
module conv_128_32 ( clk, reset, s_valid_x, s_valid_f, m_ready_y, s_data_in_x, 
        s_data_in_f, s_ready_f, s_ready_x, m_valid_y, m_data_out_y );
  input [7:0] s_data_in_x;
  input [7:0] s_data_in_f;
  output [20:0] m_data_out_y;
  input clk, reset, s_valid_x, s_valid_f, m_ready_y;
  output s_ready_f, s_ready_x, m_valid_y;
  wire   \xmem_data[127][7] , \xmem_data[127][6] , \xmem_data[127][5] ,
         \xmem_data[127][4] , \xmem_data[127][3] , \xmem_data[127][2] ,
         \xmem_data[127][1] , \xmem_data[127][0] , \xmem_data[126][7] ,
         \xmem_data[126][6] , \xmem_data[126][5] , \xmem_data[126][4] ,
         \xmem_data[126][3] , \xmem_data[126][2] , \xmem_data[126][1] ,
         \xmem_data[126][0] , \xmem_data[125][7] , \xmem_data[125][6] ,
         \xmem_data[125][5] , \xmem_data[125][4] , \xmem_data[125][3] ,
         \xmem_data[125][2] , \xmem_data[125][1] , \xmem_data[125][0] ,
         \xmem_data[124][7] , \xmem_data[124][6] , \xmem_data[124][5] ,
         \xmem_data[124][4] , \xmem_data[124][3] , \xmem_data[124][2] ,
         \xmem_data[124][1] , \xmem_data[124][0] , \xmem_data[123][7] ,
         \xmem_data[123][6] , \xmem_data[123][5] , \xmem_data[123][4] ,
         \xmem_data[123][3] , \xmem_data[123][2] , \xmem_data[123][1] ,
         \xmem_data[123][0] , \xmem_data[122][7] , \xmem_data[122][6] ,
         \xmem_data[122][5] , \xmem_data[122][4] , \xmem_data[122][3] ,
         \xmem_data[122][2] , \xmem_data[122][1] , \xmem_data[122][0] ,
         \xmem_data[121][7] , \xmem_data[121][6] , \xmem_data[121][5] ,
         \xmem_data[121][4] , \xmem_data[121][3] , \xmem_data[121][2] ,
         \xmem_data[121][1] , \xmem_data[121][0] , \xmem_data[120][7] ,
         \xmem_data[120][6] , \xmem_data[120][5] , \xmem_data[120][4] ,
         \xmem_data[120][3] , \xmem_data[120][2] , \xmem_data[120][1] ,
         \xmem_data[120][0] , \xmem_data[119][7] , \xmem_data[119][6] ,
         \xmem_data[119][5] , \xmem_data[119][4] , \xmem_data[119][3] ,
         \xmem_data[119][2] , \xmem_data[119][1] , \xmem_data[119][0] ,
         \xmem_data[118][7] , \xmem_data[118][6] , \xmem_data[118][5] ,
         \xmem_data[118][4] , \xmem_data[118][3] , \xmem_data[118][2] ,
         \xmem_data[118][1] , \xmem_data[118][0] , \xmem_data[117][7] ,
         \xmem_data[117][6] , \xmem_data[117][5] , \xmem_data[117][4] ,
         \xmem_data[117][3] , \xmem_data[117][2] , \xmem_data[117][1] ,
         \xmem_data[117][0] , \xmem_data[116][7] , \xmem_data[116][6] ,
         \xmem_data[116][5] , \xmem_data[116][4] , \xmem_data[116][3] ,
         \xmem_data[116][2] , \xmem_data[116][1] , \xmem_data[116][0] ,
         \xmem_data[115][7] , \xmem_data[115][6] , \xmem_data[115][5] ,
         \xmem_data[115][4] , \xmem_data[115][3] , \xmem_data[115][2] ,
         \xmem_data[115][1] , \xmem_data[115][0] , \xmem_data[114][7] ,
         \xmem_data[114][6] , \xmem_data[114][5] , \xmem_data[114][4] ,
         \xmem_data[114][3] , \xmem_data[114][2] , \xmem_data[114][1] ,
         \xmem_data[114][0] , \xmem_data[113][7] , \xmem_data[113][6] ,
         \xmem_data[113][5] , \xmem_data[113][4] , \xmem_data[113][3] ,
         \xmem_data[113][2] , \xmem_data[113][1] , \xmem_data[113][0] ,
         \xmem_data[112][7] , \xmem_data[112][6] , \xmem_data[112][5] ,
         \xmem_data[112][4] , \xmem_data[112][3] , \xmem_data[112][2] ,
         \xmem_data[112][1] , \xmem_data[112][0] , \xmem_data[111][7] ,
         \xmem_data[111][6] , \xmem_data[111][5] , \xmem_data[111][4] ,
         \xmem_data[111][3] , \xmem_data[111][2] , \xmem_data[111][1] ,
         \xmem_data[111][0] , \xmem_data[110][7] , \xmem_data[110][6] ,
         \xmem_data[110][5] , \xmem_data[110][4] , \xmem_data[110][3] ,
         \xmem_data[110][2] , \xmem_data[110][1] , \xmem_data[110][0] ,
         \xmem_data[109][7] , \xmem_data[109][6] , \xmem_data[109][5] ,
         \xmem_data[109][4] , \xmem_data[109][3] , \xmem_data[109][2] ,
         \xmem_data[109][1] , \xmem_data[109][0] , \xmem_data[108][7] ,
         \xmem_data[108][6] , \xmem_data[108][5] , \xmem_data[108][4] ,
         \xmem_data[108][3] , \xmem_data[108][2] , \xmem_data[108][1] ,
         \xmem_data[108][0] , \xmem_data[107][7] , \xmem_data[107][6] ,
         \xmem_data[107][5] , \xmem_data[107][4] , \xmem_data[107][3] ,
         \xmem_data[107][2] , \xmem_data[107][1] , \xmem_data[107][0] ,
         \xmem_data[106][7] , \xmem_data[106][6] , \xmem_data[106][5] ,
         \xmem_data[106][4] , \xmem_data[106][3] , \xmem_data[106][2] ,
         \xmem_data[106][1] , \xmem_data[106][0] , \xmem_data[105][7] ,
         \xmem_data[105][6] , \xmem_data[105][5] , \xmem_data[105][4] ,
         \xmem_data[105][3] , \xmem_data[105][2] , \xmem_data[105][1] ,
         \xmem_data[105][0] , \xmem_data[104][7] , \xmem_data[104][6] ,
         \xmem_data[104][5] , \xmem_data[104][4] , \xmem_data[104][3] ,
         \xmem_data[104][2] , \xmem_data[104][1] , \xmem_data[104][0] ,
         \xmem_data[103][7] , \xmem_data[103][6] , \xmem_data[103][5] ,
         \xmem_data[103][4] , \xmem_data[103][3] , \xmem_data[103][2] ,
         \xmem_data[103][1] , \xmem_data[103][0] , \xmem_data[102][7] ,
         \xmem_data[102][6] , \xmem_data[102][5] , \xmem_data[102][4] ,
         \xmem_data[102][3] , \xmem_data[102][2] , \xmem_data[102][1] ,
         \xmem_data[102][0] , \xmem_data[101][7] , \xmem_data[101][6] ,
         \xmem_data[101][5] , \xmem_data[101][4] , \xmem_data[101][3] ,
         \xmem_data[101][2] , \xmem_data[101][1] , \xmem_data[101][0] ,
         \xmem_data[100][7] , \xmem_data[100][6] , \xmem_data[100][5] ,
         \xmem_data[100][4] , \xmem_data[100][3] , \xmem_data[100][2] ,
         \xmem_data[100][1] , \xmem_data[100][0] , \xmem_data[99][7] ,
         \xmem_data[99][6] , \xmem_data[99][5] , \xmem_data[99][4] ,
         \xmem_data[99][3] , \xmem_data[99][2] , \xmem_data[99][1] ,
         \xmem_data[99][0] , \xmem_data[98][7] , \xmem_data[98][6] ,
         \xmem_data[98][5] , \xmem_data[98][4] , \xmem_data[98][3] ,
         \xmem_data[98][2] , \xmem_data[98][1] , \xmem_data[98][0] ,
         \xmem_data[97][7] , \xmem_data[97][6] , \xmem_data[97][5] ,
         \xmem_data[97][4] , \xmem_data[97][3] , \xmem_data[97][2] ,
         \xmem_data[97][1] , \xmem_data[97][0] , \xmem_data[96][7] ,
         \xmem_data[96][6] , \xmem_data[96][5] , \xmem_data[96][4] ,
         \xmem_data[96][3] , \xmem_data[96][2] , \xmem_data[96][1] ,
         \xmem_data[96][0] , \xmem_data[95][7] , \xmem_data[95][6] ,
         \xmem_data[95][5] , \xmem_data[95][4] , \xmem_data[95][3] ,
         \xmem_data[95][2] , \xmem_data[95][1] , \xmem_data[95][0] ,
         \xmem_data[94][7] , \xmem_data[94][6] , \xmem_data[94][5] ,
         \xmem_data[94][4] , \xmem_data[94][3] , \xmem_data[94][2] ,
         \xmem_data[94][1] , \xmem_data[94][0] , \xmem_data[93][7] ,
         \xmem_data[93][6] , \xmem_data[93][5] , \xmem_data[93][4] ,
         \xmem_data[93][3] , \xmem_data[93][2] , \xmem_data[93][1] ,
         \xmem_data[93][0] , \xmem_data[92][7] , \xmem_data[92][6] ,
         \xmem_data[92][5] , \xmem_data[92][4] , \xmem_data[92][3] ,
         \xmem_data[92][2] , \xmem_data[92][1] , \xmem_data[92][0] ,
         \xmem_data[91][7] , \xmem_data[91][6] , \xmem_data[91][5] ,
         \xmem_data[91][4] , \xmem_data[91][3] , \xmem_data[91][2] ,
         \xmem_data[91][1] , \xmem_data[91][0] , \xmem_data[90][7] ,
         \xmem_data[90][6] , \xmem_data[90][5] , \xmem_data[90][4] ,
         \xmem_data[90][3] , \xmem_data[90][2] , \xmem_data[90][1] ,
         \xmem_data[90][0] , \xmem_data[89][7] , \xmem_data[89][6] ,
         \xmem_data[89][5] , \xmem_data[89][4] , \xmem_data[89][3] ,
         \xmem_data[89][2] , \xmem_data[89][1] , \xmem_data[89][0] ,
         \xmem_data[88][7] , \xmem_data[88][6] , \xmem_data[88][5] ,
         \xmem_data[88][4] , \xmem_data[88][3] , \xmem_data[88][2] ,
         \xmem_data[88][1] , \xmem_data[88][0] , \xmem_data[87][7] ,
         \xmem_data[87][6] , \xmem_data[87][5] , \xmem_data[87][4] ,
         \xmem_data[87][3] , \xmem_data[87][2] , \xmem_data[87][1] ,
         \xmem_data[87][0] , \xmem_data[86][7] , \xmem_data[86][6] ,
         \xmem_data[86][5] , \xmem_data[86][4] , \xmem_data[86][3] ,
         \xmem_data[86][2] , \xmem_data[86][1] , \xmem_data[86][0] ,
         \xmem_data[85][7] , \xmem_data[85][6] , \xmem_data[85][5] ,
         \xmem_data[85][4] , \xmem_data[85][3] , \xmem_data[85][2] ,
         \xmem_data[85][1] , \xmem_data[85][0] , \xmem_data[84][7] ,
         \xmem_data[84][6] , \xmem_data[84][5] , \xmem_data[84][4] ,
         \xmem_data[84][3] , \xmem_data[84][2] , \xmem_data[84][1] ,
         \xmem_data[84][0] , \xmem_data[83][7] , \xmem_data[83][6] ,
         \xmem_data[83][5] , \xmem_data[83][4] , \xmem_data[83][3] ,
         \xmem_data[83][2] , \xmem_data[83][1] , \xmem_data[83][0] ,
         \xmem_data[82][7] , \xmem_data[82][6] , \xmem_data[82][5] ,
         \xmem_data[82][4] , \xmem_data[82][3] , \xmem_data[82][2] ,
         \xmem_data[82][1] , \xmem_data[82][0] , \xmem_data[81][7] ,
         \xmem_data[81][6] , \xmem_data[81][5] , \xmem_data[81][4] ,
         \xmem_data[81][3] , \xmem_data[81][2] , \xmem_data[81][1] ,
         \xmem_data[81][0] , \xmem_data[80][7] , \xmem_data[80][6] ,
         \xmem_data[80][5] , \xmem_data[80][4] , \xmem_data[80][3] ,
         \xmem_data[80][2] , \xmem_data[80][1] , \xmem_data[80][0] ,
         \xmem_data[79][7] , \xmem_data[79][6] , \xmem_data[79][5] ,
         \xmem_data[79][4] , \xmem_data[79][3] , \xmem_data[79][2] ,
         \xmem_data[79][1] , \xmem_data[79][0] , \xmem_data[78][7] ,
         \xmem_data[78][6] , \xmem_data[78][5] , \xmem_data[78][4] ,
         \xmem_data[78][3] , \xmem_data[78][2] , \xmem_data[78][1] ,
         \xmem_data[78][0] , \xmem_data[77][7] , \xmem_data[77][6] ,
         \xmem_data[77][5] , \xmem_data[77][4] , \xmem_data[77][3] ,
         \xmem_data[77][2] , \xmem_data[77][1] , \xmem_data[77][0] ,
         \xmem_data[76][7] , \xmem_data[76][6] , \xmem_data[76][5] ,
         \xmem_data[76][4] , \xmem_data[76][3] , \xmem_data[76][2] ,
         \xmem_data[76][1] , \xmem_data[76][0] , \xmem_data[75][7] ,
         \xmem_data[75][6] , \xmem_data[75][5] , \xmem_data[75][4] ,
         \xmem_data[75][3] , \xmem_data[75][2] , \xmem_data[75][1] ,
         \xmem_data[75][0] , \xmem_data[74][7] , \xmem_data[74][6] ,
         \xmem_data[74][5] , \xmem_data[74][4] , \xmem_data[74][3] ,
         \xmem_data[74][2] , \xmem_data[74][1] , \xmem_data[74][0] ,
         \xmem_data[73][7] , \xmem_data[73][6] , \xmem_data[73][5] ,
         \xmem_data[73][4] , \xmem_data[73][3] , \xmem_data[73][2] ,
         \xmem_data[73][1] , \xmem_data[73][0] , \xmem_data[72][7] ,
         \xmem_data[72][6] , \xmem_data[72][5] , \xmem_data[72][4] ,
         \xmem_data[72][3] , \xmem_data[72][2] , \xmem_data[72][1] ,
         \xmem_data[72][0] , \xmem_data[71][7] , \xmem_data[71][6] ,
         \xmem_data[71][5] , \xmem_data[71][4] , \xmem_data[71][3] ,
         \xmem_data[71][2] , \xmem_data[71][1] , \xmem_data[71][0] ,
         \xmem_data[70][7] , \xmem_data[70][6] , \xmem_data[70][5] ,
         \xmem_data[70][4] , \xmem_data[70][3] , \xmem_data[70][2] ,
         \xmem_data[70][1] , \xmem_data[70][0] , \xmem_data[69][7] ,
         \xmem_data[69][6] , \xmem_data[69][5] , \xmem_data[69][4] ,
         \xmem_data[69][3] , \xmem_data[69][2] , \xmem_data[69][1] ,
         \xmem_data[69][0] , \xmem_data[68][7] , \xmem_data[68][6] ,
         \xmem_data[68][5] , \xmem_data[68][4] , \xmem_data[68][3] ,
         \xmem_data[68][2] , \xmem_data[68][1] , \xmem_data[68][0] ,
         \xmem_data[67][7] , \xmem_data[67][6] , \xmem_data[67][5] ,
         \xmem_data[67][4] , \xmem_data[67][3] , \xmem_data[67][2] ,
         \xmem_data[67][1] , \xmem_data[67][0] , \xmem_data[66][7] ,
         \xmem_data[66][6] , \xmem_data[66][5] , \xmem_data[66][4] ,
         \xmem_data[66][3] , \xmem_data[66][2] , \xmem_data[66][1] ,
         \xmem_data[66][0] , \xmem_data[65][7] , \xmem_data[65][6] ,
         \xmem_data[65][5] , \xmem_data[65][4] , \xmem_data[65][3] ,
         \xmem_data[65][2] , \xmem_data[65][1] , \xmem_data[65][0] ,
         \xmem_data[64][7] , \xmem_data[64][6] , \xmem_data[64][5] ,
         \xmem_data[64][4] , \xmem_data[64][3] , \xmem_data[64][2] ,
         \xmem_data[64][1] , \xmem_data[64][0] , \xmem_data[63][7] ,
         \xmem_data[63][6] , \xmem_data[63][5] , \xmem_data[63][4] ,
         \xmem_data[63][3] , \xmem_data[63][2] , \xmem_data[63][1] ,
         \xmem_data[63][0] , \xmem_data[62][7] , \xmem_data[62][6] ,
         \xmem_data[62][5] , \xmem_data[62][4] , \xmem_data[62][3] ,
         \xmem_data[62][2] , \xmem_data[62][1] , \xmem_data[62][0] ,
         \xmem_data[61][7] , \xmem_data[61][6] , \xmem_data[61][5] ,
         \xmem_data[61][4] , \xmem_data[61][3] , \xmem_data[61][2] ,
         \xmem_data[61][1] , \xmem_data[61][0] , \xmem_data[60][7] ,
         \xmem_data[60][6] , \xmem_data[60][5] , \xmem_data[60][4] ,
         \xmem_data[60][3] , \xmem_data[60][2] , \xmem_data[60][1] ,
         \xmem_data[60][0] , \xmem_data[59][7] , \xmem_data[59][6] ,
         \xmem_data[59][5] , \xmem_data[59][4] , \xmem_data[59][3] ,
         \xmem_data[59][2] , \xmem_data[59][1] , \xmem_data[59][0] ,
         \xmem_data[58][7] , \xmem_data[58][6] , \xmem_data[58][5] ,
         \xmem_data[58][4] , \xmem_data[58][3] , \xmem_data[58][2] ,
         \xmem_data[58][1] , \xmem_data[58][0] , \xmem_data[57][7] ,
         \xmem_data[57][6] , \xmem_data[57][5] , \xmem_data[57][4] ,
         \xmem_data[57][3] , \xmem_data[57][2] , \xmem_data[57][1] ,
         \xmem_data[57][0] , \xmem_data[56][7] , \xmem_data[56][6] ,
         \xmem_data[56][5] , \xmem_data[56][4] , \xmem_data[56][3] ,
         \xmem_data[56][2] , \xmem_data[56][1] , \xmem_data[56][0] ,
         \xmem_data[55][7] , \xmem_data[55][6] , \xmem_data[55][5] ,
         \xmem_data[55][4] , \xmem_data[55][3] , \xmem_data[55][2] ,
         \xmem_data[55][1] , \xmem_data[55][0] , \xmem_data[54][7] ,
         \xmem_data[54][6] , \xmem_data[54][5] , \xmem_data[54][4] ,
         \xmem_data[54][3] , \xmem_data[54][2] , \xmem_data[54][1] ,
         \xmem_data[54][0] , \xmem_data[53][7] , \xmem_data[53][6] ,
         \xmem_data[53][5] , \xmem_data[53][4] , \xmem_data[53][3] ,
         \xmem_data[53][2] , \xmem_data[53][1] , \xmem_data[53][0] ,
         \xmem_data[52][7] , \xmem_data[52][6] , \xmem_data[52][5] ,
         \xmem_data[52][4] , \xmem_data[52][3] , \xmem_data[52][2] ,
         \xmem_data[52][1] , \xmem_data[52][0] , \xmem_data[51][7] ,
         \xmem_data[51][6] , \xmem_data[51][5] , \xmem_data[51][4] ,
         \xmem_data[51][3] , \xmem_data[51][2] , \xmem_data[51][1] ,
         \xmem_data[51][0] , \xmem_data[50][7] , \xmem_data[50][6] ,
         \xmem_data[50][5] , \xmem_data[50][4] , \xmem_data[50][3] ,
         \xmem_data[50][2] , \xmem_data[50][1] , \xmem_data[50][0] ,
         \xmem_data[49][7] , \xmem_data[49][6] , \xmem_data[49][5] ,
         \xmem_data[49][4] , \xmem_data[49][3] , \xmem_data[49][2] ,
         \xmem_data[49][1] , \xmem_data[49][0] , \xmem_data[48][7] ,
         \xmem_data[48][6] , \xmem_data[48][5] , \xmem_data[48][4] ,
         \xmem_data[48][3] , \xmem_data[48][2] , \xmem_data[48][1] ,
         \xmem_data[48][0] , \xmem_data[47][7] , \xmem_data[47][6] ,
         \xmem_data[47][5] , \xmem_data[47][4] , \xmem_data[47][3] ,
         \xmem_data[47][2] , \xmem_data[47][1] , \xmem_data[47][0] ,
         \xmem_data[46][7] , \xmem_data[46][6] , \xmem_data[46][5] ,
         \xmem_data[46][4] , \xmem_data[46][3] , \xmem_data[46][2] ,
         \xmem_data[46][1] , \xmem_data[46][0] , \xmem_data[45][7] ,
         \xmem_data[45][6] , \xmem_data[45][5] , \xmem_data[45][4] ,
         \xmem_data[45][3] , \xmem_data[45][2] , \xmem_data[45][1] ,
         \xmem_data[45][0] , \xmem_data[44][7] , \xmem_data[44][6] ,
         \xmem_data[44][5] , \xmem_data[44][4] , \xmem_data[44][3] ,
         \xmem_data[44][2] , \xmem_data[44][1] , \xmem_data[44][0] ,
         \xmem_data[43][7] , \xmem_data[43][6] , \xmem_data[43][5] ,
         \xmem_data[43][4] , \xmem_data[43][3] , \xmem_data[43][2] ,
         \xmem_data[43][1] , \xmem_data[43][0] , \xmem_data[42][7] ,
         \xmem_data[42][6] , \xmem_data[42][5] , \xmem_data[42][4] ,
         \xmem_data[42][3] , \xmem_data[42][2] , \xmem_data[42][1] ,
         \xmem_data[42][0] , \xmem_data[41][7] , \xmem_data[41][6] ,
         \xmem_data[41][5] , \xmem_data[41][4] , \xmem_data[41][3] ,
         \xmem_data[41][2] , \xmem_data[41][1] , \xmem_data[41][0] ,
         \xmem_data[40][7] , \xmem_data[40][6] , \xmem_data[40][5] ,
         \xmem_data[40][4] , \xmem_data[40][3] , \xmem_data[40][2] ,
         \xmem_data[40][1] , \xmem_data[40][0] , \xmem_data[39][7] ,
         \xmem_data[39][6] , \xmem_data[39][5] , \xmem_data[39][4] ,
         \xmem_data[39][3] , \xmem_data[39][2] , \xmem_data[39][1] ,
         \xmem_data[39][0] , \xmem_data[38][7] , \xmem_data[38][6] ,
         \xmem_data[38][5] , \xmem_data[38][4] , \xmem_data[38][3] ,
         \xmem_data[38][2] , \xmem_data[38][1] , \xmem_data[38][0] ,
         \xmem_data[37][7] , \xmem_data[37][6] , \xmem_data[37][5] ,
         \xmem_data[37][4] , \xmem_data[37][3] , \xmem_data[37][2] ,
         \xmem_data[37][1] , \xmem_data[37][0] , \xmem_data[36][7] ,
         \xmem_data[36][6] , \xmem_data[36][5] , \xmem_data[36][4] ,
         \xmem_data[36][3] , \xmem_data[36][2] , \xmem_data[36][1] ,
         \xmem_data[36][0] , \xmem_data[35][7] , \xmem_data[35][6] ,
         \xmem_data[35][5] , \xmem_data[35][4] , \xmem_data[35][3] ,
         \xmem_data[35][2] , \xmem_data[35][1] , \xmem_data[35][0] ,
         \xmem_data[34][7] , \xmem_data[34][6] , \xmem_data[34][5] ,
         \xmem_data[34][4] , \xmem_data[34][3] , \xmem_data[34][2] ,
         \xmem_data[34][1] , \xmem_data[34][0] , \xmem_data[33][7] ,
         \xmem_data[33][6] , \xmem_data[33][5] , \xmem_data[33][4] ,
         \xmem_data[33][3] , \xmem_data[33][2] , \xmem_data[33][1] ,
         \xmem_data[33][0] , \xmem_data[32][7] , \xmem_data[32][6] ,
         \xmem_data[32][5] , \xmem_data[32][4] , \xmem_data[32][3] ,
         \xmem_data[32][2] , \xmem_data[32][1] , \xmem_data[32][0] ,
         \xmem_data[31][7] , \xmem_data[31][6] , \xmem_data[31][5] ,
         \xmem_data[31][4] , \xmem_data[31][3] , \xmem_data[31][2] ,
         \xmem_data[31][1] , \xmem_data[31][0] , \xmem_data[30][7] ,
         \xmem_data[30][6] , \xmem_data[30][5] , \xmem_data[30][4] ,
         \xmem_data[30][3] , \xmem_data[30][2] , \xmem_data[30][1] ,
         \xmem_data[30][0] , \xmem_data[29][7] , \xmem_data[29][6] ,
         \xmem_data[29][5] , \xmem_data[29][4] , \xmem_data[29][3] ,
         \xmem_data[29][2] , \xmem_data[29][1] , \xmem_data[29][0] ,
         \xmem_data[28][7] , \xmem_data[28][6] , \xmem_data[28][5] ,
         \xmem_data[28][4] , \xmem_data[28][3] , \xmem_data[28][2] ,
         \xmem_data[28][1] , \xmem_data[28][0] , \xmem_data[27][7] ,
         \xmem_data[27][6] , \xmem_data[27][5] , \xmem_data[27][4] ,
         \xmem_data[27][3] , \xmem_data[27][2] , \xmem_data[27][1] ,
         \xmem_data[27][0] , \xmem_data[26][7] , \xmem_data[26][6] ,
         \xmem_data[26][5] , \xmem_data[26][4] , \xmem_data[26][3] ,
         \xmem_data[26][2] , \xmem_data[26][1] , \xmem_data[26][0] ,
         \xmem_data[25][7] , \xmem_data[25][6] , \xmem_data[25][5] ,
         \xmem_data[25][4] , \xmem_data[25][3] , \xmem_data[25][2] ,
         \xmem_data[25][1] , \xmem_data[25][0] , \xmem_data[24][7] ,
         \xmem_data[24][6] , \xmem_data[24][5] , \xmem_data[24][4] ,
         \xmem_data[24][3] , \xmem_data[24][2] , \xmem_data[24][1] ,
         \xmem_data[24][0] , \xmem_data[23][7] , \xmem_data[23][6] ,
         \xmem_data[23][5] , \xmem_data[23][4] , \xmem_data[23][3] ,
         \xmem_data[23][2] , \xmem_data[23][1] , \xmem_data[23][0] ,
         \xmem_data[22][7] , \xmem_data[22][6] , \xmem_data[22][5] ,
         \xmem_data[22][4] , \xmem_data[22][3] , \xmem_data[22][2] ,
         \xmem_data[22][1] , \xmem_data[22][0] , \xmem_data[21][7] ,
         \xmem_data[21][6] , \xmem_data[21][5] , \xmem_data[21][4] ,
         \xmem_data[21][3] , \xmem_data[21][2] , \xmem_data[21][1] ,
         \xmem_data[21][0] , \xmem_data[20][7] , \xmem_data[20][6] ,
         \xmem_data[20][5] , \xmem_data[20][4] , \xmem_data[20][3] ,
         \xmem_data[20][2] , \xmem_data[20][1] , \xmem_data[20][0] ,
         \xmem_data[19][7] , \xmem_data[19][6] , \xmem_data[19][5] ,
         \xmem_data[19][4] , \xmem_data[19][3] , \xmem_data[19][2] ,
         \xmem_data[19][1] , \xmem_data[19][0] , \xmem_data[18][7] ,
         \xmem_data[18][6] , \xmem_data[18][5] , \xmem_data[18][4] ,
         \xmem_data[18][3] , \xmem_data[18][2] , \xmem_data[18][1] ,
         \xmem_data[18][0] , \xmem_data[17][7] , \xmem_data[17][6] ,
         \xmem_data[17][5] , \xmem_data[17][4] , \xmem_data[17][3] ,
         \xmem_data[17][2] , \xmem_data[17][1] , \xmem_data[17][0] ,
         \xmem_data[16][7] , \xmem_data[16][6] , \xmem_data[16][5] ,
         \xmem_data[16][4] , \xmem_data[16][3] , \xmem_data[16][2] ,
         \xmem_data[16][1] , \xmem_data[16][0] , \xmem_data[15][7] ,
         \xmem_data[15][6] , \xmem_data[15][5] , \xmem_data[15][4] ,
         \xmem_data[15][3] , \xmem_data[15][2] , \xmem_data[15][1] ,
         \xmem_data[15][0] , \xmem_data[14][7] , \xmem_data[14][6] ,
         \xmem_data[14][5] , \xmem_data[14][4] , \xmem_data[14][3] ,
         \xmem_data[14][2] , \xmem_data[14][1] , \xmem_data[14][0] ,
         \xmem_data[13][7] , \xmem_data[13][6] , \xmem_data[13][5] ,
         \xmem_data[13][4] , \xmem_data[13][3] , \xmem_data[13][2] ,
         \xmem_data[13][1] , \xmem_data[13][0] , \xmem_data[12][7] ,
         \xmem_data[12][6] , \xmem_data[12][5] , \xmem_data[12][4] ,
         \xmem_data[12][3] , \xmem_data[12][2] , \xmem_data[12][1] ,
         \xmem_data[12][0] , \xmem_data[11][7] , \xmem_data[11][6] ,
         \xmem_data[11][5] , \xmem_data[11][4] , \xmem_data[11][3] ,
         \xmem_data[11][2] , \xmem_data[11][1] , \xmem_data[11][0] ,
         \xmem_data[10][7] , \xmem_data[10][6] , \xmem_data[10][5] ,
         \xmem_data[10][4] , \xmem_data[10][3] , \xmem_data[10][2] ,
         \xmem_data[10][1] , \xmem_data[10][0] , \xmem_data[9][7] ,
         \xmem_data[9][6] , \xmem_data[9][5] , \xmem_data[9][4] ,
         \xmem_data[9][3] , \xmem_data[9][2] , \xmem_data[9][1] ,
         \xmem_data[9][0] , \xmem_data[8][7] , \xmem_data[8][6] ,
         \xmem_data[8][5] , \xmem_data[8][4] , \xmem_data[8][3] ,
         \xmem_data[8][2] , \xmem_data[8][1] , \xmem_data[8][0] ,
         \xmem_data[7][7] , \xmem_data[7][6] , \xmem_data[7][5] ,
         \xmem_data[7][4] , \xmem_data[7][3] , \xmem_data[7][2] ,
         \xmem_data[7][1] , \xmem_data[7][0] , \xmem_data[6][7] ,
         \xmem_data[6][6] , \xmem_data[6][5] , \xmem_data[6][4] ,
         \xmem_data[6][3] , \xmem_data[6][2] , \xmem_data[6][1] ,
         \xmem_data[6][0] , \xmem_data[5][7] , \xmem_data[5][6] ,
         \xmem_data[5][5] , \xmem_data[5][4] , \xmem_data[5][3] ,
         \xmem_data[5][2] , \xmem_data[5][1] , \xmem_data[5][0] ,
         \xmem_data[4][7] , \xmem_data[4][6] , \xmem_data[4][5] ,
         \xmem_data[4][4] , \xmem_data[4][3] , \xmem_data[4][2] ,
         \xmem_data[4][1] , \xmem_data[4][0] , \xmem_data[3][7] ,
         \xmem_data[3][6] , \xmem_data[3][5] , \xmem_data[3][4] ,
         \xmem_data[3][3] , \xmem_data[3][2] , \xmem_data[3][1] ,
         \xmem_data[3][0] , \xmem_data[2][7] , \xmem_data[2][6] ,
         \xmem_data[2][5] , \xmem_data[2][4] , \xmem_data[2][3] ,
         \xmem_data[2][2] , \xmem_data[2][1] , \xmem_data[2][0] ,
         \xmem_data[1][7] , \xmem_data[1][6] , \xmem_data[1][5] ,
         \xmem_data[1][4] , \xmem_data[1][3] , \xmem_data[1][2] ,
         \xmem_data[1][1] , \xmem_data[1][0] , \xmem_data[0][7] ,
         \xmem_data[0][6] , \xmem_data[0][5] , \xmem_data[0][4] ,
         \xmem_data[0][3] , \xmem_data[0][2] , \xmem_data[0][1] ,
         \xmem_data[0][0] , \fmem_data[31][7] , \fmem_data[31][6] ,
         \fmem_data[31][5] , \fmem_data[31][4] , \fmem_data[31][3] ,
         \fmem_data[31][2] , \fmem_data[31][1] , \fmem_data[30][7] ,
         \fmem_data[30][6] , \fmem_data[30][5] , \fmem_data[30][4] ,
         \fmem_data[30][3] , \fmem_data[30][2] , \fmem_data[30][1] ,
         \fmem_data[30][0] , \fmem_data[29][7] , \fmem_data[29][6] ,
         \fmem_data[29][5] , \fmem_data[29][4] , \fmem_data[29][3] ,
         \fmem_data[29][2] , \fmem_data[29][1] , \fmem_data[29][0] ,
         \fmem_data[28][7] , \fmem_data[28][6] , \fmem_data[28][5] ,
         \fmem_data[28][4] , \fmem_data[28][3] , \fmem_data[28][2] ,
         \fmem_data[28][1] , \fmem_data[28][0] , \fmem_data[27][7] ,
         \fmem_data[27][6] , \fmem_data[27][5] , \fmem_data[27][4] ,
         \fmem_data[27][3] , \fmem_data[27][2] , \fmem_data[27][1] ,
         \fmem_data[27][0] , \fmem_data[26][7] , \fmem_data[26][6] ,
         \fmem_data[26][5] , \fmem_data[26][4] , \fmem_data[26][3] ,
         \fmem_data[26][2] , \fmem_data[26][1] , \fmem_data[26][0] ,
         \fmem_data[25][7] , \fmem_data[25][6] , \fmem_data[25][5] ,
         \fmem_data[25][4] , \fmem_data[25][3] , \fmem_data[25][2] ,
         \fmem_data[25][1] , \fmem_data[25][0] , \fmem_data[24][7] ,
         \fmem_data[24][6] , \fmem_data[24][5] , \fmem_data[24][4] ,
         \fmem_data[24][3] , \fmem_data[24][2] , \fmem_data[24][1] ,
         \fmem_data[24][0] , \fmem_data[23][7] , \fmem_data[23][6] ,
         \fmem_data[23][5] , \fmem_data[23][4] , \fmem_data[23][3] ,
         \fmem_data[23][2] , \fmem_data[23][1] , \fmem_data[23][0] ,
         \fmem_data[22][7] , \fmem_data[22][6] , \fmem_data[22][5] ,
         \fmem_data[22][4] , \fmem_data[22][3] , \fmem_data[22][2] ,
         \fmem_data[22][1] , \fmem_data[22][0] , \fmem_data[21][7] ,
         \fmem_data[21][6] , \fmem_data[21][5] , \fmem_data[21][4] ,
         \fmem_data[21][3] , \fmem_data[21][2] , \fmem_data[21][1] ,
         \fmem_data[21][0] , \fmem_data[20][7] , \fmem_data[20][6] ,
         \fmem_data[20][5] , \fmem_data[20][4] , \fmem_data[20][3] ,
         \fmem_data[20][2] , \fmem_data[20][1] , \fmem_data[20][0] ,
         \fmem_data[19][7] , \fmem_data[19][6] , \fmem_data[19][5] ,
         \fmem_data[19][4] , \fmem_data[19][3] , \fmem_data[19][2] ,
         \fmem_data[19][1] , \fmem_data[19][0] , \fmem_data[18][7] ,
         \fmem_data[18][6] , \fmem_data[18][5] , \fmem_data[18][4] ,
         \fmem_data[18][3] , \fmem_data[18][2] , \fmem_data[18][1] ,
         \fmem_data[18][0] , \fmem_data[17][7] , \fmem_data[17][6] ,
         \fmem_data[17][5] , \fmem_data[17][4] , \fmem_data[17][3] ,
         \fmem_data[17][2] , \fmem_data[17][1] , \fmem_data[17][0] ,
         \fmem_data[16][7] , \fmem_data[16][6] , \fmem_data[16][5] ,
         \fmem_data[16][4] , \fmem_data[16][3] , \fmem_data[16][2] ,
         \fmem_data[16][1] , \fmem_data[16][0] , \fmem_data[15][7] ,
         \fmem_data[15][6] , \fmem_data[15][5] , \fmem_data[15][4] ,
         \fmem_data[15][3] , \fmem_data[15][2] , \fmem_data[15][1] ,
         \fmem_data[15][0] , \fmem_data[14][7] , \fmem_data[14][6] ,
         \fmem_data[14][5] , \fmem_data[14][4] , \fmem_data[14][3] ,
         \fmem_data[14][2] , \fmem_data[14][1] , \fmem_data[14][0] ,
         \fmem_data[13][7] , \fmem_data[13][6] , \fmem_data[13][5] ,
         \fmem_data[13][4] , \fmem_data[13][3] , \fmem_data[13][2] ,
         \fmem_data[13][1] , \fmem_data[13][0] , \fmem_data[12][7] ,
         \fmem_data[12][6] , \fmem_data[12][5] , \fmem_data[12][4] ,
         \fmem_data[12][3] , \fmem_data[12][2] , \fmem_data[12][1] ,
         \fmem_data[12][0] , \fmem_data[11][7] , \fmem_data[11][6] ,
         \fmem_data[11][5] , \fmem_data[11][4] , \fmem_data[11][3] ,
         \fmem_data[11][2] , \fmem_data[11][1] , \fmem_data[11][0] ,
         \fmem_data[10][7] , \fmem_data[10][6] , \fmem_data[10][5] ,
         \fmem_data[10][4] , \fmem_data[10][3] , \fmem_data[10][2] ,
         \fmem_data[10][1] , \fmem_data[10][0] , \fmem_data[9][7] ,
         \fmem_data[9][6] , \fmem_data[9][5] , \fmem_data[9][4] ,
         \fmem_data[9][3] , \fmem_data[9][2] , \fmem_data[9][1] ,
         \fmem_data[9][0] , \fmem_data[8][7] , \fmem_data[8][6] ,
         \fmem_data[8][5] , \fmem_data[8][4] , \fmem_data[8][3] ,
         \fmem_data[8][2] , \fmem_data[8][1] , \fmem_data[8][0] ,
         \fmem_data[7][7] , \fmem_data[7][6] , \fmem_data[7][5] ,
         \fmem_data[7][4] , \fmem_data[7][3] , \fmem_data[7][2] ,
         \fmem_data[7][1] , \fmem_data[7][0] , \fmem_data[6][7] ,
         \fmem_data[6][6] , \fmem_data[6][5] , \fmem_data[6][4] ,
         \fmem_data[6][3] , \fmem_data[6][2] , \fmem_data[6][1] ,
         \fmem_data[6][0] , \fmem_data[5][7] , \fmem_data[5][6] ,
         \fmem_data[5][5] , \fmem_data[5][4] , \fmem_data[5][3] ,
         \fmem_data[5][2] , \fmem_data[5][1] , \fmem_data[5][0] ,
         \fmem_data[4][7] , \fmem_data[4][6] , \fmem_data[4][5] ,
         \fmem_data[4][4] , \fmem_data[4][3] , \fmem_data[4][2] ,
         \fmem_data[4][1] , \fmem_data[4][0] , \fmem_data[3][7] ,
         \fmem_data[3][6] , \fmem_data[3][5] , \fmem_data[3][4] ,
         \fmem_data[3][3] , \fmem_data[3][2] , \fmem_data[3][1] ,
         \fmem_data[3][0] , \fmem_data[2][7] , \fmem_data[2][6] ,
         \fmem_data[2][5] , \fmem_data[2][4] , \fmem_data[2][3] ,
         \fmem_data[2][2] , \fmem_data[2][1] , \fmem_data[2][0] ,
         \fmem_data[1][7] , \fmem_data[1][6] , \fmem_data[1][5] ,
         \fmem_data[1][4] , \fmem_data[1][3] , \fmem_data[1][2] ,
         \fmem_data[1][1] , \fmem_data[1][0] , \fmem_data[0][7] ,
         \fmem_data[0][6] , \fmem_data[0][5] , \fmem_data[0][4] ,
         \fmem_data[0][3] , \fmem_data[0][2] , \fmem_data[0][1] ,
         \fmem_data[0][0] , conv_pre_start, N229, N284, N345, N466,
         \xmem_inst/mem[127][7] , \xmem_inst/mem[127][6] ,
         \xmem_inst/mem[127][5] , \xmem_inst/mem[127][4] ,
         \xmem_inst/mem[127][3] , \xmem_inst/mem[127][2] ,
         \xmem_inst/mem[127][1] , \xmem_inst/mem[127][0] ,
         \xmem_inst/mem[126][7] , \xmem_inst/mem[126][6] ,
         \xmem_inst/mem[126][5] , \xmem_inst/mem[126][4] ,
         \xmem_inst/mem[126][3] , \xmem_inst/mem[126][2] ,
         \xmem_inst/mem[126][1] , \xmem_inst/mem[126][0] ,
         \xmem_inst/mem[125][7] , \xmem_inst/mem[125][6] ,
         \xmem_inst/mem[125][5] , \xmem_inst/mem[125][4] ,
         \xmem_inst/mem[125][3] , \xmem_inst/mem[125][2] ,
         \xmem_inst/mem[125][1] , \xmem_inst/mem[125][0] ,
         \xmem_inst/mem[124][7] , \xmem_inst/mem[124][6] ,
         \xmem_inst/mem[124][5] , \xmem_inst/mem[124][4] ,
         \xmem_inst/mem[124][3] , \xmem_inst/mem[124][2] ,
         \xmem_inst/mem[124][1] , \xmem_inst/mem[124][0] ,
         \xmem_inst/mem[123][7] , \xmem_inst/mem[123][6] ,
         \xmem_inst/mem[123][5] , \xmem_inst/mem[123][4] ,
         \xmem_inst/mem[123][3] , \xmem_inst/mem[123][2] ,
         \xmem_inst/mem[123][1] , \xmem_inst/mem[123][0] ,
         \xmem_inst/mem[122][7] , \xmem_inst/mem[122][6] ,
         \xmem_inst/mem[122][5] , \xmem_inst/mem[122][4] ,
         \xmem_inst/mem[122][3] , \xmem_inst/mem[122][2] ,
         \xmem_inst/mem[122][1] , \xmem_inst/mem[122][0] ,
         \xmem_inst/mem[121][7] , \xmem_inst/mem[121][6] ,
         \xmem_inst/mem[121][5] , \xmem_inst/mem[121][4] ,
         \xmem_inst/mem[121][3] , \xmem_inst/mem[121][2] ,
         \xmem_inst/mem[121][1] , \xmem_inst/mem[121][0] ,
         \xmem_inst/mem[120][7] , \xmem_inst/mem[120][6] ,
         \xmem_inst/mem[120][5] , \xmem_inst/mem[120][4] ,
         \xmem_inst/mem[120][3] , \xmem_inst/mem[120][2] ,
         \xmem_inst/mem[120][1] , \xmem_inst/mem[120][0] ,
         \xmem_inst/mem[119][7] , \xmem_inst/mem[119][6] ,
         \xmem_inst/mem[119][5] , \xmem_inst/mem[119][4] ,
         \xmem_inst/mem[119][3] , \xmem_inst/mem[119][2] ,
         \xmem_inst/mem[119][1] , \xmem_inst/mem[119][0] ,
         \xmem_inst/mem[118][7] , \xmem_inst/mem[118][6] ,
         \xmem_inst/mem[118][5] , \xmem_inst/mem[118][4] ,
         \xmem_inst/mem[118][3] , \xmem_inst/mem[118][2] ,
         \xmem_inst/mem[118][1] , \xmem_inst/mem[118][0] ,
         \xmem_inst/mem[117][7] , \xmem_inst/mem[117][6] ,
         \xmem_inst/mem[117][5] , \xmem_inst/mem[117][4] ,
         \xmem_inst/mem[117][3] , \xmem_inst/mem[117][2] ,
         \xmem_inst/mem[117][1] , \xmem_inst/mem[117][0] ,
         \xmem_inst/mem[116][7] , \xmem_inst/mem[116][6] ,
         \xmem_inst/mem[116][5] , \xmem_inst/mem[116][4] ,
         \xmem_inst/mem[116][3] , \xmem_inst/mem[116][2] ,
         \xmem_inst/mem[116][1] , \xmem_inst/mem[116][0] ,
         \xmem_inst/mem[115][7] , \xmem_inst/mem[115][6] ,
         \xmem_inst/mem[115][5] , \xmem_inst/mem[115][4] ,
         \xmem_inst/mem[115][3] , \xmem_inst/mem[115][2] ,
         \xmem_inst/mem[115][1] , \xmem_inst/mem[115][0] ,
         \xmem_inst/mem[114][7] , \xmem_inst/mem[114][6] ,
         \xmem_inst/mem[114][5] , \xmem_inst/mem[114][4] ,
         \xmem_inst/mem[114][3] , \xmem_inst/mem[114][2] ,
         \xmem_inst/mem[114][1] , \xmem_inst/mem[114][0] ,
         \xmem_inst/mem[113][7] , \xmem_inst/mem[113][6] ,
         \xmem_inst/mem[113][5] , \xmem_inst/mem[113][4] ,
         \xmem_inst/mem[113][3] , \xmem_inst/mem[113][2] ,
         \xmem_inst/mem[113][1] , \xmem_inst/mem[113][0] ,
         \xmem_inst/mem[112][7] , \xmem_inst/mem[112][6] ,
         \xmem_inst/mem[112][5] , \xmem_inst/mem[112][4] ,
         \xmem_inst/mem[112][3] , \xmem_inst/mem[112][2] ,
         \xmem_inst/mem[112][1] , \xmem_inst/mem[112][0] ,
         \xmem_inst/mem[111][7] , \xmem_inst/mem[111][6] ,
         \xmem_inst/mem[111][5] , \xmem_inst/mem[111][4] ,
         \xmem_inst/mem[111][3] , \xmem_inst/mem[111][2] ,
         \xmem_inst/mem[111][1] , \xmem_inst/mem[111][0] ,
         \xmem_inst/mem[110][7] , \xmem_inst/mem[110][6] ,
         \xmem_inst/mem[110][5] , \xmem_inst/mem[110][4] ,
         \xmem_inst/mem[110][3] , \xmem_inst/mem[110][2] ,
         \xmem_inst/mem[110][1] , \xmem_inst/mem[110][0] ,
         \xmem_inst/mem[109][7] , \xmem_inst/mem[109][6] ,
         \xmem_inst/mem[109][5] , \xmem_inst/mem[109][4] ,
         \xmem_inst/mem[109][3] , \xmem_inst/mem[109][2] ,
         \xmem_inst/mem[109][1] , \xmem_inst/mem[109][0] ,
         \xmem_inst/mem[108][7] , \xmem_inst/mem[108][6] ,
         \xmem_inst/mem[108][5] , \xmem_inst/mem[108][4] ,
         \xmem_inst/mem[108][3] , \xmem_inst/mem[108][2] ,
         \xmem_inst/mem[108][1] , \xmem_inst/mem[108][0] ,
         \xmem_inst/mem[107][7] , \xmem_inst/mem[107][6] ,
         \xmem_inst/mem[107][5] , \xmem_inst/mem[107][4] ,
         \xmem_inst/mem[107][3] , \xmem_inst/mem[107][2] ,
         \xmem_inst/mem[107][1] , \xmem_inst/mem[107][0] ,
         \xmem_inst/mem[106][7] , \xmem_inst/mem[106][6] ,
         \xmem_inst/mem[106][5] , \xmem_inst/mem[106][4] ,
         \xmem_inst/mem[106][3] , \xmem_inst/mem[106][2] ,
         \xmem_inst/mem[106][1] , \xmem_inst/mem[106][0] ,
         \xmem_inst/mem[105][7] , \xmem_inst/mem[105][6] ,
         \xmem_inst/mem[105][5] , \xmem_inst/mem[105][4] ,
         \xmem_inst/mem[105][3] , \xmem_inst/mem[105][2] ,
         \xmem_inst/mem[105][1] , \xmem_inst/mem[105][0] ,
         \xmem_inst/mem[104][7] , \xmem_inst/mem[104][6] ,
         \xmem_inst/mem[104][5] , \xmem_inst/mem[104][4] ,
         \xmem_inst/mem[104][3] , \xmem_inst/mem[104][2] ,
         \xmem_inst/mem[104][1] , \xmem_inst/mem[104][0] ,
         \xmem_inst/mem[103][7] , \xmem_inst/mem[103][6] ,
         \xmem_inst/mem[103][5] , \xmem_inst/mem[103][4] ,
         \xmem_inst/mem[103][3] , \xmem_inst/mem[103][2] ,
         \xmem_inst/mem[103][1] , \xmem_inst/mem[103][0] ,
         \xmem_inst/mem[102][7] , \xmem_inst/mem[102][6] ,
         \xmem_inst/mem[102][5] , \xmem_inst/mem[102][4] ,
         \xmem_inst/mem[102][3] , \xmem_inst/mem[102][2] ,
         \xmem_inst/mem[102][1] , \xmem_inst/mem[102][0] ,
         \xmem_inst/mem[101][7] , \xmem_inst/mem[101][6] ,
         \xmem_inst/mem[101][5] , \xmem_inst/mem[101][4] ,
         \xmem_inst/mem[101][3] , \xmem_inst/mem[101][2] ,
         \xmem_inst/mem[101][1] , \xmem_inst/mem[101][0] ,
         \xmem_inst/mem[100][7] , \xmem_inst/mem[100][6] ,
         \xmem_inst/mem[100][5] , \xmem_inst/mem[100][4] ,
         \xmem_inst/mem[100][3] , \xmem_inst/mem[100][2] ,
         \xmem_inst/mem[100][1] , \xmem_inst/mem[100][0] ,
         \xmem_inst/mem[99][7] , \xmem_inst/mem[99][6] ,
         \xmem_inst/mem[99][5] , \xmem_inst/mem[99][4] ,
         \xmem_inst/mem[99][3] , \xmem_inst/mem[99][2] ,
         \xmem_inst/mem[99][1] , \xmem_inst/mem[99][0] ,
         \xmem_inst/mem[98][7] , \xmem_inst/mem[98][6] ,
         \xmem_inst/mem[98][5] , \xmem_inst/mem[98][4] ,
         \xmem_inst/mem[98][3] , \xmem_inst/mem[98][2] ,
         \xmem_inst/mem[98][1] , \xmem_inst/mem[98][0] ,
         \xmem_inst/mem[97][7] , \xmem_inst/mem[97][6] ,
         \xmem_inst/mem[97][5] , \xmem_inst/mem[97][4] ,
         \xmem_inst/mem[97][3] , \xmem_inst/mem[97][2] ,
         \xmem_inst/mem[97][1] , \xmem_inst/mem[97][0] ,
         \xmem_inst/mem[96][7] , \xmem_inst/mem[96][6] ,
         \xmem_inst/mem[96][5] , \xmem_inst/mem[96][4] ,
         \xmem_inst/mem[96][3] , \xmem_inst/mem[96][2] ,
         \xmem_inst/mem[96][1] , \xmem_inst/mem[96][0] ,
         \xmem_inst/mem[95][7] , \xmem_inst/mem[95][6] ,
         \xmem_inst/mem[95][5] , \xmem_inst/mem[95][4] ,
         \xmem_inst/mem[95][3] , \xmem_inst/mem[95][2] ,
         \xmem_inst/mem[95][1] , \xmem_inst/mem[95][0] ,
         \xmem_inst/mem[94][7] , \xmem_inst/mem[94][6] ,
         \xmem_inst/mem[94][5] , \xmem_inst/mem[94][4] ,
         \xmem_inst/mem[94][3] , \xmem_inst/mem[94][2] ,
         \xmem_inst/mem[94][1] , \xmem_inst/mem[94][0] ,
         \xmem_inst/mem[93][7] , \xmem_inst/mem[93][6] ,
         \xmem_inst/mem[93][5] , \xmem_inst/mem[93][4] ,
         \xmem_inst/mem[93][3] , \xmem_inst/mem[93][2] ,
         \xmem_inst/mem[93][1] , \xmem_inst/mem[93][0] ,
         \xmem_inst/mem[92][7] , \xmem_inst/mem[92][6] ,
         \xmem_inst/mem[92][5] , \xmem_inst/mem[92][4] ,
         \xmem_inst/mem[92][3] , \xmem_inst/mem[92][2] ,
         \xmem_inst/mem[92][1] , \xmem_inst/mem[92][0] ,
         \xmem_inst/mem[91][7] , \xmem_inst/mem[91][6] ,
         \xmem_inst/mem[91][5] , \xmem_inst/mem[91][4] ,
         \xmem_inst/mem[91][3] , \xmem_inst/mem[91][2] ,
         \xmem_inst/mem[91][1] , \xmem_inst/mem[91][0] ,
         \xmem_inst/mem[90][7] , \xmem_inst/mem[90][6] ,
         \xmem_inst/mem[90][5] , \xmem_inst/mem[90][4] ,
         \xmem_inst/mem[90][3] , \xmem_inst/mem[90][2] ,
         \xmem_inst/mem[90][1] , \xmem_inst/mem[90][0] ,
         \xmem_inst/mem[89][7] , \xmem_inst/mem[89][6] ,
         \xmem_inst/mem[89][5] , \xmem_inst/mem[89][4] ,
         \xmem_inst/mem[89][3] , \xmem_inst/mem[89][2] ,
         \xmem_inst/mem[89][1] , \xmem_inst/mem[89][0] ,
         \xmem_inst/mem[88][7] , \xmem_inst/mem[88][6] ,
         \xmem_inst/mem[88][5] , \xmem_inst/mem[88][4] ,
         \xmem_inst/mem[88][3] , \xmem_inst/mem[88][2] ,
         \xmem_inst/mem[88][1] , \xmem_inst/mem[88][0] ,
         \xmem_inst/mem[87][7] , \xmem_inst/mem[87][6] ,
         \xmem_inst/mem[87][5] , \xmem_inst/mem[87][4] ,
         \xmem_inst/mem[87][3] , \xmem_inst/mem[87][2] ,
         \xmem_inst/mem[87][1] , \xmem_inst/mem[87][0] ,
         \xmem_inst/mem[86][7] , \xmem_inst/mem[86][6] ,
         \xmem_inst/mem[86][5] , \xmem_inst/mem[86][4] ,
         \xmem_inst/mem[86][3] , \xmem_inst/mem[86][2] ,
         \xmem_inst/mem[86][1] , \xmem_inst/mem[86][0] ,
         \xmem_inst/mem[85][7] , \xmem_inst/mem[85][6] ,
         \xmem_inst/mem[85][5] , \xmem_inst/mem[85][4] ,
         \xmem_inst/mem[85][3] , \xmem_inst/mem[85][2] ,
         \xmem_inst/mem[85][1] , \xmem_inst/mem[85][0] ,
         \xmem_inst/mem[84][7] , \xmem_inst/mem[84][6] ,
         \xmem_inst/mem[84][5] , \xmem_inst/mem[84][4] ,
         \xmem_inst/mem[84][3] , \xmem_inst/mem[84][2] ,
         \xmem_inst/mem[84][1] , \xmem_inst/mem[84][0] ,
         \xmem_inst/mem[83][7] , \xmem_inst/mem[83][6] ,
         \xmem_inst/mem[83][5] , \xmem_inst/mem[83][4] ,
         \xmem_inst/mem[83][3] , \xmem_inst/mem[83][2] ,
         \xmem_inst/mem[83][1] , \xmem_inst/mem[83][0] ,
         \xmem_inst/mem[82][7] , \xmem_inst/mem[82][6] ,
         \xmem_inst/mem[82][5] , \xmem_inst/mem[82][4] ,
         \xmem_inst/mem[82][3] , \xmem_inst/mem[82][2] ,
         \xmem_inst/mem[82][1] , \xmem_inst/mem[82][0] ,
         \xmem_inst/mem[81][7] , \xmem_inst/mem[81][6] ,
         \xmem_inst/mem[81][5] , \xmem_inst/mem[81][4] ,
         \xmem_inst/mem[81][3] , \xmem_inst/mem[81][2] ,
         \xmem_inst/mem[81][1] , \xmem_inst/mem[81][0] ,
         \xmem_inst/mem[80][7] , \xmem_inst/mem[80][6] ,
         \xmem_inst/mem[80][5] , \xmem_inst/mem[80][4] ,
         \xmem_inst/mem[80][3] , \xmem_inst/mem[80][2] ,
         \xmem_inst/mem[80][1] , \xmem_inst/mem[80][0] ,
         \xmem_inst/mem[79][7] , \xmem_inst/mem[79][6] ,
         \xmem_inst/mem[79][5] , \xmem_inst/mem[79][4] ,
         \xmem_inst/mem[79][3] , \xmem_inst/mem[79][2] ,
         \xmem_inst/mem[79][1] , \xmem_inst/mem[79][0] ,
         \xmem_inst/mem[78][7] , \xmem_inst/mem[78][6] ,
         \xmem_inst/mem[78][5] , \xmem_inst/mem[78][4] ,
         \xmem_inst/mem[78][3] , \xmem_inst/mem[78][2] ,
         \xmem_inst/mem[78][1] , \xmem_inst/mem[78][0] ,
         \xmem_inst/mem[77][7] , \xmem_inst/mem[77][6] ,
         \xmem_inst/mem[77][5] , \xmem_inst/mem[77][4] ,
         \xmem_inst/mem[77][3] , \xmem_inst/mem[77][2] ,
         \xmem_inst/mem[77][1] , \xmem_inst/mem[77][0] ,
         \xmem_inst/mem[76][7] , \xmem_inst/mem[76][6] ,
         \xmem_inst/mem[76][5] , \xmem_inst/mem[76][4] ,
         \xmem_inst/mem[76][3] , \xmem_inst/mem[76][2] ,
         \xmem_inst/mem[76][1] , \xmem_inst/mem[76][0] ,
         \xmem_inst/mem[75][7] , \xmem_inst/mem[75][6] ,
         \xmem_inst/mem[75][5] , \xmem_inst/mem[75][4] ,
         \xmem_inst/mem[75][3] , \xmem_inst/mem[75][2] ,
         \xmem_inst/mem[75][1] , \xmem_inst/mem[75][0] ,
         \xmem_inst/mem[74][7] , \xmem_inst/mem[74][6] ,
         \xmem_inst/mem[74][5] , \xmem_inst/mem[74][4] ,
         \xmem_inst/mem[74][3] , \xmem_inst/mem[74][2] ,
         \xmem_inst/mem[74][1] , \xmem_inst/mem[74][0] ,
         \xmem_inst/mem[73][7] , \xmem_inst/mem[73][6] ,
         \xmem_inst/mem[73][5] , \xmem_inst/mem[73][4] ,
         \xmem_inst/mem[73][3] , \xmem_inst/mem[73][2] ,
         \xmem_inst/mem[73][1] , \xmem_inst/mem[73][0] ,
         \xmem_inst/mem[72][7] , \xmem_inst/mem[72][6] ,
         \xmem_inst/mem[72][5] , \xmem_inst/mem[72][4] ,
         \xmem_inst/mem[72][3] , \xmem_inst/mem[72][2] ,
         \xmem_inst/mem[72][1] , \xmem_inst/mem[72][0] ,
         \xmem_inst/mem[71][7] , \xmem_inst/mem[71][6] ,
         \xmem_inst/mem[71][5] , \xmem_inst/mem[71][4] ,
         \xmem_inst/mem[71][3] , \xmem_inst/mem[71][2] ,
         \xmem_inst/mem[71][1] , \xmem_inst/mem[71][0] ,
         \xmem_inst/mem[70][7] , \xmem_inst/mem[70][6] ,
         \xmem_inst/mem[70][5] , \xmem_inst/mem[70][4] ,
         \xmem_inst/mem[70][3] , \xmem_inst/mem[70][2] ,
         \xmem_inst/mem[70][1] , \xmem_inst/mem[70][0] ,
         \xmem_inst/mem[69][7] , \xmem_inst/mem[69][6] ,
         \xmem_inst/mem[69][5] , \xmem_inst/mem[69][4] ,
         \xmem_inst/mem[69][3] , \xmem_inst/mem[69][2] ,
         \xmem_inst/mem[69][1] , \xmem_inst/mem[69][0] ,
         \xmem_inst/mem[68][7] , \xmem_inst/mem[68][6] ,
         \xmem_inst/mem[68][5] , \xmem_inst/mem[68][4] ,
         \xmem_inst/mem[68][3] , \xmem_inst/mem[68][2] ,
         \xmem_inst/mem[68][1] , \xmem_inst/mem[68][0] ,
         \xmem_inst/mem[67][7] , \xmem_inst/mem[67][6] ,
         \xmem_inst/mem[67][5] , \xmem_inst/mem[67][4] ,
         \xmem_inst/mem[67][3] , \xmem_inst/mem[67][2] ,
         \xmem_inst/mem[67][1] , \xmem_inst/mem[67][0] ,
         \xmem_inst/mem[66][7] , \xmem_inst/mem[66][6] ,
         \xmem_inst/mem[66][5] , \xmem_inst/mem[66][4] ,
         \xmem_inst/mem[66][3] , \xmem_inst/mem[66][2] ,
         \xmem_inst/mem[66][1] , \xmem_inst/mem[66][0] ,
         \xmem_inst/mem[65][7] , \xmem_inst/mem[65][6] ,
         \xmem_inst/mem[65][5] , \xmem_inst/mem[65][4] ,
         \xmem_inst/mem[65][3] , \xmem_inst/mem[65][2] ,
         \xmem_inst/mem[65][1] , \xmem_inst/mem[65][0] ,
         \xmem_inst/mem[64][7] , \xmem_inst/mem[64][6] ,
         \xmem_inst/mem[64][5] , \xmem_inst/mem[64][4] ,
         \xmem_inst/mem[64][3] , \xmem_inst/mem[64][2] ,
         \xmem_inst/mem[64][1] , \xmem_inst/mem[64][0] ,
         \xmem_inst/mem[63][7] , \xmem_inst/mem[63][6] ,
         \xmem_inst/mem[63][5] , \xmem_inst/mem[63][4] ,
         \xmem_inst/mem[63][3] , \xmem_inst/mem[63][2] ,
         \xmem_inst/mem[63][1] , \xmem_inst/mem[63][0] ,
         \xmem_inst/mem[62][7] , \xmem_inst/mem[62][6] ,
         \xmem_inst/mem[62][5] , \xmem_inst/mem[62][4] ,
         \xmem_inst/mem[62][3] , \xmem_inst/mem[62][2] ,
         \xmem_inst/mem[62][1] , \xmem_inst/mem[62][0] ,
         \xmem_inst/mem[61][7] , \xmem_inst/mem[61][6] ,
         \xmem_inst/mem[61][5] , \xmem_inst/mem[61][4] ,
         \xmem_inst/mem[61][3] , \xmem_inst/mem[61][2] ,
         \xmem_inst/mem[61][1] , \xmem_inst/mem[61][0] ,
         \xmem_inst/mem[60][7] , \xmem_inst/mem[60][6] ,
         \xmem_inst/mem[60][5] , \xmem_inst/mem[60][4] ,
         \xmem_inst/mem[60][3] , \xmem_inst/mem[60][2] ,
         \xmem_inst/mem[60][1] , \xmem_inst/mem[60][0] ,
         \xmem_inst/mem[59][7] , \xmem_inst/mem[59][6] ,
         \xmem_inst/mem[59][5] , \xmem_inst/mem[59][4] ,
         \xmem_inst/mem[59][3] , \xmem_inst/mem[59][2] ,
         \xmem_inst/mem[59][1] , \xmem_inst/mem[59][0] ,
         \xmem_inst/mem[58][7] , \xmem_inst/mem[58][6] ,
         \xmem_inst/mem[58][5] , \xmem_inst/mem[58][4] ,
         \xmem_inst/mem[58][3] , \xmem_inst/mem[58][2] ,
         \xmem_inst/mem[58][1] , \xmem_inst/mem[58][0] ,
         \xmem_inst/mem[57][7] , \xmem_inst/mem[57][6] ,
         \xmem_inst/mem[57][5] , \xmem_inst/mem[57][4] ,
         \xmem_inst/mem[57][3] , \xmem_inst/mem[57][2] ,
         \xmem_inst/mem[57][1] , \xmem_inst/mem[57][0] ,
         \xmem_inst/mem[56][7] , \xmem_inst/mem[56][6] ,
         \xmem_inst/mem[56][5] , \xmem_inst/mem[56][4] ,
         \xmem_inst/mem[56][3] , \xmem_inst/mem[56][2] ,
         \xmem_inst/mem[56][1] , \xmem_inst/mem[56][0] ,
         \xmem_inst/mem[55][7] , \xmem_inst/mem[55][6] ,
         \xmem_inst/mem[55][5] , \xmem_inst/mem[55][4] ,
         \xmem_inst/mem[55][3] , \xmem_inst/mem[55][2] ,
         \xmem_inst/mem[55][1] , \xmem_inst/mem[55][0] ,
         \xmem_inst/mem[54][7] , \xmem_inst/mem[54][6] ,
         \xmem_inst/mem[54][5] , \xmem_inst/mem[54][4] ,
         \xmem_inst/mem[54][3] , \xmem_inst/mem[54][2] ,
         \xmem_inst/mem[54][1] , \xmem_inst/mem[54][0] ,
         \xmem_inst/mem[53][7] , \xmem_inst/mem[53][6] ,
         \xmem_inst/mem[53][5] , \xmem_inst/mem[53][4] ,
         \xmem_inst/mem[53][3] , \xmem_inst/mem[53][2] ,
         \xmem_inst/mem[53][1] , \xmem_inst/mem[53][0] ,
         \xmem_inst/mem[52][7] , \xmem_inst/mem[52][6] ,
         \xmem_inst/mem[52][5] , \xmem_inst/mem[52][4] ,
         \xmem_inst/mem[52][3] , \xmem_inst/mem[52][2] ,
         \xmem_inst/mem[52][1] , \xmem_inst/mem[52][0] ,
         \xmem_inst/mem[51][7] , \xmem_inst/mem[51][6] ,
         \xmem_inst/mem[51][5] , \xmem_inst/mem[51][4] ,
         \xmem_inst/mem[51][3] , \xmem_inst/mem[51][2] ,
         \xmem_inst/mem[51][1] , \xmem_inst/mem[51][0] ,
         \xmem_inst/mem[50][7] , \xmem_inst/mem[50][6] ,
         \xmem_inst/mem[50][5] , \xmem_inst/mem[50][4] ,
         \xmem_inst/mem[50][3] , \xmem_inst/mem[50][2] ,
         \xmem_inst/mem[50][1] , \xmem_inst/mem[50][0] ,
         \xmem_inst/mem[49][7] , \xmem_inst/mem[49][6] ,
         \xmem_inst/mem[49][5] , \xmem_inst/mem[49][4] ,
         \xmem_inst/mem[49][3] , \xmem_inst/mem[49][2] ,
         \xmem_inst/mem[49][1] , \xmem_inst/mem[49][0] ,
         \xmem_inst/mem[48][7] , \xmem_inst/mem[48][6] ,
         \xmem_inst/mem[48][5] , \xmem_inst/mem[48][4] ,
         \xmem_inst/mem[48][3] , \xmem_inst/mem[48][2] ,
         \xmem_inst/mem[48][1] , \xmem_inst/mem[48][0] ,
         \xmem_inst/mem[47][7] , \xmem_inst/mem[47][6] ,
         \xmem_inst/mem[47][5] , \xmem_inst/mem[47][4] ,
         \xmem_inst/mem[47][3] , \xmem_inst/mem[47][2] ,
         \xmem_inst/mem[47][1] , \xmem_inst/mem[47][0] ,
         \xmem_inst/mem[46][7] , \xmem_inst/mem[46][6] ,
         \xmem_inst/mem[46][5] , \xmem_inst/mem[46][4] ,
         \xmem_inst/mem[46][3] , \xmem_inst/mem[46][2] ,
         \xmem_inst/mem[46][1] , \xmem_inst/mem[46][0] ,
         \xmem_inst/mem[45][7] , \xmem_inst/mem[45][6] ,
         \xmem_inst/mem[45][5] , \xmem_inst/mem[45][4] ,
         \xmem_inst/mem[45][3] , \xmem_inst/mem[45][2] ,
         \xmem_inst/mem[45][1] , \xmem_inst/mem[45][0] ,
         \xmem_inst/mem[44][7] , \xmem_inst/mem[44][6] ,
         \xmem_inst/mem[44][5] , \xmem_inst/mem[44][4] ,
         \xmem_inst/mem[44][3] , \xmem_inst/mem[44][2] ,
         \xmem_inst/mem[44][1] , \xmem_inst/mem[44][0] ,
         \xmem_inst/mem[43][7] , \xmem_inst/mem[43][6] ,
         \xmem_inst/mem[43][5] , \xmem_inst/mem[43][4] ,
         \xmem_inst/mem[43][3] , \xmem_inst/mem[43][2] ,
         \xmem_inst/mem[43][1] , \xmem_inst/mem[43][0] ,
         \xmem_inst/mem[42][7] , \xmem_inst/mem[42][6] ,
         \xmem_inst/mem[42][5] , \xmem_inst/mem[42][4] ,
         \xmem_inst/mem[42][3] , \xmem_inst/mem[42][2] ,
         \xmem_inst/mem[42][1] , \xmem_inst/mem[42][0] ,
         \xmem_inst/mem[41][7] , \xmem_inst/mem[41][6] ,
         \xmem_inst/mem[41][5] , \xmem_inst/mem[41][4] ,
         \xmem_inst/mem[41][3] , \xmem_inst/mem[41][2] ,
         \xmem_inst/mem[41][1] , \xmem_inst/mem[41][0] ,
         \xmem_inst/mem[40][7] , \xmem_inst/mem[40][6] ,
         \xmem_inst/mem[40][5] , \xmem_inst/mem[40][4] ,
         \xmem_inst/mem[40][3] , \xmem_inst/mem[40][2] ,
         \xmem_inst/mem[40][1] , \xmem_inst/mem[40][0] ,
         \xmem_inst/mem[39][7] , \xmem_inst/mem[39][6] ,
         \xmem_inst/mem[39][5] , \xmem_inst/mem[39][4] ,
         \xmem_inst/mem[39][3] , \xmem_inst/mem[39][2] ,
         \xmem_inst/mem[39][1] , \xmem_inst/mem[39][0] ,
         \xmem_inst/mem[38][7] , \xmem_inst/mem[38][6] ,
         \xmem_inst/mem[38][5] , \xmem_inst/mem[38][4] ,
         \xmem_inst/mem[38][3] , \xmem_inst/mem[38][2] ,
         \xmem_inst/mem[38][1] , \xmem_inst/mem[38][0] ,
         \xmem_inst/mem[37][7] , \xmem_inst/mem[37][6] ,
         \xmem_inst/mem[37][5] , \xmem_inst/mem[37][4] ,
         \xmem_inst/mem[37][3] , \xmem_inst/mem[37][2] ,
         \xmem_inst/mem[37][1] , \xmem_inst/mem[37][0] ,
         \xmem_inst/mem[36][7] , \xmem_inst/mem[36][6] ,
         \xmem_inst/mem[36][5] , \xmem_inst/mem[36][4] ,
         \xmem_inst/mem[36][3] , \xmem_inst/mem[36][2] ,
         \xmem_inst/mem[36][1] , \xmem_inst/mem[36][0] ,
         \xmem_inst/mem[35][7] , \xmem_inst/mem[35][6] ,
         \xmem_inst/mem[35][5] , \xmem_inst/mem[35][4] ,
         \xmem_inst/mem[35][3] , \xmem_inst/mem[35][2] ,
         \xmem_inst/mem[35][1] , \xmem_inst/mem[35][0] ,
         \xmem_inst/mem[34][7] , \xmem_inst/mem[34][6] ,
         \xmem_inst/mem[34][5] , \xmem_inst/mem[34][4] ,
         \xmem_inst/mem[34][3] , \xmem_inst/mem[34][2] ,
         \xmem_inst/mem[34][1] , \xmem_inst/mem[34][0] ,
         \xmem_inst/mem[33][7] , \xmem_inst/mem[33][6] ,
         \xmem_inst/mem[33][5] , \xmem_inst/mem[33][4] ,
         \xmem_inst/mem[33][3] , \xmem_inst/mem[33][2] ,
         \xmem_inst/mem[33][1] , \xmem_inst/mem[33][0] ,
         \xmem_inst/mem[32][7] , \xmem_inst/mem[32][6] ,
         \xmem_inst/mem[32][5] , \xmem_inst/mem[32][4] ,
         \xmem_inst/mem[32][3] , \xmem_inst/mem[32][2] ,
         \xmem_inst/mem[32][1] , \xmem_inst/mem[32][0] ,
         \xmem_inst/mem[31][7] , \xmem_inst/mem[31][6] ,
         \xmem_inst/mem[31][5] , \xmem_inst/mem[31][4] ,
         \xmem_inst/mem[31][3] , \xmem_inst/mem[31][2] ,
         \xmem_inst/mem[31][1] , \xmem_inst/mem[31][0] ,
         \xmem_inst/mem[30][7] , \xmem_inst/mem[30][6] ,
         \xmem_inst/mem[30][5] , \xmem_inst/mem[30][4] ,
         \xmem_inst/mem[30][3] , \xmem_inst/mem[30][2] ,
         \xmem_inst/mem[30][1] , \xmem_inst/mem[30][0] ,
         \xmem_inst/mem[29][7] , \xmem_inst/mem[29][6] ,
         \xmem_inst/mem[29][5] , \xmem_inst/mem[29][4] ,
         \xmem_inst/mem[29][3] , \xmem_inst/mem[29][2] ,
         \xmem_inst/mem[29][1] , \xmem_inst/mem[29][0] ,
         \xmem_inst/mem[28][7] , \xmem_inst/mem[28][6] ,
         \xmem_inst/mem[28][5] , \xmem_inst/mem[28][4] ,
         \xmem_inst/mem[28][3] , \xmem_inst/mem[28][2] ,
         \xmem_inst/mem[28][1] , \xmem_inst/mem[28][0] ,
         \xmem_inst/mem[27][7] , \xmem_inst/mem[27][6] ,
         \xmem_inst/mem[27][5] , \xmem_inst/mem[27][4] ,
         \xmem_inst/mem[27][3] , \xmem_inst/mem[27][2] ,
         \xmem_inst/mem[27][1] , \xmem_inst/mem[27][0] ,
         \xmem_inst/mem[26][7] , \xmem_inst/mem[26][6] ,
         \xmem_inst/mem[26][5] , \xmem_inst/mem[26][4] ,
         \xmem_inst/mem[26][3] , \xmem_inst/mem[26][2] ,
         \xmem_inst/mem[26][1] , \xmem_inst/mem[26][0] ,
         \xmem_inst/mem[25][7] , \xmem_inst/mem[25][6] ,
         \xmem_inst/mem[25][5] , \xmem_inst/mem[25][4] ,
         \xmem_inst/mem[25][3] , \xmem_inst/mem[25][2] ,
         \xmem_inst/mem[25][1] , \xmem_inst/mem[25][0] ,
         \xmem_inst/mem[24][7] , \xmem_inst/mem[24][6] ,
         \xmem_inst/mem[24][5] , \xmem_inst/mem[24][4] ,
         \xmem_inst/mem[24][3] , \xmem_inst/mem[24][2] ,
         \xmem_inst/mem[24][1] , \xmem_inst/mem[24][0] ,
         \xmem_inst/mem[23][7] , \xmem_inst/mem[23][6] ,
         \xmem_inst/mem[23][5] , \xmem_inst/mem[23][4] ,
         \xmem_inst/mem[23][3] , \xmem_inst/mem[23][2] ,
         \xmem_inst/mem[23][1] , \xmem_inst/mem[23][0] ,
         \xmem_inst/mem[22][7] , \xmem_inst/mem[22][6] ,
         \xmem_inst/mem[22][5] , \xmem_inst/mem[22][4] ,
         \xmem_inst/mem[22][3] , \xmem_inst/mem[22][2] ,
         \xmem_inst/mem[22][1] , \xmem_inst/mem[22][0] ,
         \xmem_inst/mem[21][7] , \xmem_inst/mem[21][6] ,
         \xmem_inst/mem[21][5] , \xmem_inst/mem[21][4] ,
         \xmem_inst/mem[21][3] , \xmem_inst/mem[21][2] ,
         \xmem_inst/mem[21][1] , \xmem_inst/mem[21][0] ,
         \xmem_inst/mem[20][7] , \xmem_inst/mem[20][6] ,
         \xmem_inst/mem[20][5] , \xmem_inst/mem[20][4] ,
         \xmem_inst/mem[20][3] , \xmem_inst/mem[20][2] ,
         \xmem_inst/mem[20][1] , \xmem_inst/mem[20][0] ,
         \xmem_inst/mem[19][7] , \xmem_inst/mem[19][6] ,
         \xmem_inst/mem[19][5] , \xmem_inst/mem[19][4] ,
         \xmem_inst/mem[19][3] , \xmem_inst/mem[19][2] ,
         \xmem_inst/mem[19][1] , \xmem_inst/mem[19][0] ,
         \xmem_inst/mem[18][7] , \xmem_inst/mem[18][6] ,
         \xmem_inst/mem[18][5] , \xmem_inst/mem[18][4] ,
         \xmem_inst/mem[18][3] , \xmem_inst/mem[18][2] ,
         \xmem_inst/mem[18][1] , \xmem_inst/mem[18][0] ,
         \xmem_inst/mem[17][7] , \xmem_inst/mem[17][6] ,
         \xmem_inst/mem[17][5] , \xmem_inst/mem[17][4] ,
         \xmem_inst/mem[17][3] , \xmem_inst/mem[17][2] ,
         \xmem_inst/mem[17][1] , \xmem_inst/mem[17][0] ,
         \xmem_inst/mem[16][7] , \xmem_inst/mem[16][6] ,
         \xmem_inst/mem[16][5] , \xmem_inst/mem[16][4] ,
         \xmem_inst/mem[16][3] , \xmem_inst/mem[16][2] ,
         \xmem_inst/mem[16][1] , \xmem_inst/mem[16][0] ,
         \xmem_inst/mem[15][7] , \xmem_inst/mem[15][6] ,
         \xmem_inst/mem[15][5] , \xmem_inst/mem[15][4] ,
         \xmem_inst/mem[15][3] , \xmem_inst/mem[15][2] ,
         \xmem_inst/mem[15][1] , \xmem_inst/mem[15][0] ,
         \xmem_inst/mem[14][7] , \xmem_inst/mem[14][6] ,
         \xmem_inst/mem[14][5] , \xmem_inst/mem[14][4] ,
         \xmem_inst/mem[14][3] , \xmem_inst/mem[14][2] ,
         \xmem_inst/mem[14][1] , \xmem_inst/mem[14][0] ,
         \xmem_inst/mem[13][7] , \xmem_inst/mem[13][6] ,
         \xmem_inst/mem[13][5] , \xmem_inst/mem[13][4] ,
         \xmem_inst/mem[13][3] , \xmem_inst/mem[13][2] ,
         \xmem_inst/mem[13][1] , \xmem_inst/mem[13][0] ,
         \xmem_inst/mem[12][7] , \xmem_inst/mem[12][6] ,
         \xmem_inst/mem[12][5] , \xmem_inst/mem[12][4] ,
         \xmem_inst/mem[12][3] , \xmem_inst/mem[12][2] ,
         \xmem_inst/mem[12][1] , \xmem_inst/mem[12][0] ,
         \xmem_inst/mem[11][7] , \xmem_inst/mem[11][6] ,
         \xmem_inst/mem[11][5] , \xmem_inst/mem[11][4] ,
         \xmem_inst/mem[11][3] , \xmem_inst/mem[11][2] ,
         \xmem_inst/mem[11][1] , \xmem_inst/mem[11][0] ,
         \xmem_inst/mem[10][7] , \xmem_inst/mem[10][6] ,
         \xmem_inst/mem[10][5] , \xmem_inst/mem[10][4] ,
         \xmem_inst/mem[10][3] , \xmem_inst/mem[10][2] ,
         \xmem_inst/mem[10][1] , \xmem_inst/mem[10][0] , \xmem_inst/mem[9][7] ,
         \xmem_inst/mem[9][6] , \xmem_inst/mem[9][5] , \xmem_inst/mem[9][4] ,
         \xmem_inst/mem[9][3] , \xmem_inst/mem[9][2] , \xmem_inst/mem[9][1] ,
         \xmem_inst/mem[9][0] , \xmem_inst/mem[8][7] , \xmem_inst/mem[8][6] ,
         \xmem_inst/mem[8][5] , \xmem_inst/mem[8][4] , \xmem_inst/mem[8][3] ,
         \xmem_inst/mem[8][2] , \xmem_inst/mem[8][1] , \xmem_inst/mem[8][0] ,
         \xmem_inst/mem[7][7] , \xmem_inst/mem[7][6] , \xmem_inst/mem[7][5] ,
         \xmem_inst/mem[7][4] , \xmem_inst/mem[7][3] , \xmem_inst/mem[7][2] ,
         \xmem_inst/mem[7][1] , \xmem_inst/mem[7][0] , \xmem_inst/mem[6][7] ,
         \xmem_inst/mem[6][6] , \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] ,
         \xmem_inst/mem[6][3] , \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] ,
         \xmem_inst/mem[6][0] , \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] ,
         \xmem_inst/mem[5][5] , \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] ,
         \xmem_inst/mem[5][2] , \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] ,
         \xmem_inst/mem[4][7] , \xmem_inst/mem[4][6] , \xmem_inst/mem[4][5] ,
         \xmem_inst/mem[4][4] , \xmem_inst/mem[4][3] , \xmem_inst/mem[4][2] ,
         \xmem_inst/mem[4][1] , \xmem_inst/mem[4][0] , \xmem_inst/mem[3][7] ,
         \xmem_inst/mem[3][6] , \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] ,
         \xmem_inst/mem[3][3] , \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] ,
         \xmem_inst/mem[3][0] , \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] ,
         \xmem_inst/mem[2][5] , \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] ,
         \xmem_inst/mem[2][2] , \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] ,
         \xmem_inst/mem[1][7] , \xmem_inst/mem[1][6] , \xmem_inst/mem[1][5] ,
         \xmem_inst/mem[1][4] , \xmem_inst/mem[1][3] , \xmem_inst/mem[1][2] ,
         \xmem_inst/mem[1][1] , \xmem_inst/mem[1][0] , \xmem_inst/mem[0][7] ,
         \xmem_inst/mem[0][6] , \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] ,
         \xmem_inst/mem[0][3] , \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] ,
         \xmem_inst/mem[0][0] , \fmem_inst/mem[31][7] , \fmem_inst/mem[31][6] ,
         \fmem_inst/mem[31][5] , \fmem_inst/mem[31][4] ,
         \fmem_inst/mem[31][3] , \fmem_inst/mem[31][2] ,
         \fmem_inst/mem[31][1] , \fmem_inst/mem[31][0] ,
         \fmem_inst/mem[30][7] , \fmem_inst/mem[30][6] ,
         \fmem_inst/mem[30][5] , \fmem_inst/mem[30][4] ,
         \fmem_inst/mem[30][3] , \fmem_inst/mem[30][2] ,
         \fmem_inst/mem[30][1] , \fmem_inst/mem[30][0] ,
         \fmem_inst/mem[29][7] , \fmem_inst/mem[29][6] ,
         \fmem_inst/mem[29][5] , \fmem_inst/mem[29][4] ,
         \fmem_inst/mem[29][3] , \fmem_inst/mem[29][2] ,
         \fmem_inst/mem[29][1] , \fmem_inst/mem[29][0] ,
         \fmem_inst/mem[28][7] , \fmem_inst/mem[28][6] ,
         \fmem_inst/mem[28][5] , \fmem_inst/mem[28][4] ,
         \fmem_inst/mem[28][3] , \fmem_inst/mem[28][2] ,
         \fmem_inst/mem[28][1] , \fmem_inst/mem[28][0] ,
         \fmem_inst/mem[27][7] , \fmem_inst/mem[27][6] ,
         \fmem_inst/mem[27][5] , \fmem_inst/mem[27][4] ,
         \fmem_inst/mem[27][3] , \fmem_inst/mem[27][2] ,
         \fmem_inst/mem[27][1] , \fmem_inst/mem[27][0] ,
         \fmem_inst/mem[26][7] , \fmem_inst/mem[26][6] ,
         \fmem_inst/mem[26][5] , \fmem_inst/mem[26][4] ,
         \fmem_inst/mem[26][3] , \fmem_inst/mem[26][2] ,
         \fmem_inst/mem[26][1] , \fmem_inst/mem[26][0] ,
         \fmem_inst/mem[25][7] , \fmem_inst/mem[25][6] ,
         \fmem_inst/mem[25][5] , \fmem_inst/mem[25][4] ,
         \fmem_inst/mem[25][3] , \fmem_inst/mem[25][2] ,
         \fmem_inst/mem[25][1] , \fmem_inst/mem[25][0] ,
         \fmem_inst/mem[24][7] , \fmem_inst/mem[24][6] ,
         \fmem_inst/mem[24][5] , \fmem_inst/mem[24][4] ,
         \fmem_inst/mem[24][3] , \fmem_inst/mem[24][2] ,
         \fmem_inst/mem[24][1] , \fmem_inst/mem[24][0] ,
         \fmem_inst/mem[23][7] , \fmem_inst/mem[23][6] ,
         \fmem_inst/mem[23][5] , \fmem_inst/mem[23][4] ,
         \fmem_inst/mem[23][3] , \fmem_inst/mem[23][2] ,
         \fmem_inst/mem[23][1] , \fmem_inst/mem[23][0] ,
         \fmem_inst/mem[22][7] , \fmem_inst/mem[22][6] ,
         \fmem_inst/mem[22][5] , \fmem_inst/mem[22][4] ,
         \fmem_inst/mem[22][3] , \fmem_inst/mem[22][2] ,
         \fmem_inst/mem[22][1] , \fmem_inst/mem[22][0] ,
         \fmem_inst/mem[21][7] , \fmem_inst/mem[21][6] ,
         \fmem_inst/mem[21][5] , \fmem_inst/mem[21][4] ,
         \fmem_inst/mem[21][3] , \fmem_inst/mem[21][2] ,
         \fmem_inst/mem[21][1] , \fmem_inst/mem[21][0] ,
         \fmem_inst/mem[20][7] , \fmem_inst/mem[20][6] ,
         \fmem_inst/mem[20][5] , \fmem_inst/mem[20][4] ,
         \fmem_inst/mem[20][3] , \fmem_inst/mem[20][2] ,
         \fmem_inst/mem[20][1] , \fmem_inst/mem[20][0] ,
         \fmem_inst/mem[19][7] , \fmem_inst/mem[19][6] ,
         \fmem_inst/mem[19][5] , \fmem_inst/mem[19][4] ,
         \fmem_inst/mem[19][3] , \fmem_inst/mem[19][2] ,
         \fmem_inst/mem[19][1] , \fmem_inst/mem[19][0] ,
         \fmem_inst/mem[18][7] , \fmem_inst/mem[18][6] ,
         \fmem_inst/mem[18][5] , \fmem_inst/mem[18][4] ,
         \fmem_inst/mem[18][3] , \fmem_inst/mem[18][2] ,
         \fmem_inst/mem[18][1] , \fmem_inst/mem[18][0] ,
         \fmem_inst/mem[17][7] , \fmem_inst/mem[17][6] ,
         \fmem_inst/mem[17][5] , \fmem_inst/mem[17][4] ,
         \fmem_inst/mem[17][3] , \fmem_inst/mem[17][2] ,
         \fmem_inst/mem[17][1] , \fmem_inst/mem[17][0] ,
         \fmem_inst/mem[16][7] , \fmem_inst/mem[16][6] ,
         \fmem_inst/mem[16][5] , \fmem_inst/mem[16][4] ,
         \fmem_inst/mem[16][3] , \fmem_inst/mem[16][2] ,
         \fmem_inst/mem[16][1] , \fmem_inst/mem[16][0] ,
         \fmem_inst/mem[15][7] , \fmem_inst/mem[15][6] ,
         \fmem_inst/mem[15][5] , \fmem_inst/mem[15][4] ,
         \fmem_inst/mem[15][3] , \fmem_inst/mem[15][2] ,
         \fmem_inst/mem[15][1] , \fmem_inst/mem[15][0] ,
         \fmem_inst/mem[14][7] , \fmem_inst/mem[14][6] ,
         \fmem_inst/mem[14][5] , \fmem_inst/mem[14][4] ,
         \fmem_inst/mem[14][3] , \fmem_inst/mem[14][2] ,
         \fmem_inst/mem[14][1] , \fmem_inst/mem[14][0] ,
         \fmem_inst/mem[13][7] , \fmem_inst/mem[13][6] ,
         \fmem_inst/mem[13][5] , \fmem_inst/mem[13][4] ,
         \fmem_inst/mem[13][3] , \fmem_inst/mem[13][2] ,
         \fmem_inst/mem[13][1] , \fmem_inst/mem[13][0] ,
         \fmem_inst/mem[12][7] , \fmem_inst/mem[12][6] ,
         \fmem_inst/mem[12][5] , \fmem_inst/mem[12][4] ,
         \fmem_inst/mem[12][3] , \fmem_inst/mem[12][2] ,
         \fmem_inst/mem[12][1] , \fmem_inst/mem[12][0] ,
         \fmem_inst/mem[11][7] , \fmem_inst/mem[11][6] ,
         \fmem_inst/mem[11][5] , \fmem_inst/mem[11][4] ,
         \fmem_inst/mem[11][3] , \fmem_inst/mem[11][2] ,
         \fmem_inst/mem[11][1] , \fmem_inst/mem[11][0] ,
         \fmem_inst/mem[10][7] , \fmem_inst/mem[10][6] ,
         \fmem_inst/mem[10][5] , \fmem_inst/mem[10][4] ,
         \fmem_inst/mem[10][3] , \fmem_inst/mem[10][2] ,
         \fmem_inst/mem[10][1] , \fmem_inst/mem[10][0] , \fmem_inst/mem[9][7] ,
         \fmem_inst/mem[9][6] , \fmem_inst/mem[9][5] , \fmem_inst/mem[9][4] ,
         \fmem_inst/mem[9][3] , \fmem_inst/mem[9][2] , \fmem_inst/mem[9][1] ,
         \fmem_inst/mem[9][0] , \fmem_inst/mem[8][7] , \fmem_inst/mem[8][6] ,
         \fmem_inst/mem[8][5] , \fmem_inst/mem[8][4] , \fmem_inst/mem[8][3] ,
         \fmem_inst/mem[8][2] , \fmem_inst/mem[8][1] , \fmem_inst/mem[8][0] ,
         \fmem_inst/mem[7][7] , \fmem_inst/mem[7][6] , \fmem_inst/mem[7][5] ,
         \fmem_inst/mem[7][4] , \fmem_inst/mem[7][3] , \fmem_inst/mem[7][2] ,
         \fmem_inst/mem[7][1] , \fmem_inst/mem[7][0] , \fmem_inst/mem[6][7] ,
         \fmem_inst/mem[6][6] , \fmem_inst/mem[6][5] , \fmem_inst/mem[6][4] ,
         \fmem_inst/mem[6][3] , \fmem_inst/mem[6][2] , \fmem_inst/mem[6][1] ,
         \fmem_inst/mem[6][0] , \fmem_inst/mem[5][7] , \fmem_inst/mem[5][6] ,
         \fmem_inst/mem[5][5] , \fmem_inst/mem[5][4] , \fmem_inst/mem[5][3] ,
         \fmem_inst/mem[5][2] , \fmem_inst/mem[5][1] , \fmem_inst/mem[5][0] ,
         \fmem_inst/mem[4][7] , \fmem_inst/mem[4][6] , \fmem_inst/mem[4][5] ,
         \fmem_inst/mem[4][4] , \fmem_inst/mem[4][3] , \fmem_inst/mem[4][2] ,
         \fmem_inst/mem[4][1] , \fmem_inst/mem[4][0] , \fmem_inst/mem[3][7] ,
         \fmem_inst/mem[3][6] , \fmem_inst/mem[3][5] , \fmem_inst/mem[3][4] ,
         \fmem_inst/mem[3][3] , \fmem_inst/mem[3][2] , \fmem_inst/mem[3][1] ,
         \fmem_inst/mem[3][0] , \fmem_inst/mem[2][7] , \fmem_inst/mem[2][6] ,
         \fmem_inst/mem[2][5] , \fmem_inst/mem[2][4] , \fmem_inst/mem[2][3] ,
         \fmem_inst/mem[2][2] , \fmem_inst/mem[2][1] , \fmem_inst/mem[2][0] ,
         \fmem_inst/mem[1][7] , \fmem_inst/mem[1][6] , \fmem_inst/mem[1][5] ,
         \fmem_inst/mem[1][4] , \fmem_inst/mem[1][3] , \fmem_inst/mem[1][2] ,
         \fmem_inst/mem[1][1] , \fmem_inst/mem[1][0] , \fmem_inst/mem[0][7] ,
         \fmem_inst/mem[0][6] , \fmem_inst/mem[0][5] , \fmem_inst/mem[0][4] ,
         \fmem_inst/mem[0][3] , \fmem_inst/mem[0][2] , \fmem_inst/mem[0][1] ,
         \fmem_inst/mem[0][0] , \ctrl_conv_output_inst/N7 ,
         \ctrl_conv_output_inst/conv_start_reg , n1814, n1815, n1816, n1817,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, \add_x_2/A[0] ,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
         n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
         n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
         n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
         n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836,
         n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
         n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
         n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
         n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
         n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
         n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
         n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
         n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
         n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908,
         n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
         n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
         n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
         n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
         n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
         n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
         n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
         n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
         n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
         n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
         n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
         n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
         n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
         n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
         n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
         n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100,
         n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
         n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
         n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
         n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
         n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
         n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
         n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
         n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
         n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
         n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
         n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
         n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
         n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220,
         n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
         n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236,
         n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
         n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
         n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
         n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
         n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
         n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
         n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292,
         n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
         n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308,
         n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
         n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324,
         n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
         n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
         n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
         n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
         n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364,
         n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
         n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
         n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
         n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
         n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
         n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
         n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
         n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
         n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436,
         n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
         n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452,
         n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
         n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468,
         n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
         n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
         n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492,
         n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
         n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508,
         n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
         n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524,
         n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
         n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540,
         n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
         n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
         n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
         n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
         n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
         n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
         n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
         n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
         n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
         n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
         n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652,
         n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
         n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
         n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
         n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
         n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
         n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
         n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
         n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
         n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724,
         n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
         n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
         n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
         n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
         n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
         n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
         n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
         n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
         n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796,
         n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
         n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
         n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
         n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
         n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
         n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844,
         n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
         n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
         n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
         n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
         n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900,
         n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
         n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
         n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
         n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
         n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940,
         n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
         n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
         n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
         n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036,
         n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
         n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
         n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
         n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
         n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
         n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
         n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132,
         n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
         n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
         n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156,
         n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
         n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
         n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180,
         n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
         n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
         n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204,
         n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
         n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228,
         n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
         n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
         n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252,
         n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
         n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
         n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276,
         n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284,
         n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
         n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300,
         n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
         n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
         n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324,
         n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
         n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
         n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348,
         n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356,
         n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
         n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372,
         n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
         n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
         n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396,
         n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
         n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
         n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420,
         n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
         n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
         n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
         n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
         n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492,
         n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500,
         n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
         n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516,
         n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
         n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
         n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540,
         n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
         n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
         n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564,
         n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
         n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
         n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588,
         n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
         n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
         n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612,
         n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
         n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
         n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
         n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
         n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
         n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
         n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708,
         n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716,
         n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
         n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
         n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
         n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
         n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
         n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
         n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
         n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
         n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
         n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
         n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
         n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
         n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
         n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116,
         n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
         n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
         n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140,
         n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148,
         n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
         n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164,
         n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
         n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
         n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188,
         n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
         n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
         n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212,
         n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
         n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
         n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236,
         n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
         n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
         n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260,
         n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
         n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
         n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284,
         n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292,
         n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
         n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308,
         n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
         n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
         n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332,
         n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340,
         n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
         n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364,
         n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
         n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380,
         n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
         n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396,
         n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404,
         n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412,
         n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
         n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
         n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436,
         n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
         n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
         n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
         n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
         n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476,
         n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
         n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
         n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
         n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508,
         n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
         n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
         n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
         n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
         n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548,
         n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
         n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
         n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
         n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
         n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
         n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
         n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
         n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
         n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
         n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
         n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
         n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668,
         n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
         n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
         n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692,
         n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
         n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
         n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
         n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
         n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
         n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740,
         n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
         n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
         n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
         n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
         n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
         n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
         n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
         n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
         n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812,
         n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
         n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
         n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
         n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
         n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
         n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
         n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
         n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884,
         n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
         n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
         n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
         n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
         n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
         n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
         n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
         n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
         n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
         n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
         n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
         n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
         n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
         n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
         n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
         n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
         n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
         n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028,
         n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
         n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
         n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052,
         n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060,
         n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
         n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
         n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084,
         n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
         n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
         n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
         n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
         n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124,
         n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
         n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
         n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
         n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156,
         n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
         n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172,
         n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
         n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
         n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
         n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
         n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
         n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
         n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228,
         n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
         n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
         n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
         n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
         n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268,
         n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
         n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
         n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300,
         n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
         n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
         n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
         n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
         n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340,
         n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
         n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
         n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
         n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
         n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
         n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388,
         n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412,
         n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
         n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
         n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
         n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
         n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
         n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
         n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
         n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
         n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
         n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
         n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
         n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
         n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
         n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580,
         n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
         n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
         n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
         n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
         n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
         n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
         n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
         n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
         n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
         n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
         n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
         n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
         n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
         n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
         n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
         n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
         n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
         n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
         n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
         n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
         n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
         n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
         n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
         n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
         n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
         n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
         n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
         n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
         n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
         n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
         n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
         n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
         n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
         n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
         n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
         n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
         n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
         n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
         n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
         n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
         n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
         n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
         n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
         n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
         n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
         n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
         n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
         n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
         n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
         n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
         n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
         n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
         n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
         n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
         n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
         n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
         n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
         n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
         n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
         n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
         n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
         n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
         n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
         n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
         n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
         n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
         n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
         n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
         n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
         n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
         n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
         n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
         n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
         n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
         n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
         n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
         n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
         n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
         n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
         n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
         n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
         n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
         n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
         n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
         n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
         n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
         n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
         n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
         n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
         n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
         n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
         n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
         n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
         n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
         n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308,
         n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
         n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
         n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
         n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
         n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
         n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
         n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
         n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
         n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380,
         n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
         n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
         n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
         n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
         n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
         n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
         n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
         n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460,
         n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
         n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
         n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
         n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
         n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500,
         n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
         n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
         n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524,
         n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
         n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
         n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
         n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
         n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
         n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
         n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
         n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
         n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
         n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
         n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
         n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
         n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
         n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
         n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
         n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
         n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
         n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
         n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
         n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
         n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
         n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748,
         n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
         n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
         n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
         n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
         n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788,
         n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
         n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
         n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
         n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
         n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
         n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
         n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
         n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860,
         n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
         n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
         n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
         n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892,
         n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
         n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
         n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
         n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
         n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004,
         n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
         n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
         n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
         n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068,
         n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076,
         n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
         n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
         n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100,
         n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108,
         n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
         n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
         n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
         n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
         n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148,
         n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
         n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164,
         n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172,
         n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180,
         n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
         n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196,
         n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204,
         n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
         n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220,
         n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
         n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236,
         n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244,
         n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252,
         n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
         n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
         n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
         n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284,
         n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292,
         n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
         n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308,
         n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316,
         n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324,
         n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
         n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340,
         n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
         n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356,
         n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364,
         n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372,
         n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380,
         n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388,
         n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396,
         n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
         n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412,
         n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420,
         n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428,
         n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436,
         n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444,
         n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452,
         n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460,
         n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468,
         n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
         n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484,
         n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492,
         n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500,
         n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508,
         n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
         n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524,
         n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532,
         n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
         n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
         n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556,
         n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
         n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
         n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580,
         n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
         n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596,
         n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
         n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612,
         n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
         n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628,
         n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636,
         n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644,
         n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652,
         n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
         n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
         n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
         n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684,
         n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
         n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700,
         n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708,
         n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716,
         n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724,
         n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732,
         n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740,
         n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748,
         n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756,
         n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
         n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772,
         n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
         n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788,
         n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796,
         n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804,
         n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812,
         n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820,
         n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828,
         n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
         n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844,
         n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852,
         n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860,
         n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868,
         n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876,
         n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884,
         n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892,
         n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900,
         n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
         n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916,
         n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924,
         n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932,
         n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940,
         n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948,
         n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956,
         n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964,
         n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972,
         n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980,
         n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988,
         n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996,
         n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004,
         n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012,
         n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020,
         n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028,
         n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036,
         n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044,
         n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
         n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
         n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
         n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
         n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084,
         n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
         n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100,
         n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
         n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116,
         n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
         n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132,
         n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
         n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148,
         n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156,
         n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
         n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172,
         n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180,
         n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188,
         n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
         n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204,
         n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212,
         n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220,
         n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228,
         n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236,
         n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244,
         n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252,
         n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260,
         n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
         n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276,
         n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284,
         n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292,
         n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300,
         n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308,
         n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316,
         n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324,
         n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332,
         n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
         n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348,
         n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356,
         n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364,
         n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372,
         n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380,
         n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388,
         n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396,
         n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404,
         n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412,
         n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420,
         n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428,
         n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436,
         n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444,
         n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452,
         n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
         n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468,
         n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476,
         n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
         n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492,
         n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
         n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
         n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516,
         n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
         n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
         n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
         n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548,
         n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
         n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564,
         n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572,
         n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580,
         n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588,
         n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
         n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604,
         n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612,
         n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620,
         n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
         n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636,
         n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644,
         n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652,
         n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660,
         n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
         n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676,
         n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684,
         n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692,
         n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
         n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708,
         n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716,
         n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724,
         n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732,
         n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740,
         n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
         n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756,
         n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764,
         n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
         n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780,
         n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
         n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796,
         n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804,
         n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812,
         n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820,
         n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828,
         n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836,
         n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
         n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852,
         n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860,
         n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868,
         n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876,
         n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884,
         n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892,
         n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900,
         n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908,
         n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
         n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924,
         n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
         n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940,
         n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948,
         n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956,
         n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964,
         n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972,
         n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980,
         n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
         n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996,
         n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
         n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012,
         n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020,
         n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028,
         n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
         n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
         n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052,
         n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
         n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068,
         n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
         n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
         n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
         n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
         n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
         n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
         n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124,
         n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
         n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140,
         n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
         n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
         n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164,
         n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
         n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
         n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188,
         n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196,
         n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
         n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212,
         n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
         n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
         n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236,
         n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244,
         n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
         n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260,
         n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
         n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
         n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284,
         n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
         n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
         n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308,
         n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
         n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324,
         n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332,
         n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340,
         n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
         n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
         n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
         n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
         n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380,
         n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
         n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
         n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428,
         n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
         n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
         n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452,
         n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
         n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
         n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476,
         n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484,
         n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
         n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500,
         n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
         n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516,
         n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524,
         n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
         n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
         n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548,
         n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
         n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
         n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
         n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
         n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
         n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596,
         n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
         n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
         n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
         n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
         n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
         n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644,
         n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
         n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
         n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668,
         n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
         n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
         n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
         n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
         n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
         n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
         n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740,
         n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
         n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
         n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764,
         n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
         n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
         n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
         n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
         n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
         n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
         n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
         n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
         n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
         n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
         n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
         n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
         n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
         n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
         n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
         n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908,
         n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
         n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
         n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
         n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
         n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
         n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
         n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
         n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
         n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980,
         n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
         n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
         n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
         n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
         n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
         n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
         n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
         n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052,
         n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
         n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
         n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
         n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
         n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092,
         n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
         n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108,
         n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116,
         n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124,
         n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132,
         n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
         n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148,
         n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
         n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
         n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
         n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196,
         n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204,
         n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
         n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220,
         n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
         n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236,
         n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244,
         n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
         n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260,
         n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
         n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
         n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
         n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
         n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
         n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
         n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316,
         n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324,
         n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332,
         n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340,
         n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348,
         n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
         n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364,
         n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
         n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
         n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388,
         n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396,
         n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404,
         n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412,
         n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
         n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
         n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436,
         n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
         n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
         n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460,
         n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
         n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
         n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484,
         n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
         n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
         n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508,
         n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
         n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
         n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532,
         n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540,
         n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
         n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556,
         n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
         n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
         n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580,
         n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
         n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
         n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604,
         n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
         n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620,
         n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
         n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
         n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
         n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652,
         n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
         n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
         n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676,
         n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684,
         n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692,
         n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700,
         n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
         n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
         n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724,
         n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
         n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740,
         n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748,
         n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756,
         n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764,
         n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772,
         n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780,
         n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
         n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796,
         n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
         n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812,
         n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820,
         n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
         n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836,
         n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844,
         n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852,
         n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
         n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868,
         n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
         n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884,
         n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892,
         n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900,
         n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908,
         n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916,
         n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924,
         n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
         n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940,
         n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
         n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956,
         n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964,
         n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972,
         n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980,
         n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
         n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
         n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
         n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012,
         n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
         n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028,
         n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036,
         n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044,
         n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
         n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
         n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068,
         n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
         n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084,
         n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
         n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100,
         n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108,
         n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
         n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
         n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132,
         n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140,
         n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
         n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156,
         n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
         n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
         n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180,
         n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
         n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212,
         n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
         n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
         n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
         n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
         n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300,
         n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
         n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
         n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324,
         n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
         n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
         n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
         n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
         n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
         n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
         n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
         n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
         n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
         n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
         n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444,
         n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
         n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
         n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468,
         n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
         n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
         n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
         n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
         n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
         n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516,
         n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
         n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
         n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540,
         n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
         n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
         n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
         n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572,
         n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
         n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588,
         n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
         n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604,
         n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612,
         n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
         n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628,
         n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636,
         n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644,
         n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
         n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660,
         n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
         n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
         n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684,
         n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
         n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700,
         n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708,
         n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716,
         n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
         n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732,
         n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
         n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748,
         n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756,
         n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
         n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772,
         n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780,
         n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788,
         n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
         n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804,
         n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
         n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820,
         n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828,
         n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
         n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
         n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852,
         n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860,
         n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
         n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876,
         n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
         n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
         n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
         n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
         n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916,
         n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
         n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932,
         n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
         n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948,
         n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
         n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
         n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972,
         n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
         n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
         n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
         n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004,
         n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
         n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
         n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
         n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044,
         n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
         n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
         n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068,
         n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076,
         n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
         n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092,
         n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
         n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108,
         n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116,
         n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
         n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
         n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140,
         n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148,
         n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
         n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164,
         n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
         n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
         n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188,
         n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
         n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
         n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212,
         n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220,
         n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
         n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236,
         n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
         n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
         n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260,
         n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
         n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
         n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284,
         n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292,
         n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
         n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308,
         n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
         n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
         n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332,
         n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
         n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348,
         n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356,
         n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
         n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
         n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380,
         n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
         n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
         n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404,
         n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
         n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420,
         n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428,
         n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
         n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
         n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452,
         n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
         n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
         n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476,
         n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
         n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492,
         n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500,
         n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508,
         n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
         n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524,
         n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
         n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540,
         n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548,
         n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
         n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564,
         n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572,
         n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580,
         n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
         n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596,
         n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
         n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612,
         n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
         n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628,
         n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636,
         n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644,
         n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652,
         n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
         n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668,
         n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
         n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684,
         n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692,
         n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700,
         n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708,
         n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716,
         n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724,
         n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732,
         n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740,
         n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
         n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756,
         n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764,
         n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772,
         n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780,
         n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788,
         n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796,
         n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804,
         n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812,
         n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
         n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828,
         n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836,
         n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844,
         n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852,
         n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860,
         n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868,
         n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876,
         n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884,
         n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892,
         n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900,
         n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908,
         n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
         n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924,
         n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932,
         n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940,
         n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948,
         n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956,
         n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964,
         n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972,
         n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980,
         n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
         n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996,
         n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004,
         n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012,
         n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020,
         n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028,
         n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036,
         n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044,
         n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052,
         n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060,
         n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068,
         n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076,
         n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084,
         n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092,
         n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100,
         n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
         n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116,
         n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124,
         n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132,
         n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140,
         n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148,
         n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156,
         n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164,
         n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172,
         n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180,
         n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188,
         n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196,
         n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204,
         n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212,
         n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220,
         n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228,
         n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
         n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244,
         n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
         n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260,
         n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268,
         n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276,
         n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284,
         n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292,
         n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300,
         n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
         n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316,
         n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324,
         n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332,
         n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340,
         n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
         n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356,
         n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364,
         n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372,
         n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
         n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388,
         n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
         n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
         n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412,
         n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
         n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
         n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436,
         n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444,
         n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
         n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460,
         n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468,
         n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476,
         n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484,
         n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492,
         n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500,
         n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508,
         n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516,
         n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
         n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532,
         n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
         n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548,
         n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556,
         n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564,
         n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572,
         n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580,
         n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588,
         n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
         n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604,
         n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
         n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620,
         n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628,
         n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
         n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644,
         n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652,
         n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660,
         n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668,
         n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676,
         n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
         n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692,
         n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700,
         n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708,
         n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716,
         n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724,
         n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732,
         n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
         n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748,
         n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756,
         n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764,
         n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772,
         n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780,
         n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788,
         n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796,
         n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
         n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812,
         n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820,
         n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
         n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836,
         n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844,
         n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852,
         n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860,
         n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868,
         n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876,
         n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884,
         n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892,
         n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900,
         n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908,
         n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916,
         n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924,
         n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932,
         n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940,
         n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948,
         n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956,
         n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964,
         n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972,
         n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980,
         n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988,
         n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996,
         n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
         n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012,
         n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020,
         n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028,
         n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036,
         n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044,
         n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052,
         n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060,
         n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068,
         n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076,
         n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084,
         n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092,
         n36093, n36094, n36095, n36096, n36098, n36099, n36100, n36101,
         n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109,
         n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117,
         n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125,
         n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133,
         n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141,
         n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149,
         n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157,
         n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165,
         n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173,
         n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181,
         n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189,
         n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197,
         n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205,
         n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213,
         n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221,
         n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229,
         n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237,
         n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245,
         n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253,
         n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261,
         n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269,
         n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277,
         n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285,
         n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293,
         n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301,
         n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309,
         n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317,
         n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325,
         n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333,
         n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341,
         n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349,
         n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357,
         n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365,
         n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373,
         n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381,
         n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389,
         n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397,
         n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405,
         n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413,
         n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421,
         n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429,
         n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437,
         n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445,
         n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453,
         n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461,
         n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469,
         n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477,
         n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485,
         n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493,
         n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501,
         n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509,
         n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517,
         n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525,
         n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533,
         n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541,
         n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549,
         n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557,
         n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565,
         n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573,
         n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581,
         n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589,
         n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597,
         n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605,
         n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613,
         n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621,
         n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629,
         n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637,
         n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645,
         n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653,
         n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661,
         n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669,
         n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677,
         n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685,
         n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693,
         n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701,
         n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709,
         n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717,
         n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725,
         n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733,
         n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741,
         n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749,
         n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757,
         n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765,
         n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773,
         n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781,
         n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789,
         n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797,
         n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805,
         n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813,
         n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821,
         n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829,
         n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837,
         n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845,
         n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853,
         n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861,
         n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869,
         n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877,
         n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885,
         n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893,
         n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
         n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909,
         n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917,
         n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925,
         n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933,
         n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941,
         n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949,
         n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957,
         n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965,
         n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973,
         n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981,
         n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989,
         n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997,
         n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005,
         n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013,
         n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021,
         n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029,
         n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037,
         n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
         n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053,
         n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061,
         n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069,
         n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077,
         n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085,
         n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093,
         n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101,
         n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109,
         n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
         n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125,
         n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133,
         n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141,
         n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149,
         n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157,
         n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165,
         n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173,
         n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181,
         n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189,
         n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197,
         n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205,
         n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213,
         n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221,
         n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229,
         n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237,
         n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245,
         n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253,
         n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261,
         n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269,
         n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277,
         n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285,
         n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293,
         n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301,
         n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309,
         n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317,
         n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325,
         n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333,
         n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341,
         n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349,
         n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357,
         n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365,
         n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373,
         n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381,
         n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389,
         n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397,
         n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405,
         n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413,
         n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421,
         n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429,
         n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437,
         n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445,
         n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453,
         n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461,
         n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469,
         n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477,
         n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485,
         n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493,
         n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501,
         n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509,
         n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517,
         n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525,
         n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533,
         n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541,
         n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549,
         n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557,
         n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565,
         n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573,
         n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581,
         n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589,
         n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597,
         n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605,
         n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613,
         n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621,
         n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629,
         n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637,
         n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645,
         n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653,
         n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661,
         n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669,
         n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677,
         n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685,
         n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693,
         n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701,
         n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709,
         n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717,
         n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725,
         n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733,
         n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741,
         n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749,
         n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757,
         n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765,
         n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773,
         n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781,
         n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789,
         n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797,
         n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805,
         n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813,
         n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821,
         n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829,
         n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837,
         n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845,
         n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853,
         n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861,
         n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869,
         n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877,
         n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885,
         n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893,
         n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901,
         n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909,
         n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917,
         n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925,
         n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933,
         n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941,
         n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949,
         n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957,
         n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965,
         n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973,
         n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981,
         n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989,
         n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997,
         n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005,
         n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013,
         n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021,
         n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029,
         n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037,
         n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045,
         n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053,
         n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061,
         n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069,
         n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077,
         n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085,
         n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093,
         n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101,
         n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109,
         n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117,
         n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125,
         n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133,
         n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141,
         n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149,
         n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157,
         n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165,
         n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173,
         n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181,
         n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189,
         n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197,
         n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205,
         n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213,
         n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221,
         n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229,
         n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237,
         n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245,
         n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253,
         n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261,
         n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269,
         n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277,
         n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285,
         n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293,
         n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301,
         n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309,
         n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317,
         n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325,
         n38326, n38327, n38328, n38329, n38330, n38331, n38332, n38333,
         n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341,
         n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349,
         n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357,
         n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365,
         n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373,
         n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381,
         n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389,
         n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397,
         n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405,
         n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413,
         n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421,
         n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429,
         n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437,
         n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445,
         n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453,
         n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461,
         n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469,
         n38470, n38471, n38472, n38473, n38474, n38475, n38476, n38477,
         n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485,
         n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493,
         n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501,
         n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509,
         n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517,
         n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525,
         n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533,
         n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541,
         n38542, n38543, n38544, n38545, n38546, n38547, n38548, n38549,
         n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
         n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565,
         n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573,
         n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581,
         n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589,
         n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597,
         n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605,
         n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613,
         n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621,
         n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629,
         n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637,
         n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645,
         n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653,
         n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661,
         n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669,
         n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677,
         n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685,
         n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693,
         n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701,
         n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709,
         n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717,
         n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725,
         n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733,
         n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741,
         n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749,
         n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757,
         n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765,
         n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
         n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781,
         n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789,
         n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797,
         n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805,
         n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813,
         n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821,
         n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829,
         n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837,
         n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845,
         n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853,
         n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861,
         n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869,
         n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877,
         n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885,
         n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893,
         n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901,
         n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909,
         n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917,
         n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925,
         n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933,
         n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941,
         n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949,
         n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957,
         n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965,
         n38966, n38967, n38968, n38969, n38970, n38971, n38972, n38973,
         n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981,
         n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989,
         n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997,
         n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005,
         n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013,
         n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021,
         n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029,
         n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037,
         n39038, n39039, n39040, n39041, n39042, n39043, n39044, n39045,
         n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053,
         n39054;
  wire   [6:0] xmem_addr;
  wire   [4:0] fmem_addr;
  wire   [6:0] load_xaddr_val;

  DFF_X1 \ctrl_conv_output_inst/conv_start_reg_reg  ( .D(
        \ctrl_conv_output_inst/N7 ), .CK(clk), .Q(
        \ctrl_conv_output_inst/conv_start_reg ) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n2850), .CK(clk), .Q(
        xmem_addr[0]), .QN(n39048) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n2849), .CK(clk), .Q(
        xmem_addr[1]), .QN(n39049) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n2848), .CK(clk), .Q(
        xmem_addr[2]), .QN(n38999) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[3]  ( .D(n2847), .CK(clk), .Q(
        xmem_addr[3]), .QN(n39044) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[4]  ( .D(n2846), .CK(clk), .Q(
        xmem_addr[4]), .QN(n39042) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[5]  ( .D(n2845), .CK(clk), .Q(
        xmem_addr[5]), .QN(n38998) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[6]  ( .D(n2844), .CK(clk), .Q(
        xmem_addr[6]), .QN(n39043) );
  DFF_X1 \xmem_inst/mem_reg[112][0]  ( .D(n1947), .CK(clk), .Q(
        \xmem_inst/mem[112][0] ) );
  DFF_X1 \xmem_inst/mem_reg[112][1]  ( .D(n1946), .CK(clk), .Q(
        \xmem_inst/mem[112][1] ) );
  DFF_X1 \xmem_inst/mem_reg[112][2]  ( .D(n1945), .CK(clk), .Q(
        \xmem_inst/mem[112][2] ) );
  DFF_X1 \xmem_inst/mem_reg[112][3]  ( .D(n1944), .CK(clk), .Q(
        \xmem_inst/mem[112][3] ) );
  DFF_X1 \xmem_inst/mem_reg[112][4]  ( .D(n1943), .CK(clk), .Q(
        \xmem_inst/mem[112][4] ) );
  DFF_X1 \xmem_inst/mem_reg[112][5]  ( .D(n1942), .CK(clk), .Q(
        \xmem_inst/mem[112][5] ) );
  DFF_X1 \xmem_inst/mem_reg[112][6]  ( .D(n1941), .CK(clk), .Q(
        \xmem_inst/mem[112][6] ) );
  DFF_X1 \xmem_inst/mem_reg[112][7]  ( .D(n1940), .CK(clk), .Q(
        \xmem_inst/mem[112][7] ) );
  DFF_X1 \xmem_inst/mem_reg[113][0]  ( .D(n1939), .CK(clk), .Q(
        \xmem_inst/mem[113][0] ) );
  DFF_X1 \xmem_inst/mem_reg[113][1]  ( .D(n1938), .CK(clk), .Q(
        \xmem_inst/mem[113][1] ) );
  DFF_X1 \xmem_inst/mem_reg[113][2]  ( .D(n1937), .CK(clk), .Q(
        \xmem_inst/mem[113][2] ) );
  DFF_X1 \xmem_inst/mem_reg[113][3]  ( .D(n1936), .CK(clk), .Q(
        \xmem_inst/mem[113][3] ) );
  DFF_X1 \xmem_inst/mem_reg[113][4]  ( .D(n1935), .CK(clk), .Q(
        \xmem_inst/mem[113][4] ) );
  DFF_X1 \xmem_inst/mem_reg[113][5]  ( .D(n1934), .CK(clk), .Q(
        \xmem_inst/mem[113][5] ) );
  DFF_X1 \xmem_inst/mem_reg[113][6]  ( .D(n1933), .CK(clk), .Q(
        \xmem_inst/mem[113][6] ) );
  DFF_X1 \xmem_inst/mem_reg[113][7]  ( .D(n1932), .CK(clk), .Q(
        \xmem_inst/mem[113][7] ) );
  DFF_X1 \xmem_inst/mem_reg[114][0]  ( .D(n1931), .CK(clk), .Q(
        \xmem_inst/mem[114][0] ) );
  DFF_X1 \xmem_inst/mem_reg[114][1]  ( .D(n1930), .CK(clk), .Q(
        \xmem_inst/mem[114][1] ) );
  DFF_X1 \xmem_inst/mem_reg[114][2]  ( .D(n1929), .CK(clk), .Q(
        \xmem_inst/mem[114][2] ) );
  DFF_X1 \xmem_inst/mem_reg[114][3]  ( .D(n1928), .CK(clk), .Q(
        \xmem_inst/mem[114][3] ) );
  DFF_X1 \xmem_inst/mem_reg[114][4]  ( .D(n1927), .CK(clk), .Q(
        \xmem_inst/mem[114][4] ) );
  DFF_X1 \xmem_inst/mem_reg[114][5]  ( .D(n1926), .CK(clk), .Q(
        \xmem_inst/mem[114][5] ) );
  DFF_X1 \xmem_inst/mem_reg[114][6]  ( .D(n1925), .CK(clk), .Q(
        \xmem_inst/mem[114][6] ) );
  DFF_X1 \xmem_inst/mem_reg[114][7]  ( .D(n1924), .CK(clk), .Q(
        \xmem_inst/mem[114][7] ) );
  DFF_X1 \xmem_inst/mem_reg[115][0]  ( .D(n1923), .CK(clk), .Q(
        \xmem_inst/mem[115][0] ) );
  DFF_X1 \xmem_inst/mem_reg[115][1]  ( .D(n1922), .CK(clk), .Q(
        \xmem_inst/mem[115][1] ) );
  DFF_X1 \xmem_inst/mem_reg[115][2]  ( .D(n1921), .CK(clk), .Q(
        \xmem_inst/mem[115][2] ) );
  DFF_X1 \xmem_inst/mem_reg[115][3]  ( .D(n1920), .CK(clk), .Q(
        \xmem_inst/mem[115][3] ) );
  DFF_X1 \xmem_inst/mem_reg[115][4]  ( .D(n1919), .CK(clk), .Q(
        \xmem_inst/mem[115][4] ) );
  DFF_X1 \xmem_inst/mem_reg[115][5]  ( .D(n1918), .CK(clk), .Q(
        \xmem_inst/mem[115][5] ) );
  DFF_X1 \xmem_inst/mem_reg[115][6]  ( .D(n1917), .CK(clk), .Q(
        \xmem_inst/mem[115][6] ) );
  DFF_X1 \xmem_inst/mem_reg[115][7]  ( .D(n1916), .CK(clk), .Q(
        \xmem_inst/mem[115][7] ) );
  DFF_X1 \xmem_inst/mem_reg[116][0]  ( .D(n1915), .CK(clk), .Q(
        \xmem_inst/mem[116][0] ) );
  DFF_X1 \xmem_inst/mem_reg[116][1]  ( .D(n1914), .CK(clk), .Q(
        \xmem_inst/mem[116][1] ) );
  DFF_X1 \xmem_inst/mem_reg[116][2]  ( .D(n1913), .CK(clk), .Q(
        \xmem_inst/mem[116][2] ) );
  DFF_X1 \xmem_inst/mem_reg[116][3]  ( .D(n1912), .CK(clk), .Q(
        \xmem_inst/mem[116][3] ) );
  DFF_X1 \xmem_inst/mem_reg[116][4]  ( .D(n1911), .CK(clk), .Q(
        \xmem_inst/mem[116][4] ) );
  DFF_X1 \xmem_inst/mem_reg[116][5]  ( .D(n1910), .CK(clk), .Q(
        \xmem_inst/mem[116][5] ) );
  DFF_X1 \xmem_inst/mem_reg[116][6]  ( .D(n1909), .CK(clk), .Q(
        \xmem_inst/mem[116][6] ) );
  DFF_X1 \xmem_inst/mem_reg[116][7]  ( .D(n1908), .CK(clk), .Q(
        \xmem_inst/mem[116][7] ) );
  DFF_X1 \xmem_inst/mem_reg[117][0]  ( .D(n1907), .CK(clk), .Q(
        \xmem_inst/mem[117][0] ) );
  DFF_X1 \xmem_inst/mem_reg[117][1]  ( .D(n1906), .CK(clk), .Q(
        \xmem_inst/mem[117][1] ) );
  DFF_X1 \xmem_inst/mem_reg[117][2]  ( .D(n1905), .CK(clk), .Q(
        \xmem_inst/mem[117][2] ) );
  DFF_X1 \xmem_inst/mem_reg[117][3]  ( .D(n1904), .CK(clk), .Q(
        \xmem_inst/mem[117][3] ) );
  DFF_X1 \xmem_inst/mem_reg[117][4]  ( .D(n1903), .CK(clk), .Q(
        \xmem_inst/mem[117][4] ) );
  DFF_X1 \xmem_inst/mem_reg[117][5]  ( .D(n1902), .CK(clk), .Q(
        \xmem_inst/mem[117][5] ) );
  DFF_X1 \xmem_inst/mem_reg[117][6]  ( .D(n1901), .CK(clk), .Q(
        \xmem_inst/mem[117][6] ) );
  DFF_X1 \xmem_inst/mem_reg[117][7]  ( .D(n1900), .CK(clk), .Q(
        \xmem_inst/mem[117][7] ) );
  DFF_X1 \xmem_inst/mem_reg[118][0]  ( .D(n1899), .CK(clk), .Q(
        \xmem_inst/mem[118][0] ) );
  DFF_X1 \xmem_inst/mem_reg[118][1]  ( .D(n1898), .CK(clk), .Q(
        \xmem_inst/mem[118][1] ) );
  DFF_X1 \xmem_inst/mem_reg[118][2]  ( .D(n1897), .CK(clk), .Q(
        \xmem_inst/mem[118][2] ) );
  DFF_X1 \xmem_inst/mem_reg[118][3]  ( .D(n1896), .CK(clk), .Q(
        \xmem_inst/mem[118][3] ) );
  DFF_X1 \xmem_inst/mem_reg[118][4]  ( .D(n1895), .CK(clk), .Q(
        \xmem_inst/mem[118][4] ) );
  DFF_X1 \xmem_inst/mem_reg[118][5]  ( .D(n1894), .CK(clk), .Q(
        \xmem_inst/mem[118][5] ) );
  DFF_X1 \xmem_inst/mem_reg[118][6]  ( .D(n1893), .CK(clk), .Q(
        \xmem_inst/mem[118][6] ) );
  DFF_X1 \xmem_inst/mem_reg[118][7]  ( .D(n1892), .CK(clk), .Q(
        \xmem_inst/mem[118][7] ) );
  DFF_X1 \xmem_inst/mem_reg[119][0]  ( .D(n1891), .CK(clk), .Q(
        \xmem_inst/mem[119][0] ) );
  DFF_X1 \xmem_inst/mem_reg[119][1]  ( .D(n1890), .CK(clk), .Q(
        \xmem_inst/mem[119][1] ) );
  DFF_X1 \xmem_inst/mem_reg[119][2]  ( .D(n1889), .CK(clk), .Q(
        \xmem_inst/mem[119][2] ) );
  DFF_X1 \xmem_inst/mem_reg[119][3]  ( .D(n1888), .CK(clk), .Q(
        \xmem_inst/mem[119][3] ) );
  DFF_X1 \xmem_inst/mem_reg[119][4]  ( .D(n1887), .CK(clk), .Q(
        \xmem_inst/mem[119][4] ) );
  DFF_X1 \xmem_inst/mem_reg[119][5]  ( .D(n1886), .CK(clk), .Q(
        \xmem_inst/mem[119][5] ) );
  DFF_X1 \xmem_inst/mem_reg[119][6]  ( .D(n1885), .CK(clk), .Q(
        \xmem_inst/mem[119][6] ) );
  DFF_X1 \xmem_inst/mem_reg[119][7]  ( .D(n1884), .CK(clk), .Q(
        \xmem_inst/mem[119][7] ) );
  DFF_X1 \xmem_inst/mem_reg[120][0]  ( .D(n1883), .CK(clk), .Q(
        \xmem_inst/mem[120][0] ) );
  DFF_X1 \xmem_inst/mem_reg[120][1]  ( .D(n1882), .CK(clk), .Q(
        \xmem_inst/mem[120][1] ) );
  DFF_X1 \xmem_inst/mem_reg[120][2]  ( .D(n1881), .CK(clk), .Q(
        \xmem_inst/mem[120][2] ) );
  DFF_X1 \xmem_inst/mem_reg[120][3]  ( .D(n1880), .CK(clk), .Q(
        \xmem_inst/mem[120][3] ) );
  DFF_X1 \xmem_inst/mem_reg[120][4]  ( .D(n1879), .CK(clk), .Q(
        \xmem_inst/mem[120][4] ) );
  DFF_X1 \xmem_inst/mem_reg[120][5]  ( .D(n1878), .CK(clk), .Q(
        \xmem_inst/mem[120][5] ) );
  DFF_X1 \xmem_inst/mem_reg[120][6]  ( .D(n1877), .CK(clk), .Q(
        \xmem_inst/mem[120][6] ) );
  DFF_X1 \xmem_inst/mem_reg[120][7]  ( .D(n1876), .CK(clk), .Q(
        \xmem_inst/mem[120][7] ) );
  DFF_X1 \xmem_inst/mem_reg[121][0]  ( .D(n1875), .CK(clk), .Q(
        \xmem_inst/mem[121][0] ) );
  DFF_X1 \xmem_inst/mem_reg[121][1]  ( .D(n1874), .CK(clk), .Q(
        \xmem_inst/mem[121][1] ) );
  DFF_X1 \xmem_inst/mem_reg[121][2]  ( .D(n1873), .CK(clk), .Q(
        \xmem_inst/mem[121][2] ) );
  DFF_X1 \xmem_inst/mem_reg[121][3]  ( .D(n1872), .CK(clk), .Q(
        \xmem_inst/mem[121][3] ) );
  DFF_X1 \xmem_inst/mem_reg[121][4]  ( .D(n1871), .CK(clk), .Q(
        \xmem_inst/mem[121][4] ) );
  DFF_X1 \xmem_inst/mem_reg[121][5]  ( .D(n1870), .CK(clk), .Q(
        \xmem_inst/mem[121][5] ) );
  DFF_X1 \xmem_inst/mem_reg[121][6]  ( .D(n1869), .CK(clk), .Q(
        \xmem_inst/mem[121][6] ) );
  DFF_X1 \xmem_inst/mem_reg[121][7]  ( .D(n1868), .CK(clk), .Q(
        \xmem_inst/mem[121][7] ) );
  DFF_X1 \xmem_inst/mem_reg[122][0]  ( .D(n1867), .CK(clk), .Q(
        \xmem_inst/mem[122][0] ) );
  DFF_X1 \xmem_inst/mem_reg[122][1]  ( .D(n1866), .CK(clk), .Q(
        \xmem_inst/mem[122][1] ) );
  DFF_X1 \xmem_inst/mem_reg[122][2]  ( .D(n1865), .CK(clk), .Q(
        \xmem_inst/mem[122][2] ) );
  DFF_X1 \xmem_inst/mem_reg[122][3]  ( .D(n1864), .CK(clk), .Q(
        \xmem_inst/mem[122][3] ) );
  DFF_X1 \xmem_inst/mem_reg[122][4]  ( .D(n1863), .CK(clk), .Q(
        \xmem_inst/mem[122][4] ) );
  DFF_X1 \xmem_inst/mem_reg[122][5]  ( .D(n1862), .CK(clk), .Q(
        \xmem_inst/mem[122][5] ) );
  DFF_X1 \xmem_inst/mem_reg[122][6]  ( .D(n1861), .CK(clk), .Q(
        \xmem_inst/mem[122][6] ) );
  DFF_X1 \xmem_inst/mem_reg[122][7]  ( .D(n1860), .CK(clk), .Q(
        \xmem_inst/mem[122][7] ) );
  DFF_X1 \xmem_inst/mem_reg[123][0]  ( .D(n1859), .CK(clk), .Q(
        \xmem_inst/mem[123][0] ) );
  DFF_X1 \xmem_inst/mem_reg[123][1]  ( .D(n1858), .CK(clk), .Q(
        \xmem_inst/mem[123][1] ) );
  DFF_X1 \xmem_inst/mem_reg[123][2]  ( .D(n1857), .CK(clk), .Q(
        \xmem_inst/mem[123][2] ) );
  DFF_X1 \xmem_inst/mem_reg[123][3]  ( .D(n1856), .CK(clk), .Q(
        \xmem_inst/mem[123][3] ) );
  DFF_X1 \xmem_inst/mem_reg[123][4]  ( .D(n1855), .CK(clk), .Q(
        \xmem_inst/mem[123][4] ) );
  DFF_X1 \xmem_inst/mem_reg[123][5]  ( .D(n1854), .CK(clk), .Q(
        \xmem_inst/mem[123][5] ) );
  DFF_X1 \xmem_inst/mem_reg[123][6]  ( .D(n1853), .CK(clk), .Q(
        \xmem_inst/mem[123][6] ) );
  DFF_X1 \xmem_inst/mem_reg[123][7]  ( .D(n1852), .CK(clk), .Q(
        \xmem_inst/mem[123][7] ) );
  DFF_X1 \xmem_inst/mem_reg[124][0]  ( .D(n1851), .CK(clk), .Q(
        \xmem_inst/mem[124][0] ) );
  DFF_X1 \xmem_inst/mem_reg[124][1]  ( .D(n1850), .CK(clk), .Q(
        \xmem_inst/mem[124][1] ) );
  DFF_X1 \xmem_inst/mem_reg[124][2]  ( .D(n1849), .CK(clk), .Q(
        \xmem_inst/mem[124][2] ) );
  DFF_X1 \xmem_inst/mem_reg[124][3]  ( .D(n1848), .CK(clk), .Q(
        \xmem_inst/mem[124][3] ) );
  DFF_X1 \xmem_inst/mem_reg[124][4]  ( .D(n1847), .CK(clk), .Q(
        \xmem_inst/mem[124][4] ) );
  DFF_X1 \xmem_inst/mem_reg[124][5]  ( .D(n1846), .CK(clk), .Q(
        \xmem_inst/mem[124][5] ) );
  DFF_X1 \xmem_inst/mem_reg[124][6]  ( .D(n1845), .CK(clk), .Q(
        \xmem_inst/mem[124][6] ) );
  DFF_X1 \xmem_inst/mem_reg[124][7]  ( .D(n1844), .CK(clk), .Q(
        \xmem_inst/mem[124][7] ) );
  DFF_X1 \xmem_inst/mem_reg[125][0]  ( .D(n1843), .CK(clk), .Q(
        \xmem_inst/mem[125][0] ) );
  DFF_X1 \xmem_inst/mem_reg[125][1]  ( .D(n1842), .CK(clk), .Q(
        \xmem_inst/mem[125][1] ) );
  DFF_X1 \xmem_inst/mem_reg[125][2]  ( .D(n1841), .CK(clk), .Q(
        \xmem_inst/mem[125][2] ) );
  DFF_X1 \xmem_inst/mem_reg[125][3]  ( .D(n1840), .CK(clk), .Q(
        \xmem_inst/mem[125][3] ) );
  DFF_X1 \xmem_inst/mem_reg[125][4]  ( .D(n1839), .CK(clk), .Q(
        \xmem_inst/mem[125][4] ) );
  DFF_X1 \xmem_inst/mem_reg[125][5]  ( .D(n1838), .CK(clk), .Q(
        \xmem_inst/mem[125][5] ) );
  DFF_X1 \xmem_inst/mem_reg[125][6]  ( .D(n1837), .CK(clk), .Q(
        \xmem_inst/mem[125][6] ) );
  DFF_X1 \xmem_inst/mem_reg[125][7]  ( .D(n1836), .CK(clk), .Q(
        \xmem_inst/mem[125][7] ) );
  DFF_X1 \xmem_inst/mem_reg[126][0]  ( .D(n1835), .CK(clk), .Q(
        \xmem_inst/mem[126][0] ) );
  DFF_X1 \xmem_inst/mem_reg[126][1]  ( .D(n1834), .CK(clk), .Q(
        \xmem_inst/mem[126][1] ) );
  DFF_X1 \xmem_inst/mem_reg[126][2]  ( .D(n1833), .CK(clk), .Q(
        \xmem_inst/mem[126][2] ) );
  DFF_X1 \xmem_inst/mem_reg[126][3]  ( .D(n1832), .CK(clk), .Q(
        \xmem_inst/mem[126][3] ) );
  DFF_X1 \xmem_inst/mem_reg[126][4]  ( .D(n1831), .CK(clk), .Q(
        \xmem_inst/mem[126][4] ) );
  DFF_X1 \xmem_inst/mem_reg[126][5]  ( .D(n1830), .CK(clk), .Q(
        \xmem_inst/mem[126][5] ) );
  DFF_X1 \xmem_inst/mem_reg[126][6]  ( .D(n1829), .CK(clk), .Q(
        \xmem_inst/mem[126][6] ) );
  DFF_X1 \xmem_inst/mem_reg[126][7]  ( .D(n1828), .CK(clk), .Q(
        \xmem_inst/mem[126][7] ) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n2851), .CK(clk), .Q(
        s_ready_x), .QN(n39051) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n2843), .CK(clk), .Q(
        \xmem_inst/mem[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n2842), .CK(clk), .Q(
        \xmem_inst/mem[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n2841), .CK(clk), .Q(
        \xmem_inst/mem[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n2840), .CK(clk), .Q(
        \xmem_inst/mem[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n2839), .CK(clk), .Q(
        \xmem_inst/mem[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n2838), .CK(clk), .Q(
        \xmem_inst/mem[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n2837), .CK(clk), .Q(
        \xmem_inst/mem[0][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n2836), .CK(clk), .Q(
        \xmem_inst/mem[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n2835), .CK(clk), .Q(
        \xmem_inst/mem[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n2834), .CK(clk), .Q(
        \xmem_inst/mem[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n2833), .CK(clk), .Q(
        \xmem_inst/mem[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n2832), .CK(clk), .Q(
        \xmem_inst/mem[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n2831), .CK(clk), .Q(
        \xmem_inst/mem[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n2830), .CK(clk), .Q(
        \xmem_inst/mem[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n2829), .CK(clk), .Q(
        \xmem_inst/mem[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n2828), .CK(clk), .Q(
        \xmem_inst/mem[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n2827), .CK(clk), .Q(
        \xmem_inst/mem[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n2826), .CK(clk), .Q(
        \xmem_inst/mem[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n2825), .CK(clk), .Q(
        \xmem_inst/mem[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n2824), .CK(clk), .Q(
        \xmem_inst/mem[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n2823), .CK(clk), .Q(
        \xmem_inst/mem[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n2822), .CK(clk), .Q(
        \xmem_inst/mem[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n2821), .CK(clk), .Q(
        \xmem_inst/mem[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n2820), .CK(clk), .Q(
        \xmem_inst/mem[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n2819), .CK(clk), .Q(
        \xmem_inst/mem[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n2818), .CK(clk), .Q(
        \xmem_inst/mem[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n2817), .CK(clk), .Q(
        \xmem_inst/mem[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n2816), .CK(clk), .Q(
        \xmem_inst/mem[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n2815), .CK(clk), .Q(
        \xmem_inst/mem[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n2814), .CK(clk), .Q(
        \xmem_inst/mem[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n2813), .CK(clk), .Q(
        \xmem_inst/mem[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n2812), .CK(clk), .Q(
        \xmem_inst/mem[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n2811), .CK(clk), .Q(
        \xmem_inst/mem[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n2810), .CK(clk), .Q(
        \xmem_inst/mem[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n2809), .CK(clk), .Q(
        \xmem_inst/mem[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n2808), .CK(clk), .Q(
        \xmem_inst/mem[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n2807), .CK(clk), .Q(
        \xmem_inst/mem[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n2806), .CK(clk), .Q(
        \xmem_inst/mem[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n2805), .CK(clk), .Q(
        \xmem_inst/mem[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n2804), .CK(clk), .Q(
        \xmem_inst/mem[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n2803), .CK(clk), .Q(
        \xmem_inst/mem[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n2802), .CK(clk), .Q(
        \xmem_inst/mem[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n2801), .CK(clk), .Q(
        \xmem_inst/mem[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n2800), .CK(clk), .Q(
        \xmem_inst/mem[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n2799), .CK(clk), .Q(
        \xmem_inst/mem[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n2798), .CK(clk), .Q(
        \xmem_inst/mem[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n2797), .CK(clk), .Q(
        \xmem_inst/mem[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n2796), .CK(clk), .Q(
        \xmem_inst/mem[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n2795), .CK(clk), .Q(
        \xmem_inst/mem[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n2794), .CK(clk), .Q(
        \xmem_inst/mem[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n2793), .CK(clk), .Q(
        \xmem_inst/mem[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n2792), .CK(clk), .Q(
        \xmem_inst/mem[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n2791), .CK(clk), .Q(
        \xmem_inst/mem[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n2790), .CK(clk), .Q(
        \xmem_inst/mem[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n2789), .CK(clk), .Q(
        \xmem_inst/mem[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n2788), .CK(clk), .Q(
        \xmem_inst/mem[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n2787), .CK(clk), .Q(
        \xmem_inst/mem[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n2786), .CK(clk), .Q(
        \xmem_inst/mem[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n2785), .CK(clk), .Q(
        \xmem_inst/mem[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n2784), .CK(clk), .Q(
        \xmem_inst/mem[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n2783), .CK(clk), .Q(
        \xmem_inst/mem[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n2782), .CK(clk), .Q(
        \xmem_inst/mem[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n2781), .CK(clk), .Q(
        \xmem_inst/mem[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n2780), .CK(clk), .Q(
        \xmem_inst/mem[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n2779), .CK(clk), .Q(
        \xmem_inst/mem[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n2778), .CK(clk), .Q(
        \xmem_inst/mem[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n2777), .CK(clk), .Q(
        \xmem_inst/mem[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n2776), .CK(clk), .Q(
        \xmem_inst/mem[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n2775), .CK(clk), .Q(
        \xmem_inst/mem[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n2774), .CK(clk), .Q(
        \xmem_inst/mem[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n2773), .CK(clk), .Q(
        \xmem_inst/mem[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n2772), .CK(clk), .Q(
        \xmem_inst/mem[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n2771), .CK(clk), .Q(
        \xmem_inst/mem[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n2770), .CK(clk), .Q(
        \xmem_inst/mem[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n2769), .CK(clk), .Q(
        \xmem_inst/mem[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n2768), .CK(clk), .Q(
        \xmem_inst/mem[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n2767), .CK(clk), .Q(
        \xmem_inst/mem[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n2766), .CK(clk), .Q(
        \xmem_inst/mem[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n2765), .CK(clk), .Q(
        \xmem_inst/mem[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n2764), .CK(clk), .Q(
        \xmem_inst/mem[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n2763), .CK(clk), .Q(
        \xmem_inst/mem[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n2762), .CK(clk), .Q(
        \xmem_inst/mem[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n2761), .CK(clk), .Q(
        \xmem_inst/mem[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n2760), .CK(clk), .Q(
        \xmem_inst/mem[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n2759), .CK(clk), .Q(
        \xmem_inst/mem[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n2758), .CK(clk), .Q(
        \xmem_inst/mem[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n2757), .CK(clk), .Q(
        \xmem_inst/mem[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n2756), .CK(clk), .Q(
        \xmem_inst/mem[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n2755), .CK(clk), .Q(
        \xmem_inst/mem[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n2754), .CK(clk), .Q(
        \xmem_inst/mem[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n2753), .CK(clk), .Q(
        \xmem_inst/mem[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n2752), .CK(clk), .Q(
        \xmem_inst/mem[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n2751), .CK(clk), .Q(
        \xmem_inst/mem[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n2750), .CK(clk), .Q(
        \xmem_inst/mem[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n2749), .CK(clk), .Q(
        \xmem_inst/mem[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n2748), .CK(clk), .Q(
        \xmem_inst/mem[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n2747), .CK(clk), .Q(
        \xmem_inst/mem[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n2746), .CK(clk), .Q(
        \xmem_inst/mem[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n2745), .CK(clk), .Q(
        \xmem_inst/mem[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n2744), .CK(clk), .Q(
        \xmem_inst/mem[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n2743), .CK(clk), .Q(
        \xmem_inst/mem[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n2742), .CK(clk), .Q(
        \xmem_inst/mem[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n2741), .CK(clk), .Q(
        \xmem_inst/mem[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n2740), .CK(clk), .Q(
        \xmem_inst/mem[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n2739), .CK(clk), .Q(
        \xmem_inst/mem[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n2738), .CK(clk), .Q(
        \xmem_inst/mem[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n2737), .CK(clk), .Q(
        \xmem_inst/mem[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n2736), .CK(clk), .Q(
        \xmem_inst/mem[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n2735), .CK(clk), .Q(
        \xmem_inst/mem[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n2734), .CK(clk), .Q(
        \xmem_inst/mem[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n2733), .CK(clk), .Q(
        \xmem_inst/mem[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n2732), .CK(clk), .Q(
        \xmem_inst/mem[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n2731), .CK(clk), .Q(
        \xmem_inst/mem[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n2730), .CK(clk), .Q(
        \xmem_inst/mem[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n2729), .CK(clk), .Q(
        \xmem_inst/mem[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n2728), .CK(clk), .Q(
        \xmem_inst/mem[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n2727), .CK(clk), .Q(
        \xmem_inst/mem[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n2726), .CK(clk), .Q(
        \xmem_inst/mem[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n2725), .CK(clk), .Q(
        \xmem_inst/mem[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n2724), .CK(clk), .Q(
        \xmem_inst/mem[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n2723), .CK(clk), .Q(
        \xmem_inst/mem[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n2722), .CK(clk), .Q(
        \xmem_inst/mem[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n2721), .CK(clk), .Q(
        \xmem_inst/mem[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n2720), .CK(clk), .Q(
        \xmem_inst/mem[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n2719), .CK(clk), .Q(
        \xmem_inst/mem[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n2718), .CK(clk), .Q(
        \xmem_inst/mem[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n2717), .CK(clk), .Q(
        \xmem_inst/mem[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n2716), .CK(clk), .Q(
        \xmem_inst/mem[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n2715), .CK(clk), .Q(
        \xmem_inst/mem[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n2714), .CK(clk), .Q(
        \xmem_inst/mem[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n2713), .CK(clk), .Q(
        \xmem_inst/mem[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n2712), .CK(clk), .Q(
        \xmem_inst/mem[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n2711), .CK(clk), .Q(
        \xmem_inst/mem[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n2710), .CK(clk), .Q(
        \xmem_inst/mem[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n2709), .CK(clk), .Q(
        \xmem_inst/mem[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n2708), .CK(clk), .Q(
        \xmem_inst/mem[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n2707), .CK(clk), .Q(
        \xmem_inst/mem[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n2706), .CK(clk), .Q(
        \xmem_inst/mem[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n2705), .CK(clk), .Q(
        \xmem_inst/mem[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n2704), .CK(clk), .Q(
        \xmem_inst/mem[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n2703), .CK(clk), .Q(
        \xmem_inst/mem[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n2702), .CK(clk), .Q(
        \xmem_inst/mem[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n2701), .CK(clk), .Q(
        \xmem_inst/mem[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n2700), .CK(clk), .Q(
        \xmem_inst/mem[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n2699), .CK(clk), .Q(
        \xmem_inst/mem[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n2698), .CK(clk), .Q(
        \xmem_inst/mem[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n2697), .CK(clk), .Q(
        \xmem_inst/mem[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n2696), .CK(clk), .Q(
        \xmem_inst/mem[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n2695), .CK(clk), .Q(
        \xmem_inst/mem[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n2694), .CK(clk), .Q(
        \xmem_inst/mem[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n2693), .CK(clk), .Q(
        \xmem_inst/mem[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n2692), .CK(clk), .Q(
        \xmem_inst/mem[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n2691), .CK(clk), .Q(
        \xmem_inst/mem[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n2690), .CK(clk), .Q(
        \xmem_inst/mem[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n2689), .CK(clk), .Q(
        \xmem_inst/mem[19][2] ) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n2688), .CK(clk), .Q(
        \xmem_inst/mem[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n2687), .CK(clk), .Q(
        \xmem_inst/mem[19][4] ) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n2686), .CK(clk), .Q(
        \xmem_inst/mem[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n2685), .CK(clk), .Q(
        \xmem_inst/mem[19][6] ) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n2684), .CK(clk), .Q(
        \xmem_inst/mem[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[20][0]  ( .D(n2683), .CK(clk), .Q(
        \xmem_inst/mem[20][0] ) );
  DFF_X1 \xmem_inst/mem_reg[20][1]  ( .D(n2682), .CK(clk), .Q(
        \xmem_inst/mem[20][1] ) );
  DFF_X1 \xmem_inst/mem_reg[20][2]  ( .D(n2681), .CK(clk), .Q(
        \xmem_inst/mem[20][2] ) );
  DFF_X1 \xmem_inst/mem_reg[20][3]  ( .D(n2680), .CK(clk), .Q(
        \xmem_inst/mem[20][3] ) );
  DFF_X1 \xmem_inst/mem_reg[20][4]  ( .D(n2679), .CK(clk), .Q(
        \xmem_inst/mem[20][4] ) );
  DFF_X1 \xmem_inst/mem_reg[20][5]  ( .D(n2678), .CK(clk), .Q(
        \xmem_inst/mem[20][5] ) );
  DFF_X1 \xmem_inst/mem_reg[20][6]  ( .D(n2677), .CK(clk), .Q(
        \xmem_inst/mem[20][6] ) );
  DFF_X1 \xmem_inst/mem_reg[20][7]  ( .D(n2676), .CK(clk), .Q(
        \xmem_inst/mem[20][7] ) );
  DFF_X1 \xmem_inst/mem_reg[21][0]  ( .D(n2675), .CK(clk), .Q(
        \xmem_inst/mem[21][0] ) );
  DFF_X1 \xmem_inst/mem_reg[21][1]  ( .D(n2674), .CK(clk), .Q(
        \xmem_inst/mem[21][1] ) );
  DFF_X1 \xmem_inst/mem_reg[21][2]  ( .D(n2673), .CK(clk), .Q(
        \xmem_inst/mem[21][2] ) );
  DFF_X1 \xmem_inst/mem_reg[21][3]  ( .D(n2672), .CK(clk), .Q(
        \xmem_inst/mem[21][3] ) );
  DFF_X1 \xmem_inst/mem_reg[21][4]  ( .D(n2671), .CK(clk), .Q(
        \xmem_inst/mem[21][4] ) );
  DFF_X1 \xmem_inst/mem_reg[21][5]  ( .D(n2670), .CK(clk), .Q(
        \xmem_inst/mem[21][5] ) );
  DFF_X1 \xmem_inst/mem_reg[21][6]  ( .D(n2669), .CK(clk), .Q(
        \xmem_inst/mem[21][6] ) );
  DFF_X1 \xmem_inst/mem_reg[21][7]  ( .D(n2668), .CK(clk), .Q(
        \xmem_inst/mem[21][7] ) );
  DFF_X1 \xmem_inst/mem_reg[22][0]  ( .D(n2667), .CK(clk), .Q(
        \xmem_inst/mem[22][0] ) );
  DFF_X1 \xmem_inst/mem_reg[22][1]  ( .D(n2666), .CK(clk), .Q(
        \xmem_inst/mem[22][1] ) );
  DFF_X1 \xmem_inst/mem_reg[22][2]  ( .D(n2665), .CK(clk), .Q(
        \xmem_inst/mem[22][2] ) );
  DFF_X1 \xmem_inst/mem_reg[22][3]  ( .D(n2664), .CK(clk), .Q(
        \xmem_inst/mem[22][3] ) );
  DFF_X1 \xmem_inst/mem_reg[22][4]  ( .D(n2663), .CK(clk), .Q(
        \xmem_inst/mem[22][4] ) );
  DFF_X1 \xmem_inst/mem_reg[22][5]  ( .D(n2662), .CK(clk), .Q(
        \xmem_inst/mem[22][5] ) );
  DFF_X1 \xmem_inst/mem_reg[22][6]  ( .D(n2661), .CK(clk), .Q(
        \xmem_inst/mem[22][6] ) );
  DFF_X1 \xmem_inst/mem_reg[22][7]  ( .D(n2660), .CK(clk), .Q(
        \xmem_inst/mem[22][7] ) );
  DFF_X1 \xmem_inst/mem_reg[23][0]  ( .D(n2659), .CK(clk), .Q(
        \xmem_inst/mem[23][0] ) );
  DFF_X1 \xmem_inst/mem_reg[23][1]  ( .D(n2658), .CK(clk), .Q(
        \xmem_inst/mem[23][1] ) );
  DFF_X1 \xmem_inst/mem_reg[23][2]  ( .D(n2657), .CK(clk), .Q(
        \xmem_inst/mem[23][2] ) );
  DFF_X1 \xmem_inst/mem_reg[23][3]  ( .D(n2656), .CK(clk), .Q(
        \xmem_inst/mem[23][3] ) );
  DFF_X1 \xmem_inst/mem_reg[23][4]  ( .D(n2655), .CK(clk), .Q(
        \xmem_inst/mem[23][4] ) );
  DFF_X1 \xmem_inst/mem_reg[23][5]  ( .D(n2654), .CK(clk), .Q(
        \xmem_inst/mem[23][5] ) );
  DFF_X1 \xmem_inst/mem_reg[23][6]  ( .D(n2653), .CK(clk), .Q(
        \xmem_inst/mem[23][6] ) );
  DFF_X1 \xmem_inst/mem_reg[23][7]  ( .D(n2652), .CK(clk), .Q(
        \xmem_inst/mem[23][7] ) );
  DFF_X1 \xmem_inst/mem_reg[24][0]  ( .D(n2651), .CK(clk), .Q(
        \xmem_inst/mem[24][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][1]  ( .D(n2650), .CK(clk), .Q(
        \xmem_inst/mem[24][1] ) );
  DFF_X1 \xmem_inst/mem_reg[24][2]  ( .D(n2649), .CK(clk), .Q(
        \xmem_inst/mem[24][2] ) );
  DFF_X1 \xmem_inst/mem_reg[24][3]  ( .D(n2648), .CK(clk), .Q(
        \xmem_inst/mem[24][3] ) );
  DFF_X1 \xmem_inst/mem_reg[24][4]  ( .D(n2647), .CK(clk), .Q(
        \xmem_inst/mem[24][4] ) );
  DFF_X1 \xmem_inst/mem_reg[24][5]  ( .D(n2646), .CK(clk), .Q(
        \xmem_inst/mem[24][5] ) );
  DFF_X1 \xmem_inst/mem_reg[24][6]  ( .D(n2645), .CK(clk), .Q(
        \xmem_inst/mem[24][6] ) );
  DFF_X1 \xmem_inst/mem_reg[24][7]  ( .D(n2644), .CK(clk), .Q(
        \xmem_inst/mem[24][7] ) );
  DFF_X1 \xmem_inst/mem_reg[25][0]  ( .D(n2643), .CK(clk), .Q(
        \xmem_inst/mem[25][0] ) );
  DFF_X1 \xmem_inst/mem_reg[25][1]  ( .D(n2642), .CK(clk), .Q(
        \xmem_inst/mem[25][1] ) );
  DFF_X1 \xmem_inst/mem_reg[25][2]  ( .D(n2641), .CK(clk), .Q(
        \xmem_inst/mem[25][2] ) );
  DFF_X1 \xmem_inst/mem_reg[25][3]  ( .D(n2640), .CK(clk), .Q(
        \xmem_inst/mem[25][3] ) );
  DFF_X1 \xmem_inst/mem_reg[25][4]  ( .D(n2639), .CK(clk), .Q(
        \xmem_inst/mem[25][4] ) );
  DFF_X1 \xmem_inst/mem_reg[25][5]  ( .D(n2638), .CK(clk), .Q(
        \xmem_inst/mem[25][5] ) );
  DFF_X1 \xmem_inst/mem_reg[25][6]  ( .D(n2637), .CK(clk), .Q(
        \xmem_inst/mem[25][6] ) );
  DFF_X1 \xmem_inst/mem_reg[25][7]  ( .D(n2636), .CK(clk), .Q(
        \xmem_inst/mem[25][7] ) );
  DFF_X1 \xmem_inst/mem_reg[26][0]  ( .D(n2635), .CK(clk), .Q(
        \xmem_inst/mem[26][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][1]  ( .D(n2634), .CK(clk), .Q(
        \xmem_inst/mem[26][1] ) );
  DFF_X1 \xmem_inst/mem_reg[26][2]  ( .D(n2633), .CK(clk), .Q(
        \xmem_inst/mem[26][2] ) );
  DFF_X1 \xmem_inst/mem_reg[26][3]  ( .D(n2632), .CK(clk), .Q(
        \xmem_inst/mem[26][3] ) );
  DFF_X1 \xmem_inst/mem_reg[26][4]  ( .D(n2631), .CK(clk), .Q(
        \xmem_inst/mem[26][4] ) );
  DFF_X1 \xmem_inst/mem_reg[26][5]  ( .D(n2630), .CK(clk), .Q(
        \xmem_inst/mem[26][5] ) );
  DFF_X1 \xmem_inst/mem_reg[26][6]  ( .D(n2629), .CK(clk), .Q(
        \xmem_inst/mem[26][6] ) );
  DFF_X1 \xmem_inst/mem_reg[26][7]  ( .D(n2628), .CK(clk), .Q(
        \xmem_inst/mem[26][7] ) );
  DFF_X1 \xmem_inst/mem_reg[27][0]  ( .D(n2627), .CK(clk), .Q(
        \xmem_inst/mem[27][0] ) );
  DFF_X1 \xmem_inst/mem_reg[27][1]  ( .D(n2626), .CK(clk), .Q(
        \xmem_inst/mem[27][1] ) );
  DFF_X1 \xmem_inst/mem_reg[27][2]  ( .D(n2625), .CK(clk), .Q(
        \xmem_inst/mem[27][2] ) );
  DFF_X1 \xmem_inst/mem_reg[27][3]  ( .D(n2624), .CK(clk), .Q(
        \xmem_inst/mem[27][3] ) );
  DFF_X1 \xmem_inst/mem_reg[27][4]  ( .D(n2623), .CK(clk), .Q(
        \xmem_inst/mem[27][4] ) );
  DFF_X1 \xmem_inst/mem_reg[27][5]  ( .D(n2622), .CK(clk), .Q(
        \xmem_inst/mem[27][5] ) );
  DFF_X1 \xmem_inst/mem_reg[27][6]  ( .D(n2621), .CK(clk), .Q(
        \xmem_inst/mem[27][6] ) );
  DFF_X1 \xmem_inst/mem_reg[27][7]  ( .D(n2620), .CK(clk), .Q(
        \xmem_inst/mem[27][7] ) );
  DFF_X1 \xmem_inst/mem_reg[28][0]  ( .D(n2619), .CK(clk), .Q(
        \xmem_inst/mem[28][0] ) );
  DFF_X1 \xmem_inst/mem_reg[28][1]  ( .D(n2618), .CK(clk), .Q(
        \xmem_inst/mem[28][1] ) );
  DFF_X1 \xmem_inst/mem_reg[28][2]  ( .D(n2617), .CK(clk), .Q(
        \xmem_inst/mem[28][2] ) );
  DFF_X1 \xmem_inst/mem_reg[28][3]  ( .D(n2616), .CK(clk), .Q(
        \xmem_inst/mem[28][3] ) );
  DFF_X1 \xmem_inst/mem_reg[28][4]  ( .D(n2615), .CK(clk), .Q(
        \xmem_inst/mem[28][4] ) );
  DFF_X1 \xmem_inst/mem_reg[28][5]  ( .D(n2614), .CK(clk), .Q(
        \xmem_inst/mem[28][5] ) );
  DFF_X1 \xmem_inst/mem_reg[28][6]  ( .D(n2613), .CK(clk), .Q(
        \xmem_inst/mem[28][6] ) );
  DFF_X1 \xmem_inst/mem_reg[28][7]  ( .D(n2612), .CK(clk), .Q(
        \xmem_inst/mem[28][7] ) );
  DFF_X1 \xmem_inst/mem_reg[29][0]  ( .D(n2611), .CK(clk), .Q(
        \xmem_inst/mem[29][0] ) );
  DFF_X1 \xmem_inst/mem_reg[29][1]  ( .D(n2610), .CK(clk), .Q(
        \xmem_inst/mem[29][1] ) );
  DFF_X1 \xmem_inst/mem_reg[29][2]  ( .D(n2609), .CK(clk), .Q(
        \xmem_inst/mem[29][2] ) );
  DFF_X1 \xmem_inst/mem_reg[29][3]  ( .D(n2608), .CK(clk), .Q(
        \xmem_inst/mem[29][3] ) );
  DFF_X1 \xmem_inst/mem_reg[29][4]  ( .D(n2607), .CK(clk), .Q(
        \xmem_inst/mem[29][4] ) );
  DFF_X1 \xmem_inst/mem_reg[29][5]  ( .D(n2606), .CK(clk), .Q(
        \xmem_inst/mem[29][5] ) );
  DFF_X1 \xmem_inst/mem_reg[29][6]  ( .D(n2605), .CK(clk), .Q(
        \xmem_inst/mem[29][6] ) );
  DFF_X1 \xmem_inst/mem_reg[29][7]  ( .D(n2604), .CK(clk), .Q(
        \xmem_inst/mem[29][7] ) );
  DFF_X1 \xmem_inst/mem_reg[30][0]  ( .D(n2603), .CK(clk), .Q(
        \xmem_inst/mem[30][0] ) );
  DFF_X1 \xmem_inst/mem_reg[30][1]  ( .D(n2602), .CK(clk), .Q(
        \xmem_inst/mem[30][1] ) );
  DFF_X1 \xmem_inst/mem_reg[30][2]  ( .D(n2601), .CK(clk), .Q(
        \xmem_inst/mem[30][2] ) );
  DFF_X1 \xmem_inst/mem_reg[30][3]  ( .D(n2600), .CK(clk), .Q(
        \xmem_inst/mem[30][3] ) );
  DFF_X1 \xmem_inst/mem_reg[30][4]  ( .D(n2599), .CK(clk), .Q(
        \xmem_inst/mem[30][4] ) );
  DFF_X1 \xmem_inst/mem_reg[30][5]  ( .D(n2598), .CK(clk), .Q(
        \xmem_inst/mem[30][5] ) );
  DFF_X1 \xmem_inst/mem_reg[30][6]  ( .D(n2597), .CK(clk), .Q(
        \xmem_inst/mem[30][6] ) );
  DFF_X1 \xmem_inst/mem_reg[30][7]  ( .D(n2596), .CK(clk), .Q(
        \xmem_inst/mem[30][7] ) );
  DFF_X1 \xmem_inst/mem_reg[31][0]  ( .D(n2595), .CK(clk), .Q(
        \xmem_inst/mem[31][0] ) );
  DFF_X1 \xmem_inst/mem_reg[31][1]  ( .D(n2594), .CK(clk), .Q(
        \xmem_inst/mem[31][1] ) );
  DFF_X1 \xmem_inst/mem_reg[31][2]  ( .D(n2593), .CK(clk), .Q(
        \xmem_inst/mem[31][2] ) );
  DFF_X1 \xmem_inst/mem_reg[31][3]  ( .D(n2592), .CK(clk), .Q(
        \xmem_inst/mem[31][3] ) );
  DFF_X1 \xmem_inst/mem_reg[31][4]  ( .D(n2591), .CK(clk), .Q(
        \xmem_inst/mem[31][4] ) );
  DFF_X1 \xmem_inst/mem_reg[31][5]  ( .D(n2590), .CK(clk), .Q(
        \xmem_inst/mem[31][5] ) );
  DFF_X1 \xmem_inst/mem_reg[31][6]  ( .D(n2589), .CK(clk), .Q(
        \xmem_inst/mem[31][6] ) );
  DFF_X1 \xmem_inst/mem_reg[31][7]  ( .D(n2588), .CK(clk), .Q(
        \xmem_inst/mem[31][7] ) );
  DFF_X1 \xmem_inst/mem_reg[32][0]  ( .D(n2587), .CK(clk), .Q(
        \xmem_inst/mem[32][0] ) );
  DFF_X1 \xmem_inst/mem_reg[32][1]  ( .D(n2586), .CK(clk), .Q(
        \xmem_inst/mem[32][1] ) );
  DFF_X1 \xmem_inst/mem_reg[32][2]  ( .D(n2585), .CK(clk), .Q(
        \xmem_inst/mem[32][2] ) );
  DFF_X1 \xmem_inst/mem_reg[32][3]  ( .D(n2584), .CK(clk), .Q(
        \xmem_inst/mem[32][3] ) );
  DFF_X1 \xmem_inst/mem_reg[32][4]  ( .D(n2583), .CK(clk), .Q(
        \xmem_inst/mem[32][4] ) );
  DFF_X1 \xmem_inst/mem_reg[32][5]  ( .D(n2582), .CK(clk), .Q(
        \xmem_inst/mem[32][5] ) );
  DFF_X1 \xmem_inst/mem_reg[32][6]  ( .D(n2581), .CK(clk), .Q(
        \xmem_inst/mem[32][6] ) );
  DFF_X1 \xmem_inst/mem_reg[32][7]  ( .D(n2580), .CK(clk), .Q(
        \xmem_inst/mem[32][7] ) );
  DFF_X1 \xmem_inst/mem_reg[33][0]  ( .D(n2579), .CK(clk), .Q(
        \xmem_inst/mem[33][0] ) );
  DFF_X1 \xmem_inst/mem_reg[33][1]  ( .D(n2578), .CK(clk), .Q(
        \xmem_inst/mem[33][1] ) );
  DFF_X1 \xmem_inst/mem_reg[33][2]  ( .D(n2577), .CK(clk), .Q(
        \xmem_inst/mem[33][2] ) );
  DFF_X1 \xmem_inst/mem_reg[33][3]  ( .D(n2576), .CK(clk), .Q(
        \xmem_inst/mem[33][3] ) );
  DFF_X1 \xmem_inst/mem_reg[33][4]  ( .D(n2575), .CK(clk), .Q(
        \xmem_inst/mem[33][4] ) );
  DFF_X1 \xmem_inst/mem_reg[33][5]  ( .D(n2574), .CK(clk), .Q(
        \xmem_inst/mem[33][5] ) );
  DFF_X1 \xmem_inst/mem_reg[33][6]  ( .D(n2573), .CK(clk), .Q(
        \xmem_inst/mem[33][6] ) );
  DFF_X1 \xmem_inst/mem_reg[33][7]  ( .D(n2572), .CK(clk), .Q(
        \xmem_inst/mem[33][7] ) );
  DFF_X1 \xmem_inst/mem_reg[34][0]  ( .D(n2571), .CK(clk), .Q(
        \xmem_inst/mem[34][0] ) );
  DFF_X1 \xmem_inst/mem_reg[34][1]  ( .D(n2570), .CK(clk), .Q(
        \xmem_inst/mem[34][1] ) );
  DFF_X1 \xmem_inst/mem_reg[34][2]  ( .D(n2569), .CK(clk), .Q(
        \xmem_inst/mem[34][2] ) );
  DFF_X1 \xmem_inst/mem_reg[34][3]  ( .D(n2568), .CK(clk), .Q(
        \xmem_inst/mem[34][3] ) );
  DFF_X1 \xmem_inst/mem_reg[34][4]  ( .D(n2567), .CK(clk), .Q(
        \xmem_inst/mem[34][4] ) );
  DFF_X1 \xmem_inst/mem_reg[34][5]  ( .D(n2566), .CK(clk), .Q(
        \xmem_inst/mem[34][5] ) );
  DFF_X1 \xmem_inst/mem_reg[34][6]  ( .D(n2565), .CK(clk), .Q(
        \xmem_inst/mem[34][6] ) );
  DFF_X1 \xmem_inst/mem_reg[34][7]  ( .D(n2564), .CK(clk), .Q(
        \xmem_inst/mem[34][7] ) );
  DFF_X1 \xmem_inst/mem_reg[35][0]  ( .D(n2563), .CK(clk), .Q(
        \xmem_inst/mem[35][0] ) );
  DFF_X1 \xmem_inst/mem_reg[35][1]  ( .D(n2562), .CK(clk), .Q(
        \xmem_inst/mem[35][1] ) );
  DFF_X1 \xmem_inst/mem_reg[35][2]  ( .D(n2561), .CK(clk), .Q(
        \xmem_inst/mem[35][2] ) );
  DFF_X1 \xmem_inst/mem_reg[35][3]  ( .D(n2560), .CK(clk), .Q(
        \xmem_inst/mem[35][3] ) );
  DFF_X1 \xmem_inst/mem_reg[35][4]  ( .D(n2559), .CK(clk), .Q(
        \xmem_inst/mem[35][4] ) );
  DFF_X1 \xmem_inst/mem_reg[35][5]  ( .D(n2558), .CK(clk), .Q(
        \xmem_inst/mem[35][5] ) );
  DFF_X1 \xmem_inst/mem_reg[35][6]  ( .D(n2557), .CK(clk), .Q(
        \xmem_inst/mem[35][6] ) );
  DFF_X1 \xmem_inst/mem_reg[35][7]  ( .D(n2556), .CK(clk), .Q(
        \xmem_inst/mem[35][7] ) );
  DFF_X1 \xmem_inst/mem_reg[36][0]  ( .D(n2555), .CK(clk), .Q(
        \xmem_inst/mem[36][0] ) );
  DFF_X1 \xmem_inst/mem_reg[36][1]  ( .D(n2554), .CK(clk), .Q(
        \xmem_inst/mem[36][1] ) );
  DFF_X1 \xmem_inst/mem_reg[36][2]  ( .D(n2553), .CK(clk), .Q(
        \xmem_inst/mem[36][2] ) );
  DFF_X1 \xmem_inst/mem_reg[36][3]  ( .D(n2552), .CK(clk), .Q(
        \xmem_inst/mem[36][3] ) );
  DFF_X1 \xmem_inst/mem_reg[36][4]  ( .D(n2551), .CK(clk), .Q(
        \xmem_inst/mem[36][4] ) );
  DFF_X1 \xmem_inst/mem_reg[36][5]  ( .D(n2550), .CK(clk), .Q(
        \xmem_inst/mem[36][5] ) );
  DFF_X1 \xmem_inst/mem_reg[36][6]  ( .D(n2549), .CK(clk), .Q(
        \xmem_inst/mem[36][6] ) );
  DFF_X1 \xmem_inst/mem_reg[36][7]  ( .D(n2548), .CK(clk), .Q(
        \xmem_inst/mem[36][7] ) );
  DFF_X1 \xmem_inst/mem_reg[37][0]  ( .D(n2547), .CK(clk), .Q(
        \xmem_inst/mem[37][0] ) );
  DFF_X1 \xmem_inst/mem_reg[37][1]  ( .D(n2546), .CK(clk), .Q(
        \xmem_inst/mem[37][1] ) );
  DFF_X1 \xmem_inst/mem_reg[37][2]  ( .D(n2545), .CK(clk), .Q(
        \xmem_inst/mem[37][2] ) );
  DFF_X1 \xmem_inst/mem_reg[37][3]  ( .D(n2544), .CK(clk), .Q(
        \xmem_inst/mem[37][3] ) );
  DFF_X1 \xmem_inst/mem_reg[37][4]  ( .D(n2543), .CK(clk), .Q(
        \xmem_inst/mem[37][4] ) );
  DFF_X1 \xmem_inst/mem_reg[37][5]  ( .D(n2542), .CK(clk), .Q(
        \xmem_inst/mem[37][5] ) );
  DFF_X1 \xmem_inst/mem_reg[37][6]  ( .D(n2541), .CK(clk), .Q(
        \xmem_inst/mem[37][6] ) );
  DFF_X1 \xmem_inst/mem_reg[37][7]  ( .D(n2540), .CK(clk), .Q(
        \xmem_inst/mem[37][7] ) );
  DFF_X1 \xmem_inst/mem_reg[38][0]  ( .D(n2539), .CK(clk), .Q(
        \xmem_inst/mem[38][0] ) );
  DFF_X1 \xmem_inst/mem_reg[38][1]  ( .D(n2538), .CK(clk), .Q(
        \xmem_inst/mem[38][1] ) );
  DFF_X1 \xmem_inst/mem_reg[38][2]  ( .D(n2537), .CK(clk), .Q(
        \xmem_inst/mem[38][2] ) );
  DFF_X1 \xmem_inst/mem_reg[38][3]  ( .D(n2536), .CK(clk), .Q(
        \xmem_inst/mem[38][3] ) );
  DFF_X1 \xmem_inst/mem_reg[38][4]  ( .D(n2535), .CK(clk), .Q(
        \xmem_inst/mem[38][4] ) );
  DFF_X1 \xmem_inst/mem_reg[38][5]  ( .D(n2534), .CK(clk), .Q(
        \xmem_inst/mem[38][5] ) );
  DFF_X1 \xmem_inst/mem_reg[38][6]  ( .D(n2533), .CK(clk), .Q(
        \xmem_inst/mem[38][6] ) );
  DFF_X1 \xmem_inst/mem_reg[38][7]  ( .D(n2532), .CK(clk), .Q(
        \xmem_inst/mem[38][7] ) );
  DFF_X1 \xmem_inst/mem_reg[39][0]  ( .D(n2531), .CK(clk), .Q(
        \xmem_inst/mem[39][0] ) );
  DFF_X1 \xmem_inst/mem_reg[39][1]  ( .D(n2530), .CK(clk), .Q(
        \xmem_inst/mem[39][1] ) );
  DFF_X1 \xmem_inst/mem_reg[39][2]  ( .D(n2529), .CK(clk), .Q(
        \xmem_inst/mem[39][2] ) );
  DFF_X1 \xmem_inst/mem_reg[39][3]  ( .D(n2528), .CK(clk), .Q(
        \xmem_inst/mem[39][3] ) );
  DFF_X1 \xmem_inst/mem_reg[39][4]  ( .D(n2527), .CK(clk), .Q(
        \xmem_inst/mem[39][4] ) );
  DFF_X1 \xmem_inst/mem_reg[39][5]  ( .D(n2526), .CK(clk), .Q(
        \xmem_inst/mem[39][5] ) );
  DFF_X1 \xmem_inst/mem_reg[39][6]  ( .D(n2525), .CK(clk), .Q(
        \xmem_inst/mem[39][6] ) );
  DFF_X1 \xmem_inst/mem_reg[39][7]  ( .D(n2524), .CK(clk), .Q(
        \xmem_inst/mem[39][7] ) );
  DFF_X1 \xmem_inst/mem_reg[40][0]  ( .D(n2523), .CK(clk), .Q(
        \xmem_inst/mem[40][0] ) );
  DFF_X1 \xmem_inst/mem_reg[40][1]  ( .D(n2522), .CK(clk), .Q(
        \xmem_inst/mem[40][1] ) );
  DFF_X1 \xmem_inst/mem_reg[40][2]  ( .D(n2521), .CK(clk), .Q(
        \xmem_inst/mem[40][2] ) );
  DFF_X1 \xmem_inst/mem_reg[40][3]  ( .D(n2520), .CK(clk), .Q(
        \xmem_inst/mem[40][3] ) );
  DFF_X1 \xmem_inst/mem_reg[40][4]  ( .D(n2519), .CK(clk), .Q(
        \xmem_inst/mem[40][4] ) );
  DFF_X1 \xmem_inst/mem_reg[40][5]  ( .D(n2518), .CK(clk), .Q(
        \xmem_inst/mem[40][5] ) );
  DFF_X1 \xmem_inst/mem_reg[40][6]  ( .D(n2517), .CK(clk), .Q(
        \xmem_inst/mem[40][6] ) );
  DFF_X1 \xmem_inst/mem_reg[40][7]  ( .D(n2516), .CK(clk), .Q(
        \xmem_inst/mem[40][7] ) );
  DFF_X1 \xmem_inst/mem_reg[41][0]  ( .D(n2515), .CK(clk), .Q(
        \xmem_inst/mem[41][0] ) );
  DFF_X1 \xmem_inst/mem_reg[41][1]  ( .D(n2514), .CK(clk), .Q(
        \xmem_inst/mem[41][1] ) );
  DFF_X1 \xmem_inst/mem_reg[41][2]  ( .D(n2513), .CK(clk), .Q(
        \xmem_inst/mem[41][2] ) );
  DFF_X1 \xmem_inst/mem_reg[41][3]  ( .D(n2512), .CK(clk), .Q(
        \xmem_inst/mem[41][3] ) );
  DFF_X1 \xmem_inst/mem_reg[41][4]  ( .D(n2511), .CK(clk), .Q(
        \xmem_inst/mem[41][4] ) );
  DFF_X1 \xmem_inst/mem_reg[41][5]  ( .D(n2510), .CK(clk), .Q(
        \xmem_inst/mem[41][5] ) );
  DFF_X1 \xmem_inst/mem_reg[41][6]  ( .D(n2509), .CK(clk), .Q(
        \xmem_inst/mem[41][6] ) );
  DFF_X1 \xmem_inst/mem_reg[41][7]  ( .D(n2508), .CK(clk), .Q(
        \xmem_inst/mem[41][7] ) );
  DFF_X1 \xmem_inst/mem_reg[42][0]  ( .D(n2507), .CK(clk), .Q(
        \xmem_inst/mem[42][0] ) );
  DFF_X1 \xmem_inst/mem_reg[42][1]  ( .D(n2506), .CK(clk), .Q(
        \xmem_inst/mem[42][1] ) );
  DFF_X1 \xmem_inst/mem_reg[42][2]  ( .D(n2505), .CK(clk), .Q(
        \xmem_inst/mem[42][2] ) );
  DFF_X1 \xmem_inst/mem_reg[42][3]  ( .D(n2504), .CK(clk), .Q(
        \xmem_inst/mem[42][3] ) );
  DFF_X1 \xmem_inst/mem_reg[42][4]  ( .D(n2503), .CK(clk), .Q(
        \xmem_inst/mem[42][4] ) );
  DFF_X1 \xmem_inst/mem_reg[42][5]  ( .D(n2502), .CK(clk), .Q(
        \xmem_inst/mem[42][5] ) );
  DFF_X1 \xmem_inst/mem_reg[42][6]  ( .D(n2501), .CK(clk), .Q(
        \xmem_inst/mem[42][6] ) );
  DFF_X1 \xmem_inst/mem_reg[42][7]  ( .D(n2500), .CK(clk), .Q(
        \xmem_inst/mem[42][7] ) );
  DFF_X1 \xmem_inst/mem_reg[43][0]  ( .D(n2499), .CK(clk), .Q(
        \xmem_inst/mem[43][0] ) );
  DFF_X1 \xmem_inst/mem_reg[43][1]  ( .D(n2498), .CK(clk), .Q(
        \xmem_inst/mem[43][1] ) );
  DFF_X1 \xmem_inst/mem_reg[43][2]  ( .D(n2497), .CK(clk), .Q(
        \xmem_inst/mem[43][2] ) );
  DFF_X1 \xmem_inst/mem_reg[43][3]  ( .D(n2496), .CK(clk), .Q(
        \xmem_inst/mem[43][3] ) );
  DFF_X1 \xmem_inst/mem_reg[43][4]  ( .D(n2495), .CK(clk), .Q(
        \xmem_inst/mem[43][4] ) );
  DFF_X1 \xmem_inst/mem_reg[43][5]  ( .D(n2494), .CK(clk), .Q(
        \xmem_inst/mem[43][5] ) );
  DFF_X1 \xmem_inst/mem_reg[43][6]  ( .D(n2493), .CK(clk), .Q(
        \xmem_inst/mem[43][6] ) );
  DFF_X1 \xmem_inst/mem_reg[43][7]  ( .D(n2492), .CK(clk), .Q(
        \xmem_inst/mem[43][7] ) );
  DFF_X1 \xmem_inst/mem_reg[44][0]  ( .D(n2491), .CK(clk), .Q(
        \xmem_inst/mem[44][0] ) );
  DFF_X1 \xmem_inst/mem_reg[44][1]  ( .D(n2490), .CK(clk), .Q(
        \xmem_inst/mem[44][1] ) );
  DFF_X1 \xmem_inst/mem_reg[44][2]  ( .D(n2489), .CK(clk), .Q(
        \xmem_inst/mem[44][2] ) );
  DFF_X1 \xmem_inst/mem_reg[44][3]  ( .D(n2488), .CK(clk), .Q(
        \xmem_inst/mem[44][3] ) );
  DFF_X1 \xmem_inst/mem_reg[44][4]  ( .D(n2487), .CK(clk), .Q(
        \xmem_inst/mem[44][4] ) );
  DFF_X1 \xmem_inst/mem_reg[44][5]  ( .D(n2486), .CK(clk), .Q(
        \xmem_inst/mem[44][5] ) );
  DFF_X1 \xmem_inst/mem_reg[44][6]  ( .D(n2485), .CK(clk), .Q(
        \xmem_inst/mem[44][6] ) );
  DFF_X1 \xmem_inst/mem_reg[44][7]  ( .D(n2484), .CK(clk), .Q(
        \xmem_inst/mem[44][7] ) );
  DFF_X1 \xmem_inst/mem_reg[45][0]  ( .D(n2483), .CK(clk), .Q(
        \xmem_inst/mem[45][0] ) );
  DFF_X1 \xmem_inst/mem_reg[45][1]  ( .D(n2482), .CK(clk), .Q(
        \xmem_inst/mem[45][1] ) );
  DFF_X1 \xmem_inst/mem_reg[45][2]  ( .D(n2481), .CK(clk), .Q(
        \xmem_inst/mem[45][2] ) );
  DFF_X1 \xmem_inst/mem_reg[45][3]  ( .D(n2480), .CK(clk), .Q(
        \xmem_inst/mem[45][3] ) );
  DFF_X1 \xmem_inst/mem_reg[45][4]  ( .D(n2479), .CK(clk), .Q(
        \xmem_inst/mem[45][4] ) );
  DFF_X1 \xmem_inst/mem_reg[45][5]  ( .D(n2478), .CK(clk), .Q(
        \xmem_inst/mem[45][5] ) );
  DFF_X1 \xmem_inst/mem_reg[45][6]  ( .D(n2477), .CK(clk), .Q(
        \xmem_inst/mem[45][6] ) );
  DFF_X1 \xmem_inst/mem_reg[45][7]  ( .D(n2476), .CK(clk), .Q(
        \xmem_inst/mem[45][7] ) );
  DFF_X1 \xmem_inst/mem_reg[46][0]  ( .D(n2475), .CK(clk), .Q(
        \xmem_inst/mem[46][0] ) );
  DFF_X1 \xmem_inst/mem_reg[46][1]  ( .D(n2474), .CK(clk), .Q(
        \xmem_inst/mem[46][1] ) );
  DFF_X1 \xmem_inst/mem_reg[46][2]  ( .D(n2473), .CK(clk), .Q(
        \xmem_inst/mem[46][2] ) );
  DFF_X1 \xmem_inst/mem_reg[46][3]  ( .D(n2472), .CK(clk), .Q(
        \xmem_inst/mem[46][3] ) );
  DFF_X1 \xmem_inst/mem_reg[46][4]  ( .D(n2471), .CK(clk), .Q(
        \xmem_inst/mem[46][4] ) );
  DFF_X1 \xmem_inst/mem_reg[46][5]  ( .D(n2470), .CK(clk), .Q(
        \xmem_inst/mem[46][5] ) );
  DFF_X1 \xmem_inst/mem_reg[46][6]  ( .D(n2469), .CK(clk), .Q(
        \xmem_inst/mem[46][6] ) );
  DFF_X1 \xmem_inst/mem_reg[46][7]  ( .D(n2468), .CK(clk), .Q(
        \xmem_inst/mem[46][7] ) );
  DFF_X1 \xmem_inst/mem_reg[47][0]  ( .D(n2467), .CK(clk), .Q(
        \xmem_inst/mem[47][0] ) );
  DFF_X1 \xmem_inst/mem_reg[47][1]  ( .D(n2466), .CK(clk), .Q(
        \xmem_inst/mem[47][1] ) );
  DFF_X1 \xmem_inst/mem_reg[47][2]  ( .D(n2465), .CK(clk), .Q(
        \xmem_inst/mem[47][2] ) );
  DFF_X1 \xmem_inst/mem_reg[47][3]  ( .D(n2464), .CK(clk), .Q(
        \xmem_inst/mem[47][3] ) );
  DFF_X1 \xmem_inst/mem_reg[47][4]  ( .D(n2463), .CK(clk), .Q(
        \xmem_inst/mem[47][4] ) );
  DFF_X1 \xmem_inst/mem_reg[47][5]  ( .D(n2462), .CK(clk), .Q(
        \xmem_inst/mem[47][5] ) );
  DFF_X1 \xmem_inst/mem_reg[47][6]  ( .D(n2461), .CK(clk), .Q(
        \xmem_inst/mem[47][6] ) );
  DFF_X1 \xmem_inst/mem_reg[47][7]  ( .D(n2460), .CK(clk), .Q(
        \xmem_inst/mem[47][7] ) );
  DFF_X1 \xmem_inst/mem_reg[48][0]  ( .D(n2459), .CK(clk), .Q(
        \xmem_inst/mem[48][0] ) );
  DFF_X1 \xmem_inst/mem_reg[48][1]  ( .D(n2458), .CK(clk), .Q(
        \xmem_inst/mem[48][1] ) );
  DFF_X1 \xmem_inst/mem_reg[48][2]  ( .D(n2457), .CK(clk), .Q(
        \xmem_inst/mem[48][2] ) );
  DFF_X1 \xmem_inst/mem_reg[48][3]  ( .D(n2456), .CK(clk), .Q(
        \xmem_inst/mem[48][3] ) );
  DFF_X1 \xmem_inst/mem_reg[48][4]  ( .D(n2455), .CK(clk), .Q(
        \xmem_inst/mem[48][4] ) );
  DFF_X1 \xmem_inst/mem_reg[48][5]  ( .D(n2454), .CK(clk), .Q(
        \xmem_inst/mem[48][5] ) );
  DFF_X1 \xmem_inst/mem_reg[48][6]  ( .D(n2453), .CK(clk), .Q(
        \xmem_inst/mem[48][6] ) );
  DFF_X1 \xmem_inst/mem_reg[48][7]  ( .D(n2452), .CK(clk), .Q(
        \xmem_inst/mem[48][7] ) );
  DFF_X1 \xmem_inst/mem_reg[49][0]  ( .D(n2451), .CK(clk), .Q(
        \xmem_inst/mem[49][0] ) );
  DFF_X1 \xmem_inst/mem_reg[49][1]  ( .D(n2450), .CK(clk), .Q(
        \xmem_inst/mem[49][1] ) );
  DFF_X1 \xmem_inst/mem_reg[49][2]  ( .D(n2449), .CK(clk), .Q(
        \xmem_inst/mem[49][2] ) );
  DFF_X1 \xmem_inst/mem_reg[49][3]  ( .D(n2448), .CK(clk), .Q(
        \xmem_inst/mem[49][3] ) );
  DFF_X1 \xmem_inst/mem_reg[49][4]  ( .D(n2447), .CK(clk), .Q(
        \xmem_inst/mem[49][4] ) );
  DFF_X1 \xmem_inst/mem_reg[49][5]  ( .D(n2446), .CK(clk), .Q(
        \xmem_inst/mem[49][5] ) );
  DFF_X1 \xmem_inst/mem_reg[49][6]  ( .D(n2445), .CK(clk), .Q(
        \xmem_inst/mem[49][6] ) );
  DFF_X1 \xmem_inst/mem_reg[49][7]  ( .D(n2444), .CK(clk), .Q(
        \xmem_inst/mem[49][7] ) );
  DFF_X1 \xmem_inst/mem_reg[50][0]  ( .D(n2443), .CK(clk), .Q(
        \xmem_inst/mem[50][0] ) );
  DFF_X1 \xmem_inst/mem_reg[50][1]  ( .D(n2442), .CK(clk), .Q(
        \xmem_inst/mem[50][1] ) );
  DFF_X1 \xmem_inst/mem_reg[50][2]  ( .D(n2441), .CK(clk), .Q(
        \xmem_inst/mem[50][2] ) );
  DFF_X1 \xmem_inst/mem_reg[50][3]  ( .D(n2440), .CK(clk), .Q(
        \xmem_inst/mem[50][3] ) );
  DFF_X1 \xmem_inst/mem_reg[50][4]  ( .D(n2439), .CK(clk), .Q(
        \xmem_inst/mem[50][4] ) );
  DFF_X1 \xmem_inst/mem_reg[50][5]  ( .D(n2438), .CK(clk), .Q(
        \xmem_inst/mem[50][5] ) );
  DFF_X1 \xmem_inst/mem_reg[50][6]  ( .D(n2437), .CK(clk), .Q(
        \xmem_inst/mem[50][6] ) );
  DFF_X1 \xmem_inst/mem_reg[50][7]  ( .D(n2436), .CK(clk), .Q(
        \xmem_inst/mem[50][7] ) );
  DFF_X1 \xmem_inst/mem_reg[51][0]  ( .D(n2435), .CK(clk), .Q(
        \xmem_inst/mem[51][0] ) );
  DFF_X1 \xmem_inst/mem_reg[51][1]  ( .D(n2434), .CK(clk), .Q(
        \xmem_inst/mem[51][1] ) );
  DFF_X1 \xmem_inst/mem_reg[51][2]  ( .D(n2433), .CK(clk), .Q(
        \xmem_inst/mem[51][2] ) );
  DFF_X1 \xmem_inst/mem_reg[51][3]  ( .D(n2432), .CK(clk), .Q(
        \xmem_inst/mem[51][3] ) );
  DFF_X1 \xmem_inst/mem_reg[51][4]  ( .D(n2431), .CK(clk), .Q(
        \xmem_inst/mem[51][4] ) );
  DFF_X1 \xmem_inst/mem_reg[51][5]  ( .D(n2430), .CK(clk), .Q(
        \xmem_inst/mem[51][5] ) );
  DFF_X1 \xmem_inst/mem_reg[51][6]  ( .D(n2429), .CK(clk), .Q(
        \xmem_inst/mem[51][6] ) );
  DFF_X1 \xmem_inst/mem_reg[51][7]  ( .D(n2428), .CK(clk), .Q(
        \xmem_inst/mem[51][7] ) );
  DFF_X1 \xmem_inst/mem_reg[52][0]  ( .D(n2427), .CK(clk), .Q(
        \xmem_inst/mem[52][0] ) );
  DFF_X1 \xmem_inst/mem_reg[52][1]  ( .D(n2426), .CK(clk), .Q(
        \xmem_inst/mem[52][1] ) );
  DFF_X1 \xmem_inst/mem_reg[52][2]  ( .D(n2425), .CK(clk), .Q(
        \xmem_inst/mem[52][2] ) );
  DFF_X1 \xmem_inst/mem_reg[52][3]  ( .D(n2424), .CK(clk), .Q(
        \xmem_inst/mem[52][3] ) );
  DFF_X1 \xmem_inst/mem_reg[52][4]  ( .D(n2423), .CK(clk), .Q(
        \xmem_inst/mem[52][4] ) );
  DFF_X1 \xmem_inst/mem_reg[52][5]  ( .D(n2422), .CK(clk), .Q(
        \xmem_inst/mem[52][5] ) );
  DFF_X1 \xmem_inst/mem_reg[52][6]  ( .D(n2421), .CK(clk), .Q(
        \xmem_inst/mem[52][6] ) );
  DFF_X1 \xmem_inst/mem_reg[52][7]  ( .D(n2420), .CK(clk), .Q(
        \xmem_inst/mem[52][7] ) );
  DFF_X1 \xmem_inst/mem_reg[53][0]  ( .D(n2419), .CK(clk), .Q(
        \xmem_inst/mem[53][0] ) );
  DFF_X1 \xmem_inst/mem_reg[53][1]  ( .D(n2418), .CK(clk), .Q(
        \xmem_inst/mem[53][1] ) );
  DFF_X1 \xmem_inst/mem_reg[53][2]  ( .D(n2417), .CK(clk), .Q(
        \xmem_inst/mem[53][2] ) );
  DFF_X1 \xmem_inst/mem_reg[53][3]  ( .D(n2416), .CK(clk), .Q(
        \xmem_inst/mem[53][3] ) );
  DFF_X1 \xmem_inst/mem_reg[53][4]  ( .D(n2415), .CK(clk), .Q(
        \xmem_inst/mem[53][4] ) );
  DFF_X1 \xmem_inst/mem_reg[53][5]  ( .D(n2414), .CK(clk), .Q(
        \xmem_inst/mem[53][5] ) );
  DFF_X1 \xmem_inst/mem_reg[53][6]  ( .D(n2413), .CK(clk), .Q(
        \xmem_inst/mem[53][6] ) );
  DFF_X1 \xmem_inst/mem_reg[53][7]  ( .D(n2412), .CK(clk), .Q(
        \xmem_inst/mem[53][7] ) );
  DFF_X1 \xmem_inst/mem_reg[54][0]  ( .D(n2411), .CK(clk), .Q(
        \xmem_inst/mem[54][0] ) );
  DFF_X1 \xmem_inst/mem_reg[54][1]  ( .D(n2410), .CK(clk), .Q(
        \xmem_inst/mem[54][1] ) );
  DFF_X1 \xmem_inst/mem_reg[54][2]  ( .D(n2409), .CK(clk), .Q(
        \xmem_inst/mem[54][2] ) );
  DFF_X1 \xmem_inst/mem_reg[54][3]  ( .D(n2408), .CK(clk), .Q(
        \xmem_inst/mem[54][3] ) );
  DFF_X1 \xmem_inst/mem_reg[54][4]  ( .D(n2407), .CK(clk), .Q(
        \xmem_inst/mem[54][4] ) );
  DFF_X1 \xmem_inst/mem_reg[54][5]  ( .D(n2406), .CK(clk), .Q(
        \xmem_inst/mem[54][5] ) );
  DFF_X1 \xmem_inst/mem_reg[54][6]  ( .D(n2405), .CK(clk), .Q(
        \xmem_inst/mem[54][6] ) );
  DFF_X1 \xmem_inst/mem_reg[54][7]  ( .D(n2404), .CK(clk), .Q(
        \xmem_inst/mem[54][7] ) );
  DFF_X1 \xmem_inst/mem_reg[55][0]  ( .D(n2403), .CK(clk), .Q(
        \xmem_inst/mem[55][0] ) );
  DFF_X1 \xmem_inst/mem_reg[55][1]  ( .D(n2402), .CK(clk), .Q(
        \xmem_inst/mem[55][1] ) );
  DFF_X1 \xmem_inst/mem_reg[55][2]  ( .D(n2401), .CK(clk), .Q(
        \xmem_inst/mem[55][2] ) );
  DFF_X1 \xmem_inst/mem_reg[55][3]  ( .D(n2400), .CK(clk), .Q(
        \xmem_inst/mem[55][3] ) );
  DFF_X1 \xmem_inst/mem_reg[55][4]  ( .D(n2399), .CK(clk), .Q(
        \xmem_inst/mem[55][4] ) );
  DFF_X1 \xmem_inst/mem_reg[55][5]  ( .D(n2398), .CK(clk), .Q(
        \xmem_inst/mem[55][5] ) );
  DFF_X1 \xmem_inst/mem_reg[55][6]  ( .D(n2397), .CK(clk), .Q(
        \xmem_inst/mem[55][6] ) );
  DFF_X1 \xmem_inst/mem_reg[55][7]  ( .D(n2396), .CK(clk), .Q(
        \xmem_inst/mem[55][7] ) );
  DFF_X1 \xmem_inst/mem_reg[56][0]  ( .D(n2395), .CK(clk), .Q(
        \xmem_inst/mem[56][0] ) );
  DFF_X1 \xmem_inst/mem_reg[56][1]  ( .D(n2394), .CK(clk), .Q(
        \xmem_inst/mem[56][1] ) );
  DFF_X1 \xmem_inst/mem_reg[56][2]  ( .D(n2393), .CK(clk), .Q(
        \xmem_inst/mem[56][2] ) );
  DFF_X1 \xmem_inst/mem_reg[56][3]  ( .D(n2392), .CK(clk), .Q(
        \xmem_inst/mem[56][3] ) );
  DFF_X1 \xmem_inst/mem_reg[56][4]  ( .D(n2391), .CK(clk), .Q(
        \xmem_inst/mem[56][4] ) );
  DFF_X1 \xmem_inst/mem_reg[56][5]  ( .D(n2390), .CK(clk), .Q(
        \xmem_inst/mem[56][5] ) );
  DFF_X1 \xmem_inst/mem_reg[56][6]  ( .D(n2389), .CK(clk), .Q(
        \xmem_inst/mem[56][6] ) );
  DFF_X1 \xmem_inst/mem_reg[56][7]  ( .D(n2388), .CK(clk), .Q(
        \xmem_inst/mem[56][7] ) );
  DFF_X1 \xmem_inst/mem_reg[57][0]  ( .D(n2387), .CK(clk), .Q(
        \xmem_inst/mem[57][0] ) );
  DFF_X1 \xmem_inst/mem_reg[57][1]  ( .D(n2386), .CK(clk), .Q(
        \xmem_inst/mem[57][1] ) );
  DFF_X1 \xmem_inst/mem_reg[57][2]  ( .D(n2385), .CK(clk), .Q(
        \xmem_inst/mem[57][2] ) );
  DFF_X1 \xmem_inst/mem_reg[57][3]  ( .D(n2384), .CK(clk), .Q(
        \xmem_inst/mem[57][3] ) );
  DFF_X1 \xmem_inst/mem_reg[57][4]  ( .D(n2383), .CK(clk), .Q(
        \xmem_inst/mem[57][4] ) );
  DFF_X1 \xmem_inst/mem_reg[57][5]  ( .D(n2382), .CK(clk), .Q(
        \xmem_inst/mem[57][5] ) );
  DFF_X1 \xmem_inst/mem_reg[57][6]  ( .D(n2381), .CK(clk), .Q(
        \xmem_inst/mem[57][6] ) );
  DFF_X1 \xmem_inst/mem_reg[57][7]  ( .D(n2380), .CK(clk), .Q(
        \xmem_inst/mem[57][7] ) );
  DFF_X1 \xmem_inst/mem_reg[58][0]  ( .D(n2379), .CK(clk), .Q(
        \xmem_inst/mem[58][0] ) );
  DFF_X1 \xmem_inst/mem_reg[58][1]  ( .D(n2378), .CK(clk), .Q(
        \xmem_inst/mem[58][1] ) );
  DFF_X1 \xmem_inst/mem_reg[58][2]  ( .D(n2377), .CK(clk), .Q(
        \xmem_inst/mem[58][2] ) );
  DFF_X1 \xmem_inst/mem_reg[58][3]  ( .D(n2376), .CK(clk), .Q(
        \xmem_inst/mem[58][3] ) );
  DFF_X1 \xmem_inst/mem_reg[58][4]  ( .D(n2375), .CK(clk), .Q(
        \xmem_inst/mem[58][4] ) );
  DFF_X1 \xmem_inst/mem_reg[58][5]  ( .D(n2374), .CK(clk), .Q(
        \xmem_inst/mem[58][5] ) );
  DFF_X1 \xmem_inst/mem_reg[58][6]  ( .D(n2373), .CK(clk), .Q(
        \xmem_inst/mem[58][6] ) );
  DFF_X1 \xmem_inst/mem_reg[58][7]  ( .D(n2372), .CK(clk), .Q(
        \xmem_inst/mem[58][7] ) );
  DFF_X1 \xmem_inst/mem_reg[59][0]  ( .D(n2371), .CK(clk), .Q(
        \xmem_inst/mem[59][0] ) );
  DFF_X1 \xmem_inst/mem_reg[59][1]  ( .D(n2370), .CK(clk), .Q(
        \xmem_inst/mem[59][1] ) );
  DFF_X1 \xmem_inst/mem_reg[59][2]  ( .D(n2369), .CK(clk), .Q(
        \xmem_inst/mem[59][2] ) );
  DFF_X1 \xmem_inst/mem_reg[59][3]  ( .D(n2368), .CK(clk), .Q(
        \xmem_inst/mem[59][3] ) );
  DFF_X1 \xmem_inst/mem_reg[59][4]  ( .D(n2367), .CK(clk), .Q(
        \xmem_inst/mem[59][4] ) );
  DFF_X1 \xmem_inst/mem_reg[59][5]  ( .D(n2366), .CK(clk), .Q(
        \xmem_inst/mem[59][5] ) );
  DFF_X1 \xmem_inst/mem_reg[59][6]  ( .D(n2365), .CK(clk), .Q(
        \xmem_inst/mem[59][6] ) );
  DFF_X1 \xmem_inst/mem_reg[59][7]  ( .D(n2364), .CK(clk), .Q(
        \xmem_inst/mem[59][7] ) );
  DFF_X1 \xmem_inst/mem_reg[60][0]  ( .D(n2363), .CK(clk), .Q(
        \xmem_inst/mem[60][0] ) );
  DFF_X1 \xmem_inst/mem_reg[60][1]  ( .D(n2362), .CK(clk), .Q(
        \xmem_inst/mem[60][1] ) );
  DFF_X1 \xmem_inst/mem_reg[60][2]  ( .D(n2361), .CK(clk), .Q(
        \xmem_inst/mem[60][2] ) );
  DFF_X1 \xmem_inst/mem_reg[60][3]  ( .D(n2360), .CK(clk), .Q(
        \xmem_inst/mem[60][3] ) );
  DFF_X1 \xmem_inst/mem_reg[60][4]  ( .D(n2359), .CK(clk), .Q(
        \xmem_inst/mem[60][4] ) );
  DFF_X1 \xmem_inst/mem_reg[60][5]  ( .D(n2358), .CK(clk), .Q(
        \xmem_inst/mem[60][5] ) );
  DFF_X1 \xmem_inst/mem_reg[60][6]  ( .D(n2357), .CK(clk), .Q(
        \xmem_inst/mem[60][6] ) );
  DFF_X1 \xmem_inst/mem_reg[60][7]  ( .D(n2356), .CK(clk), .Q(
        \xmem_inst/mem[60][7] ) );
  DFF_X1 \xmem_inst/mem_reg[61][0]  ( .D(n2355), .CK(clk), .Q(
        \xmem_inst/mem[61][0] ) );
  DFF_X1 \xmem_inst/mem_reg[61][1]  ( .D(n2354), .CK(clk), .Q(
        \xmem_inst/mem[61][1] ) );
  DFF_X1 \xmem_inst/mem_reg[61][2]  ( .D(n2353), .CK(clk), .Q(
        \xmem_inst/mem[61][2] ) );
  DFF_X1 \xmem_inst/mem_reg[61][3]  ( .D(n2352), .CK(clk), .Q(
        \xmem_inst/mem[61][3] ) );
  DFF_X1 \xmem_inst/mem_reg[61][4]  ( .D(n2351), .CK(clk), .Q(
        \xmem_inst/mem[61][4] ) );
  DFF_X1 \xmem_inst/mem_reg[61][5]  ( .D(n2350), .CK(clk), .Q(
        \xmem_inst/mem[61][5] ) );
  DFF_X1 \xmem_inst/mem_reg[61][6]  ( .D(n2349), .CK(clk), .Q(
        \xmem_inst/mem[61][6] ) );
  DFF_X1 \xmem_inst/mem_reg[61][7]  ( .D(n2348), .CK(clk), .Q(
        \xmem_inst/mem[61][7] ) );
  DFF_X1 \xmem_inst/mem_reg[62][0]  ( .D(n2347), .CK(clk), .Q(
        \xmem_inst/mem[62][0] ) );
  DFF_X1 \xmem_inst/mem_reg[62][1]  ( .D(n2346), .CK(clk), .Q(
        \xmem_inst/mem[62][1] ) );
  DFF_X1 \xmem_inst/mem_reg[62][2]  ( .D(n2345), .CK(clk), .Q(
        \xmem_inst/mem[62][2] ) );
  DFF_X1 \xmem_inst/mem_reg[62][3]  ( .D(n2344), .CK(clk), .Q(
        \xmem_inst/mem[62][3] ) );
  DFF_X1 \xmem_inst/mem_reg[62][4]  ( .D(n2343), .CK(clk), .Q(
        \xmem_inst/mem[62][4] ) );
  DFF_X1 \xmem_inst/mem_reg[62][5]  ( .D(n2342), .CK(clk), .Q(
        \xmem_inst/mem[62][5] ) );
  DFF_X1 \xmem_inst/mem_reg[62][6]  ( .D(n2341), .CK(clk), .Q(
        \xmem_inst/mem[62][6] ) );
  DFF_X1 \xmem_inst/mem_reg[62][7]  ( .D(n2340), .CK(clk), .Q(
        \xmem_inst/mem[62][7] ) );
  DFF_X1 \xmem_inst/mem_reg[63][0]  ( .D(n2339), .CK(clk), .Q(
        \xmem_inst/mem[63][0] ) );
  DFF_X1 \xmem_inst/mem_reg[63][1]  ( .D(n2338), .CK(clk), .Q(
        \xmem_inst/mem[63][1] ) );
  DFF_X1 \xmem_inst/mem_reg[63][2]  ( .D(n2337), .CK(clk), .Q(
        \xmem_inst/mem[63][2] ) );
  DFF_X1 \xmem_inst/mem_reg[63][3]  ( .D(n2336), .CK(clk), .Q(
        \xmem_inst/mem[63][3] ) );
  DFF_X1 \xmem_inst/mem_reg[63][4]  ( .D(n2335), .CK(clk), .Q(
        \xmem_inst/mem[63][4] ) );
  DFF_X1 \xmem_inst/mem_reg[63][5]  ( .D(n2334), .CK(clk), .Q(
        \xmem_inst/mem[63][5] ) );
  DFF_X1 \xmem_inst/mem_reg[63][6]  ( .D(n2333), .CK(clk), .Q(
        \xmem_inst/mem[63][6] ) );
  DFF_X1 \xmem_inst/mem_reg[63][7]  ( .D(n2332), .CK(clk), .Q(
        \xmem_inst/mem[63][7] ) );
  DFF_X1 \xmem_inst/mem_reg[64][0]  ( .D(n2331), .CK(clk), .Q(
        \xmem_inst/mem[64][0] ) );
  DFF_X1 \xmem_inst/mem_reg[64][1]  ( .D(n2330), .CK(clk), .Q(
        \xmem_inst/mem[64][1] ) );
  DFF_X1 \xmem_inst/mem_reg[64][2]  ( .D(n2329), .CK(clk), .Q(
        \xmem_inst/mem[64][2] ) );
  DFF_X1 \xmem_inst/mem_reg[64][3]  ( .D(n2328), .CK(clk), .Q(
        \xmem_inst/mem[64][3] ) );
  DFF_X1 \xmem_inst/mem_reg[64][4]  ( .D(n2327), .CK(clk), .Q(
        \xmem_inst/mem[64][4] ) );
  DFF_X1 \xmem_inst/mem_reg[64][5]  ( .D(n2326), .CK(clk), .Q(
        \xmem_inst/mem[64][5] ) );
  DFF_X1 \xmem_inst/mem_reg[64][6]  ( .D(n2325), .CK(clk), .Q(
        \xmem_inst/mem[64][6] ) );
  DFF_X1 \xmem_inst/mem_reg[64][7]  ( .D(n2324), .CK(clk), .Q(
        \xmem_inst/mem[64][7] ) );
  DFF_X1 \xmem_inst/mem_reg[65][0]  ( .D(n2323), .CK(clk), .Q(
        \xmem_inst/mem[65][0] ) );
  DFF_X1 \xmem_inst/mem_reg[65][1]  ( .D(n2322), .CK(clk), .Q(
        \xmem_inst/mem[65][1] ) );
  DFF_X1 \xmem_inst/mem_reg[65][2]  ( .D(n2321), .CK(clk), .Q(
        \xmem_inst/mem[65][2] ) );
  DFF_X1 \xmem_inst/mem_reg[65][3]  ( .D(n2320), .CK(clk), .Q(
        \xmem_inst/mem[65][3] ) );
  DFF_X1 \xmem_inst/mem_reg[65][4]  ( .D(n2319), .CK(clk), .Q(
        \xmem_inst/mem[65][4] ) );
  DFF_X1 \xmem_inst/mem_reg[65][5]  ( .D(n2318), .CK(clk), .Q(
        \xmem_inst/mem[65][5] ) );
  DFF_X1 \xmem_inst/mem_reg[65][6]  ( .D(n2317), .CK(clk), .Q(
        \xmem_inst/mem[65][6] ) );
  DFF_X1 \xmem_inst/mem_reg[65][7]  ( .D(n2316), .CK(clk), .Q(
        \xmem_inst/mem[65][7] ) );
  DFF_X1 \xmem_inst/mem_reg[66][0]  ( .D(n2315), .CK(clk), .Q(
        \xmem_inst/mem[66][0] ) );
  DFF_X1 \xmem_inst/mem_reg[66][1]  ( .D(n2314), .CK(clk), .Q(
        \xmem_inst/mem[66][1] ) );
  DFF_X1 \xmem_inst/mem_reg[66][2]  ( .D(n2313), .CK(clk), .Q(
        \xmem_inst/mem[66][2] ) );
  DFF_X1 \xmem_inst/mem_reg[66][3]  ( .D(n2312), .CK(clk), .Q(
        \xmem_inst/mem[66][3] ) );
  DFF_X1 \xmem_inst/mem_reg[66][4]  ( .D(n2311), .CK(clk), .Q(
        \xmem_inst/mem[66][4] ) );
  DFF_X1 \xmem_inst/mem_reg[66][5]  ( .D(n2310), .CK(clk), .Q(
        \xmem_inst/mem[66][5] ) );
  DFF_X1 \xmem_inst/mem_reg[66][6]  ( .D(n2309), .CK(clk), .Q(
        \xmem_inst/mem[66][6] ) );
  DFF_X1 \xmem_inst/mem_reg[66][7]  ( .D(n2308), .CK(clk), .Q(
        \xmem_inst/mem[66][7] ) );
  DFF_X1 \xmem_inst/mem_reg[67][0]  ( .D(n2307), .CK(clk), .Q(
        \xmem_inst/mem[67][0] ) );
  DFF_X1 \xmem_inst/mem_reg[67][1]  ( .D(n2306), .CK(clk), .Q(
        \xmem_inst/mem[67][1] ) );
  DFF_X1 \xmem_inst/mem_reg[67][2]  ( .D(n2305), .CK(clk), .Q(
        \xmem_inst/mem[67][2] ) );
  DFF_X1 \xmem_inst/mem_reg[67][3]  ( .D(n2304), .CK(clk), .Q(
        \xmem_inst/mem[67][3] ) );
  DFF_X1 \xmem_inst/mem_reg[67][4]  ( .D(n2303), .CK(clk), .Q(
        \xmem_inst/mem[67][4] ) );
  DFF_X1 \xmem_inst/mem_reg[67][5]  ( .D(n2302), .CK(clk), .Q(
        \xmem_inst/mem[67][5] ) );
  DFF_X1 \xmem_inst/mem_reg[67][6]  ( .D(n2301), .CK(clk), .Q(
        \xmem_inst/mem[67][6] ) );
  DFF_X1 \xmem_inst/mem_reg[67][7]  ( .D(n2300), .CK(clk), .Q(
        \xmem_inst/mem[67][7] ) );
  DFF_X1 \xmem_inst/mem_reg[68][0]  ( .D(n2299), .CK(clk), .Q(
        \xmem_inst/mem[68][0] ) );
  DFF_X1 \xmem_inst/mem_reg[68][1]  ( .D(n2298), .CK(clk), .Q(
        \xmem_inst/mem[68][1] ) );
  DFF_X1 \xmem_inst/mem_reg[68][2]  ( .D(n2297), .CK(clk), .Q(
        \xmem_inst/mem[68][2] ) );
  DFF_X1 \xmem_inst/mem_reg[68][3]  ( .D(n2296), .CK(clk), .Q(
        \xmem_inst/mem[68][3] ) );
  DFF_X1 \xmem_inst/mem_reg[68][4]  ( .D(n2295), .CK(clk), .Q(
        \xmem_inst/mem[68][4] ) );
  DFF_X1 \xmem_inst/mem_reg[68][5]  ( .D(n2294), .CK(clk), .Q(
        \xmem_inst/mem[68][5] ) );
  DFF_X1 \xmem_inst/mem_reg[68][6]  ( .D(n2293), .CK(clk), .Q(
        \xmem_inst/mem[68][6] ) );
  DFF_X1 \xmem_inst/mem_reg[68][7]  ( .D(n2292), .CK(clk), .Q(
        \xmem_inst/mem[68][7] ) );
  DFF_X1 \xmem_inst/mem_reg[69][0]  ( .D(n2291), .CK(clk), .Q(
        \xmem_inst/mem[69][0] ) );
  DFF_X1 \xmem_inst/mem_reg[69][1]  ( .D(n2290), .CK(clk), .Q(
        \xmem_inst/mem[69][1] ) );
  DFF_X1 \xmem_inst/mem_reg[69][2]  ( .D(n2289), .CK(clk), .Q(
        \xmem_inst/mem[69][2] ) );
  DFF_X1 \xmem_inst/mem_reg[69][3]  ( .D(n2288), .CK(clk), .Q(
        \xmem_inst/mem[69][3] ) );
  DFF_X1 \xmem_inst/mem_reg[69][4]  ( .D(n2287), .CK(clk), .Q(
        \xmem_inst/mem[69][4] ) );
  DFF_X1 \xmem_inst/mem_reg[69][5]  ( .D(n2286), .CK(clk), .Q(
        \xmem_inst/mem[69][5] ) );
  DFF_X1 \xmem_inst/mem_reg[69][6]  ( .D(n2285), .CK(clk), .Q(
        \xmem_inst/mem[69][6] ) );
  DFF_X1 \xmem_inst/mem_reg[69][7]  ( .D(n2284), .CK(clk), .Q(
        \xmem_inst/mem[69][7] ) );
  DFF_X1 \xmem_inst/mem_reg[70][0]  ( .D(n2283), .CK(clk), .Q(
        \xmem_inst/mem[70][0] ) );
  DFF_X1 \xmem_inst/mem_reg[70][1]  ( .D(n2282), .CK(clk), .Q(
        \xmem_inst/mem[70][1] ) );
  DFF_X1 \xmem_inst/mem_reg[70][2]  ( .D(n2281), .CK(clk), .Q(
        \xmem_inst/mem[70][2] ) );
  DFF_X1 \xmem_inst/mem_reg[70][3]  ( .D(n2280), .CK(clk), .Q(
        \xmem_inst/mem[70][3] ) );
  DFF_X1 \xmem_inst/mem_reg[70][4]  ( .D(n2279), .CK(clk), .Q(
        \xmem_inst/mem[70][4] ) );
  DFF_X1 \xmem_inst/mem_reg[70][5]  ( .D(n2278), .CK(clk), .Q(
        \xmem_inst/mem[70][5] ) );
  DFF_X1 \xmem_inst/mem_reg[70][6]  ( .D(n2277), .CK(clk), .Q(
        \xmem_inst/mem[70][6] ) );
  DFF_X1 \xmem_inst/mem_reg[70][7]  ( .D(n2276), .CK(clk), .Q(
        \xmem_inst/mem[70][7] ) );
  DFF_X1 \xmem_inst/mem_reg[71][0]  ( .D(n2275), .CK(clk), .Q(
        \xmem_inst/mem[71][0] ) );
  DFF_X1 \xmem_inst/mem_reg[71][1]  ( .D(n2274), .CK(clk), .Q(
        \xmem_inst/mem[71][1] ) );
  DFF_X1 \xmem_inst/mem_reg[71][2]  ( .D(n2273), .CK(clk), .Q(
        \xmem_inst/mem[71][2] ) );
  DFF_X1 \xmem_inst/mem_reg[71][3]  ( .D(n2272), .CK(clk), .Q(
        \xmem_inst/mem[71][3] ) );
  DFF_X1 \xmem_inst/mem_reg[71][4]  ( .D(n2271), .CK(clk), .Q(
        \xmem_inst/mem[71][4] ) );
  DFF_X1 \xmem_inst/mem_reg[71][5]  ( .D(n2270), .CK(clk), .Q(
        \xmem_inst/mem[71][5] ) );
  DFF_X1 \xmem_inst/mem_reg[71][6]  ( .D(n2269), .CK(clk), .Q(
        \xmem_inst/mem[71][6] ) );
  DFF_X1 \xmem_inst/mem_reg[71][7]  ( .D(n2268), .CK(clk), .Q(
        \xmem_inst/mem[71][7] ) );
  DFF_X1 \xmem_inst/mem_reg[72][0]  ( .D(n2267), .CK(clk), .Q(
        \xmem_inst/mem[72][0] ) );
  DFF_X1 \xmem_inst/mem_reg[72][1]  ( .D(n2266), .CK(clk), .Q(
        \xmem_inst/mem[72][1] ) );
  DFF_X1 \xmem_inst/mem_reg[72][2]  ( .D(n2265), .CK(clk), .Q(
        \xmem_inst/mem[72][2] ) );
  DFF_X1 \xmem_inst/mem_reg[72][3]  ( .D(n2264), .CK(clk), .Q(
        \xmem_inst/mem[72][3] ) );
  DFF_X1 \xmem_inst/mem_reg[72][4]  ( .D(n2263), .CK(clk), .Q(
        \xmem_inst/mem[72][4] ) );
  DFF_X1 \xmem_inst/mem_reg[72][5]  ( .D(n2262), .CK(clk), .Q(
        \xmem_inst/mem[72][5] ) );
  DFF_X1 \xmem_inst/mem_reg[72][6]  ( .D(n2261), .CK(clk), .Q(
        \xmem_inst/mem[72][6] ) );
  DFF_X1 \xmem_inst/mem_reg[72][7]  ( .D(n2260), .CK(clk), .Q(
        \xmem_inst/mem[72][7] ) );
  DFF_X1 \xmem_inst/mem_reg[73][0]  ( .D(n2259), .CK(clk), .Q(
        \xmem_inst/mem[73][0] ) );
  DFF_X1 \xmem_inst/mem_reg[73][1]  ( .D(n2258), .CK(clk), .Q(
        \xmem_inst/mem[73][1] ) );
  DFF_X1 \xmem_inst/mem_reg[73][2]  ( .D(n2257), .CK(clk), .Q(
        \xmem_inst/mem[73][2] ) );
  DFF_X1 \xmem_inst/mem_reg[73][3]  ( .D(n2256), .CK(clk), .Q(
        \xmem_inst/mem[73][3] ) );
  DFF_X1 \xmem_inst/mem_reg[73][4]  ( .D(n2255), .CK(clk), .Q(
        \xmem_inst/mem[73][4] ) );
  DFF_X1 \xmem_inst/mem_reg[73][5]  ( .D(n2254), .CK(clk), .Q(
        \xmem_inst/mem[73][5] ) );
  DFF_X1 \xmem_inst/mem_reg[73][6]  ( .D(n2253), .CK(clk), .Q(
        \xmem_inst/mem[73][6] ) );
  DFF_X1 \xmem_inst/mem_reg[73][7]  ( .D(n2252), .CK(clk), .Q(
        \xmem_inst/mem[73][7] ) );
  DFF_X1 \xmem_inst/mem_reg[74][0]  ( .D(n2251), .CK(clk), .Q(
        \xmem_inst/mem[74][0] ) );
  DFF_X1 \xmem_inst/mem_reg[74][1]  ( .D(n2250), .CK(clk), .Q(
        \xmem_inst/mem[74][1] ) );
  DFF_X1 \xmem_inst/mem_reg[74][2]  ( .D(n2249), .CK(clk), .Q(
        \xmem_inst/mem[74][2] ) );
  DFF_X1 \xmem_inst/mem_reg[74][3]  ( .D(n2248), .CK(clk), .Q(
        \xmem_inst/mem[74][3] ) );
  DFF_X1 \xmem_inst/mem_reg[74][4]  ( .D(n2247), .CK(clk), .Q(
        \xmem_inst/mem[74][4] ) );
  DFF_X1 \xmem_inst/mem_reg[74][5]  ( .D(n2246), .CK(clk), .Q(
        \xmem_inst/mem[74][5] ) );
  DFF_X1 \xmem_inst/mem_reg[74][6]  ( .D(n2245), .CK(clk), .Q(
        \xmem_inst/mem[74][6] ) );
  DFF_X1 \xmem_inst/mem_reg[74][7]  ( .D(n2244), .CK(clk), .Q(
        \xmem_inst/mem[74][7] ) );
  DFF_X1 \xmem_inst/mem_reg[75][0]  ( .D(n2243), .CK(clk), .Q(
        \xmem_inst/mem[75][0] ) );
  DFF_X1 \xmem_inst/mem_reg[75][1]  ( .D(n2242), .CK(clk), .Q(
        \xmem_inst/mem[75][1] ) );
  DFF_X1 \xmem_inst/mem_reg[75][2]  ( .D(n2241), .CK(clk), .Q(
        \xmem_inst/mem[75][2] ) );
  DFF_X1 \xmem_inst/mem_reg[75][3]  ( .D(n2240), .CK(clk), .Q(
        \xmem_inst/mem[75][3] ) );
  DFF_X1 \xmem_inst/mem_reg[75][4]  ( .D(n2239), .CK(clk), .Q(
        \xmem_inst/mem[75][4] ) );
  DFF_X1 \xmem_inst/mem_reg[75][5]  ( .D(n2238), .CK(clk), .Q(
        \xmem_inst/mem[75][5] ) );
  DFF_X1 \xmem_inst/mem_reg[75][6]  ( .D(n2237), .CK(clk), .Q(
        \xmem_inst/mem[75][6] ) );
  DFF_X1 \xmem_inst/mem_reg[75][7]  ( .D(n2236), .CK(clk), .Q(
        \xmem_inst/mem[75][7] ) );
  DFF_X1 \xmem_inst/mem_reg[76][0]  ( .D(n2235), .CK(clk), .Q(
        \xmem_inst/mem[76][0] ) );
  DFF_X1 \xmem_inst/mem_reg[76][1]  ( .D(n2234), .CK(clk), .Q(
        \xmem_inst/mem[76][1] ) );
  DFF_X1 \xmem_inst/mem_reg[76][2]  ( .D(n2233), .CK(clk), .Q(
        \xmem_inst/mem[76][2] ) );
  DFF_X1 \xmem_inst/mem_reg[76][3]  ( .D(n2232), .CK(clk), .Q(
        \xmem_inst/mem[76][3] ) );
  DFF_X1 \xmem_inst/mem_reg[76][4]  ( .D(n2231), .CK(clk), .Q(
        \xmem_inst/mem[76][4] ) );
  DFF_X1 \xmem_inst/mem_reg[76][5]  ( .D(n2230), .CK(clk), .Q(
        \xmem_inst/mem[76][5] ) );
  DFF_X1 \xmem_inst/mem_reg[76][6]  ( .D(n2229), .CK(clk), .Q(
        \xmem_inst/mem[76][6] ) );
  DFF_X1 \xmem_inst/mem_reg[76][7]  ( .D(n2228), .CK(clk), .Q(
        \xmem_inst/mem[76][7] ) );
  DFF_X1 \xmem_inst/mem_reg[77][0]  ( .D(n2227), .CK(clk), .Q(
        \xmem_inst/mem[77][0] ) );
  DFF_X1 \xmem_inst/mem_reg[77][1]  ( .D(n2226), .CK(clk), .Q(
        \xmem_inst/mem[77][1] ) );
  DFF_X1 \xmem_inst/mem_reg[77][2]  ( .D(n2225), .CK(clk), .Q(
        \xmem_inst/mem[77][2] ) );
  DFF_X1 \xmem_inst/mem_reg[77][3]  ( .D(n2224), .CK(clk), .Q(
        \xmem_inst/mem[77][3] ) );
  DFF_X1 \xmem_inst/mem_reg[77][4]  ( .D(n2223), .CK(clk), .Q(
        \xmem_inst/mem[77][4] ) );
  DFF_X1 \xmem_inst/mem_reg[77][5]  ( .D(n2222), .CK(clk), .Q(
        \xmem_inst/mem[77][5] ) );
  DFF_X1 \xmem_inst/mem_reg[77][6]  ( .D(n2221), .CK(clk), .Q(
        \xmem_inst/mem[77][6] ) );
  DFF_X1 \xmem_inst/mem_reg[77][7]  ( .D(n2220), .CK(clk), .Q(
        \xmem_inst/mem[77][7] ) );
  DFF_X1 \xmem_inst/mem_reg[78][0]  ( .D(n2219), .CK(clk), .Q(
        \xmem_inst/mem[78][0] ) );
  DFF_X1 \xmem_inst/mem_reg[78][1]  ( .D(n2218), .CK(clk), .Q(
        \xmem_inst/mem[78][1] ) );
  DFF_X1 \xmem_inst/mem_reg[78][2]  ( .D(n2217), .CK(clk), .Q(
        \xmem_inst/mem[78][2] ) );
  DFF_X1 \xmem_inst/mem_reg[78][3]  ( .D(n2216), .CK(clk), .Q(
        \xmem_inst/mem[78][3] ) );
  DFF_X1 \xmem_inst/mem_reg[78][4]  ( .D(n2215), .CK(clk), .Q(
        \xmem_inst/mem[78][4] ) );
  DFF_X1 \xmem_inst/mem_reg[78][5]  ( .D(n2214), .CK(clk), .Q(
        \xmem_inst/mem[78][5] ) );
  DFF_X1 \xmem_inst/mem_reg[78][6]  ( .D(n2213), .CK(clk), .Q(
        \xmem_inst/mem[78][6] ) );
  DFF_X1 \xmem_inst/mem_reg[78][7]  ( .D(n2212), .CK(clk), .Q(
        \xmem_inst/mem[78][7] ) );
  DFF_X1 \xmem_inst/mem_reg[79][0]  ( .D(n2211), .CK(clk), .Q(
        \xmem_inst/mem[79][0] ) );
  DFF_X1 \xmem_inst/mem_reg[79][1]  ( .D(n2210), .CK(clk), .Q(
        \xmem_inst/mem[79][1] ) );
  DFF_X1 \xmem_inst/mem_reg[79][2]  ( .D(n2209), .CK(clk), .Q(
        \xmem_inst/mem[79][2] ) );
  DFF_X1 \xmem_inst/mem_reg[79][3]  ( .D(n2208), .CK(clk), .Q(
        \xmem_inst/mem[79][3] ) );
  DFF_X1 \xmem_inst/mem_reg[79][4]  ( .D(n2207), .CK(clk), .Q(
        \xmem_inst/mem[79][4] ) );
  DFF_X1 \xmem_inst/mem_reg[79][5]  ( .D(n2206), .CK(clk), .Q(
        \xmem_inst/mem[79][5] ) );
  DFF_X1 \xmem_inst/mem_reg[79][6]  ( .D(n2205), .CK(clk), .Q(
        \xmem_inst/mem[79][6] ) );
  DFF_X1 \xmem_inst/mem_reg[79][7]  ( .D(n2204), .CK(clk), .Q(
        \xmem_inst/mem[79][7] ) );
  DFF_X1 \xmem_inst/mem_reg[80][0]  ( .D(n2203), .CK(clk), .Q(
        \xmem_inst/mem[80][0] ) );
  DFF_X1 \xmem_inst/mem_reg[80][1]  ( .D(n2202), .CK(clk), .Q(
        \xmem_inst/mem[80][1] ) );
  DFF_X1 \xmem_inst/mem_reg[80][2]  ( .D(n2201), .CK(clk), .Q(
        \xmem_inst/mem[80][2] ) );
  DFF_X1 \xmem_inst/mem_reg[80][3]  ( .D(n2200), .CK(clk), .Q(
        \xmem_inst/mem[80][3] ) );
  DFF_X1 \xmem_inst/mem_reg[80][4]  ( .D(n2199), .CK(clk), .Q(
        \xmem_inst/mem[80][4] ) );
  DFF_X1 \xmem_inst/mem_reg[80][5]  ( .D(n2198), .CK(clk), .Q(
        \xmem_inst/mem[80][5] ) );
  DFF_X1 \xmem_inst/mem_reg[80][6]  ( .D(n2197), .CK(clk), .Q(
        \xmem_inst/mem[80][6] ) );
  DFF_X1 \xmem_inst/mem_reg[80][7]  ( .D(n2196), .CK(clk), .Q(
        \xmem_inst/mem[80][7] ) );
  DFF_X1 \xmem_inst/mem_reg[81][0]  ( .D(n2195), .CK(clk), .Q(
        \xmem_inst/mem[81][0] ) );
  DFF_X1 \xmem_inst/mem_reg[81][1]  ( .D(n2194), .CK(clk), .Q(
        \xmem_inst/mem[81][1] ) );
  DFF_X1 \xmem_inst/mem_reg[81][2]  ( .D(n2193), .CK(clk), .Q(
        \xmem_inst/mem[81][2] ) );
  DFF_X1 \xmem_inst/mem_reg[81][3]  ( .D(n2192), .CK(clk), .Q(
        \xmem_inst/mem[81][3] ) );
  DFF_X1 \xmem_inst/mem_reg[81][4]  ( .D(n2191), .CK(clk), .Q(
        \xmem_inst/mem[81][4] ) );
  DFF_X1 \xmem_inst/mem_reg[81][5]  ( .D(n2190), .CK(clk), .Q(
        \xmem_inst/mem[81][5] ) );
  DFF_X1 \xmem_inst/mem_reg[81][6]  ( .D(n2189), .CK(clk), .Q(
        \xmem_inst/mem[81][6] ) );
  DFF_X1 \xmem_inst/mem_reg[81][7]  ( .D(n2188), .CK(clk), .Q(
        \xmem_inst/mem[81][7] ) );
  DFF_X1 \xmem_inst/mem_reg[82][0]  ( .D(n2187), .CK(clk), .Q(
        \xmem_inst/mem[82][0] ) );
  DFF_X1 \xmem_inst/mem_reg[82][1]  ( .D(n2186), .CK(clk), .Q(
        \xmem_inst/mem[82][1] ) );
  DFF_X1 \xmem_inst/mem_reg[82][2]  ( .D(n2185), .CK(clk), .Q(
        \xmem_inst/mem[82][2] ) );
  DFF_X1 \xmem_inst/mem_reg[82][3]  ( .D(n2184), .CK(clk), .Q(
        \xmem_inst/mem[82][3] ) );
  DFF_X1 \xmem_inst/mem_reg[82][4]  ( .D(n2183), .CK(clk), .Q(
        \xmem_inst/mem[82][4] ) );
  DFF_X1 \xmem_inst/mem_reg[82][5]  ( .D(n2182), .CK(clk), .Q(
        \xmem_inst/mem[82][5] ) );
  DFF_X1 \xmem_inst/mem_reg[82][6]  ( .D(n2181), .CK(clk), .Q(
        \xmem_inst/mem[82][6] ) );
  DFF_X1 \xmem_inst/mem_reg[82][7]  ( .D(n2180), .CK(clk), .Q(
        \xmem_inst/mem[82][7] ) );
  DFF_X1 \xmem_inst/mem_reg[83][0]  ( .D(n2179), .CK(clk), .Q(
        \xmem_inst/mem[83][0] ) );
  DFF_X1 \xmem_inst/mem_reg[83][1]  ( .D(n2178), .CK(clk), .Q(
        \xmem_inst/mem[83][1] ) );
  DFF_X1 \xmem_inst/mem_reg[83][2]  ( .D(n2177), .CK(clk), .Q(
        \xmem_inst/mem[83][2] ) );
  DFF_X1 \xmem_inst/mem_reg[83][3]  ( .D(n2176), .CK(clk), .Q(
        \xmem_inst/mem[83][3] ) );
  DFF_X1 \xmem_inst/mem_reg[83][4]  ( .D(n2175), .CK(clk), .Q(
        \xmem_inst/mem[83][4] ) );
  DFF_X1 \xmem_inst/mem_reg[83][5]  ( .D(n2174), .CK(clk), .Q(
        \xmem_inst/mem[83][5] ) );
  DFF_X1 \xmem_inst/mem_reg[83][6]  ( .D(n2173), .CK(clk), .Q(
        \xmem_inst/mem[83][6] ) );
  DFF_X1 \xmem_inst/mem_reg[83][7]  ( .D(n2172), .CK(clk), .Q(
        \xmem_inst/mem[83][7] ) );
  DFF_X1 \xmem_inst/mem_reg[84][0]  ( .D(n2171), .CK(clk), .Q(
        \xmem_inst/mem[84][0] ) );
  DFF_X1 \xmem_inst/mem_reg[84][1]  ( .D(n2170), .CK(clk), .Q(
        \xmem_inst/mem[84][1] ) );
  DFF_X1 \xmem_inst/mem_reg[84][2]  ( .D(n2169), .CK(clk), .Q(
        \xmem_inst/mem[84][2] ) );
  DFF_X1 \xmem_inst/mem_reg[84][3]  ( .D(n2168), .CK(clk), .Q(
        \xmem_inst/mem[84][3] ) );
  DFF_X1 \xmem_inst/mem_reg[84][4]  ( .D(n2167), .CK(clk), .Q(
        \xmem_inst/mem[84][4] ) );
  DFF_X1 \xmem_inst/mem_reg[84][5]  ( .D(n2166), .CK(clk), .Q(
        \xmem_inst/mem[84][5] ) );
  DFF_X1 \xmem_inst/mem_reg[84][6]  ( .D(n2165), .CK(clk), .Q(
        \xmem_inst/mem[84][6] ) );
  DFF_X1 \xmem_inst/mem_reg[84][7]  ( .D(n2164), .CK(clk), .Q(
        \xmem_inst/mem[84][7] ) );
  DFF_X1 \xmem_inst/mem_reg[85][0]  ( .D(n2163), .CK(clk), .Q(
        \xmem_inst/mem[85][0] ) );
  DFF_X1 \xmem_inst/mem_reg[85][1]  ( .D(n2162), .CK(clk), .Q(
        \xmem_inst/mem[85][1] ) );
  DFF_X1 \xmem_inst/mem_reg[85][2]  ( .D(n2161), .CK(clk), .Q(
        \xmem_inst/mem[85][2] ) );
  DFF_X1 \xmem_inst/mem_reg[85][3]  ( .D(n2160), .CK(clk), .Q(
        \xmem_inst/mem[85][3] ) );
  DFF_X1 \xmem_inst/mem_reg[85][4]  ( .D(n2159), .CK(clk), .Q(
        \xmem_inst/mem[85][4] ) );
  DFF_X1 \xmem_inst/mem_reg[85][5]  ( .D(n2158), .CK(clk), .Q(
        \xmem_inst/mem[85][5] ) );
  DFF_X1 \xmem_inst/mem_reg[85][6]  ( .D(n2157), .CK(clk), .Q(
        \xmem_inst/mem[85][6] ) );
  DFF_X1 \xmem_inst/mem_reg[85][7]  ( .D(n2156), .CK(clk), .Q(
        \xmem_inst/mem[85][7] ) );
  DFF_X1 \xmem_inst/mem_reg[86][0]  ( .D(n2155), .CK(clk), .Q(
        \xmem_inst/mem[86][0] ) );
  DFF_X1 \xmem_inst/mem_reg[86][1]  ( .D(n2154), .CK(clk), .Q(
        \xmem_inst/mem[86][1] ) );
  DFF_X1 \xmem_inst/mem_reg[86][2]  ( .D(n2153), .CK(clk), .Q(
        \xmem_inst/mem[86][2] ) );
  DFF_X1 \xmem_inst/mem_reg[86][3]  ( .D(n2152), .CK(clk), .Q(
        \xmem_inst/mem[86][3] ) );
  DFF_X1 \xmem_inst/mem_reg[86][4]  ( .D(n2151), .CK(clk), .Q(
        \xmem_inst/mem[86][4] ) );
  DFF_X1 \xmem_inst/mem_reg[86][5]  ( .D(n2150), .CK(clk), .Q(
        \xmem_inst/mem[86][5] ) );
  DFF_X1 \xmem_inst/mem_reg[86][6]  ( .D(n2149), .CK(clk), .Q(
        \xmem_inst/mem[86][6] ) );
  DFF_X1 \xmem_inst/mem_reg[86][7]  ( .D(n2148), .CK(clk), .Q(
        \xmem_inst/mem[86][7] ) );
  DFF_X1 \xmem_inst/mem_reg[87][0]  ( .D(n2147), .CK(clk), .Q(
        \xmem_inst/mem[87][0] ) );
  DFF_X1 \xmem_inst/mem_reg[87][1]  ( .D(n2146), .CK(clk), .Q(
        \xmem_inst/mem[87][1] ) );
  DFF_X1 \xmem_inst/mem_reg[87][2]  ( .D(n2145), .CK(clk), .Q(
        \xmem_inst/mem[87][2] ) );
  DFF_X1 \xmem_inst/mem_reg[87][3]  ( .D(n2144), .CK(clk), .Q(
        \xmem_inst/mem[87][3] ) );
  DFF_X1 \xmem_inst/mem_reg[87][4]  ( .D(n2143), .CK(clk), .Q(
        \xmem_inst/mem[87][4] ) );
  DFF_X1 \xmem_inst/mem_reg[87][5]  ( .D(n2142), .CK(clk), .Q(
        \xmem_inst/mem[87][5] ) );
  DFF_X1 \xmem_inst/mem_reg[87][6]  ( .D(n2141), .CK(clk), .Q(
        \xmem_inst/mem[87][6] ) );
  DFF_X1 \xmem_inst/mem_reg[87][7]  ( .D(n2140), .CK(clk), .Q(
        \xmem_inst/mem[87][7] ) );
  DFF_X1 \xmem_inst/mem_reg[88][0]  ( .D(n2139), .CK(clk), .Q(
        \xmem_inst/mem[88][0] ) );
  DFF_X1 \xmem_inst/mem_reg[88][1]  ( .D(n2138), .CK(clk), .Q(
        \xmem_inst/mem[88][1] ) );
  DFF_X1 \xmem_inst/mem_reg[88][2]  ( .D(n2137), .CK(clk), .Q(
        \xmem_inst/mem[88][2] ) );
  DFF_X1 \xmem_inst/mem_reg[88][3]  ( .D(n2136), .CK(clk), .Q(
        \xmem_inst/mem[88][3] ) );
  DFF_X1 \xmem_inst/mem_reg[88][4]  ( .D(n2135), .CK(clk), .Q(
        \xmem_inst/mem[88][4] ) );
  DFF_X1 \xmem_inst/mem_reg[88][5]  ( .D(n2134), .CK(clk), .Q(
        \xmem_inst/mem[88][5] ) );
  DFF_X1 \xmem_inst/mem_reg[88][6]  ( .D(n2133), .CK(clk), .Q(
        \xmem_inst/mem[88][6] ) );
  DFF_X1 \xmem_inst/mem_reg[88][7]  ( .D(n2132), .CK(clk), .Q(
        \xmem_inst/mem[88][7] ) );
  DFF_X1 \xmem_inst/mem_reg[89][0]  ( .D(n2131), .CK(clk), .Q(
        \xmem_inst/mem[89][0] ) );
  DFF_X1 \xmem_inst/mem_reg[89][1]  ( .D(n2130), .CK(clk), .Q(
        \xmem_inst/mem[89][1] ) );
  DFF_X1 \xmem_inst/mem_reg[89][2]  ( .D(n2129), .CK(clk), .Q(
        \xmem_inst/mem[89][2] ) );
  DFF_X1 \xmem_inst/mem_reg[89][3]  ( .D(n2128), .CK(clk), .Q(
        \xmem_inst/mem[89][3] ) );
  DFF_X1 \xmem_inst/mem_reg[89][4]  ( .D(n2127), .CK(clk), .Q(
        \xmem_inst/mem[89][4] ) );
  DFF_X1 \xmem_inst/mem_reg[89][5]  ( .D(n2126), .CK(clk), .Q(
        \xmem_inst/mem[89][5] ) );
  DFF_X1 \xmem_inst/mem_reg[89][6]  ( .D(n2125), .CK(clk), .Q(
        \xmem_inst/mem[89][6] ) );
  DFF_X1 \xmem_inst/mem_reg[89][7]  ( .D(n2124), .CK(clk), .Q(
        \xmem_inst/mem[89][7] ) );
  DFF_X1 \xmem_inst/mem_reg[90][0]  ( .D(n2123), .CK(clk), .Q(
        \xmem_inst/mem[90][0] ) );
  DFF_X1 \xmem_inst/mem_reg[90][1]  ( .D(n2122), .CK(clk), .Q(
        \xmem_inst/mem[90][1] ) );
  DFF_X1 \xmem_inst/mem_reg[90][2]  ( .D(n2121), .CK(clk), .Q(
        \xmem_inst/mem[90][2] ) );
  DFF_X1 \xmem_inst/mem_reg[90][3]  ( .D(n2120), .CK(clk), .Q(
        \xmem_inst/mem[90][3] ) );
  DFF_X1 \xmem_inst/mem_reg[90][4]  ( .D(n2119), .CK(clk), .Q(
        \xmem_inst/mem[90][4] ) );
  DFF_X1 \xmem_inst/mem_reg[90][5]  ( .D(n2118), .CK(clk), .Q(
        \xmem_inst/mem[90][5] ) );
  DFF_X1 \xmem_inst/mem_reg[90][6]  ( .D(n2117), .CK(clk), .Q(
        \xmem_inst/mem[90][6] ) );
  DFF_X1 \xmem_inst/mem_reg[90][7]  ( .D(n2116), .CK(clk), .Q(
        \xmem_inst/mem[90][7] ) );
  DFF_X1 \xmem_inst/mem_reg[91][0]  ( .D(n2115), .CK(clk), .Q(
        \xmem_inst/mem[91][0] ) );
  DFF_X1 \xmem_inst/mem_reg[91][1]  ( .D(n2114), .CK(clk), .Q(
        \xmem_inst/mem[91][1] ) );
  DFF_X1 \xmem_inst/mem_reg[91][2]  ( .D(n2113), .CK(clk), .Q(
        \xmem_inst/mem[91][2] ) );
  DFF_X1 \xmem_inst/mem_reg[91][3]  ( .D(n2112), .CK(clk), .Q(
        \xmem_inst/mem[91][3] ) );
  DFF_X1 \xmem_inst/mem_reg[91][4]  ( .D(n2111), .CK(clk), .Q(
        \xmem_inst/mem[91][4] ) );
  DFF_X1 \xmem_inst/mem_reg[91][5]  ( .D(n2110), .CK(clk), .Q(
        \xmem_inst/mem[91][5] ) );
  DFF_X1 \xmem_inst/mem_reg[91][6]  ( .D(n2109), .CK(clk), .Q(
        \xmem_inst/mem[91][6] ) );
  DFF_X1 \xmem_inst/mem_reg[91][7]  ( .D(n2108), .CK(clk), .Q(
        \xmem_inst/mem[91][7] ) );
  DFF_X1 \xmem_inst/mem_reg[92][0]  ( .D(n2107), .CK(clk), .Q(
        \xmem_inst/mem[92][0] ) );
  DFF_X1 \xmem_inst/mem_reg[92][1]  ( .D(n2106), .CK(clk), .Q(
        \xmem_inst/mem[92][1] ) );
  DFF_X1 \xmem_inst/mem_reg[92][2]  ( .D(n2105), .CK(clk), .Q(
        \xmem_inst/mem[92][2] ) );
  DFF_X1 \xmem_inst/mem_reg[92][3]  ( .D(n2104), .CK(clk), .Q(
        \xmem_inst/mem[92][3] ) );
  DFF_X1 \xmem_inst/mem_reg[92][4]  ( .D(n2103), .CK(clk), .Q(
        \xmem_inst/mem[92][4] ) );
  DFF_X1 \xmem_inst/mem_reg[92][5]  ( .D(n2102), .CK(clk), .Q(
        \xmem_inst/mem[92][5] ) );
  DFF_X1 \xmem_inst/mem_reg[92][6]  ( .D(n2101), .CK(clk), .Q(
        \xmem_inst/mem[92][6] ) );
  DFF_X1 \xmem_inst/mem_reg[92][7]  ( .D(n2100), .CK(clk), .Q(
        \xmem_inst/mem[92][7] ) );
  DFF_X1 \xmem_inst/mem_reg[93][0]  ( .D(n2099), .CK(clk), .Q(
        \xmem_inst/mem[93][0] ) );
  DFF_X1 \xmem_inst/mem_reg[93][1]  ( .D(n2098), .CK(clk), .Q(
        \xmem_inst/mem[93][1] ) );
  DFF_X1 \xmem_inst/mem_reg[93][2]  ( .D(n2097), .CK(clk), .Q(
        \xmem_inst/mem[93][2] ) );
  DFF_X1 \xmem_inst/mem_reg[93][3]  ( .D(n2096), .CK(clk), .Q(
        \xmem_inst/mem[93][3] ) );
  DFF_X1 \xmem_inst/mem_reg[93][4]  ( .D(n2095), .CK(clk), .Q(
        \xmem_inst/mem[93][4] ) );
  DFF_X1 \xmem_inst/mem_reg[93][5]  ( .D(n2094), .CK(clk), .Q(
        \xmem_inst/mem[93][5] ) );
  DFF_X1 \xmem_inst/mem_reg[93][6]  ( .D(n2093), .CK(clk), .Q(
        \xmem_inst/mem[93][6] ) );
  DFF_X1 \xmem_inst/mem_reg[93][7]  ( .D(n2092), .CK(clk), .Q(
        \xmem_inst/mem[93][7] ) );
  DFF_X1 \xmem_inst/mem_reg[94][0]  ( .D(n2091), .CK(clk), .Q(
        \xmem_inst/mem[94][0] ) );
  DFF_X1 \xmem_inst/mem_reg[94][1]  ( .D(n2090), .CK(clk), .Q(
        \xmem_inst/mem[94][1] ) );
  DFF_X1 \xmem_inst/mem_reg[94][2]  ( .D(n2089), .CK(clk), .Q(
        \xmem_inst/mem[94][2] ) );
  DFF_X1 \xmem_inst/mem_reg[94][3]  ( .D(n2088), .CK(clk), .Q(
        \xmem_inst/mem[94][3] ) );
  DFF_X1 \xmem_inst/mem_reg[94][4]  ( .D(n2087), .CK(clk), .Q(
        \xmem_inst/mem[94][4] ) );
  DFF_X1 \xmem_inst/mem_reg[94][5]  ( .D(n2086), .CK(clk), .Q(
        \xmem_inst/mem[94][5] ) );
  DFF_X1 \xmem_inst/mem_reg[94][6]  ( .D(n2085), .CK(clk), .Q(
        \xmem_inst/mem[94][6] ) );
  DFF_X1 \xmem_inst/mem_reg[94][7]  ( .D(n2084), .CK(clk), .Q(
        \xmem_inst/mem[94][7] ) );
  DFF_X1 \xmem_inst/mem_reg[95][0]  ( .D(n2083), .CK(clk), .Q(
        \xmem_inst/mem[95][0] ) );
  DFF_X1 \xmem_inst/mem_reg[95][1]  ( .D(n2082), .CK(clk), .Q(
        \xmem_inst/mem[95][1] ) );
  DFF_X1 \xmem_inst/mem_reg[95][2]  ( .D(n2081), .CK(clk), .Q(
        \xmem_inst/mem[95][2] ) );
  DFF_X1 \xmem_inst/mem_reg[95][3]  ( .D(n2080), .CK(clk), .Q(
        \xmem_inst/mem[95][3] ) );
  DFF_X1 \xmem_inst/mem_reg[95][4]  ( .D(n2079), .CK(clk), .Q(
        \xmem_inst/mem[95][4] ) );
  DFF_X1 \xmem_inst/mem_reg[95][5]  ( .D(n2078), .CK(clk), .Q(
        \xmem_inst/mem[95][5] ) );
  DFF_X1 \xmem_inst/mem_reg[95][6]  ( .D(n2077), .CK(clk), .Q(
        \xmem_inst/mem[95][6] ) );
  DFF_X1 \xmem_inst/mem_reg[95][7]  ( .D(n2076), .CK(clk), .Q(
        \xmem_inst/mem[95][7] ) );
  DFF_X1 \xmem_inst/mem_reg[96][0]  ( .D(n2075), .CK(clk), .Q(
        \xmem_inst/mem[96][0] ) );
  DFF_X1 \xmem_inst/mem_reg[96][1]  ( .D(n2074), .CK(clk), .Q(
        \xmem_inst/mem[96][1] ) );
  DFF_X1 \xmem_inst/mem_reg[96][2]  ( .D(n2073), .CK(clk), .Q(
        \xmem_inst/mem[96][2] ) );
  DFF_X1 \xmem_inst/mem_reg[96][3]  ( .D(n2072), .CK(clk), .Q(
        \xmem_inst/mem[96][3] ) );
  DFF_X1 \xmem_inst/mem_reg[96][4]  ( .D(n2071), .CK(clk), .Q(
        \xmem_inst/mem[96][4] ) );
  DFF_X1 \xmem_inst/mem_reg[96][5]  ( .D(n2070), .CK(clk), .Q(
        \xmem_inst/mem[96][5] ) );
  DFF_X1 \xmem_inst/mem_reg[96][6]  ( .D(n2069), .CK(clk), .Q(
        \xmem_inst/mem[96][6] ) );
  DFF_X1 \xmem_inst/mem_reg[96][7]  ( .D(n2068), .CK(clk), .Q(
        \xmem_inst/mem[96][7] ) );
  DFF_X1 \xmem_inst/mem_reg[97][0]  ( .D(n2067), .CK(clk), .Q(
        \xmem_inst/mem[97][0] ) );
  DFF_X1 \xmem_inst/mem_reg[97][1]  ( .D(n2066), .CK(clk), .Q(
        \xmem_inst/mem[97][1] ) );
  DFF_X1 \xmem_inst/mem_reg[97][2]  ( .D(n2065), .CK(clk), .Q(
        \xmem_inst/mem[97][2] ) );
  DFF_X1 \xmem_inst/mem_reg[97][3]  ( .D(n2064), .CK(clk), .Q(
        \xmem_inst/mem[97][3] ) );
  DFF_X1 \xmem_inst/mem_reg[97][4]  ( .D(n2063), .CK(clk), .Q(
        \xmem_inst/mem[97][4] ) );
  DFF_X1 \xmem_inst/mem_reg[97][5]  ( .D(n2062), .CK(clk), .Q(
        \xmem_inst/mem[97][5] ) );
  DFF_X1 \xmem_inst/mem_reg[97][6]  ( .D(n2061), .CK(clk), .Q(
        \xmem_inst/mem[97][6] ) );
  DFF_X1 \xmem_inst/mem_reg[97][7]  ( .D(n2060), .CK(clk), .Q(
        \xmem_inst/mem[97][7] ) );
  DFF_X1 \xmem_inst/mem_reg[98][0]  ( .D(n2059), .CK(clk), .Q(
        \xmem_inst/mem[98][0] ) );
  DFF_X1 \xmem_inst/mem_reg[98][1]  ( .D(n2058), .CK(clk), .Q(
        \xmem_inst/mem[98][1] ) );
  DFF_X1 \xmem_inst/mem_reg[98][2]  ( .D(n2057), .CK(clk), .Q(
        \xmem_inst/mem[98][2] ) );
  DFF_X1 \xmem_inst/mem_reg[98][3]  ( .D(n2056), .CK(clk), .Q(
        \xmem_inst/mem[98][3] ) );
  DFF_X1 \xmem_inst/mem_reg[98][4]  ( .D(n2055), .CK(clk), .Q(
        \xmem_inst/mem[98][4] ) );
  DFF_X1 \xmem_inst/mem_reg[98][5]  ( .D(n2054), .CK(clk), .Q(
        \xmem_inst/mem[98][5] ) );
  DFF_X1 \xmem_inst/mem_reg[98][6]  ( .D(n2053), .CK(clk), .Q(
        \xmem_inst/mem[98][6] ) );
  DFF_X1 \xmem_inst/mem_reg[98][7]  ( .D(n2052), .CK(clk), .Q(
        \xmem_inst/mem[98][7] ) );
  DFF_X1 \xmem_inst/mem_reg[99][0]  ( .D(n2051), .CK(clk), .Q(
        \xmem_inst/mem[99][0] ) );
  DFF_X1 \xmem_inst/mem_reg[99][1]  ( .D(n2050), .CK(clk), .Q(
        \xmem_inst/mem[99][1] ) );
  DFF_X1 \xmem_inst/mem_reg[99][2]  ( .D(n2049), .CK(clk), .Q(
        \xmem_inst/mem[99][2] ) );
  DFF_X1 \xmem_inst/mem_reg[99][3]  ( .D(n2048), .CK(clk), .Q(
        \xmem_inst/mem[99][3] ) );
  DFF_X1 \xmem_inst/mem_reg[99][4]  ( .D(n2047), .CK(clk), .Q(
        \xmem_inst/mem[99][4] ) );
  DFF_X1 \xmem_inst/mem_reg[99][5]  ( .D(n2046), .CK(clk), .Q(
        \xmem_inst/mem[99][5] ) );
  DFF_X1 \xmem_inst/mem_reg[99][6]  ( .D(n2045), .CK(clk), .Q(
        \xmem_inst/mem[99][6] ) );
  DFF_X1 \xmem_inst/mem_reg[99][7]  ( .D(n2044), .CK(clk), .Q(
        \xmem_inst/mem[99][7] ) );
  DFF_X1 \xmem_inst/mem_reg[100][0]  ( .D(n2043), .CK(clk), .Q(
        \xmem_inst/mem[100][0] ) );
  DFF_X1 \xmem_inst/mem_reg[100][1]  ( .D(n2042), .CK(clk), .Q(
        \xmem_inst/mem[100][1] ) );
  DFF_X1 \xmem_inst/mem_reg[100][2]  ( .D(n2041), .CK(clk), .Q(
        \xmem_inst/mem[100][2] ) );
  DFF_X1 \xmem_inst/mem_reg[100][3]  ( .D(n2040), .CK(clk), .Q(
        \xmem_inst/mem[100][3] ) );
  DFF_X1 \xmem_inst/mem_reg[100][4]  ( .D(n2039), .CK(clk), .Q(
        \xmem_inst/mem[100][4] ) );
  DFF_X1 \xmem_inst/mem_reg[100][5]  ( .D(n2038), .CK(clk), .Q(
        \xmem_inst/mem[100][5] ) );
  DFF_X1 \xmem_inst/mem_reg[100][6]  ( .D(n2037), .CK(clk), .Q(
        \xmem_inst/mem[100][6] ) );
  DFF_X1 \xmem_inst/mem_reg[100][7]  ( .D(n2036), .CK(clk), .Q(
        \xmem_inst/mem[100][7] ) );
  DFF_X1 \xmem_inst/mem_reg[101][0]  ( .D(n2035), .CK(clk), .Q(
        \xmem_inst/mem[101][0] ) );
  DFF_X1 \xmem_inst/mem_reg[101][1]  ( .D(n2034), .CK(clk), .Q(
        \xmem_inst/mem[101][1] ) );
  DFF_X1 \xmem_inst/mem_reg[101][2]  ( .D(n2033), .CK(clk), .Q(
        \xmem_inst/mem[101][2] ) );
  DFF_X1 \xmem_inst/mem_reg[101][3]  ( .D(n2032), .CK(clk), .Q(
        \xmem_inst/mem[101][3] ) );
  DFF_X1 \xmem_inst/mem_reg[101][4]  ( .D(n2031), .CK(clk), .Q(
        \xmem_inst/mem[101][4] ) );
  DFF_X1 \xmem_inst/mem_reg[101][5]  ( .D(n2030), .CK(clk), .Q(
        \xmem_inst/mem[101][5] ) );
  DFF_X1 \xmem_inst/mem_reg[101][6]  ( .D(n2029), .CK(clk), .Q(
        \xmem_inst/mem[101][6] ) );
  DFF_X1 \xmem_inst/mem_reg[101][7]  ( .D(n2028), .CK(clk), .Q(
        \xmem_inst/mem[101][7] ) );
  DFF_X1 \xmem_inst/mem_reg[102][0]  ( .D(n2027), .CK(clk), .Q(
        \xmem_inst/mem[102][0] ) );
  DFF_X1 \xmem_inst/mem_reg[102][1]  ( .D(n2026), .CK(clk), .Q(
        \xmem_inst/mem[102][1] ) );
  DFF_X1 \xmem_inst/mem_reg[102][2]  ( .D(n2025), .CK(clk), .Q(
        \xmem_inst/mem[102][2] ) );
  DFF_X1 \xmem_inst/mem_reg[102][3]  ( .D(n2024), .CK(clk), .Q(
        \xmem_inst/mem[102][3] ) );
  DFF_X1 \xmem_inst/mem_reg[102][4]  ( .D(n2023), .CK(clk), .Q(
        \xmem_inst/mem[102][4] ) );
  DFF_X1 \xmem_inst/mem_reg[102][5]  ( .D(n2022), .CK(clk), .Q(
        \xmem_inst/mem[102][5] ) );
  DFF_X1 \xmem_inst/mem_reg[102][6]  ( .D(n2021), .CK(clk), .Q(
        \xmem_inst/mem[102][6] ) );
  DFF_X1 \xmem_inst/mem_reg[102][7]  ( .D(n2020), .CK(clk), .Q(
        \xmem_inst/mem[102][7] ) );
  DFF_X1 \xmem_inst/mem_reg[103][0]  ( .D(n2019), .CK(clk), .Q(
        \xmem_inst/mem[103][0] ) );
  DFF_X1 \xmem_inst/mem_reg[103][1]  ( .D(n2018), .CK(clk), .Q(
        \xmem_inst/mem[103][1] ) );
  DFF_X1 \xmem_inst/mem_reg[103][2]  ( .D(n2017), .CK(clk), .Q(
        \xmem_inst/mem[103][2] ) );
  DFF_X1 \xmem_inst/mem_reg[103][3]  ( .D(n2016), .CK(clk), .Q(
        \xmem_inst/mem[103][3] ) );
  DFF_X1 \xmem_inst/mem_reg[103][4]  ( .D(n2015), .CK(clk), .Q(
        \xmem_inst/mem[103][4] ) );
  DFF_X1 \xmem_inst/mem_reg[103][5]  ( .D(n2014), .CK(clk), .Q(
        \xmem_inst/mem[103][5] ) );
  DFF_X1 \xmem_inst/mem_reg[103][6]  ( .D(n2013), .CK(clk), .Q(
        \xmem_inst/mem[103][6] ) );
  DFF_X1 \xmem_inst/mem_reg[103][7]  ( .D(n2012), .CK(clk), .Q(
        \xmem_inst/mem[103][7] ) );
  DFF_X1 \xmem_inst/mem_reg[104][0]  ( .D(n2011), .CK(clk), .Q(
        \xmem_inst/mem[104][0] ) );
  DFF_X1 \xmem_inst/mem_reg[104][1]  ( .D(n2010), .CK(clk), .Q(
        \xmem_inst/mem[104][1] ) );
  DFF_X1 \xmem_inst/mem_reg[104][2]  ( .D(n2009), .CK(clk), .Q(
        \xmem_inst/mem[104][2] ) );
  DFF_X1 \xmem_inst/mem_reg[104][3]  ( .D(n2008), .CK(clk), .Q(
        \xmem_inst/mem[104][3] ) );
  DFF_X1 \xmem_inst/mem_reg[104][4]  ( .D(n2007), .CK(clk), .Q(
        \xmem_inst/mem[104][4] ) );
  DFF_X1 \xmem_inst/mem_reg[104][5]  ( .D(n2006), .CK(clk), .Q(
        \xmem_inst/mem[104][5] ) );
  DFF_X1 \xmem_inst/mem_reg[104][6]  ( .D(n2005), .CK(clk), .Q(
        \xmem_inst/mem[104][6] ) );
  DFF_X1 \xmem_inst/mem_reg[104][7]  ( .D(n2004), .CK(clk), .Q(
        \xmem_inst/mem[104][7] ) );
  DFF_X1 \xmem_inst/mem_reg[105][0]  ( .D(n2003), .CK(clk), .Q(
        \xmem_inst/mem[105][0] ) );
  DFF_X1 \xmem_inst/mem_reg[105][1]  ( .D(n2002), .CK(clk), .Q(
        \xmem_inst/mem[105][1] ) );
  DFF_X1 \xmem_inst/mem_reg[105][2]  ( .D(n2001), .CK(clk), .Q(
        \xmem_inst/mem[105][2] ) );
  DFF_X1 \xmem_inst/mem_reg[105][3]  ( .D(n2000), .CK(clk), .Q(
        \xmem_inst/mem[105][3] ) );
  DFF_X1 \xmem_inst/mem_reg[105][4]  ( .D(n1999), .CK(clk), .Q(
        \xmem_inst/mem[105][4] ) );
  DFF_X1 \xmem_inst/mem_reg[105][5]  ( .D(n1998), .CK(clk), .Q(
        \xmem_inst/mem[105][5] ) );
  DFF_X1 \xmem_inst/mem_reg[105][6]  ( .D(n1997), .CK(clk), .Q(
        \xmem_inst/mem[105][6] ) );
  DFF_X1 \xmem_inst/mem_reg[105][7]  ( .D(n1996), .CK(clk), .Q(
        \xmem_inst/mem[105][7] ) );
  DFF_X1 \xmem_inst/mem_reg[106][0]  ( .D(n1995), .CK(clk), .Q(
        \xmem_inst/mem[106][0] ) );
  DFF_X1 \xmem_inst/mem_reg[106][1]  ( .D(n1994), .CK(clk), .Q(
        \xmem_inst/mem[106][1] ) );
  DFF_X1 \xmem_inst/mem_reg[106][2]  ( .D(n1993), .CK(clk), .Q(
        \xmem_inst/mem[106][2] ) );
  DFF_X1 \xmem_inst/mem_reg[106][3]  ( .D(n1992), .CK(clk), .Q(
        \xmem_inst/mem[106][3] ) );
  DFF_X1 \xmem_inst/mem_reg[106][4]  ( .D(n1991), .CK(clk), .Q(
        \xmem_inst/mem[106][4] ) );
  DFF_X1 \xmem_inst/mem_reg[106][5]  ( .D(n1990), .CK(clk), .Q(
        \xmem_inst/mem[106][5] ) );
  DFF_X1 \xmem_inst/mem_reg[106][6]  ( .D(n1989), .CK(clk), .Q(
        \xmem_inst/mem[106][6] ) );
  DFF_X1 \xmem_inst/mem_reg[106][7]  ( .D(n1988), .CK(clk), .Q(
        \xmem_inst/mem[106][7] ) );
  DFF_X1 \xmem_inst/mem_reg[107][0]  ( .D(n1987), .CK(clk), .Q(
        \xmem_inst/mem[107][0] ) );
  DFF_X1 \xmem_inst/mem_reg[107][1]  ( .D(n1986), .CK(clk), .Q(
        \xmem_inst/mem[107][1] ) );
  DFF_X1 \xmem_inst/mem_reg[107][2]  ( .D(n1985), .CK(clk), .Q(
        \xmem_inst/mem[107][2] ) );
  DFF_X1 \xmem_inst/mem_reg[107][3]  ( .D(n1984), .CK(clk), .Q(
        \xmem_inst/mem[107][3] ) );
  DFF_X1 \xmem_inst/mem_reg[107][4]  ( .D(n1983), .CK(clk), .Q(
        \xmem_inst/mem[107][4] ) );
  DFF_X1 \xmem_inst/mem_reg[107][5]  ( .D(n1982), .CK(clk), .Q(
        \xmem_inst/mem[107][5] ) );
  DFF_X1 \xmem_inst/mem_reg[107][6]  ( .D(n1981), .CK(clk), .Q(
        \xmem_inst/mem[107][6] ) );
  DFF_X1 \xmem_inst/mem_reg[107][7]  ( .D(n1980), .CK(clk), .Q(
        \xmem_inst/mem[107][7] ) );
  DFF_X1 \xmem_inst/mem_reg[108][0]  ( .D(n1979), .CK(clk), .Q(
        \xmem_inst/mem[108][0] ) );
  DFF_X1 \xmem_inst/mem_reg[108][1]  ( .D(n1978), .CK(clk), .Q(
        \xmem_inst/mem[108][1] ) );
  DFF_X1 \xmem_inst/mem_reg[108][2]  ( .D(n1977), .CK(clk), .Q(
        \xmem_inst/mem[108][2] ) );
  DFF_X1 \xmem_inst/mem_reg[108][3]  ( .D(n1976), .CK(clk), .Q(
        \xmem_inst/mem[108][3] ) );
  DFF_X1 \xmem_inst/mem_reg[108][4]  ( .D(n1975), .CK(clk), .Q(
        \xmem_inst/mem[108][4] ) );
  DFF_X1 \xmem_inst/mem_reg[108][5]  ( .D(n1974), .CK(clk), .Q(
        \xmem_inst/mem[108][5] ) );
  DFF_X1 \xmem_inst/mem_reg[108][6]  ( .D(n1973), .CK(clk), .Q(
        \xmem_inst/mem[108][6] ) );
  DFF_X1 \xmem_inst/mem_reg[108][7]  ( .D(n1972), .CK(clk), .Q(
        \xmem_inst/mem[108][7] ) );
  DFF_X1 \xmem_inst/mem_reg[109][0]  ( .D(n1971), .CK(clk), .Q(
        \xmem_inst/mem[109][0] ) );
  DFF_X1 \xmem_inst/mem_reg[109][1]  ( .D(n1970), .CK(clk), .Q(
        \xmem_inst/mem[109][1] ) );
  DFF_X1 \xmem_inst/mem_reg[109][2]  ( .D(n1969), .CK(clk), .Q(
        \xmem_inst/mem[109][2] ) );
  DFF_X1 \xmem_inst/mem_reg[109][3]  ( .D(n1968), .CK(clk), .Q(
        \xmem_inst/mem[109][3] ) );
  DFF_X1 \xmem_inst/mem_reg[109][4]  ( .D(n1967), .CK(clk), .Q(
        \xmem_inst/mem[109][4] ) );
  DFF_X1 \xmem_inst/mem_reg[109][5]  ( .D(n1966), .CK(clk), .Q(
        \xmem_inst/mem[109][5] ) );
  DFF_X1 \xmem_inst/mem_reg[109][6]  ( .D(n1965), .CK(clk), .Q(
        \xmem_inst/mem[109][6] ) );
  DFF_X1 \xmem_inst/mem_reg[109][7]  ( .D(n1964), .CK(clk), .Q(
        \xmem_inst/mem[109][7] ) );
  DFF_X1 \xmem_inst/mem_reg[110][0]  ( .D(n1963), .CK(clk), .Q(
        \xmem_inst/mem[110][0] ) );
  DFF_X1 \xmem_inst/mem_reg[110][1]  ( .D(n1962), .CK(clk), .Q(
        \xmem_inst/mem[110][1] ) );
  DFF_X1 \xmem_inst/mem_reg[110][2]  ( .D(n1961), .CK(clk), .Q(
        \xmem_inst/mem[110][2] ) );
  DFF_X1 \xmem_inst/mem_reg[110][3]  ( .D(n1960), .CK(clk), .Q(
        \xmem_inst/mem[110][3] ) );
  DFF_X1 \xmem_inst/mem_reg[110][4]  ( .D(n1959), .CK(clk), .Q(
        \xmem_inst/mem[110][4] ) );
  DFF_X1 \xmem_inst/mem_reg[110][5]  ( .D(n1958), .CK(clk), .Q(
        \xmem_inst/mem[110][5] ) );
  DFF_X1 \xmem_inst/mem_reg[110][6]  ( .D(n1957), .CK(clk), .Q(
        \xmem_inst/mem[110][6] ) );
  DFF_X1 \xmem_inst/mem_reg[110][7]  ( .D(n1956), .CK(clk), .Q(
        \xmem_inst/mem[110][7] ) );
  DFF_X1 \xmem_inst/mem_reg[111][0]  ( .D(n1955), .CK(clk), .Q(
        \xmem_inst/mem[111][0] ) );
  DFF_X1 \xmem_inst/mem_reg[111][1]  ( .D(n1954), .CK(clk), .Q(
        \xmem_inst/mem[111][1] ) );
  DFF_X1 \xmem_inst/mem_reg[111][2]  ( .D(n1953), .CK(clk), .Q(
        \xmem_inst/mem[111][2] ) );
  DFF_X1 \xmem_inst/mem_reg[111][3]  ( .D(n1952), .CK(clk), .Q(
        \xmem_inst/mem[111][3] ) );
  DFF_X1 \xmem_inst/mem_reg[111][4]  ( .D(n1951), .CK(clk), .Q(
        \xmem_inst/mem[111][4] ) );
  DFF_X1 \xmem_inst/mem_reg[111][5]  ( .D(n1950), .CK(clk), .Q(
        \xmem_inst/mem[111][5] ) );
  DFF_X1 \xmem_inst/mem_reg[111][6]  ( .D(n1949), .CK(clk), .Q(
        \xmem_inst/mem[111][6] ) );
  DFF_X1 \xmem_inst/mem_reg[111][7]  ( .D(n1948), .CK(clk), .Q(
        \xmem_inst/mem[111][7] ) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[0]  ( .D(n3112), .CK(clk), .Q(
        fmem_addr[0]), .QN(n39046) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[1]  ( .D(n3111), .CK(clk), .Q(
        fmem_addr[1]), .QN(n39047) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[2]  ( .D(n3110), .CK(clk), .Q(
        fmem_addr[2]), .QN(n39000) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[3]  ( .D(n3109), .CK(clk), .Q(
        fmem_addr[3]) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[4]  ( .D(n3108), .CK(clk), .Q(
        fmem_addr[4]), .QN(n39045) );
  DFF_X1 \fmem_inst/mem_reg[24][0]  ( .D(n2915), .CK(clk), .Q(
        \fmem_inst/mem[24][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][0]  ( .D(\fmem_inst/mem[24][0] ), .CK(clk), .Q(\fmem_data[24][0] ), .QN(n3565) );
  DFF_X1 \fmem_inst/mem_reg[24][1]  ( .D(n2914), .CK(clk), .Q(
        \fmem_inst/mem[24][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][1]  ( .D(\fmem_inst/mem[24][1] ), .CK(clk), .Q(\fmem_data[24][1] ), .QN(n3670) );
  DFF_X1 \fmem_inst/mem_reg[24][2]  ( .D(n2913), .CK(clk), .Q(
        \fmem_inst/mem[24][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][2]  ( .D(\fmem_inst/mem[24][2] ), .CK(clk), .Q(\fmem_data[24][2] ) );
  DFF_X1 \fmem_inst/mem_reg[24][3]  ( .D(n2912), .CK(clk), .Q(
        \fmem_inst/mem[24][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][3]  ( .D(\fmem_inst/mem[24][3] ), .CK(clk), .Q(\fmem_data[24][3] ), .QN(n3605) );
  DFF_X1 \fmem_inst/mem_reg[24][4]  ( .D(n2911), .CK(clk), .Q(
        \fmem_inst/mem[24][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][4]  ( .D(\fmem_inst/mem[24][4] ), .CK(clk), .Q(\fmem_data[24][4] ) );
  DFF_X1 \fmem_inst/mem_reg[24][5]  ( .D(n2910), .CK(clk), .Q(
        \fmem_inst/mem[24][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][5]  ( .D(\fmem_inst/mem[24][5] ), .CK(clk), .Q(\fmem_data[24][5] ), .QN(n3651) );
  DFF_X1 \fmem_inst/mem_reg[24][6]  ( .D(n2909), .CK(clk), .Q(
        \fmem_inst/mem[24][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][6]  ( .D(\fmem_inst/mem[24][6] ), .CK(clk), .Q(\fmem_data[24][6] ) );
  DFF_X1 \fmem_inst/mem_reg[24][7]  ( .D(n2908), .CK(clk), .Q(
        \fmem_inst/mem[24][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[24][7]  ( .D(\fmem_inst/mem[24][7] ), .CK(clk), .Q(\fmem_data[24][7] ), .QN(n3599) );
  DFF_X1 \fmem_inst/mem_reg[25][0]  ( .D(n2907), .CK(clk), .Q(
        \fmem_inst/mem[25][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][0]  ( .D(\fmem_inst/mem[25][0] ), .CK(clk), .Q(\fmem_data[25][0] ), .QN(n3483) );
  DFF_X1 \fmem_inst/mem_reg[25][1]  ( .D(n2906), .CK(clk), .Q(
        \fmem_inst/mem[25][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][1]  ( .D(\fmem_inst/mem[25][1] ), .CK(clk), .Q(\fmem_data[25][1] ), .QN(n3679) );
  DFF_X1 \fmem_inst/mem_reg[25][2]  ( .D(n2905), .CK(clk), .Q(
        \fmem_inst/mem[25][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][2]  ( .D(\fmem_inst/mem[25][2] ), .CK(clk), .Q(\fmem_data[25][2] ) );
  DFF_X1 \fmem_inst/mem_reg[25][3]  ( .D(n2904), .CK(clk), .Q(
        \fmem_inst/mem[25][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][3]  ( .D(\fmem_inst/mem[25][3] ), .CK(clk), .Q(\fmem_data[25][3] ), .QN(n3634) );
  DFF_X1 \fmem_inst/mem_reg[25][4]  ( .D(n2903), .CK(clk), .Q(
        \fmem_inst/mem[25][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][4]  ( .D(\fmem_inst/mem[25][4] ), .CK(clk), .Q(\fmem_data[25][4] ) );
  DFF_X1 \fmem_inst/mem_reg[25][5]  ( .D(n2902), .CK(clk), .Q(
        \fmem_inst/mem[25][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][5]  ( .D(\fmem_inst/mem[25][5] ), .CK(clk), .Q(\fmem_data[25][5] ), .QN(n3644) );
  DFF_X1 \fmem_inst/mem_reg[25][6]  ( .D(n2901), .CK(clk), .Q(
        \fmem_inst/mem[25][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][6]  ( .D(\fmem_inst/mem[25][6] ), .CK(clk), .Q(\fmem_data[25][6] ) );
  DFF_X1 \fmem_inst/mem_reg[25][7]  ( .D(n2900), .CK(clk), .Q(
        \fmem_inst/mem[25][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[25][7]  ( .D(\fmem_inst/mem[25][7] ), .CK(clk), .Q(\fmem_data[25][7] ), .QN(n3622) );
  DFF_X1 \fmem_inst/mem_reg[26][0]  ( .D(n2899), .CK(clk), .Q(
        \fmem_inst/mem[26][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][0]  ( .D(\fmem_inst/mem[26][0] ), .CK(clk), .Q(\fmem_data[26][0] ), .QN(n3678) );
  DFF_X1 \fmem_inst/mem_reg[26][1]  ( .D(n2898), .CK(clk), .Q(
        \fmem_inst/mem[26][1] ) );
  DFF_X1 \fmem_inst/mem_reg[26][2]  ( .D(n2897), .CK(clk), .Q(
        \fmem_inst/mem[26][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][2]  ( .D(\fmem_inst/mem[26][2] ), .CK(clk), .Q(\fmem_data[26][2] ) );
  DFF_X1 \fmem_inst/mem_reg[26][3]  ( .D(n2896), .CK(clk), .Q(
        \fmem_inst/mem[26][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][3]  ( .D(\fmem_inst/mem[26][3] ), .CK(clk), .Q(\fmem_data[26][3] ), .QN(n3658) );
  DFF_X1 \fmem_inst/mem_reg[26][4]  ( .D(n2895), .CK(clk), .Q(
        \fmem_inst/mem[26][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][4]  ( .D(\fmem_inst/mem[26][4] ), .CK(clk), .Q(\fmem_data[26][4] ) );
  DFF_X1 \fmem_inst/mem_reg[26][5]  ( .D(n2894), .CK(clk), .Q(
        \fmem_inst/mem[26][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][5]  ( .D(\fmem_inst/mem[26][5] ), .CK(clk), .Q(\fmem_data[26][5] ), .QN(n3677) );
  DFF_X1 \fmem_inst/mem_reg[26][6]  ( .D(n2893), .CK(clk), .Q(
        \fmem_inst/mem[26][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][6]  ( .D(\fmem_inst/mem[26][6] ), .CK(clk), .Q(\fmem_data[26][6] ) );
  DFF_X1 \fmem_inst/mem_reg[26][7]  ( .D(n2892), .CK(clk), .Q(
        \fmem_inst/mem[26][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[26][7]  ( .D(\fmem_inst/mem[26][7] ), .CK(clk), .Q(\fmem_data[26][7] ), .QN(n3655) );
  DFF_X1 \fmem_inst/mem_reg[27][0]  ( .D(n2891), .CK(clk), .Q(
        \fmem_inst/mem[27][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][0]  ( .D(\fmem_inst/mem[27][0] ), .CK(clk), .Q(\fmem_data[27][0] ), .QN(n3482) );
  DFF_X1 \fmem_inst/mem_reg[27][1]  ( .D(n2890), .CK(clk), .Q(
        \fmem_inst/mem[27][1] ) );
  DFF_X1 \fmem_inst/mem_reg[27][2]  ( .D(n2889), .CK(clk), .Q(
        \fmem_inst/mem[27][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][2]  ( .D(\fmem_inst/mem[27][2] ), .CK(clk), .Q(\fmem_data[27][2] ) );
  DFF_X1 \fmem_inst/mem_reg[27][3]  ( .D(n2888), .CK(clk), .Q(
        \fmem_inst/mem[27][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][3]  ( .D(\fmem_inst/mem[27][3] ), .CK(clk), .Q(\fmem_data[27][3] ), .QN(n3643) );
  DFF_X1 \fmem_inst/mem_reg[27][4]  ( .D(n2887), .CK(clk), .Q(
        \fmem_inst/mem[27][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][4]  ( .D(\fmem_inst/mem[27][4] ), .CK(clk), .Q(\fmem_data[27][4] ) );
  DFF_X1 \fmem_inst/mem_reg[27][5]  ( .D(n2886), .CK(clk), .Q(
        \fmem_inst/mem[27][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][5]  ( .D(\fmem_inst/mem[27][5] ), .CK(clk), .Q(\fmem_data[27][5] ), .QN(n3636) );
  DFF_X1 \fmem_inst/mem_reg[27][6]  ( .D(n2885), .CK(clk), .Q(
        \fmem_inst/mem[27][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][6]  ( .D(\fmem_inst/mem[27][6] ), .CK(clk), .Q(\fmem_data[27][6] ) );
  DFF_X1 \fmem_inst/mem_reg[27][7]  ( .D(n2884), .CK(clk), .Q(
        \fmem_inst/mem[27][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[27][7]  ( .D(\fmem_inst/mem[27][7] ), .CK(clk), .Q(\fmem_data[27][7] ), .QN(n3698) );
  DFF_X1 \fmem_inst/mem_reg[28][0]  ( .D(n2883), .CK(clk), .Q(
        \fmem_inst/mem[28][0] ) );
  DFF_X1 \fmem_inst/mem_reg[28][1]  ( .D(n2882), .CK(clk), .Q(
        \fmem_inst/mem[28][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][1]  ( .D(\fmem_inst/mem[28][1] ), .CK(clk), .Q(\fmem_data[28][1] ), .QN(n3671) );
  DFF_X1 \fmem_inst/mem_reg[28][2]  ( .D(n2881), .CK(clk), .Q(
        \fmem_inst/mem[28][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][2]  ( .D(\fmem_inst/mem[28][2] ), .CK(clk), .Q(\fmem_data[28][2] ) );
  DFF_X1 \fmem_inst/mem_reg[28][3]  ( .D(n2880), .CK(clk), .Q(
        \fmem_inst/mem[28][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][3]  ( .D(\fmem_inst/mem[28][3] ), .CK(clk), .Q(\fmem_data[28][3] ), .QN(n3604) );
  DFF_X1 \fmem_inst/mem_reg[28][4]  ( .D(n2879), .CK(clk), .Q(
        \fmem_inst/mem[28][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][4]  ( .D(\fmem_inst/mem[28][4] ), .CK(clk), .Q(\fmem_data[28][4] ) );
  DFF_X1 \fmem_inst/mem_reg[28][5]  ( .D(n2878), .CK(clk), .Q(
        \fmem_inst/mem[28][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][5]  ( .D(\fmem_inst/mem[28][5] ), .CK(clk), .Q(\fmem_data[28][5] ), .QN(n3650) );
  DFF_X1 \fmem_inst/mem_reg[28][6]  ( .D(n2877), .CK(clk), .Q(
        \fmem_inst/mem[28][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][6]  ( .D(\fmem_inst/mem[28][6] ), .CK(clk), .Q(\fmem_data[28][6] ) );
  DFF_X1 \fmem_inst/mem_reg[28][7]  ( .D(n2876), .CK(clk), .Q(
        \fmem_inst/mem[28][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[28][7]  ( .D(\fmem_inst/mem[28][7] ), .CK(clk), .Q(\fmem_data[28][7] ), .QN(n3659) );
  DFF_X1 \fmem_inst/mem_reg[29][0]  ( .D(n2875), .CK(clk), .Q(
        \fmem_inst/mem[29][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][0]  ( .D(\fmem_inst/mem[29][0] ), .CK(clk), .Q(\fmem_data[29][0] ), .QN(n3575) );
  DFF_X1 \fmem_inst/mem_reg[29][1]  ( .D(n2874), .CK(clk), .Q(
        \fmem_inst/mem[29][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][1]  ( .D(\fmem_inst/mem[29][1] ), .CK(clk), .Q(\fmem_data[29][1] ), .QN(n3660) );
  DFF_X1 \fmem_inst/mem_reg[29][2]  ( .D(n2873), .CK(clk), .Q(
        \fmem_inst/mem[29][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][2]  ( .D(\fmem_inst/mem[29][2] ), .CK(clk), .Q(\fmem_data[29][2] ) );
  DFF_X1 \fmem_inst/mem_reg[29][3]  ( .D(n2872), .CK(clk), .Q(
        \fmem_inst/mem[29][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][3]  ( .D(\fmem_inst/mem[29][3] ), .CK(clk), .Q(\fmem_data[29][3] ), .QN(n3587) );
  DFF_X1 \fmem_inst/mem_reg[29][4]  ( .D(n2871), .CK(clk), .Q(
        \fmem_inst/mem[29][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][4]  ( .D(\fmem_inst/mem[29][4] ), .CK(clk), .Q(\fmem_data[29][4] ) );
  DFF_X1 \fmem_inst/mem_reg[29][5]  ( .D(n2870), .CK(clk), .Q(
        \fmem_inst/mem[29][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][5]  ( .D(\fmem_inst/mem[29][5] ), .CK(clk), .Q(\fmem_data[29][5] ), .QN(n3588) );
  DFF_X1 \fmem_inst/mem_reg[29][6]  ( .D(n2869), .CK(clk), .Q(
        \fmem_inst/mem[29][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][6]  ( .D(\fmem_inst/mem[29][6] ), .CK(clk), .Q(\fmem_data[29][6] ) );
  DFF_X1 \fmem_inst/mem_reg[29][7]  ( .D(n2868), .CK(clk), .Q(
        \fmem_inst/mem[29][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[29][7]  ( .D(\fmem_inst/mem[29][7] ), .CK(clk), .Q(\fmem_data[29][7] ), .QN(n3602) );
  DFF_X1 \fmem_inst/mem_reg[30][0]  ( .D(n2867), .CK(clk), .Q(
        \fmem_inst/mem[30][0] ) );
  DFF_X1 \fmem_inst/mem_reg[30][1]  ( .D(n2866), .CK(clk), .Q(
        \fmem_inst/mem[30][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][1]  ( .D(\fmem_inst/mem[30][1] ), .CK(clk), .Q(\fmem_data[30][1] ), .QN(n3672) );
  DFF_X1 \fmem_inst/mem_reg[30][2]  ( .D(n2865), .CK(clk), .Q(
        \fmem_inst/mem[30][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][2]  ( .D(\fmem_inst/mem[30][2] ), .CK(clk), .Q(\fmem_data[30][2] ) );
  DFF_X1 \fmem_inst/mem_reg[30][3]  ( .D(n2864), .CK(clk), .Q(
        \fmem_inst/mem[30][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][3]  ( .D(\fmem_inst/mem[30][3] ), .CK(clk), .Q(\fmem_data[30][3] ), .QN(n3592) );
  DFF_X1 \fmem_inst/mem_reg[30][4]  ( .D(n2863), .CK(clk), .Q(
        \fmem_inst/mem[30][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][4]  ( .D(\fmem_inst/mem[30][4] ), .CK(clk), .Q(\fmem_data[30][4] ) );
  DFF_X1 \fmem_inst/mem_reg[30][5]  ( .D(n2862), .CK(clk), .Q(
        \fmem_inst/mem[30][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][5]  ( .D(\fmem_inst/mem[30][5] ), .CK(clk), .Q(\fmem_data[30][5] ), .QN(n3597) );
  DFF_X1 \fmem_inst/mem_reg[30][6]  ( .D(n2861), .CK(clk), .Q(
        \fmem_inst/mem[30][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][6]  ( .D(\fmem_inst/mem[30][6] ), .CK(clk), .Q(\fmem_data[30][6] ) );
  DFF_X1 \fmem_inst/mem_reg[30][7]  ( .D(n2860), .CK(clk), .Q(
        \fmem_inst/mem[30][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[30][7]  ( .D(\fmem_inst/mem[30][7] ), .CK(clk), .Q(\fmem_data[30][7] ), .QN(n3585) );
  DFF_X1 \ctrl_fmem_write_inst/s_ready_reg  ( .D(n3113), .CK(clk), .Q(
        s_ready_f), .QN(n39001) );
  DFF_X1 \fmem_inst/mem_reg[0][0]  ( .D(n3107), .CK(clk), .Q(
        \fmem_inst/mem[0][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][0]  ( .D(\fmem_inst/mem[0][0] ), .CK(clk), 
        .Q(\fmem_data[0][0] ), .QN(n3564) );
  DFF_X1 \fmem_inst/mem_reg[0][1]  ( .D(n3106), .CK(clk), .Q(
        \fmem_inst/mem[0][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][1]  ( .D(\fmem_inst/mem[0][1] ), .CK(clk), 
        .Q(\fmem_data[0][1] ), .QN(n4020) );
  DFF_X1 \fmem_inst/mem_reg[0][2]  ( .D(n3105), .CK(clk), .Q(
        \fmem_inst/mem[0][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][2]  ( .D(\fmem_inst/mem[0][2] ), .CK(clk), 
        .Q(\fmem_data[0][2] ) );
  DFF_X1 \fmem_inst/mem_reg[0][3]  ( .D(n3104), .CK(clk), .Q(
        \fmem_inst/mem[0][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][3]  ( .D(\fmem_inst/mem[0][3] ), .CK(clk), 
        .Q(\fmem_data[0][3] ), .QN(n3667) );
  DFF_X1 \fmem_inst/mem_reg[0][4]  ( .D(n3103), .CK(clk), .Q(
        \fmem_inst/mem[0][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][4]  ( .D(\fmem_inst/mem[0][4] ), .CK(clk), 
        .Q(\fmem_data[0][4] ) );
  DFF_X1 \fmem_inst/mem_reg[0][5]  ( .D(n3102), .CK(clk), .Q(
        \fmem_inst/mem[0][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][5]  ( .D(\fmem_inst/mem[0][5] ), .CK(clk), 
        .Q(\fmem_data[0][5] ), .QN(n3629) );
  DFF_X1 \fmem_inst/mem_reg[0][6]  ( .D(n3101), .CK(clk), .Q(
        \fmem_inst/mem[0][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][6]  ( .D(\fmem_inst/mem[0][6] ), .CK(clk), 
        .Q(\fmem_data[0][6] ) );
  DFF_X1 \fmem_inst/mem_reg[0][7]  ( .D(n3100), .CK(clk), .Q(
        \fmem_inst/mem[0][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[0][7]  ( .D(\fmem_inst/mem[0][7] ), .CK(clk), 
        .Q(\fmem_data[0][7] ), .QN(n3637) );
  DFF_X1 \fmem_inst/mem_reg[1][0]  ( .D(n3099), .CK(clk), .Q(
        \fmem_inst/mem[1][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][0]  ( .D(\fmem_inst/mem[1][0] ), .CK(clk), 
        .Q(\fmem_data[1][0] ), .QN(n3558) );
  DFF_X1 \fmem_inst/mem_reg[1][1]  ( .D(n3098), .CK(clk), .Q(
        \fmem_inst/mem[1][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][1]  ( .D(\fmem_inst/mem[1][1] ), .CK(clk), 
        .Q(\fmem_data[1][1] ), .QN(n3661) );
  DFF_X1 \fmem_inst/mem_reg[1][2]  ( .D(n3097), .CK(clk), .Q(
        \fmem_inst/mem[1][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][2]  ( .D(\fmem_inst/mem[1][2] ), .CK(clk), 
        .Q(\fmem_data[1][2] ) );
  DFF_X1 \fmem_inst/mem_reg[1][3]  ( .D(n3096), .CK(clk), .Q(
        \fmem_inst/mem[1][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][3]  ( .D(\fmem_inst/mem[1][3] ), .CK(clk), 
        .Q(\fmem_data[1][3] ), .QN(n3590) );
  DFF_X1 \fmem_inst/mem_reg[1][4]  ( .D(n3095), .CK(clk), .Q(
        \fmem_inst/mem[1][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][4]  ( .D(\fmem_inst/mem[1][4] ), .CK(clk), 
        .Q(\fmem_data[1][4] ) );
  DFF_X1 \fmem_inst/mem_reg[1][5]  ( .D(n3094), .CK(clk), .Q(
        \fmem_inst/mem[1][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][5]  ( .D(\fmem_inst/mem[1][5] ), .CK(clk), 
        .Q(\fmem_data[1][5] ), .QN(n3583) );
  DFF_X1 \fmem_inst/mem_reg[1][6]  ( .D(n3093), .CK(clk), .Q(
        \fmem_inst/mem[1][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][6]  ( .D(\fmem_inst/mem[1][6] ), .CK(clk), 
        .Q(\fmem_data[1][6] ) );
  DFF_X1 \fmem_inst/mem_reg[1][7]  ( .D(n3092), .CK(clk), .Q(
        \fmem_inst/mem[1][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[1][7]  ( .D(\fmem_inst/mem[1][7] ), .CK(clk), 
        .Q(\fmem_data[1][7] ), .QN(n3601) );
  DFF_X1 \fmem_inst/mem_reg[2][0]  ( .D(n3091), .CK(clk), .Q(
        \fmem_inst/mem[2][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][0]  ( .D(\fmem_inst/mem[2][0] ), .CK(clk), 
        .Q(\fmem_data[2][0] ), .QN(n3578) );
  DFF_X1 \fmem_inst/mem_reg[2][1]  ( .D(n3090), .CK(clk), .Q(
        \fmem_inst/mem[2][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][1]  ( .D(\fmem_inst/mem[2][1] ), .CK(clk), 
        .Q(\fmem_data[2][1] ), .QN(n3691) );
  DFF_X1 \fmem_inst/mem_reg[2][2]  ( .D(n3089), .CK(clk), .Q(
        \fmem_inst/mem[2][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][2]  ( .D(\fmem_inst/mem[2][2] ), .CK(clk), 
        .Q(\fmem_data[2][2] ) );
  DFF_X1 \fmem_inst/mem_reg[2][3]  ( .D(n3088), .CK(clk), .Q(
        \fmem_inst/mem[2][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][3]  ( .D(\fmem_inst/mem[2][3] ), .CK(clk), 
        .Q(\fmem_data[2][3] ), .QN(n3652) );
  DFF_X1 \fmem_inst/mem_reg[2][4]  ( .D(n3087), .CK(clk), .Q(
        \fmem_inst/mem[2][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][4]  ( .D(\fmem_inst/mem[2][4] ), .CK(clk), 
        .Q(\fmem_data[2][4] ) );
  DFF_X1 \fmem_inst/mem_reg[2][5]  ( .D(n3086), .CK(clk), .Q(
        \fmem_inst/mem[2][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][5]  ( .D(\fmem_inst/mem[2][5] ), .CK(clk), 
        .Q(\fmem_data[2][5] ), .QN(n3620) );
  DFF_X1 \fmem_inst/mem_reg[2][6]  ( .D(n3085), .CK(clk), .Q(
        \fmem_inst/mem[2][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][6]  ( .D(\fmem_inst/mem[2][6] ), .CK(clk), 
        .Q(\fmem_data[2][6] ) );
  DFF_X1 \fmem_inst/mem_reg[2][7]  ( .D(n3084), .CK(clk), .Q(
        \fmem_inst/mem[2][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[2][7]  ( .D(\fmem_inst/mem[2][7] ), .CK(clk), 
        .Q(\fmem_data[2][7] ), .QN(n3624) );
  DFF_X1 \fmem_inst/mem_reg[3][0]  ( .D(n3083), .CK(clk), .Q(
        \fmem_inst/mem[3][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][0]  ( .D(\fmem_inst/mem[3][0] ), .CK(clk), 
        .Q(\fmem_data[3][0] ), .QN(n3582) );
  DFF_X1 \fmem_inst/mem_reg[3][1]  ( .D(n3082), .CK(clk), .Q(
        \fmem_inst/mem[3][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][1]  ( .D(\fmem_inst/mem[3][1] ), .CK(clk), 
        .Q(\fmem_data[3][1] ), .QN(n3695) );
  DFF_X1 \fmem_inst/mem_reg[3][2]  ( .D(n3081), .CK(clk), .Q(
        \fmem_inst/mem[3][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][2]  ( .D(\fmem_inst/mem[3][2] ), .CK(clk), 
        .Q(\fmem_data[3][2] ) );
  DFF_X1 \fmem_inst/mem_reg[3][3]  ( .D(n3080), .CK(clk), .Q(
        \fmem_inst/mem[3][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][3]  ( .D(\fmem_inst/mem[3][3] ), .CK(clk), 
        .Q(\fmem_data[3][3] ), .QN(n3642) );
  DFF_X1 \fmem_inst/mem_reg[3][4]  ( .D(n3079), .CK(clk), .Q(
        \fmem_inst/mem[3][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][4]  ( .D(\fmem_inst/mem[3][4] ), .CK(clk), 
        .Q(\fmem_data[3][4] ) );
  DFF_X1 \fmem_inst/mem_reg[3][5]  ( .D(n3078), .CK(clk), .Q(
        \fmem_inst/mem[3][5] ) );
  DFF_X1 \fmem_inst/mem_reg[3][6]  ( .D(n3077), .CK(clk), .Q(
        \fmem_inst/mem[3][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][6]  ( .D(\fmem_inst/mem[3][6] ), .CK(clk), 
        .Q(\fmem_data[3][6] ) );
  DFF_X1 \fmem_inst/mem_reg[3][7]  ( .D(n3076), .CK(clk), .Q(
        \fmem_inst/mem[3][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[3][7]  ( .D(\fmem_inst/mem[3][7] ), .CK(clk), 
        .Q(\fmem_data[3][7] ), .QN(n3656) );
  DFF_X1 \fmem_inst/mem_reg[4][0]  ( .D(n3075), .CK(clk), .Q(
        \fmem_inst/mem[4][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][0]  ( .D(\fmem_inst/mem[4][0] ), .CK(clk), 
        .Q(\fmem_data[4][0] ), .QN(n3569) );
  DFF_X1 \fmem_inst/mem_reg[4][1]  ( .D(n3074), .CK(clk), .Q(
        \fmem_inst/mem[4][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][1]  ( .D(\fmem_inst/mem[4][1] ), .CK(clk), 
        .Q(\fmem_data[4][1] ) );
  DFF_X1 \fmem_inst/mem_reg[4][2]  ( .D(n3073), .CK(clk), .Q(
        \fmem_inst/mem[4][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][2]  ( .D(\fmem_inst/mem[4][2] ), .CK(clk), 
        .Q(\fmem_data[4][2] ) );
  DFF_X1 \fmem_inst/mem_reg[4][3]  ( .D(n3072), .CK(clk), .Q(
        \fmem_inst/mem[4][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][3]  ( .D(\fmem_inst/mem[4][3] ), .CK(clk), 
        .Q(\fmem_data[4][3] ), .QN(n3610) );
  DFF_X1 \fmem_inst/mem_reg[4][4]  ( .D(n3071), .CK(clk), .Q(
        \fmem_inst/mem[4][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][4]  ( .D(\fmem_inst/mem[4][4] ), .CK(clk), 
        .Q(\fmem_data[4][4] ) );
  DFF_X1 \fmem_inst/mem_reg[4][5]  ( .D(n3070), .CK(clk), .Q(
        \fmem_inst/mem[4][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][5]  ( .D(\fmem_inst/mem[4][5] ), .CK(clk), 
        .Q(\fmem_data[4][5] ), .QN(n3632) );
  DFF_X1 \fmem_inst/mem_reg[4][6]  ( .D(n3069), .CK(clk), .Q(
        \fmem_inst/mem[4][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][6]  ( .D(\fmem_inst/mem[4][6] ), .CK(clk), 
        .Q(\fmem_data[4][6] ) );
  DFF_X1 \fmem_inst/mem_reg[4][7]  ( .D(n3068), .CK(clk), .Q(
        \fmem_inst/mem[4][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[4][7]  ( .D(\fmem_inst/mem[4][7] ), .CK(clk), 
        .Q(\fmem_data[4][7] ), .QN(n3614) );
  DFF_X1 \fmem_inst/mem_reg[5][0]  ( .D(n3067), .CK(clk), .Q(
        \fmem_inst/mem[5][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][0]  ( .D(\fmem_inst/mem[5][0] ), .CK(clk), 
        .Q(\fmem_data[5][0] ), .QN(n3576) );
  DFF_X1 \fmem_inst/mem_reg[5][1]  ( .D(n3066), .CK(clk), .Q(
        \fmem_inst/mem[5][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][1]  ( .D(\fmem_inst/mem[5][1] ), .CK(clk), 
        .Q(\fmem_data[5][1] ), .QN(n3694) );
  DFF_X1 \fmem_inst/mem_reg[5][2]  ( .D(n3065), .CK(clk), .Q(
        \fmem_inst/mem[5][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][2]  ( .D(\fmem_inst/mem[5][2] ), .CK(clk), 
        .Q(\fmem_data[5][2] ) );
  DFF_X1 \fmem_inst/mem_reg[5][3]  ( .D(n3064), .CK(clk), .Q(
        \fmem_inst/mem[5][3] ) );
  DFF_X1 \fmem_inst/mem_reg[5][4]  ( .D(n3063), .CK(clk), .Q(
        \fmem_inst/mem[5][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][4]  ( .D(\fmem_inst/mem[5][4] ), .CK(clk), 
        .Q(\fmem_data[5][4] ) );
  DFF_X1 \fmem_inst/mem_reg[5][5]  ( .D(n3062), .CK(clk), .Q(
        \fmem_inst/mem[5][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][5]  ( .D(\fmem_inst/mem[5][5] ), .CK(clk), 
        .Q(\fmem_data[5][5] ), .QN(n3635) );
  DFF_X1 \fmem_inst/mem_reg[5][6]  ( .D(n3061), .CK(clk), .Q(
        \fmem_inst/mem[5][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][6]  ( .D(\fmem_inst/mem[5][6] ), .CK(clk), 
        .Q(\fmem_data[5][6] ) );
  DFF_X1 \fmem_inst/mem_reg[5][7]  ( .D(n3060), .CK(clk), .Q(
        \fmem_inst/mem[5][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[5][7]  ( .D(\fmem_inst/mem[5][7] ), .CK(clk), 
        .Q(\fmem_data[5][7] ), .QN(n3623) );
  DFF_X1 \fmem_inst/mem_reg[6][0]  ( .D(n3059), .CK(clk), .Q(
        \fmem_inst/mem[6][0] ) );
  DFF_X1 \fmem_inst/mem_reg[6][1]  ( .D(n3058), .CK(clk), .Q(
        \fmem_inst/mem[6][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][1]  ( .D(\fmem_inst/mem[6][1] ), .CK(clk), 
        .Q(\fmem_data[6][1] ), .QN(n3682) );
  DFF_X1 \fmem_inst/mem_reg[6][2]  ( .D(n3057), .CK(clk), .Q(
        \fmem_inst/mem[6][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][2]  ( .D(\fmem_inst/mem[6][2] ), .CK(clk), 
        .Q(\fmem_data[6][2] ) );
  DFF_X1 \fmem_inst/mem_reg[6][3]  ( .D(n3056), .CK(clk), .Q(
        \fmem_inst/mem[6][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][3]  ( .D(\fmem_inst/mem[6][3] ), .CK(clk), 
        .Q(\fmem_data[6][3] ), .QN(n3646) );
  DFF_X1 \fmem_inst/mem_reg[6][4]  ( .D(n3055), .CK(clk), .Q(
        \fmem_inst/mem[6][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][4]  ( .D(\fmem_inst/mem[6][4] ), .CK(clk), 
        .Q(\fmem_data[6][4] ) );
  DFF_X1 \fmem_inst/mem_reg[6][5]  ( .D(n3054), .CK(clk), .Q(
        \fmem_inst/mem[6][5] ) );
  DFF_X1 \fmem_inst/mem_reg[6][6]  ( .D(n3053), .CK(clk), .Q(
        \fmem_inst/mem[6][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][6]  ( .D(\fmem_inst/mem[6][6] ), .CK(clk), 
        .Q(\fmem_data[6][6] ) );
  DFF_X1 \fmem_inst/mem_reg[6][7]  ( .D(n3052), .CK(clk), .Q(
        \fmem_inst/mem[6][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[6][7]  ( .D(\fmem_inst/mem[6][7] ), .CK(clk), 
        .Q(\fmem_data[6][7] ), .QN(n3630) );
  DFF_X1 \fmem_inst/mem_reg[7][0]  ( .D(n3051), .CK(clk), .Q(
        \fmem_inst/mem[7][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][0]  ( .D(\fmem_inst/mem[7][0] ), .CK(clk), 
        .Q(\fmem_data[7][0] ), .QN(n3581) );
  DFF_X1 \fmem_inst/mem_reg[7][1]  ( .D(n3050), .CK(clk), .Q(
        \fmem_inst/mem[7][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][1]  ( .D(\fmem_inst/mem[7][1] ), .CK(clk), 
        .Q(\fmem_data[7][1] ), .QN(n3945) );
  DFF_X1 \fmem_inst/mem_reg[7][2]  ( .D(n3049), .CK(clk), .Q(
        \fmem_inst/mem[7][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][2]  ( .D(\fmem_inst/mem[7][2] ), .CK(clk), 
        .Q(\fmem_data[7][2] ) );
  DFF_X1 \fmem_inst/mem_reg[7][3]  ( .D(n3048), .CK(clk), .Q(
        \fmem_inst/mem[7][3] ) );
  DFF_X1 \fmem_inst/mem_reg[7][4]  ( .D(n3047), .CK(clk), .Q(
        \fmem_inst/mem[7][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][4]  ( .D(\fmem_inst/mem[7][4] ), .CK(clk), 
        .Q(\fmem_data[7][4] ) );
  DFF_X1 \fmem_inst/mem_reg[7][5]  ( .D(n3046), .CK(clk), .Q(
        \fmem_inst/mem[7][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][5]  ( .D(\fmem_inst/mem[7][5] ), .CK(clk), 
        .Q(\fmem_data[7][5] ), .QN(n3648) );
  DFF_X1 \fmem_inst/mem_reg[7][6]  ( .D(n3045), .CK(clk), .Q(
        \fmem_inst/mem[7][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][6]  ( .D(\fmem_inst/mem[7][6] ), .CK(clk), 
        .Q(\fmem_data[7][6] ) );
  DFF_X1 \fmem_inst/mem_reg[7][7]  ( .D(n3044), .CK(clk), .Q(
        \fmem_inst/mem[7][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[7][7]  ( .D(\fmem_inst/mem[7][7] ), .CK(clk), 
        .Q(\fmem_data[7][7] ), .QN(n3490) );
  DFF_X1 \fmem_inst/mem_reg[8][0]  ( .D(n3043), .CK(clk), .Q(
        \fmem_inst/mem[8][0] ) );
  DFF_X1 \fmem_inst/mem_reg[8][1]  ( .D(n3042), .CK(clk), .Q(
        \fmem_inst/mem[8][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][1]  ( .D(\fmem_inst/mem[8][1] ), .CK(clk), 
        .Q(\fmem_data[8][1] ), .QN(n3666) );
  DFF_X1 \fmem_inst/mem_reg[8][2]  ( .D(n3041), .CK(clk), .Q(
        \fmem_inst/mem[8][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][2]  ( .D(\fmem_inst/mem[8][2] ), .CK(clk), 
        .Q(\fmem_data[8][2] ) );
  DFF_X1 \fmem_inst/mem_reg[8][3]  ( .D(n3040), .CK(clk), .Q(
        \fmem_inst/mem[8][3] ) );
  DFF_X1 \fmem_inst/mem_reg[8][4]  ( .D(n3039), .CK(clk), .Q(
        \fmem_inst/mem[8][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][4]  ( .D(\fmem_inst/mem[8][4] ), .CK(clk), 
        .Q(\fmem_data[8][4] ) );
  DFF_X1 \fmem_inst/mem_reg[8][5]  ( .D(n3038), .CK(clk), .Q(
        \fmem_inst/mem[8][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][5]  ( .D(\fmem_inst/mem[8][5] ), .CK(clk), 
        .Q(\fmem_data[8][5] ), .QN(n3594) );
  DFF_X1 \fmem_inst/mem_reg[8][6]  ( .D(n3037), .CK(clk), .Q(
        \fmem_inst/mem[8][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][6]  ( .D(\fmem_inst/mem[8][6] ), .CK(clk), 
        .Q(\fmem_data[8][6] ) );
  DFF_X1 \fmem_inst/mem_reg[8][7]  ( .D(n3036), .CK(clk), .Q(
        \fmem_inst/mem[8][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[8][7]  ( .D(\fmem_inst/mem[8][7] ), .CK(clk), 
        .Q(\fmem_data[8][7] ), .QN(n3638) );
  DFF_X1 \fmem_inst/mem_reg[9][0]  ( .D(n3035), .CK(clk), .Q(
        \fmem_inst/mem[9][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][0]  ( .D(\fmem_inst/mem[9][0] ), .CK(clk), 
        .Q(\fmem_data[9][0] ), .QN(n3579) );
  DFF_X1 \fmem_inst/mem_reg[9][1]  ( .D(n3034), .CK(clk), .Q(
        \fmem_inst/mem[9][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][1]  ( .D(\fmem_inst/mem[9][1] ), .CK(clk), 
        .Q(\fmem_data[9][1] ), .QN(n3689) );
  DFF_X1 \fmem_inst/mem_reg[9][2]  ( .D(n3033), .CK(clk), .Q(
        \fmem_inst/mem[9][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][2]  ( .D(\fmem_inst/mem[9][2] ), .CK(clk), 
        .Q(\fmem_data[9][2] ) );
  DFF_X1 \fmem_inst/mem_reg[9][3]  ( .D(n3032), .CK(clk), .Q(
        \fmem_inst/mem[9][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][3]  ( .D(\fmem_inst/mem[9][3] ), .CK(clk), 
        .Q(\fmem_data[9][3] ), .QN(n3607) );
  DFF_X1 \fmem_inst/mem_reg[9][4]  ( .D(n3031), .CK(clk), .Q(
        \fmem_inst/mem[9][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][4]  ( .D(\fmem_inst/mem[9][4] ), .CK(clk), 
        .Q(\fmem_data[9][4] ) );
  DFF_X1 \fmem_inst/mem_reg[9][5]  ( .D(n3030), .CK(clk), .Q(
        \fmem_inst/mem[9][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][5]  ( .D(\fmem_inst/mem[9][5] ), .CK(clk), 
        .Q(\fmem_data[9][5] ), .QN(n3608) );
  DFF_X1 \fmem_inst/mem_reg[9][6]  ( .D(n3029), .CK(clk), .Q(
        \fmem_inst/mem[9][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][6]  ( .D(\fmem_inst/mem[9][6] ), .CK(clk), 
        .Q(\fmem_data[9][6] ) );
  DFF_X1 \fmem_inst/mem_reg[9][7]  ( .D(n3028), .CK(clk), .Q(
        \fmem_inst/mem[9][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[9][7]  ( .D(\fmem_inst/mem[9][7] ), .CK(clk), 
        .Q(\fmem_data[9][7] ), .QN(n3625) );
  DFF_X1 \fmem_inst/mem_reg[10][0]  ( .D(n3027), .CK(clk), .Q(
        \fmem_inst/mem[10][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][0]  ( .D(\fmem_inst/mem[10][0] ), .CK(clk), .Q(\fmem_data[10][0] ), .QN(n3561) );
  DFF_X1 \fmem_inst/mem_reg[10][1]  ( .D(n3026), .CK(clk), .Q(
        \fmem_inst/mem[10][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][1]  ( .D(\fmem_inst/mem[10][1] ), .CK(clk), .Q(\fmem_data[10][1] ), .QN(n3681) );
  DFF_X1 \fmem_inst/mem_reg[10][2]  ( .D(n3025), .CK(clk), .Q(
        \fmem_inst/mem[10][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][2]  ( .D(\fmem_inst/mem[10][2] ), .CK(clk), .Q(\fmem_data[10][2] ) );
  DFF_X1 \fmem_inst/mem_reg[10][3]  ( .D(n3024), .CK(clk), .Q(
        \fmem_inst/mem[10][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][3]  ( .D(\fmem_inst/mem[10][3] ), .CK(clk), .Q(\fmem_data[10][3] ), .QN(n3611) );
  DFF_X1 \fmem_inst/mem_reg[10][4]  ( .D(n3023), .CK(clk), .Q(
        \fmem_inst/mem[10][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][4]  ( .D(\fmem_inst/mem[10][4] ), .CK(clk), .Q(\fmem_data[10][4] ) );
  DFF_X1 \fmem_inst/mem_reg[10][5]  ( .D(n3022), .CK(clk), .Q(
        \fmem_inst/mem[10][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][5]  ( .D(\fmem_inst/mem[10][5] ), .CK(clk), .Q(\fmem_data[10][5] ), .QN(n3595) );
  DFF_X1 \fmem_inst/mem_reg[10][6]  ( .D(n3021), .CK(clk), .Q(
        \fmem_inst/mem[10][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][6]  ( .D(\fmem_inst/mem[10][6] ), .CK(clk), .Q(\fmem_data[10][6] ) );
  DFF_X1 \fmem_inst/mem_reg[10][7]  ( .D(n3020), .CK(clk), .Q(
        \fmem_inst/mem[10][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[10][7]  ( .D(\fmem_inst/mem[10][7] ), .CK(clk), .Q(\fmem_data[10][7] ), .QN(n3631) );
  DFF_X1 \fmem_inst/mem_reg[11][0]  ( .D(n3019), .CK(clk), .Q(
        \fmem_inst/mem[11][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][0]  ( .D(\fmem_inst/mem[11][0] ), .CK(clk), .Q(\fmem_data[11][0] ), .QN(n3577) );
  DFF_X1 \fmem_inst/mem_reg[11][1]  ( .D(n3018), .CK(clk), .Q(
        \fmem_inst/mem[11][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][1]  ( .D(\fmem_inst/mem[11][1] ), .CK(clk), .Q(\fmem_data[11][1] ), .QN(n3699) );
  DFF_X1 \fmem_inst/mem_reg[11][2]  ( .D(n3017), .CK(clk), .Q(
        \fmem_inst/mem[11][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][2]  ( .D(\fmem_inst/mem[11][2] ), .CK(clk), .Q(\fmem_data[11][2] ) );
  DFF_X1 \fmem_inst/mem_reg[11][3]  ( .D(n3016), .CK(clk), .Q(
        \fmem_inst/mem[11][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][3]  ( .D(\fmem_inst/mem[11][3] ), .CK(clk), .Q(\fmem_data[11][3] ), .QN(n3657) );
  DFF_X1 \fmem_inst/mem_reg[11][4]  ( .D(n3015), .CK(clk), .Q(
        \fmem_inst/mem[11][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][4]  ( .D(\fmem_inst/mem[11][4] ), .CK(clk), .Q(\fmem_data[11][4] ) );
  DFF_X1 \fmem_inst/mem_reg[11][5]  ( .D(n3014), .CK(clk), .Q(
        \fmem_inst/mem[11][5] ) );
  DFF_X1 \fmem_inst/mem_reg[11][6]  ( .D(n3013), .CK(clk), .Q(
        \fmem_inst/mem[11][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][6]  ( .D(\fmem_inst/mem[11][6] ), .CK(clk), .Q(\fmem_data[11][6] ) );
  DFF_X1 \fmem_inst/mem_reg[11][7]  ( .D(n3012), .CK(clk), .Q(
        \fmem_inst/mem[11][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[11][7]  ( .D(\fmem_inst/mem[11][7] ), .CK(clk), .Q(\fmem_data[11][7] ), .QN(n3663) );
  DFF_X1 \fmem_inst/mem_reg[12][0]  ( .D(n3011), .CK(clk), .Q(
        \fmem_inst/mem[12][0] ) );
  DFF_X1 \fmem_inst/mem_reg[12][1]  ( .D(n3010), .CK(clk), .Q(
        \fmem_inst/mem[12][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][1]  ( .D(\fmem_inst/mem[12][1] ), .CK(clk), .Q(\fmem_data[12][1] ), .QN(n3673) );
  DFF_X1 \fmem_inst/mem_reg[12][2]  ( .D(n3009), .CK(clk), .Q(
        \fmem_inst/mem[12][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][2]  ( .D(\fmem_inst/mem[12][2] ), .CK(clk), .Q(\fmem_data[12][2] ) );
  DFF_X1 \fmem_inst/mem_reg[12][3]  ( .D(n3008), .CK(clk), .Q(
        \fmem_inst/mem[12][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][3]  ( .D(\fmem_inst/mem[12][3] ), .CK(clk), .Q(\fmem_data[12][3] ), .QN(n3616) );
  DFF_X1 \fmem_inst/mem_reg[12][4]  ( .D(n3007), .CK(clk), .Q(
        \fmem_inst/mem[12][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][4]  ( .D(\fmem_inst/mem[12][4] ), .CK(clk), .Q(\fmem_data[12][4] ) );
  DFF_X1 \fmem_inst/mem_reg[12][5]  ( .D(n3006), .CK(clk), .Q(
        \fmem_inst/mem[12][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][5]  ( .D(\fmem_inst/mem[12][5] ), .CK(clk), .Q(\fmem_data[12][5] ), .QN(n3589) );
  DFF_X1 \fmem_inst/mem_reg[12][6]  ( .D(n3005), .CK(clk), .Q(
        \fmem_inst/mem[12][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][6]  ( .D(\fmem_inst/mem[12][6] ), .CK(clk), .Q(\fmem_data[12][6] ) );
  DFF_X1 \fmem_inst/mem_reg[12][7]  ( .D(n3004), .CK(clk), .Q(
        \fmem_inst/mem[12][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[12][7]  ( .D(\fmem_inst/mem[12][7] ), .CK(clk), .Q(\fmem_data[12][7] ), .QN(n3615) );
  DFF_X1 \fmem_inst/mem_reg[13][0]  ( .D(n3003), .CK(clk), .Q(
        \fmem_inst/mem[13][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][0]  ( .D(\fmem_inst/mem[13][0] ), .CK(clk), .Q(\fmem_data[13][0] ), .QN(n3571) );
  DFF_X1 \fmem_inst/mem_reg[13][1]  ( .D(n3002), .CK(clk), .Q(
        \fmem_inst/mem[13][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][1]  ( .D(\fmem_inst/mem[13][1] ), .CK(clk), .Q(\fmem_data[13][1] ), .QN(n3683) );
  DFF_X1 \fmem_inst/mem_reg[13][2]  ( .D(n3001), .CK(clk), .Q(
        \fmem_inst/mem[13][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][2]  ( .D(\fmem_inst/mem[13][2] ), .CK(clk), .Q(\fmem_data[13][2] ) );
  DFF_X1 \fmem_inst/mem_reg[13][3]  ( .D(n3000), .CK(clk), .Q(
        \fmem_inst/mem[13][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][3]  ( .D(\fmem_inst/mem[13][3] ), .CK(clk), .Q(\fmem_data[13][3] ), .QN(n3641) );
  DFF_X1 \fmem_inst/mem_reg[13][4]  ( .D(n2999), .CK(clk), .Q(
        \fmem_inst/mem[13][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][4]  ( .D(\fmem_inst/mem[13][4] ), .CK(clk), .Q(\fmem_data[13][4] ) );
  DFF_X1 \fmem_inst/mem_reg[13][5]  ( .D(n2998), .CK(clk), .Q(
        \fmem_inst/mem[13][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][5]  ( .D(\fmem_inst/mem[13][5] ), .CK(clk), .Q(\fmem_data[13][5] ), .QN(n3612) );
  DFF_X1 \fmem_inst/mem_reg[13][6]  ( .D(n2997), .CK(clk), .Q(
        \fmem_inst/mem[13][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][6]  ( .D(\fmem_inst/mem[13][6] ), .CK(clk), .Q(\fmem_data[13][6] ) );
  DFF_X1 \fmem_inst/mem_reg[13][7]  ( .D(n2996), .CK(clk), .Q(
        \fmem_inst/mem[13][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[13][7]  ( .D(\fmem_inst/mem[13][7] ), .CK(clk), .Q(\fmem_data[13][7] ), .QN(n3613) );
  DFF_X1 \fmem_inst/mem_reg[14][0]  ( .D(n2995), .CK(clk), .Q(
        \fmem_inst/mem[14][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][0]  ( .D(\fmem_inst/mem[14][0] ), .CK(clk), .Q(\fmem_data[14][0] ), .QN(n3563) );
  DFF_X1 \fmem_inst/mem_reg[14][1]  ( .D(n2994), .CK(clk), .Q(
        \fmem_inst/mem[14][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][1]  ( .D(\fmem_inst/mem[14][1] ), .CK(clk), .Q(\fmem_data[14][1] ), .QN(n3675) );
  DFF_X1 \fmem_inst/mem_reg[14][2]  ( .D(n2993), .CK(clk), .Q(
        \fmem_inst/mem[14][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][2]  ( .D(\fmem_inst/mem[14][2] ), .CK(clk), .Q(\fmem_data[14][2] ) );
  DFF_X1 \fmem_inst/mem_reg[14][3]  ( .D(n2992), .CK(clk), .Q(
        \fmem_inst/mem[14][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][3]  ( .D(\fmem_inst/mem[14][3] ), .CK(clk), .Q(\fmem_data[14][3] ), .QN(n3617) );
  DFF_X1 \fmem_inst/mem_reg[14][4]  ( .D(n2991), .CK(clk), .Q(
        \fmem_inst/mem[14][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][4]  ( .D(\fmem_inst/mem[14][4] ), .CK(clk), .Q(\fmem_data[14][4] ) );
  DFF_X1 \fmem_inst/mem_reg[14][5]  ( .D(n2990), .CK(clk), .Q(
        \fmem_inst/mem[14][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][5]  ( .D(\fmem_inst/mem[14][5] ), .CK(clk), .Q(\fmem_data[14][5] ), .QN(n3584) );
  DFF_X1 \fmem_inst/mem_reg[14][6]  ( .D(n2989), .CK(clk), .Q(
        \fmem_inst/mem[14][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][6]  ( .D(\fmem_inst/mem[14][6] ), .CK(clk), .Q(\fmem_data[14][6] ) );
  DFF_X1 \fmem_inst/mem_reg[14][7]  ( .D(n2988), .CK(clk), .Q(
        \fmem_inst/mem[14][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[14][7]  ( .D(\fmem_inst/mem[14][7] ), .CK(clk), .Q(\fmem_data[14][7] ), .QN(n3598) );
  DFF_X1 \fmem_inst/mem_reg[15][0]  ( .D(n2987), .CK(clk), .Q(
        \fmem_inst/mem[15][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][0]  ( .D(\fmem_inst/mem[15][0] ), .CK(clk), .Q(\fmem_data[15][0] ), .QN(n3568) );
  DFF_X1 \fmem_inst/mem_reg[15][1]  ( .D(n2986), .CK(clk), .Q(
        \fmem_inst/mem[15][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][1]  ( .D(\fmem_inst/mem[15][1] ), .CK(clk), .Q(\fmem_data[15][1] ), .QN(n3692) );
  DFF_X1 \fmem_inst/mem_reg[15][2]  ( .D(n2985), .CK(clk), .Q(
        \fmem_inst/mem[15][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][2]  ( .D(\fmem_inst/mem[15][2] ), .CK(clk), .Q(\fmem_data[15][2] ) );
  DFF_X1 \fmem_inst/mem_reg[15][3]  ( .D(n2984), .CK(clk), .Q(
        \fmem_inst/mem[15][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][3]  ( .D(\fmem_inst/mem[15][3] ), .CK(clk), .Q(\fmem_data[15][3] ), .QN(n3609) );
  DFF_X1 \fmem_inst/mem_reg[15][4]  ( .D(n2983), .CK(clk), .Q(
        \fmem_inst/mem[15][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][4]  ( .D(\fmem_inst/mem[15][4] ), .CK(clk), .Q(\fmem_data[15][4] ) );
  DFF_X1 \fmem_inst/mem_reg[15][5]  ( .D(n2982), .CK(clk), .Q(
        \fmem_inst/mem[15][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][5]  ( .D(\fmem_inst/mem[15][5] ), .CK(clk), .Q(\fmem_data[15][5] ), .QN(n3619) );
  DFF_X1 \fmem_inst/mem_reg[15][6]  ( .D(n2981), .CK(clk), .Q(
        \fmem_inst/mem[15][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][6]  ( .D(\fmem_inst/mem[15][6] ), .CK(clk), .Q(\fmem_data[15][6] ) );
  DFF_X1 \fmem_inst/mem_reg[15][7]  ( .D(n2980), .CK(clk), .Q(
        \fmem_inst/mem[15][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[15][7]  ( .D(\fmem_inst/mem[15][7] ), .CK(clk), .Q(\fmem_data[15][7] ), .QN(n3486) );
  DFF_X1 \fmem_inst/mem_reg[16][0]  ( .D(n2979), .CK(clk), .Q(
        \fmem_inst/mem[16][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][0]  ( .D(\fmem_inst/mem[16][0] ), .CK(clk), .Q(\fmem_data[16][0] ), .QN(n3573) );
  DFF_X1 \fmem_inst/mem_reg[16][1]  ( .D(n2978), .CK(clk), .Q(
        \fmem_inst/mem[16][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][1]  ( .D(\fmem_inst/mem[16][1] ), .CK(clk), .Q(\fmem_data[16][1] ), .QN(n3680) );
  DFF_X1 \fmem_inst/mem_reg[16][2]  ( .D(n2977), .CK(clk), .Q(
        \fmem_inst/mem[16][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][2]  ( .D(\fmem_inst/mem[16][2] ), .CK(clk), .Q(\fmem_data[16][2] ) );
  DFF_X1 \fmem_inst/mem_reg[16][3]  ( .D(n2976), .CK(clk), .Q(
        \fmem_inst/mem[16][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][3]  ( .D(\fmem_inst/mem[16][3] ), .CK(clk), .Q(\fmem_data[16][3] ), .QN(n3627) );
  DFF_X1 \fmem_inst/mem_reg[16][4]  ( .D(n2975), .CK(clk), .Q(
        \fmem_inst/mem[16][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][4]  ( .D(\fmem_inst/mem[16][4] ), .CK(clk), .Q(\fmem_data[16][4] ) );
  DFF_X1 \fmem_inst/mem_reg[16][5]  ( .D(n2974), .CK(clk), .Q(
        \fmem_inst/mem[16][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][5]  ( .D(\fmem_inst/mem[16][5] ), .CK(clk), .Q(\fmem_data[16][5] ), .QN(n3596) );
  DFF_X1 \fmem_inst/mem_reg[16][6]  ( .D(n2973), .CK(clk), .Q(
        \fmem_inst/mem[16][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][6]  ( .D(\fmem_inst/mem[16][6] ), .CK(clk), .Q(\fmem_data[16][6] ) );
  DFF_X1 \fmem_inst/mem_reg[16][7]  ( .D(n2972), .CK(clk), .Q(
        \fmem_inst/mem[16][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[16][7]  ( .D(\fmem_inst/mem[16][7] ), .CK(clk), .Q(\fmem_data[16][7] ), .QN(n3621) );
  DFF_X1 \fmem_inst/mem_reg[17][0]  ( .D(n2971), .CK(clk), .Q(
        \fmem_inst/mem[17][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][0]  ( .D(\fmem_inst/mem[17][0] ), .CK(clk), .Q(\fmem_data[17][0] ), .QN(n3566) );
  DFF_X1 \fmem_inst/mem_reg[17][1]  ( .D(n2970), .CK(clk), .Q(
        \fmem_inst/mem[17][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][1]  ( .D(\fmem_inst/mem[17][1] ), .CK(clk), .Q(\fmem_data[17][1] ), .QN(n3669) );
  DFF_X1 \fmem_inst/mem_reg[17][2]  ( .D(n2969), .CK(clk), .Q(
        \fmem_inst/mem[17][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][2]  ( .D(\fmem_inst/mem[17][2] ), .CK(clk), .Q(\fmem_data[17][2] ) );
  DFF_X1 \fmem_inst/mem_reg[17][3]  ( .D(n2968), .CK(clk), .Q(
        \fmem_inst/mem[17][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][3]  ( .D(\fmem_inst/mem[17][3] ), .CK(clk), .Q(\fmem_data[17][3] ), .QN(n3654) );
  DFF_X1 \fmem_inst/mem_reg[17][4]  ( .D(n2967), .CK(clk), .Q(
        \fmem_inst/mem[17][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][4]  ( .D(\fmem_inst/mem[17][4] ), .CK(clk), .Q(\fmem_data[17][4] ) );
  DFF_X1 \fmem_inst/mem_reg[17][5]  ( .D(n2966), .CK(clk), .Q(
        \fmem_inst/mem[17][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][5]  ( .D(\fmem_inst/mem[17][5] ), .CK(clk), .Q(\fmem_data[17][5] ), .QN(n3626) );
  DFF_X1 \fmem_inst/mem_reg[17][6]  ( .D(n2965), .CK(clk), .Q(
        \fmem_inst/mem[17][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][6]  ( .D(\fmem_inst/mem[17][6] ), .CK(clk), .Q(\fmem_data[17][6] ) );
  DFF_X1 \fmem_inst/mem_reg[17][7]  ( .D(n2964), .CK(clk), .Q(
        \fmem_inst/mem[17][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[17][7]  ( .D(\fmem_inst/mem[17][7] ), .CK(clk), .Q(\fmem_data[17][7] ), .QN(n3653) );
  DFF_X1 \fmem_inst/mem_reg[18][0]  ( .D(n2963), .CK(clk), .Q(
        \fmem_inst/mem[18][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][0]  ( .D(\fmem_inst/mem[18][0] ), .CK(clk), .Q(\fmem_data[18][0] ), .QN(n3580) );
  DFF_X1 \fmem_inst/mem_reg[18][1]  ( .D(n2962), .CK(clk), .Q(
        \fmem_inst/mem[18][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][1]  ( .D(\fmem_inst/mem[18][1] ), .CK(clk), .Q(\fmem_data[18][1] ), .QN(n3690) );
  DFF_X1 \fmem_inst/mem_reg[18][2]  ( .D(n2961), .CK(clk), .Q(
        \fmem_inst/mem[18][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][2]  ( .D(\fmem_inst/mem[18][2] ), .CK(clk), .Q(\fmem_data[18][2] ) );
  DFF_X1 \fmem_inst/mem_reg[18][3]  ( .D(n2960), .CK(clk), .Q(
        \fmem_inst/mem[18][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][3]  ( .D(\fmem_inst/mem[18][3] ), .CK(clk), .Q(\fmem_data[18][3] ), .QN(n3664) );
  DFF_X1 \fmem_inst/mem_reg[18][4]  ( .D(n2959), .CK(clk), .Q(
        \fmem_inst/mem[18][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][4]  ( .D(\fmem_inst/mem[18][4] ), .CK(clk), .Q(\fmem_data[18][4] ) );
  DFF_X1 \fmem_inst/mem_reg[18][5]  ( .D(n2958), .CK(clk), .Q(
        \fmem_inst/mem[18][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][5]  ( .D(\fmem_inst/mem[18][5] ), .CK(clk), .Q(\fmem_data[18][5] ), .QN(n3649) );
  DFF_X1 \fmem_inst/mem_reg[18][6]  ( .D(n2957), .CK(clk), .Q(
        \fmem_inst/mem[18][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][6]  ( .D(\fmem_inst/mem[18][6] ), .CK(clk), .Q(\fmem_data[18][6] ) );
  DFF_X1 \fmem_inst/mem_reg[18][7]  ( .D(n2956), .CK(clk), .Q(
        \fmem_inst/mem[18][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[18][7]  ( .D(\fmem_inst/mem[18][7] ), .CK(clk), .Q(\fmem_data[18][7] ), .QN(n3639) );
  DFF_X1 \fmem_inst/mem_reg[19][0]  ( .D(n2955), .CK(clk), .Q(
        \fmem_inst/mem[19][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][0]  ( .D(\fmem_inst/mem[19][0] ), .CK(clk), .Q(\fmem_data[19][0] ), .QN(n3633) );
  DFF_X1 \fmem_inst/mem_reg[19][1]  ( .D(n2954), .CK(clk), .Q(
        \fmem_inst/mem[19][1] ) );
  DFF_X1 \fmem_inst/mem_reg[19][2]  ( .D(n2953), .CK(clk), .Q(
        \fmem_inst/mem[19][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][2]  ( .D(\fmem_inst/mem[19][2] ), .CK(clk), .Q(\fmem_data[19][2] ) );
  DFF_X1 \fmem_inst/mem_reg[19][3]  ( .D(n2952), .CK(clk), .Q(
        \fmem_inst/mem[19][3] ) );
  DFF_X1 \fmem_inst/mem_reg[19][4]  ( .D(n2951), .CK(clk), .Q(
        \fmem_inst/mem[19][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][4]  ( .D(\fmem_inst/mem[19][4] ), .CK(clk), .Q(\fmem_data[19][4] ) );
  DFF_X1 \fmem_inst/mem_reg[19][5]  ( .D(n2950), .CK(clk), .Q(
        \fmem_inst/mem[19][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][5]  ( .D(\fmem_inst/mem[19][5] ), .CK(clk), .Q(\fmem_data[19][5] ), .QN(n3606) );
  DFF_X1 \fmem_inst/mem_reg[19][6]  ( .D(n2949), .CK(clk), .Q(
        \fmem_inst/mem[19][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][6]  ( .D(\fmem_inst/mem[19][6] ), .CK(clk), .Q(\fmem_data[19][6] ) );
  DFF_X1 \fmem_inst/mem_reg[19][7]  ( .D(n2948), .CK(clk), .Q(
        \fmem_inst/mem[19][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[19][7]  ( .D(\fmem_inst/mem[19][7] ), .CK(clk), .Q(\fmem_data[19][7] ), .QN(n3640) );
  DFF_X1 \fmem_inst/mem_reg[20][0]  ( .D(n2947), .CK(clk), .Q(
        \fmem_inst/mem[20][0] ) );
  DFF_X1 \fmem_inst/mem_reg[20][1]  ( .D(n2946), .CK(clk), .Q(
        \fmem_inst/mem[20][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][1]  ( .D(\fmem_inst/mem[20][1] ), .CK(clk), .Q(\fmem_data[20][1] ), .QN(n4018) );
  DFF_X1 \fmem_inst/mem_reg[20][2]  ( .D(n2945), .CK(clk), .Q(
        \fmem_inst/mem[20][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][2]  ( .D(\fmem_inst/mem[20][2] ), .CK(clk), .Q(\fmem_data[20][2] ) );
  DFF_X1 \fmem_inst/mem_reg[20][3]  ( .D(n2944), .CK(clk), .Q(
        \fmem_inst/mem[20][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][3]  ( .D(\fmem_inst/mem[20][3] ), .CK(clk), .Q(\fmem_data[20][3] ), .QN(n3593) );
  DFF_X1 \fmem_inst/mem_reg[20][4]  ( .D(n2943), .CK(clk), .Q(
        \fmem_inst/mem[20][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][4]  ( .D(\fmem_inst/mem[20][4] ), .CK(clk), .Q(\fmem_data[20][4] ) );
  DFF_X1 \fmem_inst/mem_reg[20][5]  ( .D(n2942), .CK(clk), .Q(
        \fmem_inst/mem[20][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][5]  ( .D(\fmem_inst/mem[20][5] ), .CK(clk), .Q(\fmem_data[20][5] ), .QN(n3628) );
  DFF_X1 \fmem_inst/mem_reg[20][6]  ( .D(n2941), .CK(clk), .Q(
        \fmem_inst/mem[20][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][6]  ( .D(\fmem_inst/mem[20][6] ), .CK(clk), .Q(\fmem_data[20][6] ) );
  DFF_X1 \fmem_inst/mem_reg[20][7]  ( .D(n2940), .CK(clk), .Q(
        \fmem_inst/mem[20][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[20][7]  ( .D(\fmem_inst/mem[20][7] ), .CK(clk), .Q(\fmem_data[20][7] ), .QN(n3484) );
  DFF_X1 \fmem_inst/mem_reg[21][0]  ( .D(n2939), .CK(clk), .Q(
        \fmem_inst/mem[21][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][0]  ( .D(\fmem_inst/mem[21][0] ), .CK(clk), .Q(\fmem_data[21][0] ), .QN(n3570) );
  DFF_X1 \fmem_inst/mem_reg[21][1]  ( .D(n2938), .CK(clk), .Q(
        \fmem_inst/mem[21][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][1]  ( .D(\fmem_inst/mem[21][1] ), .CK(clk), .Q(\fmem_data[21][1] ), .QN(n3999) );
  DFF_X1 \fmem_inst/mem_reg[21][2]  ( .D(n2937), .CK(clk), .Q(
        \fmem_inst/mem[21][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][2]  ( .D(\fmem_inst/mem[21][2] ), .CK(clk), .Q(\fmem_data[21][2] ) );
  DFF_X1 \fmem_inst/mem_reg[21][3]  ( .D(n2936), .CK(clk), .Q(
        \fmem_inst/mem[21][3] ) );
  DFF_X1 \fmem_inst/mem_reg[21][4]  ( .D(n2935), .CK(clk), .Q(
        \fmem_inst/mem[21][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][4]  ( .D(\fmem_inst/mem[21][4] ), .CK(clk), .Q(\fmem_data[21][4] ) );
  DFF_X1 \fmem_inst/mem_reg[21][5]  ( .D(n2934), .CK(clk), .Q(
        \fmem_inst/mem[21][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][5]  ( .D(\fmem_inst/mem[21][5] ), .CK(clk), .Q(\fmem_data[21][5] ), .QN(n3665) );
  DFF_X1 \fmem_inst/mem_reg[21][6]  ( .D(n2933), .CK(clk), .Q(
        \fmem_inst/mem[21][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][6]  ( .D(\fmem_inst/mem[21][6] ), .CK(clk), .Q(\fmem_data[21][6] ) );
  DFF_X1 \fmem_inst/mem_reg[21][7]  ( .D(n2932), .CK(clk), .Q(
        \fmem_inst/mem[21][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[21][7]  ( .D(\fmem_inst/mem[21][7] ), .CK(clk), .Q(\fmem_data[21][7] ), .QN(n3600) );
  DFF_X1 \fmem_inst/mem_reg[22][0]  ( .D(n2931), .CK(clk), .Q(
        \fmem_inst/mem[22][0] ) );
  DFF_X1 \fmem_inst/mem_reg[22][1]  ( .D(n2930), .CK(clk), .Q(
        \fmem_inst/mem[22][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][1]  ( .D(\fmem_inst/mem[22][1] ), .CK(clk), .Q(\fmem_data[22][1] ), .QN(n3693) );
  DFF_X1 \fmem_inst/mem_reg[22][2]  ( .D(n2929), .CK(clk), .Q(
        \fmem_inst/mem[22][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][2]  ( .D(\fmem_inst/mem[22][2] ), .CK(clk), .Q(\fmem_data[22][2] ) );
  DFF_X1 \fmem_inst/mem_reg[22][3]  ( .D(n2928), .CK(clk), .Q(
        \fmem_inst/mem[22][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][3]  ( .D(\fmem_inst/mem[22][3] ), .CK(clk), .Q(\fmem_data[22][3] ), .QN(n3603) );
  DFF_X1 \fmem_inst/mem_reg[22][4]  ( .D(n2927), .CK(clk), .Q(
        \fmem_inst/mem[22][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][4]  ( .D(\fmem_inst/mem[22][4] ), .CK(clk), .Q(\fmem_data[22][4] ) );
  DFF_X1 \fmem_inst/mem_reg[22][5]  ( .D(n2926), .CK(clk), .Q(
        \fmem_inst/mem[22][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][5]  ( .D(\fmem_inst/mem[22][5] ), .CK(clk), .Q(\fmem_data[22][5] ), .QN(n3591) );
  DFF_X1 \fmem_inst/mem_reg[22][6]  ( .D(n2925), .CK(clk), .Q(
        \fmem_inst/mem[22][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][6]  ( .D(\fmem_inst/mem[22][6] ), .CK(clk), .Q(\fmem_data[22][6] ) );
  DFF_X1 \fmem_inst/mem_reg[22][7]  ( .D(n2924), .CK(clk), .Q(
        \fmem_inst/mem[22][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][7]  ( .D(\fmem_inst/mem[22][7] ), .CK(clk), .Q(\fmem_data[22][7] ), .QN(n3645) );
  DFF_X1 \fmem_inst/mem_reg[23][0]  ( .D(n2923), .CK(clk), .Q(
        \fmem_inst/mem[23][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][0]  ( .D(\fmem_inst/mem[23][0] ), .CK(clk), .Q(\fmem_data[23][0] ), .QN(n3662) );
  DFF_X1 \fmem_inst/mem_reg[23][1]  ( .D(n2922), .CK(clk), .Q(
        \fmem_inst/mem[23][1] ) );
  DFF_X1 \fmem_inst/mem_reg[23][2]  ( .D(n2921), .CK(clk), .Q(
        \fmem_inst/mem[23][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][2]  ( .D(\fmem_inst/mem[23][2] ), .CK(clk), .Q(\fmem_data[23][2] ) );
  DFF_X1 \fmem_inst/mem_reg[23][3]  ( .D(n2920), .CK(clk), .Q(
        \fmem_inst/mem[23][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][3]  ( .D(\fmem_inst/mem[23][3] ), .CK(clk), .Q(\fmem_data[23][3] ), .QN(n3674) );
  DFF_X1 \fmem_inst/mem_reg[23][4]  ( .D(n2919), .CK(clk), .Q(
        \fmem_inst/mem[23][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][4]  ( .D(\fmem_inst/mem[23][4] ), .CK(clk), .Q(\fmem_data[23][4] ) );
  DFF_X1 \fmem_inst/mem_reg[23][5]  ( .D(n2918), .CK(clk), .Q(
        \fmem_inst/mem[23][5] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][5]  ( .D(\fmem_inst/mem[23][5] ), .CK(clk), .Q(\fmem_data[23][5] ), .QN(n3687) );
  DFF_X1 \fmem_inst/mem_reg[23][6]  ( .D(n2917), .CK(clk), .Q(
        \fmem_inst/mem[23][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][6]  ( .D(\fmem_inst/mem[23][6] ), .CK(clk), .Q(\fmem_data[23][6] ) );
  DFF_X1 \fmem_inst/mem_reg[23][7]  ( .D(n2916), .CK(clk), .Q(
        \fmem_inst/mem[23][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[23][7]  ( .D(\fmem_inst/mem[23][7] ), .CK(clk), .Q(\fmem_data[23][7] ), .QN(n3668) );
  DFF_X1 conv_pre_start_reg ( .D(N229), .CK(clk), .Q(conv_pre_start) );
  DFF_X1 \fmem_inst/mem_reg[31][0]  ( .D(n2859), .CK(clk), .Q(
        \fmem_inst/mem[31][0] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][0]  ( .D(\fmem_inst/mem[31][0] ), .CK(clk), .Q(n3489), .QN(n3931) );
  DFF_X1 \fmem_inst/mem_reg[31][1]  ( .D(n2858), .CK(clk), .Q(
        \fmem_inst/mem[31][1] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][1]  ( .D(\fmem_inst/mem[31][1] ), .CK(clk), .Q(\fmem_data[31][1] ) );
  DFF_X1 \fmem_inst/mem_reg[31][2]  ( .D(n2857), .CK(clk), .Q(
        \fmem_inst/mem[31][2] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][2]  ( .D(\fmem_inst/mem[31][2] ), .CK(clk), .Q(\fmem_data[31][2] ) );
  DFF_X1 \fmem_inst/mem_reg[31][3]  ( .D(n2856), .CK(clk), .Q(
        \fmem_inst/mem[31][3] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][3]  ( .D(\fmem_inst/mem[31][3] ), .CK(clk), .Q(\fmem_data[31][3] ), .QN(n3485) );
  DFF_X1 \fmem_inst/mem_reg[31][4]  ( .D(n2855), .CK(clk), .Q(
        \fmem_inst/mem[31][4] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][4]  ( .D(\fmem_inst/mem[31][4] ), .CK(clk), .Q(\fmem_data[31][4] ) );
  DFF_X1 \fmem_inst/mem_reg[31][5]  ( .D(n2854), .CK(clk), .Q(
        \fmem_inst/mem[31][5] ) );
  DFF_X1 \fmem_inst/mem_reg[31][6]  ( .D(n2853), .CK(clk), .Q(
        \fmem_inst/mem[31][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][6]  ( .D(\fmem_inst/mem[31][6] ), .CK(clk), .Q(\fmem_data[31][6] ) );
  DFF_X1 \fmem_inst/mem_reg[31][7]  ( .D(n2852), .CK(clk), .Q(
        \fmem_inst/mem[31][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][7]  ( .D(\fmem_inst/mem[31][7] ), .CK(clk), .Q(\fmem_data[31][7] ), .QN(n3487) );
  DFF_X1 \xmem_inst/mem_reg[127][0]  ( .D(n1827), .CK(clk), .Q(
        \xmem_inst/mem[127][0] ) );
  DFF_X1 \xmem_inst/mem_reg[127][1]  ( .D(n1826), .CK(clk), .Q(
        \xmem_inst/mem[127][1] ) );
  DFF_X1 \xmem_inst/mem_reg[127][2]  ( .D(n1825), .CK(clk), .Q(
        \xmem_inst/mem[127][2] ) );
  DFF_X1 \xmem_inst/mem_reg[127][3]  ( .D(n1824), .CK(clk), .Q(
        \xmem_inst/mem[127][3] ) );
  DFF_X1 \xmem_inst/mem_reg[127][4]  ( .D(n1823), .CK(clk), .Q(
        \xmem_inst/mem[127][4] ) );
  DFF_X1 \xmem_inst/mem_reg[127][5]  ( .D(n1822), .CK(clk), .Q(
        \xmem_inst/mem[127][5] ) );
  DFF_X1 \xmem_inst/mem_reg[127][6]  ( .D(n1821), .CK(clk), .Q(
        \xmem_inst/mem[127][6] ) );
  DFF_X1 \xmem_inst/mem_reg[127][7]  ( .D(n1820), .CK(clk), .Q(
        \xmem_inst/mem[127][7] ) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n3115), .CK(clk), .Q(
        m_valid_y), .QN(n39050) );
  DFF_X1 \ctrl_conv_output_inst/load_xaddr_val_reg[0]  ( .D(n1819), .CK(clk), 
        .Q(\add_x_2/A[0] ), .QN(n39052) );
  DFF_X1 \ctrl_conv_output_inst/load_xaddr_val_reg[2]  ( .D(n1817), .CK(clk), 
        .Q(N345), .QN(n39053) );
  DFF_X1 \ctrl_conv_output_inst/load_xaddr_val_reg[3]  ( .D(n1816), .CK(clk), 
        .Q(N466), .QN(n39035) );
  DFF_X1 \fmem_inst/data_out_reg[8][0]  ( .D(\fmem_inst/mem[8][0] ), .CK(clk), 
        .Q(\fmem_data[8][0] ), .QN(n3574) );
  DFF_X1 \fmem_inst/data_out_reg[6][0]  ( .D(\fmem_inst/mem[6][0] ), .CK(clk), 
        .Q(\fmem_data[6][0] ), .QN(n3559) );
  DFF_X1 \fmem_inst/data_out_reg[12][0]  ( .D(\fmem_inst/mem[12][0] ), .CK(clk), .Q(\fmem_data[12][0] ), .QN(n3572) );
  DFF_X1 \fmem_inst/data_out_reg[28][0]  ( .D(\fmem_inst/mem[28][0] ), .CK(clk), .Q(\fmem_data[28][0] ), .QN(n3562) );
  DFF_X1 \xmem_inst/data_out_reg[66][6]  ( .D(\xmem_inst/mem[66][6] ), .CK(clk), .Q(\xmem_data[66][6] ) );
  DFF_X1 \fmem_inst/data_out_reg[22][0]  ( .D(\fmem_inst/mem[22][0] ), .CK(clk), .Q(\fmem_data[22][0] ), .QN(n3567) );
  DFF_X1 \fmem_inst/data_out_reg[20][0]  ( .D(\fmem_inst/mem[20][0] ), .CK(clk), .Q(\fmem_data[20][0] ), .QN(n3647) );
  DFF_X1 \fmem_inst/data_out_reg[30][0]  ( .D(\fmem_inst/mem[30][0] ), .CK(clk), .Q(\fmem_data[30][0] ), .QN(n3560) );
  DFF_X2 \xmem_inst/data_out_reg[76][2]  ( .D(\xmem_inst/mem[76][2] ), .CK(clk), .Q(\xmem_data[76][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][2]  ( .D(\xmem_inst/mem[62][2] ), .CK(clk), .Q(\xmem_data[62][2] ) );
  DFF_X1 \ctrl_conv_output_inst/load_xaddr_val_reg[1]  ( .D(n38996), .CK(clk), 
        .Q(n39010), .QN(N284) );
  DFF_X2 \ctrl_conv_output_inst/load_xaddr_val_reg[6]  ( .D(n3114), .CK(clk), 
        .Q(load_xaddr_val[6]), .QN(n39040) );
  DFF_X1 \ctrl_conv_output_inst/load_xaddr_val_reg[4]  ( .D(n1815), .CK(clk), 
        .Q(n39054), .QN(n38997) );
  DFF_X2 \xmem_inst/data_out_reg[7][7]  ( .D(\xmem_inst/mem[7][7] ), .CK(clk), 
        .Q(\xmem_data[7][7] ) );
  DFF_X1 \fmem_inst/data_out_reg[31][5]  ( .D(\fmem_inst/mem[31][5] ), .CK(clk), .Q(\fmem_data[31][5] ), .QN(n3488) );
  DFF_X1 \fmem_inst/data_out_reg[27][1]  ( .D(\fmem_inst/mem[27][1] ), .CK(clk), .Q(\fmem_data[27][1] ), .QN(n3740) );
  DFF_X1 \fmem_inst/data_out_reg[23][1]  ( .D(\fmem_inst/mem[23][1] ), .CK(clk), .Q(\fmem_data[23][1] ), .QN(n3735) );
  DFF_X1 \fmem_inst/data_out_reg[26][1]  ( .D(\fmem_inst/mem[26][1] ), .CK(clk), .Q(\fmem_data[26][1] ), .QN(n3732) );
  DFF_X1 \fmem_inst/data_out_reg[19][1]  ( .D(\fmem_inst/mem[19][1] ), .CK(clk), .Q(\fmem_data[19][1] ), .QN(n3717) );
  DFF_X1 \fmem_inst/data_out_reg[5][3]  ( .D(\fmem_inst/mem[5][3] ), .CK(clk), 
        .Q(\fmem_data[5][3] ), .QN(n3701) );
  DFF_X1 \fmem_inst/data_out_reg[8][3]  ( .D(\fmem_inst/mem[8][3] ), .CK(clk), 
        .Q(\fmem_data[8][3] ), .QN(n3700) );
  DFF_X1 \fmem_inst/data_out_reg[11][5]  ( .D(\fmem_inst/mem[11][5] ), .CK(clk), .Q(\fmem_data[11][5] ), .QN(n3697) );
  DFF_X1 \fmem_inst/data_out_reg[6][5]  ( .D(\fmem_inst/mem[6][5] ), .CK(clk), 
        .Q(\fmem_data[6][5] ), .QN(n3696) );
  DFF_X1 \fmem_inst/data_out_reg[3][5]  ( .D(\fmem_inst/mem[3][5] ), .CK(clk), 
        .Q(\fmem_data[3][5] ), .QN(n3688) );
  DFF_X1 \fmem_inst/data_out_reg[19][3]  ( .D(\fmem_inst/mem[19][3] ), .CK(clk), .Q(\fmem_data[19][3] ), .QN(n3686) );
  DFF_X1 \fmem_inst/data_out_reg[7][3]  ( .D(\fmem_inst/mem[7][3] ), .CK(clk), 
        .Q(\fmem_data[7][3] ), .QN(n3685) );
  DFF_X1 \fmem_inst/data_out_reg[21][3]  ( .D(\fmem_inst/mem[21][3] ), .CK(clk), .Q(\fmem_data[21][3] ), .QN(n3684) );
  DFF_X2 \xmem_inst/data_out_reg[110][6]  ( .D(\xmem_inst/mem[110][6] ), .CK(
        clk), .Q(\xmem_data[110][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][5]  ( .D(\xmem_inst/mem[17][5] ), .CK(clk), .Q(\xmem_data[17][5] ), .QN(n39005) );
  DFF_X2 \xmem_inst/data_out_reg[17][3]  ( .D(\xmem_inst/mem[17][3] ), .CK(clk), .Q(\xmem_data[17][3] ), .QN(n39009) );
  DFF_X2 \xmem_inst/data_out_reg[17][2]  ( .D(\xmem_inst/mem[17][2] ), .CK(clk), .Q(\xmem_data[17][2] ), .QN(n39007) );
  DFF_X2 \xmem_inst/data_out_reg[22][1]  ( .D(\xmem_inst/mem[22][1] ), .CK(clk), .Q(\xmem_data[22][1] ), .QN(n39002) );
  DFF_X2 \xmem_inst/data_out_reg[22][3]  ( .D(\xmem_inst/mem[22][3] ), .CK(clk), .Q(\xmem_data[22][3] ), .QN(n39006) );
  DFF_X2 \xmem_inst/data_out_reg[22][2]  ( .D(\xmem_inst/mem[22][2] ), .CK(clk), .Q(\xmem_data[22][2] ), .QN(n39003) );
  DFF_X2 \xmem_inst/data_out_reg[95][1]  ( .D(\xmem_inst/mem[95][1] ), .CK(clk), .Q(\xmem_data[95][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][1]  ( .D(\xmem_inst/mem[79][1] ), .CK(clk), .Q(\xmem_data[79][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][1]  ( .D(\xmem_inst/mem[13][1] ), .CK(clk), .Q(\xmem_data[13][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][4]  ( .D(\xmem_inst/mem[45][4] ), .CK(clk), .Q(\xmem_data[45][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][4]  ( .D(\xmem_inst/mem[49][4] ), .CK(clk), .Q(\xmem_data[49][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][4]  ( .D(\xmem_inst/mem[47][4] ), .CK(clk), .Q(\xmem_data[47][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][1]  ( .D(\xmem_inst/mem[0][1] ), .CK(clk), 
        .Q(\xmem_data[0][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][7]  ( .D(\xmem_inst/mem[14][7] ), .CK(clk), .Q(\xmem_data[14][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][5]  ( .D(\xmem_inst/mem[19][5] ), .CK(clk), .Q(\xmem_data[19][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][1]  ( .D(\xmem_inst/mem[127][1] ), .CK(
        clk), .Q(\xmem_data[127][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][1]  ( .D(\xmem_inst/mem[125][1] ), .CK(
        clk), .Q(\xmem_data[125][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][1]  ( .D(\xmem_inst/mem[123][1] ), .CK(
        clk), .Q(\xmem_data[123][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][1]  ( .D(\xmem_inst/mem[117][1] ), .CK(
        clk), .Q(\xmem_data[117][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][1]  ( .D(\xmem_inst/mem[113][1] ), .CK(
        clk), .Q(\xmem_data[113][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][1]  ( .D(\xmem_inst/mem[99][1] ), .CK(clk), .Q(\xmem_data[99][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][1]  ( .D(\xmem_inst/mem[111][1] ), .CK(
        clk), .Q(\xmem_data[111][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][1]  ( .D(\xmem_inst/mem[107][1] ), .CK(
        clk), .Q(\xmem_data[107][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][1]  ( .D(\xmem_inst/mem[91][1] ), .CK(clk), .Q(\xmem_data[91][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][1]  ( .D(\xmem_inst/mem[73][1] ), .CK(clk), .Q(\xmem_data[73][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][1]  ( .D(\xmem_inst/mem[75][1] ), .CK(clk), .Q(\xmem_data[75][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][1]  ( .D(\xmem_inst/mem[77][1] ), .CK(clk), .Q(\xmem_data[77][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][1]  ( .D(\xmem_inst/mem[69][1] ), .CK(clk), .Q(\xmem_data[69][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][1]  ( .D(\xmem_inst/mem[67][1] ), .CK(clk), .Q(\xmem_data[67][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][1]  ( .D(\xmem_inst/mem[27][1] ), .CK(clk), .Q(\xmem_data[27][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][1]  ( .D(\xmem_inst/mem[9][1] ), .CK(clk), 
        .Q(\xmem_data[9][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][1]  ( .D(\xmem_inst/mem[59][1] ), .CK(clk), .Q(\xmem_data[59][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][1]  ( .D(\xmem_inst/mem[45][1] ), .CK(clk), .Q(\xmem_data[45][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][1]  ( .D(\xmem_inst/mem[41][1] ), .CK(clk), .Q(\xmem_data[41][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][2]  ( .D(\xmem_inst/mem[19][2] ), .CK(clk), .Q(\xmem_data[19][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[7][2]  ( .D(\xmem_inst/mem[7][2] ), .CK(clk), 
        .Q(\xmem_data[7][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][7]  ( .D(\xmem_inst/mem[31][7] ), .CK(clk), .Q(\xmem_data[31][7] ), .QN(n39024) );
  DFF_X2 \xmem_inst/data_out_reg[85][3]  ( .D(\xmem_inst/mem[85][3] ), .CK(clk), .Q(\xmem_data[85][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][3]  ( .D(\xmem_inst/mem[81][3] ), .CK(clk), .Q(\xmem_data[81][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][3]  ( .D(\xmem_inst/mem[117][3] ), .CK(
        clk), .Q(\xmem_data[117][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][3]  ( .D(\xmem_inst/mem[61][3] ), .CK(clk), .Q(\xmem_data[61][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][3]  ( .D(\xmem_inst/mem[49][3] ), .CK(clk), .Q(\xmem_data[49][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][3]  ( .D(\xmem_inst/mem[47][3] ), .CK(clk), .Q(\xmem_data[47][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][3]  ( .D(\xmem_inst/mem[45][3] ), .CK(clk), .Q(\xmem_data[45][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][3]  ( .D(\xmem_inst/mem[41][3] ), .CK(clk), .Q(\xmem_data[41][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][3]  ( .D(\xmem_inst/mem[39][3] ), .CK(clk), .Q(\xmem_data[39][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][3]  ( .D(\xmem_inst/mem[27][3] ), .CK(clk), .Q(\xmem_data[27][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][3]  ( .D(\xmem_inst/mem[29][3] ), .CK(clk), .Q(\xmem_data[29][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][4]  ( .D(\xmem_inst/mem[39][4] ), .CK(clk), .Q(\xmem_data[39][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][4]  ( .D(\xmem_inst/mem[59][4] ), .CK(clk), .Q(\xmem_data[59][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][4]  ( .D(\xmem_inst/mem[57][4] ), .CK(clk), .Q(\xmem_data[57][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][4]  ( .D(\xmem_inst/mem[41][4] ), .CK(clk), .Q(\xmem_data[41][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][4]  ( .D(\xmem_inst/mem[53][4] ), .CK(clk), .Q(\xmem_data[53][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][4]  ( .D(\xmem_inst/mem[101][4] ), .CK(
        clk), .Q(\xmem_data[101][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][4]  ( .D(\xmem_inst/mem[99][4] ), .CK(clk), .Q(\xmem_data[99][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][4]  ( .D(\xmem_inst/mem[127][4] ), .CK(
        clk), .Q(\xmem_data[127][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][4]  ( .D(\xmem_inst/mem[125][4] ), .CK(
        clk), .Q(\xmem_data[125][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][4]  ( .D(\xmem_inst/mem[123][4] ), .CK(
        clk), .Q(\xmem_data[123][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][4]  ( .D(\xmem_inst/mem[111][4] ), .CK(
        clk), .Q(\xmem_data[111][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][4]  ( .D(\xmem_inst/mem[109][4] ), .CK(
        clk), .Q(\xmem_data[109][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][4]  ( .D(\xmem_inst/mem[107][4] ), .CK(
        clk), .Q(\xmem_data[107][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][4]  ( .D(\xmem_inst/mem[105][4] ), .CK(
        clk), .Q(\xmem_data[105][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][4]  ( .D(\xmem_inst/mem[117][4] ), .CK(
        clk), .Q(\xmem_data[117][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][4]  ( .D(\xmem_inst/mem[113][4] ), .CK(
        clk), .Q(\xmem_data[113][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][5]  ( .D(\xmem_inst/mem[71][5] ), .CK(clk), .Q(\xmem_data[71][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][1]  ( .D(\xmem_inst/mem[81][1] ), .CK(clk), .Q(\xmem_data[81][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][1]  ( .D(\xmem_inst/mem[19][1] ), .CK(clk), .Q(\xmem_data[19][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][1]  ( .D(\xmem_inst/mem[17][1] ), .CK(clk), .Q(\xmem_data[17][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][1]  ( .D(\xmem_inst/mem[61][1] ), .CK(clk), .Q(\xmem_data[61][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][0]  ( .D(\xmem_inst/mem[23][0] ), .CK(clk), .Q(\xmem_data[23][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][1]  ( .D(\xmem_inst/mem[93][1] ), .CK(clk), .Q(\xmem_data[93][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][1]  ( .D(\xmem_inst/mem[25][1] ), .CK(clk), .Q(\xmem_data[25][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][1]  ( .D(\xmem_inst/mem[39][1] ), .CK(clk), .Q(\xmem_data[39][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][1]  ( .D(\xmem_inst/mem[57][1] ), .CK(clk), .Q(\xmem_data[57][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][4]  ( .D(\xmem_inst/mem[61][4] ), .CK(clk), .Q(\xmem_data[61][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][0]  ( .D(\xmem_inst/mem[17][0] ), .CK(clk), .Q(\xmem_data[17][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][5]  ( .D(\xmem_inst/mem[30][5] ), .CK(clk), .Q(\xmem_data[30][5] ), .QN(n39023) );
  DFF_X2 \xmem_inst/data_out_reg[24][5]  ( .D(\xmem_inst/mem[24][5] ), .CK(clk), .Q(\xmem_data[24][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][1]  ( .D(\xmem_inst/mem[30][1] ), .CK(clk), .Q(\xmem_data[30][1] ), .QN(n39014) );
  DFF_X2 \xmem_inst/data_out_reg[14][1]  ( .D(\xmem_inst/mem[14][1] ), .CK(clk), .Q(\xmem_data[14][1] ), .QN(n39015) );
  DFF_X2 \xmem_inst/data_out_reg[6][1]  ( .D(\xmem_inst/mem[6][1] ), .CK(clk), 
        .Q(\xmem_data[6][1] ), .QN(n39025) );
  DFF_X2 \xmem_inst/data_out_reg[52][1]  ( .D(\xmem_inst/mem[52][1] ), .CK(clk), .Q(\xmem_data[52][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][2]  ( .D(\xmem_inst/mem[30][2] ), .CK(clk), .Q(\xmem_data[30][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][2]  ( .D(\xmem_inst/mem[0][2] ), .CK(clk), 
        .Q(\xmem_data[0][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][7]  ( .D(\xmem_inst/mem[8][7] ), .CK(clk), 
        .Q(\xmem_data[8][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][1]  ( .D(\xmem_inst/mem[51][1] ), .CK(clk), .Q(\xmem_data[51][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][7]  ( .D(\xmem_inst/mem[28][7] ), .CK(clk), .Q(\xmem_data[28][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][0]  ( .D(\xmem_inst/mem[28][0] ), .CK(clk), .Q(\xmem_data[28][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][3]  ( .D(\xmem_inst/mem[13][3] ), .CK(clk), .Q(\xmem_data[13][3] ), .QN(n39018) );
  DFF_X2 \xmem_inst/data_out_reg[75][0]  ( .D(\xmem_inst/mem[75][0] ), .CK(clk), .Q(\xmem_data[75][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][0]  ( .D(\xmem_inst/mem[85][0] ), .CK(clk), .Q(\xmem_data[85][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][5]  ( .D(\xmem_inst/mem[14][5] ), .CK(clk), .Q(\xmem_data[14][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][3]  ( .D(\xmem_inst/mem[6][3] ), .CK(clk), 
        .Q(\xmem_data[6][3] ), .QN(n39012) );
  DFF_X2 \xmem_inst/data_out_reg[36][1]  ( .D(\xmem_inst/mem[36][1] ), .CK(clk), .Q(\xmem_data[36][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[7][4]  ( .D(\xmem_inst/mem[7][4] ), .CK(clk), 
        .Q(\xmem_data[7][4] ), .QN(n39039) );
  DFF_X2 \xmem_inst/data_out_reg[27][7]  ( .D(\xmem_inst/mem[27][7] ), .CK(clk), .Q(\xmem_data[27][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][6]  ( .D(\xmem_inst/mem[79][6] ), .CK(clk), .Q(\xmem_data[79][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][4]  ( .D(\xmem_inst/mem[86][4] ), .CK(clk), .Q(\xmem_data[86][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][0]  ( .D(\xmem_inst/mem[91][0] ), .CK(clk), .Q(\xmem_data[91][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][3]  ( .D(\xmem_inst/mem[3][3] ), .CK(clk), 
        .Q(\xmem_data[3][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][0]  ( .D(\xmem_inst/mem[39][0] ), .CK(clk), .Q(\xmem_data[39][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][4]  ( .D(\xmem_inst/mem[3][4] ), .CK(clk), 
        .Q(\xmem_data[3][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][0]  ( .D(\xmem_inst/mem[127][0] ), .CK(
        clk), .Q(\xmem_data[127][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][0]  ( .D(\xmem_inst/mem[95][0] ), .CK(clk), .Q(\xmem_data[95][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][5]  ( .D(\xmem_inst/mem[1][5] ), .CK(clk), 
        .Q(\xmem_data[1][5] ), .QN(n39030) );
  DFF_X2 \xmem_inst/data_out_reg[99][0]  ( .D(\xmem_inst/mem[99][0] ), .CK(clk), .Q(\xmem_data[99][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][0]  ( .D(\xmem_inst/mem[117][0] ), .CK(
        clk), .Q(\xmem_data[117][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][0]  ( .D(\xmem_inst/mem[113][0] ), .CK(
        clk), .Q(\xmem_data[113][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][0]  ( .D(\xmem_inst/mem[109][0] ), .CK(
        clk), .Q(\xmem_data[109][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][0]  ( .D(\xmem_inst/mem[107][0] ), .CK(
        clk), .Q(\xmem_data[107][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][0]  ( .D(\xmem_inst/mem[105][0] ), .CK(
        clk), .Q(\xmem_data[105][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][0]  ( .D(\xmem_inst/mem[125][0] ), .CK(
        clk), .Q(\xmem_data[125][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][0]  ( .D(\xmem_inst/mem[123][0] ), .CK(
        clk), .Q(\xmem_data[123][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][0]  ( .D(\xmem_inst/mem[69][0] ), .CK(clk), .Q(\xmem_data[69][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][0]  ( .D(\xmem_inst/mem[67][0] ), .CK(clk), .Q(\xmem_data[67][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][0]  ( .D(\xmem_inst/mem[81][0] ), .CK(clk), .Q(\xmem_data[81][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][0]  ( .D(\xmem_inst/mem[77][0] ), .CK(clk), .Q(\xmem_data[77][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][0]  ( .D(\xmem_inst/mem[73][0] ), .CK(clk), .Q(\xmem_data[73][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][3]  ( .D(\xmem_inst/mem[1][3] ), .CK(clk), 
        .Q(\xmem_data[1][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][7]  ( .D(\xmem_inst/mem[109][7] ), .CK(
        clk), .Q(\xmem_data[109][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][7]  ( .D(\xmem_inst/mem[107][7] ), .CK(
        clk), .Q(\xmem_data[107][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][7]  ( .D(\xmem_inst/mem[105][7] ), .CK(
        clk), .Q(\xmem_data[105][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][7]  ( .D(\xmem_inst/mem[101][7] ), .CK(
        clk), .Q(\xmem_data[101][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][7]  ( .D(\xmem_inst/mem[99][7] ), .CK(clk), .Q(\xmem_data[99][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][7]  ( .D(\xmem_inst/mem[123][7] ), .CK(
        clk), .Q(\xmem_data[123][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][3]  ( .D(\xmem_inst/mem[109][3] ), .CK(
        clk), .Q(\xmem_data[109][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][3]  ( .D(\xmem_inst/mem[107][3] ), .CK(
        clk), .Q(\xmem_data[107][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][3]  ( .D(\xmem_inst/mem[105][3] ), .CK(
        clk), .Q(\xmem_data[105][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][0]  ( .D(\xmem_inst/mem[47][0] ), .CK(clk), .Q(\xmem_data[47][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][0]  ( .D(\xmem_inst/mem[45][0] ), .CK(clk), .Q(\xmem_data[45][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][0]  ( .D(\xmem_inst/mem[55][0] ), .CK(clk), .Q(\xmem_data[55][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][0]  ( .D(\xmem_inst/mem[53][0] ), .CK(clk), .Q(\xmem_data[53][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][0]  ( .D(\xmem_inst/mem[51][0] ), .CK(clk), .Q(\xmem_data[51][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][0]  ( .D(\xmem_inst/mem[49][0] ), .CK(clk), .Q(\xmem_data[49][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][0]  ( .D(\xmem_inst/mem[57][0] ), .CK(clk), .Q(\xmem_data[57][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][3]  ( .D(\xmem_inst/mem[77][3] ), .CK(clk), .Q(\xmem_data[77][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][3]  ( .D(\xmem_inst/mem[75][3] ), .CK(clk), .Q(\xmem_data[75][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][3]  ( .D(\xmem_inst/mem[73][3] ), .CK(clk), .Q(\xmem_data[73][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][6]  ( .D(\xmem_inst/mem[9][6] ), .CK(clk), 
        .Q(\xmem_data[9][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][4]  ( .D(\xmem_inst/mem[1][4] ), .CK(clk), 
        .Q(\xmem_data[1][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][0]  ( .D(\xmem_inst/mem[13][0] ), .CK(clk), .Q(\xmem_data[13][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][7]  ( .D(\xmem_inst/mem[127][7] ), .CK(
        clk), .Q(\xmem_data[127][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][7]  ( .D(\xmem_inst/mem[125][7] ), .CK(
        clk), .Q(\xmem_data[125][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][0]  ( .D(\xmem_inst/mem[93][0] ), .CK(clk), .Q(\xmem_data[93][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][7]  ( .D(\xmem_inst/mem[113][7] ), .CK(
        clk), .Q(\xmem_data[113][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][0]  ( .D(\xmem_inst/mem[61][0] ), .CK(clk), .Q(\xmem_data[61][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][4]  ( .D(\xmem_inst/mem[84][4] ), .CK(clk), .Q(\xmem_data[84][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][4]  ( .D(\xmem_inst/mem[92][4] ), .CK(clk), .Q(\xmem_data[92][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[22][5]  ( .D(\xmem_inst/mem[22][5] ), .CK(clk), .Q(\xmem_data[22][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][4]  ( .D(\xmem_inst/mem[70][4] ), .CK(clk), .Q(\xmem_data[70][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][4]  ( .D(\xmem_inst/mem[78][4] ), .CK(clk), .Q(\xmem_data[78][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][4]  ( .D(\xmem_inst/mem[80][4] ), .CK(clk), .Q(\xmem_data[80][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][4]  ( .D(\xmem_inst/mem[90][4] ), .CK(clk), .Q(\xmem_data[90][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][4]  ( .D(\xmem_inst/mem[76][4] ), .CK(clk), .Q(\xmem_data[76][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][4]  ( .D(\xmem_inst/mem[72][4] ), .CK(clk), .Q(\xmem_data[72][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][7]  ( .D(\xmem_inst/mem[2][7] ), .CK(clk), 
        .Q(\xmem_data[2][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][3]  ( .D(\xmem_inst/mem[69][3] ), .CK(clk), .Q(\xmem_data[69][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][3]  ( .D(\xmem_inst/mem[101][3] ), .CK(
        clk), .Q(\xmem_data[101][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][3]  ( .D(\xmem_inst/mem[127][3] ), .CK(
        clk), .Q(\xmem_data[127][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][5]  ( .D(\xmem_inst/mem[87][5] ), .CK(clk), .Q(\xmem_data[87][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][0]  ( .D(\xmem_inst/mem[15][0] ), .CK(clk), .Q(\xmem_data[15][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][5]  ( .D(\xmem_inst/mem[6][5] ), .CK(clk), 
        .Q(\xmem_data[6][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][2]  ( .D(\xmem_inst/mem[86][2] ), .CK(clk), .Q(\xmem_data[86][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][2]  ( .D(\xmem_inst/mem[118][2] ), .CK(
        clk), .Q(\xmem_data[118][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][3]  ( .D(\xmem_inst/mem[67][3] ), .CK(clk), .Q(\xmem_data[67][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][3]  ( .D(\xmem_inst/mem[99][3] ), .CK(clk), .Q(\xmem_data[99][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][3]  ( .D(\xmem_inst/mem[19][3] ), .CK(clk), .Q(\xmem_data[19][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][7]  ( .D(\xmem_inst/mem[93][7] ), .CK(clk), .Q(\xmem_data[93][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][7]  ( .D(\xmem_inst/mem[81][7] ), .CK(clk), .Q(\xmem_data[81][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][7]  ( .D(\xmem_inst/mem[79][7] ), .CK(clk), .Q(\xmem_data[79][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][7]  ( .D(\xmem_inst/mem[77][7] ), .CK(clk), .Q(\xmem_data[77][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][7]  ( .D(\xmem_inst/mem[71][7] ), .CK(clk), .Q(\xmem_data[71][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][5]  ( .D(\xmem_inst/mem[9][5] ), .CK(clk), 
        .Q(\xmem_data[9][5] ), .QN(n39031) );
  DFF_X2 \xmem_inst/data_out_reg[117][5]  ( .D(\xmem_inst/mem[117][5] ), .CK(
        clk), .Q(\xmem_data[117][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][5]  ( .D(\xmem_inst/mem[113][5] ), .CK(
        clk), .Q(\xmem_data[113][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][4]  ( .D(\xmem_inst/mem[25][4] ), .CK(clk), .Q(\xmem_data[25][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][3]  ( .D(\xmem_inst/mem[59][3] ), .CK(clk), .Q(\xmem_data[59][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][3]  ( .D(\xmem_inst/mem[93][3] ), .CK(clk), .Q(\xmem_data[93][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][3]  ( .D(\xmem_inst/mem[91][3] ), .CK(clk), .Q(\xmem_data[91][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][5]  ( .D(\xmem_inst/mem[91][5] ), .CK(clk), .Q(\xmem_data[91][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][3]  ( .D(\xmem_inst/mem[113][3] ), .CK(
        clk), .Q(\xmem_data[113][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][5]  ( .D(\xmem_inst/mem[85][5] ), .CK(clk), .Q(\xmem_data[85][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][5]  ( .D(\xmem_inst/mem[81][5] ), .CK(clk), .Q(\xmem_data[81][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[22][7]  ( .D(\xmem_inst/mem[22][7] ), .CK(clk), .Q(\xmem_data[22][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][2]  ( .D(\xmem_inst/mem[15][2] ), .CK(clk), .Q(\xmem_data[15][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][2]  ( .D(\xmem_inst/mem[13][2] ), .CK(clk), .Q(\xmem_data[13][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][3]  ( .D(\xmem_inst/mem[95][3] ), .CK(clk), .Q(\xmem_data[95][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][2]  ( .D(\xmem_inst/mem[29][2] ), .CK(clk), .Q(\xmem_data[29][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][4]  ( .D(\xmem_inst/mem[29][4] ), .CK(clk), .Q(\xmem_data[29][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][5]  ( .D(\xmem_inst/mem[89][5] ), .CK(clk), .Q(\xmem_data[89][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][3]  ( .D(\xmem_inst/mem[53][3] ), .CK(clk), .Q(\xmem_data[53][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][0]  ( .D(\xmem_inst/mem[2][0] ), .CK(clk), 
        .Q(\xmem_data[2][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][2]  ( .D(\xmem_inst/mem[90][2] ), .CK(clk), .Q(\xmem_data[90][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][2]  ( .D(\xmem_inst/mem[80][2] ), .CK(clk), .Q(\xmem_data[80][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][2]  ( .D(\xmem_inst/mem[84][2] ), .CK(clk), .Q(\xmem_data[84][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][0]  ( .D(\xmem_inst/mem[18][0] ), .CK(clk), .Q(\xmem_data[18][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][7]  ( .D(\xmem_inst/mem[20][7] ), .CK(clk), .Q(\xmem_data[20][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][4]  ( .D(\xmem_inst/mem[18][4] ), .CK(clk), .Q(\xmem_data[18][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][2]  ( .D(\xmem_inst/mem[8][2] ), .CK(clk), 
        .Q(\xmem_data[8][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][4]  ( .D(\xmem_inst/mem[16][4] ), .CK(clk), .Q(\xmem_data[16][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][7]  ( .D(\xmem_inst/mem[24][7] ), .CK(clk), .Q(\xmem_data[24][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[22][4]  ( .D(\xmem_inst/mem[22][4] ), .CK(clk), .Q(\xmem_data[22][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][7]  ( .D(\xmem_inst/mem[84][7] ), .CK(clk), .Q(\xmem_data[84][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][3]  ( .D(\xmem_inst/mem[30][3] ), .CK(clk), .Q(\xmem_data[30][3] ), .QN(n39013) );
  DFF_X2 \xmem_inst/data_out_reg[26][2]  ( .D(\xmem_inst/mem[26][2] ), .CK(clk), .Q(\xmem_data[26][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][2]  ( .D(\xmem_inst/mem[24][2] ), .CK(clk), .Q(\xmem_data[24][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][2]  ( .D(\xmem_inst/mem[56][2] ), .CK(clk), .Q(\xmem_data[56][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][2]  ( .D(\xmem_inst/mem[78][2] ), .CK(clk), .Q(\xmem_data[78][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][2]  ( .D(\xmem_inst/mem[60][2] ), .CK(clk), .Q(\xmem_data[60][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][2]  ( .D(\xmem_inst/mem[46][2] ), .CK(clk), .Q(\xmem_data[46][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][2]  ( .D(\xmem_inst/mem[92][2] ), .CK(clk), .Q(\xmem_data[92][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][2]  ( .D(\xmem_inst/mem[122][2] ), .CK(
        clk), .Q(\xmem_data[122][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][2]  ( .D(\xmem_inst/mem[126][2] ), .CK(
        clk), .Q(\xmem_data[126][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][2]  ( .D(\xmem_inst/mem[94][2] ), .CK(clk), .Q(\xmem_data[94][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][2]  ( .D(\xmem_inst/mem[66][2] ), .CK(clk), .Q(\xmem_data[66][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][2]  ( .D(\xmem_inst/mem[106][2] ), .CK(
        clk), .Q(\xmem_data[106][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][7]  ( .D(\xmem_inst/mem[16][7] ), .CK(clk), .Q(\xmem_data[16][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][2]  ( .D(\xmem_inst/mem[58][2] ), .CK(clk), .Q(\xmem_data[58][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][2]  ( .D(\xmem_inst/mem[54][2] ), .CK(clk), .Q(\xmem_data[54][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][2]  ( .D(\xmem_inst/mem[52][2] ), .CK(clk), .Q(\xmem_data[52][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][2]  ( .D(\xmem_inst/mem[48][2] ), .CK(clk), .Q(\xmem_data[48][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][2]  ( .D(\xmem_inst/mem[44][2] ), .CK(clk), .Q(\xmem_data[44][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][2]  ( .D(\xmem_inst/mem[42][2] ), .CK(clk), .Q(\xmem_data[42][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][2]  ( .D(\xmem_inst/mem[40][2] ), .CK(clk), .Q(\xmem_data[40][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][2]  ( .D(\xmem_inst/mem[38][2] ), .CK(clk), .Q(\xmem_data[38][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][2]  ( .D(\xmem_inst/mem[32][2] ), .CK(clk), .Q(\xmem_data[32][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][2]  ( .D(\xmem_inst/mem[74][2] ), .CK(clk), .Q(\xmem_data[74][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][2]  ( .D(\xmem_inst/mem[72][2] ), .CK(clk), .Q(\xmem_data[72][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][2]  ( .D(\xmem_inst/mem[68][2] ), .CK(clk), .Q(\xmem_data[68][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][2]  ( .D(\xmem_inst/mem[124][2] ), .CK(
        clk), .Q(\xmem_data[124][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][2]  ( .D(\xmem_inst/mem[112][2] ), .CK(
        clk), .Q(\xmem_data[112][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][2]  ( .D(\xmem_inst/mem[110][2] ), .CK(
        clk), .Q(\xmem_data[110][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][2]  ( .D(\xmem_inst/mem[108][2] ), .CK(
        clk), .Q(\xmem_data[108][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][2]  ( .D(\xmem_inst/mem[104][2] ), .CK(
        clk), .Q(\xmem_data[104][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][2]  ( .D(\xmem_inst/mem[100][2] ), .CK(
        clk), .Q(\xmem_data[100][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][2]  ( .D(\xmem_inst/mem[98][2] ), .CK(clk), .Q(\xmem_data[98][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][7]  ( .D(\xmem_inst/mem[18][7] ), .CK(clk), .Q(\xmem_data[18][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][2]  ( .D(\xmem_inst/mem[116][2] ), .CK(
        clk), .Q(\xmem_data[116][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][5]  ( .D(\xmem_inst/mem[125][5] ), .CK(
        clk), .Q(\xmem_data[125][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][5]  ( .D(\xmem_inst/mem[123][5] ), .CK(
        clk), .Q(\xmem_data[123][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][5]  ( .D(\xmem_inst/mem[127][5] ), .CK(
        clk), .Q(\xmem_data[127][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][5]  ( .D(\xmem_inst/mem[12][5] ), .CK(clk), .Q(\xmem_data[12][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][5]  ( .D(\xmem_inst/mem[28][5] ), .CK(clk), .Q(\xmem_data[28][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][5]  ( .D(\xmem_inst/mem[78][5] ), .CK(clk), .Q(\xmem_data[78][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][5]  ( .D(\xmem_inst/mem[64][5] ), .CK(clk), .Q(\xmem_data[64][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][5]  ( .D(\xmem_inst/mem[76][5] ), .CK(clk), .Q(\xmem_data[76][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][6]  ( .D(\xmem_inst/mem[19][6] ), .CK(clk), .Q(\xmem_data[19][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][4]  ( .D(\xmem_inst/mem[30][4] ), .CK(clk), .Q(\xmem_data[30][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][5]  ( .D(\xmem_inst/mem[74][5] ), .CK(clk), .Q(\xmem_data[74][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][5]  ( .D(\xmem_inst/mem[72][5] ), .CK(clk), .Q(\xmem_data[72][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][5]  ( .D(\xmem_inst/mem[108][5] ), .CK(
        clk), .Q(\xmem_data[108][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][5]  ( .D(\xmem_inst/mem[106][5] ), .CK(
        clk), .Q(\xmem_data[106][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][5]  ( .D(\xmem_inst/mem[104][5] ), .CK(
        clk), .Q(\xmem_data[104][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][2]  ( .D(\xmem_inst/mem[2][2] ), .CK(clk), 
        .Q(\xmem_data[2][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][5]  ( .D(\xmem_inst/mem[100][5] ), .CK(
        clk), .Q(\xmem_data[100][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][5]  ( .D(\xmem_inst/mem[98][5] ), .CK(clk), .Q(\xmem_data[98][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][4]  ( .D(\xmem_inst/mem[15][4] ), .CK(clk), .Q(\xmem_data[15][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][6]  ( .D(\xmem_inst/mem[15][6] ), .CK(clk), .Q(\xmem_data[15][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][6]  ( .D(\xmem_inst/mem[3][6] ), .CK(clk), 
        .Q(\xmem_data[3][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][6]  ( .D(\xmem_inst/mem[12][6] ), .CK(clk), .Q(\xmem_data[12][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][6]  ( .D(\xmem_inst/mem[0][6] ), .CK(clk), 
        .Q(\xmem_data[0][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][7]  ( .D(\xmem_inst/mem[37][7] ), .CK(clk), .Q(\xmem_data[37][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][5]  ( .D(\xmem_inst/mem[39][5] ), .CK(clk), .Q(\xmem_data[39][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][6]  ( .D(\xmem_inst/mem[77][6] ), .CK(clk), .Q(\xmem_data[77][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][6]  ( .D(\xmem_inst/mem[107][6] ), .CK(
        clk), .Q(\xmem_data[107][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][7]  ( .D(\xmem_inst/mem[39][7] ), .CK(clk), .Q(\xmem_data[39][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][6]  ( .D(\xmem_inst/mem[91][6] ), .CK(clk), .Q(\xmem_data[91][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][6]  ( .D(\xmem_inst/mem[85][6] ), .CK(clk), .Q(\xmem_data[85][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][6]  ( .D(\xmem_inst/mem[23][6] ), .CK(clk), .Q(\xmem_data[23][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][7]  ( .D(\xmem_inst/mem[11][7] ), .CK(clk), .Q(\xmem_data[11][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][6]  ( .D(\xmem_inst/mem[20][6] ), .CK(clk), .Q(\xmem_data[20][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][0]  ( .D(\xmem_inst/mem[9][0] ), .CK(clk), 
        .Q(\xmem_data[9][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][5]  ( .D(\xmem_inst/mem[47][5] ), .CK(clk), .Q(\xmem_data[47][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][7]  ( .D(\xmem_inst/mem[61][7] ), .CK(clk), .Q(\xmem_data[61][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][7]  ( .D(\xmem_inst/mem[57][7] ), .CK(clk), .Q(\xmem_data[57][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][7]  ( .D(\xmem_inst/mem[53][7] ), .CK(clk), .Q(\xmem_data[53][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][7]  ( .D(\xmem_inst/mem[51][7] ), .CK(clk), .Q(\xmem_data[51][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][7]  ( .D(\xmem_inst/mem[49][7] ), .CK(clk), .Q(\xmem_data[49][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][7]  ( .D(\xmem_inst/mem[47][7] ), .CK(clk), .Q(\xmem_data[47][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][7]  ( .D(\xmem_inst/mem[1][7] ), .CK(clk), 
        .Q(\xmem_data[1][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][5]  ( .D(\xmem_inst/mem[57][5] ), .CK(clk), .Q(\xmem_data[57][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][5]  ( .D(\xmem_inst/mem[33][5] ), .CK(clk), .Q(\xmem_data[33][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][5]  ( .D(\xmem_inst/mem[53][5] ), .CK(clk), .Q(\xmem_data[53][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][5]  ( .D(\xmem_inst/mem[61][5] ), .CK(clk), .Q(\xmem_data[61][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][5]  ( .D(\xmem_inst/mem[59][5] ), .CK(clk), .Q(\xmem_data[59][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][6]  ( .D(\xmem_inst/mem[93][6] ), .CK(clk), .Q(\xmem_data[93][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][6]  ( .D(\xmem_inst/mem[89][6] ), .CK(clk), .Q(\xmem_data[89][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][6]  ( .D(\xmem_inst/mem[81][6] ), .CK(clk), .Q(\xmem_data[81][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][6]  ( .D(\xmem_inst/mem[71][6] ), .CK(clk), .Q(\xmem_data[71][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][6]  ( .D(\xmem_inst/mem[65][6] ), .CK(clk), .Q(\xmem_data[65][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][6]  ( .D(\xmem_inst/mem[119][6] ), .CK(
        clk), .Q(\xmem_data[119][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][6]  ( .D(\xmem_inst/mem[113][6] ), .CK(
        clk), .Q(\xmem_data[113][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][6]  ( .D(\xmem_inst/mem[109][6] ), .CK(
        clk), .Q(\xmem_data[109][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][6]  ( .D(\xmem_inst/mem[101][6] ), .CK(
        clk), .Q(\xmem_data[101][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][6]  ( .D(\xmem_inst/mem[99][6] ), .CK(clk), .Q(\xmem_data[99][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][6]  ( .D(\xmem_inst/mem[61][6] ), .CK(clk), .Q(\xmem_data[61][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][6]  ( .D(\xmem_inst/mem[57][6] ), .CK(clk), .Q(\xmem_data[57][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][6]  ( .D(\xmem_inst/mem[49][6] ), .CK(clk), .Q(\xmem_data[49][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][6]  ( .D(\xmem_inst/mem[47][6] ), .CK(clk), .Q(\xmem_data[47][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][6]  ( .D(\xmem_inst/mem[45][6] ), .CK(clk), .Q(\xmem_data[45][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][6]  ( .D(\xmem_inst/mem[39][6] ), .CK(clk), .Q(\xmem_data[39][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][6]  ( .D(\xmem_inst/mem[33][6] ), .CK(clk), .Q(\xmem_data[33][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][5]  ( .D(\xmem_inst/mem[45][5] ), .CK(clk), .Q(\xmem_data[45][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][4]  ( .D(\xmem_inst/mem[9][4] ), .CK(clk), 
        .Q(\xmem_data[9][4] ), .QN(n39038) );
  DFF_X2 \xmem_inst/data_out_reg[49][5]  ( .D(\xmem_inst/mem[49][5] ), .CK(clk), .Q(\xmem_data[49][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][6]  ( .D(\xmem_inst/mem[25][6] ), .CK(clk), .Q(\xmem_data[25][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][6]  ( .D(\xmem_inst/mem[123][6] ), .CK(
        clk), .Q(\xmem_data[123][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][6]  ( .D(\xmem_inst/mem[27][6] ), .CK(clk), .Q(\xmem_data[27][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][6]  ( .D(\xmem_inst/mem[53][6] ), .CK(clk), .Q(\xmem_data[53][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][7]  ( .D(\xmem_inst/mem[59][7] ), .CK(clk), .Q(\xmem_data[59][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][6]  ( .D(\xmem_inst/mem[117][6] ), .CK(
        clk), .Q(\xmem_data[117][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][6]  ( .D(\xmem_inst/mem[17][6] ), .CK(clk), .Q(\xmem_data[17][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][6]  ( .D(\xmem_inst/mem[29][6] ), .CK(clk), .Q(\xmem_data[29][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][7]  ( .D(\xmem_inst/mem[63][7] ), .CK(clk), .Q(\xmem_data[63][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][6]  ( .D(\xmem_inst/mem[30][6] ), .CK(clk), .Q(\xmem_data[30][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][6]  ( .D(\xmem_inst/mem[6][6] ), .CK(clk), 
        .Q(\xmem_data[6][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][6]  ( .D(\xmem_inst/mem[105][6] ), .CK(
        clk), .Q(\xmem_data[105][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][6]  ( .D(\xmem_inst/mem[59][6] ), .CK(clk), .Q(\xmem_data[59][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][3]  ( .D(\xmem_inst/mem[21][3] ), .CK(clk), .Q(\xmem_data[21][3] ), .QN(n39008) );
  DFF_X2 \xmem_inst/data_out_reg[21][5]  ( .D(\xmem_inst/mem[21][5] ), .CK(clk), .Q(\xmem_data[21][5] ), .QN(n39004) );
  DFF_X2 \xmem_inst/data_out_reg[43][1]  ( .D(\xmem_inst/mem[43][1] ), .CK(clk), .Q(\xmem_data[43][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][3]  ( .D(\xmem_inst/mem[71][3] ), .CK(clk), .Q(\xmem_data[71][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][5]  ( .D(\xmem_inst/mem[31][5] ), .CK(clk), .Q(\xmem_data[31][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][1]  ( .D(\xmem_inst/mem[37][1] ), .CK(clk), .Q(\xmem_data[37][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][4]  ( .D(\xmem_inst/mem[46][4] ), .CK(clk), .Q(\xmem_data[46][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][1]  ( .D(\xmem_inst/mem[100][1] ), .CK(
        clk), .Q(\xmem_data[100][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][4]  ( .D(\xmem_inst/mem[42][4] ), .CK(clk), .Q(\xmem_data[42][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][1]  ( .D(\xmem_inst/mem[103][1] ), .CK(
        clk), .Q(\xmem_data[103][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][1]  ( .D(\xmem_inst/mem[97][1] ), .CK(clk), .Q(\xmem_data[97][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][1]  ( .D(\xmem_inst/mem[71][1] ), .CK(clk), .Q(\xmem_data[71][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][1]  ( .D(\xmem_inst/mem[65][1] ), .CK(clk), .Q(\xmem_data[65][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][1]  ( .D(\xmem_inst/mem[3][1] ), .CK(clk), 
        .Q(\xmem_data[3][1] ), .QN(n39029) );
  DFF_X2 \xmem_inst/data_out_reg[47][1]  ( .D(\xmem_inst/mem[47][1] ), .CK(clk), .Q(\xmem_data[47][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][0]  ( .D(\xmem_inst/mem[25][0] ), .CK(clk), .Q(\xmem_data[25][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][3]  ( .D(\xmem_inst/mem[65][3] ), .CK(clk), .Q(\xmem_data[65][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][3]  ( .D(\xmem_inst/mem[97][3] ), .CK(clk), .Q(\xmem_data[97][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][3]  ( .D(\xmem_inst/mem[63][3] ), .CK(clk), .Q(\xmem_data[63][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][3]  ( .D(\xmem_inst/mem[9][3] ), .CK(clk), 
        .Q(\xmem_data[9][3] ), .QN(n39034) );
  DFF_X2 \xmem_inst/data_out_reg[37][4]  ( .D(\xmem_inst/mem[37][4] ), .CK(clk), .Q(\xmem_data[37][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][4]  ( .D(\xmem_inst/mem[63][4] ), .CK(clk), .Q(\xmem_data[63][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][4]  ( .D(\xmem_inst/mem[97][4] ), .CK(clk), .Q(\xmem_data[97][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][5]  ( .D(\xmem_inst/mem[103][5] ), .CK(
        clk), .Q(\xmem_data[103][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][1]  ( .D(\xmem_inst/mem[21][1] ), .CK(clk), .Q(\xmem_data[21][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][1]  ( .D(\xmem_inst/mem[29][1] ), .CK(clk), .Q(\xmem_data[29][1] ), .QN(n39028) );
  DFF_X2 \xmem_inst/data_out_reg[63][1]  ( .D(\xmem_inst/mem[63][1] ), .CK(clk), .Q(\xmem_data[63][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][2]  ( .D(\xmem_inst/mem[16][2] ), .CK(clk), .Q(\xmem_data[16][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][1]  ( .D(\xmem_inst/mem[94][1] ), .CK(clk), .Q(\xmem_data[94][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][1]  ( .D(\xmem_inst/mem[24][1] ), .CK(clk), .Q(\xmem_data[24][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][1]  ( .D(\xmem_inst/mem[56][1] ), .CK(clk), .Q(\xmem_data[56][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][1]  ( .D(\xmem_inst/mem[80][1] ), .CK(clk), .Q(\xmem_data[80][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][4]  ( .D(\xmem_inst/mem[48][4] ), .CK(clk), .Q(\xmem_data[48][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][1]  ( .D(\xmem_inst/mem[92][1] ), .CK(clk), .Q(\xmem_data[92][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][1]  ( .D(\xmem_inst/mem[126][1] ), .CK(
        clk), .Q(\xmem_data[126][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][1]  ( .D(\xmem_inst/mem[124][1] ), .CK(
        clk), .Q(\xmem_data[124][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][1]  ( .D(\xmem_inst/mem[98][1] ), .CK(clk), .Q(\xmem_data[98][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][1]  ( .D(\xmem_inst/mem[106][1] ), .CK(
        clk), .Q(\xmem_data[106][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][1]  ( .D(\xmem_inst/mem[68][1] ), .CK(clk), .Q(\xmem_data[68][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][1]  ( .D(\xmem_inst/mem[66][1] ), .CK(clk), .Q(\xmem_data[66][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][1]  ( .D(\xmem_inst/mem[26][1] ), .CK(clk), .Q(\xmem_data[26][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][1]  ( .D(\xmem_inst/mem[8][1] ), .CK(clk), 
        .Q(\xmem_data[8][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][1]  ( .D(\xmem_inst/mem[58][1] ), .CK(clk), .Q(\xmem_data[58][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][1]  ( .D(\xmem_inst/mem[48][1] ), .CK(clk), .Q(\xmem_data[48][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][1]  ( .D(\xmem_inst/mem[40][1] ), .CK(clk), .Q(\xmem_data[40][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][3]  ( .D(\xmem_inst/mem[80][3] ), .CK(clk), .Q(\xmem_data[80][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][3]  ( .D(\xmem_inst/mem[48][3] ), .CK(clk), .Q(\xmem_data[48][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][3]  ( .D(\xmem_inst/mem[46][3] ), .CK(clk), .Q(\xmem_data[46][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][3]  ( .D(\xmem_inst/mem[40][3] ), .CK(clk), .Q(\xmem_data[40][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][3]  ( .D(\xmem_inst/mem[38][3] ), .CK(clk), .Q(\xmem_data[38][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][3]  ( .D(\xmem_inst/mem[24][3] ), .CK(clk), .Q(\xmem_data[24][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][3]  ( .D(\xmem_inst/mem[28][3] ), .CK(clk), .Q(\xmem_data[28][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][4]  ( .D(\xmem_inst/mem[38][4] ), .CK(clk), .Q(\xmem_data[38][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][4]  ( .D(\xmem_inst/mem[58][4] ), .CK(clk), .Q(\xmem_data[58][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][4]  ( .D(\xmem_inst/mem[52][4] ), .CK(clk), .Q(\xmem_data[52][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][4]  ( .D(\xmem_inst/mem[100][4] ), .CK(
        clk), .Q(\xmem_data[100][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][4]  ( .D(\xmem_inst/mem[98][4] ), .CK(clk), .Q(\xmem_data[98][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][4]  ( .D(\xmem_inst/mem[126][4] ), .CK(
        clk), .Q(\xmem_data[126][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][4]  ( .D(\xmem_inst/mem[124][4] ), .CK(
        clk), .Q(\xmem_data[124][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][4]  ( .D(\xmem_inst/mem[106][4] ), .CK(
        clk), .Q(\xmem_data[106][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][4]  ( .D(\xmem_inst/mem[104][4] ), .CK(
        clk), .Q(\xmem_data[104][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][5]  ( .D(\xmem_inst/mem[70][5] ), .CK(clk), .Q(\xmem_data[70][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][5]  ( .D(\xmem_inst/mem[26][5] ), .CK(clk), .Q(\xmem_data[26][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][0]  ( .D(\xmem_inst/mem[21][0] ), .CK(clk), .Q(\xmem_data[21][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][1]  ( .D(\xmem_inst/mem[112][1] ), .CK(
        clk), .Q(\xmem_data[112][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][0]  ( .D(\xmem_inst/mem[102][0] ), .CK(
        clk), .Q(\xmem_data[102][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][3]  ( .D(\xmem_inst/mem[15][3] ), .CK(clk), .Q(\xmem_data[15][3] ), .QN(n39021) );
  DFF_X2 \xmem_inst/data_out_reg[38][1]  ( .D(\xmem_inst/mem[38][1] ), .CK(clk), .Q(\xmem_data[38][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][0]  ( .D(\xmem_inst/mem[0][0] ), .CK(clk), 
        .Q(\xmem_data[0][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][7]  ( .D(\xmem_inst/mem[9][7] ), .CK(clk), 
        .Q(\xmem_data[9][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][7]  ( .D(\xmem_inst/mem[15][7] ), .CK(clk), .Q(\xmem_data[15][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][5]  ( .D(\xmem_inst/mem[16][5] ), .CK(clk), .Q(\xmem_data[16][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][0]  ( .D(\xmem_inst/mem[101][0] ), .CK(
        clk), .Q(\xmem_data[101][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][0]  ( .D(\xmem_inst/mem[97][0] ), .CK(clk), .Q(\xmem_data[97][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][0]  ( .D(\xmem_inst/mem[71][0] ), .CK(clk), .Q(\xmem_data[71][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][0]  ( .D(\xmem_inst/mem[65][0] ), .CK(clk), .Q(\xmem_data[65][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][7]  ( .D(\xmem_inst/mem[103][7] ), .CK(
        clk), .Q(\xmem_data[103][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][7]  ( .D(\xmem_inst/mem[97][7] ), .CK(clk), .Q(\xmem_data[97][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][5]  ( .D(\xmem_inst/mem[25][5] ), .CK(clk), .Q(\xmem_data[25][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][0]  ( .D(\xmem_inst/mem[43][0] ), .CK(clk), .Q(\xmem_data[43][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][0]  ( .D(\xmem_inst/mem[37][0] ), .CK(clk), .Q(\xmem_data[37][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][0]  ( .D(\xmem_inst/mem[35][0] ), .CK(clk), .Q(\xmem_data[35][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][0]  ( .D(\xmem_inst/mem[59][0] ), .CK(clk), .Q(\xmem_data[59][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][0]  ( .D(\xmem_inst/mem[63][0] ), .CK(clk), .Q(\xmem_data[63][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][7]  ( .D(\xmem_inst/mem[112][7] ), .CK(
        clk), .Q(\xmem_data[112][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][2]  ( .D(\xmem_inst/mem[1][2] ), .CK(clk), 
        .Q(\xmem_data[1][2] ), .QN(n39036) );
  DFF_X2 \xmem_inst/data_out_reg[126][7]  ( .D(\xmem_inst/mem[126][7] ), .CK(
        clk), .Q(\xmem_data[126][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][0]  ( .D(\xmem_inst/mem[38][0] ), .CK(clk), .Q(\xmem_data[38][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][7]  ( .D(\xmem_inst/mem[106][7] ), .CK(
        clk), .Q(\xmem_data[106][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][7]  ( .D(\xmem_inst/mem[104][7] ), .CK(
        clk), .Q(\xmem_data[104][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][3]  ( .D(\xmem_inst/mem[104][3] ), .CK(
        clk), .Q(\xmem_data[104][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][0]  ( .D(\xmem_inst/mem[46][0] ), .CK(clk), .Q(\xmem_data[46][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][0]  ( .D(\xmem_inst/mem[54][0] ), .CK(clk), .Q(\xmem_data[54][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][0]  ( .D(\xmem_inst/mem[52][0] ), .CK(clk), .Q(\xmem_data[52][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][0]  ( .D(\xmem_inst/mem[48][0] ), .CK(clk), .Q(\xmem_data[48][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][0]  ( .D(\xmem_inst/mem[56][0] ), .CK(clk), .Q(\xmem_data[56][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][4]  ( .D(\xmem_inst/mem[66][4] ), .CK(clk), .Q(\xmem_data[66][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][4]  ( .D(\xmem_inst/mem[68][4] ), .CK(clk), .Q(\xmem_data[68][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][4]  ( .D(\xmem_inst/mem[94][4] ), .CK(clk), .Q(\xmem_data[94][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][3]  ( .D(\xmem_inst/mem[74][3] ), .CK(clk), .Q(\xmem_data[74][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][3]  ( .D(\xmem_inst/mem[72][3] ), .CK(clk), .Q(\xmem_data[72][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][7]  ( .D(\xmem_inst/mem[124][7] ), .CK(
        clk), .Q(\xmem_data[124][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][3]  ( .D(\xmem_inst/mem[37][3] ), .CK(clk), .Q(\xmem_data[37][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][4]  ( .D(\xmem_inst/mem[71][4] ), .CK(clk), .Q(\xmem_data[71][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][4]  ( .D(\xmem_inst/mem[35][4] ), .CK(clk), .Q(\xmem_data[35][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][2]  ( .D(\xmem_inst/mem[27][2] ), .CK(clk), .Q(\xmem_data[27][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][7]  ( .D(\xmem_inst/mem[87][7] ), .CK(clk), .Q(\xmem_data[87][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][4]  ( .D(\xmem_inst/mem[79][4] ), .CK(clk), .Q(\xmem_data[79][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][2]  ( .D(\xmem_inst/mem[31][2] ), .CK(clk), .Q(\xmem_data[31][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][7]  ( .D(\xmem_inst/mem[95][7] ), .CK(clk), .Q(\xmem_data[95][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][7]  ( .D(\xmem_inst/mem[91][7] ), .CK(clk), .Q(\xmem_data[91][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][7]  ( .D(\xmem_inst/mem[89][7] ), .CK(clk), .Q(\xmem_data[89][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][7]  ( .D(\xmem_inst/mem[75][7] ), .CK(clk), .Q(\xmem_data[75][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][7]  ( .D(\xmem_inst/mem[69][7] ), .CK(clk), .Q(\xmem_data[69][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][4]  ( .D(\xmem_inst/mem[81][4] ), .CK(clk), .Q(\xmem_data[81][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][4]  ( .D(\xmem_inst/mem[91][4] ), .CK(clk), .Q(\xmem_data[91][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][3]  ( .D(\xmem_inst/mem[123][3] ), .CK(
        clk), .Q(\xmem_data[123][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][0]  ( .D(\xmem_inst/mem[29][0] ), .CK(clk), .Q(\xmem_data[29][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][5]  ( .D(\xmem_inst/mem[3][5] ), .CK(clk), 
        .Q(\xmem_data[3][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][2]  ( .D(\xmem_inst/mem[3][2] ), .CK(clk), 
        .Q(\xmem_data[3][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][3]  ( .D(\xmem_inst/mem[2][3] ), .CK(clk), 
        .Q(\xmem_data[2][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][4]  ( .D(\xmem_inst/mem[85][4] ), .CK(clk), .Q(\xmem_data[85][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][5]  ( .D(\xmem_inst/mem[95][5] ), .CK(clk), .Q(\xmem_data[95][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[7][5]  ( .D(\xmem_inst/mem[7][5] ), .CK(clk), 
        .Q(\xmem_data[7][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][3]  ( .D(\xmem_inst/mem[51][3] ), .CK(clk), .Q(\xmem_data[51][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][2]  ( .D(\xmem_inst/mem[35][2] ), .CK(clk), .Q(\xmem_data[35][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][5]  ( .D(\xmem_inst/mem[8][5] ), .CK(clk), 
        .Q(\xmem_data[8][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][0]  ( .D(\xmem_inst/mem[126][0] ), .CK(
        clk), .Q(\xmem_data[126][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][0]  ( .D(\xmem_inst/mem[94][0] ), .CK(clk), .Q(\xmem_data[94][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][3]  ( .D(\xmem_inst/mem[94][3] ), .CK(clk), .Q(\xmem_data[94][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][0]  ( .D(\xmem_inst/mem[92][0] ), .CK(clk), .Q(\xmem_data[92][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][3]  ( .D(\xmem_inst/mem[126][3] ), .CK(
        clk), .Q(\xmem_data[126][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][7]  ( .D(\xmem_inst/mem[30][7] ), .CK(clk), .Q(\xmem_data[30][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][2]  ( .D(\xmem_inst/mem[28][2] ), .CK(clk), .Q(\xmem_data[28][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][3]  ( .D(\xmem_inst/mem[112][3] ), .CK(
        clk), .Q(\xmem_data[112][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][3]  ( .D(\xmem_inst/mem[90][3] ), .CK(clk), .Q(\xmem_data[90][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][3]  ( .D(\xmem_inst/mem[100][3] ), .CK(
        clk), .Q(\xmem_data[100][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][0]  ( .D(\xmem_inst/mem[112][0] ), .CK(
        clk), .Q(\xmem_data[112][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][0]  ( .D(\xmem_inst/mem[106][0] ), .CK(
        clk), .Q(\xmem_data[106][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][0]  ( .D(\xmem_inst/mem[104][0] ), .CK(
        clk), .Q(\xmem_data[104][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][0]  ( .D(\xmem_inst/mem[80][0] ), .CK(clk), .Q(\xmem_data[80][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][0]  ( .D(\xmem_inst/mem[74][0] ), .CK(clk), .Q(\xmem_data[74][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][0]  ( .D(\xmem_inst/mem[72][0] ), .CK(clk), .Q(\xmem_data[72][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][7]  ( .D(\xmem_inst/mem[80][7] ), .CK(clk), .Q(\xmem_data[80][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][7]  ( .D(\xmem_inst/mem[78][7] ), .CK(clk), .Q(\xmem_data[78][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][7]  ( .D(\xmem_inst/mem[70][7] ), .CK(clk), .Q(\xmem_data[70][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][7]  ( .D(\xmem_inst/mem[26][7] ), .CK(clk), .Q(\xmem_data[26][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][4]  ( .D(\xmem_inst/mem[56][4] ), .CK(clk), .Q(\xmem_data[56][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][3]  ( .D(\xmem_inst/mem[58][3] ), .CK(clk), .Q(\xmem_data[58][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][4]  ( .D(\xmem_inst/mem[20][4] ), .CK(clk), .Q(\xmem_data[20][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][3]  ( .D(\xmem_inst/mem[92][3] ), .CK(clk), .Q(\xmem_data[92][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][2]  ( .D(\xmem_inst/mem[6][2] ), .CK(clk), 
        .Q(\xmem_data[6][2] ), .QN(n39019) );
  DFF_X2 \xmem_inst/data_out_reg[64][2]  ( .D(\xmem_inst/mem[64][2] ), .CK(clk), .Q(\xmem_data[64][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][2]  ( .D(\xmem_inst/mem[36][2] ), .CK(clk), .Q(\xmem_data[36][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][2]  ( .D(\xmem_inst/mem[50][2] ), .CK(clk), .Q(\xmem_data[50][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][2]  ( .D(\xmem_inst/mem[102][2] ), .CK(
        clk), .Q(\xmem_data[102][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][2]  ( .D(\xmem_inst/mem[96][2] ), .CK(clk), .Q(\xmem_data[96][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][4]  ( .D(\xmem_inst/mem[26][4] ), .CK(clk), .Q(\xmem_data[26][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][7]  ( .D(\xmem_inst/mem[85][7] ), .CK(clk), .Q(\xmem_data[85][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[9][2]  ( .D(\xmem_inst/mem[9][2] ), .CK(clk), 
        .Q(\xmem_data[9][2] ), .QN(n39037) );
  DFF_X2 \xmem_inst/data_out_reg[52][3]  ( .D(\xmem_inst/mem[52][3] ), .CK(clk), .Q(\xmem_data[52][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][2]  ( .D(\xmem_inst/mem[14][2] ), .CK(clk), .Q(\xmem_data[14][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][5]  ( .D(\xmem_inst/mem[67][5] ), .CK(clk), .Q(\xmem_data[67][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][5]  ( .D(\xmem_inst/mem[29][5] ), .CK(clk), .Q(\xmem_data[29][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][5]  ( .D(\xmem_inst/mem[86][5] ), .CK(clk), .Q(\xmem_data[86][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][3]  ( .D(\xmem_inst/mem[16][3] ), .CK(clk), .Q(\xmem_data[16][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][4]  ( .D(\xmem_inst/mem[6][4] ), .CK(clk), 
        .Q(\xmem_data[6][4] ), .QN(n39032) );
  DFF_X2 \xmem_inst/data_out_reg[10][2]  ( .D(\xmem_inst/mem[10][2] ), .CK(clk), .Q(\xmem_data[10][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][5]  ( .D(\xmem_inst/mem[118][5] ), .CK(
        clk), .Q(\xmem_data[118][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][5]  ( .D(\xmem_inst/mem[126][5] ), .CK(
        clk), .Q(\xmem_data[126][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][5]  ( .D(\xmem_inst/mem[68][5] ), .CK(clk), .Q(\xmem_data[68][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[47][2]  ( .D(\xmem_inst/mem[47][2] ), .CK(clk), .Q(\xmem_data[47][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][2]  ( .D(\xmem_inst/mem[93][2] ), .CK(clk), .Q(\xmem_data[93][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][2]  ( .D(\xmem_inst/mem[69][2] ), .CK(clk), .Q(\xmem_data[69][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][2]  ( .D(\xmem_inst/mem[127][2] ), .CK(
        clk), .Q(\xmem_data[127][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][2]  ( .D(\xmem_inst/mem[53][2] ), .CK(clk), .Q(\xmem_data[53][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[59][2]  ( .D(\xmem_inst/mem[59][2] ), .CK(clk), .Q(\xmem_data[59][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][2]  ( .D(\xmem_inst/mem[55][2] ), .CK(clk), .Q(\xmem_data[55][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][2]  ( .D(\xmem_inst/mem[49][2] ), .CK(clk), .Q(\xmem_data[49][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][2]  ( .D(\xmem_inst/mem[43][2] ), .CK(clk), .Q(\xmem_data[43][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][2]  ( .D(\xmem_inst/mem[41][2] ), .CK(clk), .Q(\xmem_data[41][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[39][2]  ( .D(\xmem_inst/mem[39][2] ), .CK(clk), .Q(\xmem_data[39][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][2]  ( .D(\xmem_inst/mem[95][2] ), .CK(clk), .Q(\xmem_data[95][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][2]  ( .D(\xmem_inst/mem[75][2] ), .CK(clk), .Q(\xmem_data[75][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][2]  ( .D(\xmem_inst/mem[73][2] ), .CK(clk), .Q(\xmem_data[73][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][2]  ( .D(\xmem_inst/mem[67][2] ), .CK(clk), .Q(\xmem_data[67][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][2]  ( .D(\xmem_inst/mem[125][2] ), .CK(
        clk), .Q(\xmem_data[125][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[113][2]  ( .D(\xmem_inst/mem[113][2] ), .CK(
        clk), .Q(\xmem_data[113][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][2]  ( .D(\xmem_inst/mem[107][2] ), .CK(
        clk), .Q(\xmem_data[107][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][2]  ( .D(\xmem_inst/mem[105][2] ), .CK(
        clk), .Q(\xmem_data[105][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][2]  ( .D(\xmem_inst/mem[101][2] ), .CK(
        clk), .Q(\xmem_data[101][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][2]  ( .D(\xmem_inst/mem[99][2] ), .CK(clk), .Q(\xmem_data[99][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][2]  ( .D(\xmem_inst/mem[57][2] ), .CK(clk), .Q(\xmem_data[57][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][2]  ( .D(\xmem_inst/mem[117][2] ), .CK(
        clk), .Q(\xmem_data[117][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[81][2]  ( .D(\xmem_inst/mem[81][2] ), .CK(clk), .Q(\xmem_data[81][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][2]  ( .D(\xmem_inst/mem[87][2] ), .CK(clk), .Q(\xmem_data[87][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][2]  ( .D(\xmem_inst/mem[85][2] ), .CK(clk), .Q(\xmem_data[85][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][2]  ( .D(\xmem_inst/mem[119][2] ), .CK(
        clk), .Q(\xmem_data[119][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][5]  ( .D(\xmem_inst/mem[84][5] ), .CK(clk), .Q(\xmem_data[84][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][5]  ( .D(\xmem_inst/mem[88][5] ), .CK(clk), .Q(\xmem_data[88][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][0]  ( .D(\xmem_inst/mem[14][0] ), .CK(clk), .Q(\xmem_data[14][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][5]  ( .D(\xmem_inst/mem[112][5] ), .CK(
        clk), .Q(\xmem_data[112][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][5]  ( .D(\xmem_inst/mem[80][5] ), .CK(clk), .Q(\xmem_data[80][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][5]  ( .D(\xmem_inst/mem[90][5] ), .CK(clk), .Q(\xmem_data[90][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][5]  ( .D(\xmem_inst/mem[124][5] ), .CK(
        clk), .Q(\xmem_data[124][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][5]  ( .D(\xmem_inst/mem[122][5] ), .CK(
        clk), .Q(\xmem_data[122][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][2]  ( .D(\xmem_inst/mem[25][2] ), .CK(clk), .Q(\xmem_data[25][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][7]  ( .D(\xmem_inst/mem[17][7] ), .CK(clk), .Q(\xmem_data[17][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][7]  ( .D(\xmem_inst/mem[19][7] ), .CK(clk), .Q(\xmem_data[19][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][7]  ( .D(\xmem_inst/mem[21][7] ), .CK(clk), .Q(\xmem_data[21][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][4]  ( .D(\xmem_inst/mem[4][4] ), .CK(clk), 
        .Q(\xmem_data[4][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][6]  ( .D(\xmem_inst/mem[4][6] ), .CK(clk), 
        .Q(\xmem_data[4][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][7]  ( .D(\xmem_inst/mem[23][7] ), .CK(clk), .Q(\xmem_data[23][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][0]  ( .D(\xmem_inst/mem[3][0] ), .CK(clk), 
        .Q(\xmem_data[3][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][5]  ( .D(\xmem_inst/mem[79][5] ), .CK(clk), .Q(\xmem_data[79][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][6]  ( .D(\xmem_inst/mem[31][6] ), .CK(clk), .Q(\xmem_data[31][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][4]  ( .D(\xmem_inst/mem[8][4] ), .CK(clk), 
        .Q(\xmem_data[8][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][5]  ( .D(\xmem_inst/mem[96][5] ), .CK(clk), .Q(\xmem_data[96][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][5]  ( .D(\xmem_inst/mem[77][5] ), .CK(clk), .Q(\xmem_data[77][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][6]  ( .D(\xmem_inst/mem[95][6] ), .CK(clk), .Q(\xmem_data[95][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[127][6]  ( .D(\xmem_inst/mem[127][6] ), .CK(
        clk), .Q(\xmem_data[127][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][4]  ( .D(\xmem_inst/mem[11][4] ), .CK(clk), .Q(\xmem_data[11][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][5]  ( .D(\xmem_inst/mem[43][5] ), .CK(clk), .Q(\xmem_data[43][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][6]  ( .D(\xmem_inst/mem[21][6] ), .CK(clk), .Q(\xmem_data[21][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][4]  ( .D(\xmem_inst/mem[2][4] ), .CK(clk), 
        .Q(\xmem_data[2][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][7]  ( .D(\xmem_inst/mem[25][7] ), .CK(clk), .Q(\xmem_data[25][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][5]  ( .D(\xmem_inst/mem[41][5] ), .CK(clk), .Q(\xmem_data[41][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][7]  ( .D(\xmem_inst/mem[41][7] ), .CK(clk), .Q(\xmem_data[41][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][5]  ( .D(\xmem_inst/mem[63][5] ), .CK(clk), .Q(\xmem_data[63][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][5]  ( .D(\xmem_inst/mem[73][5] ), .CK(clk), .Q(\xmem_data[73][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][5]  ( .D(\xmem_inst/mem[101][5] ), .CK(
        clk), .Q(\xmem_data[101][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[99][5]  ( .D(\xmem_inst/mem[99][5] ), .CK(clk), .Q(\xmem_data[99][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[107][5]  ( .D(\xmem_inst/mem[107][5] ), .CK(
        clk), .Q(\xmem_data[107][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][5]  ( .D(\xmem_inst/mem[105][5] ), .CK(
        clk), .Q(\xmem_data[105][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][6]  ( .D(\xmem_inst/mem[83][6] ), .CK(clk), .Q(\xmem_data[83][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][6]  ( .D(\xmem_inst/mem[73][6] ), .CK(clk), .Q(\xmem_data[73][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][6]  ( .D(\xmem_inst/mem[103][6] ), .CK(
        clk), .Q(\xmem_data[103][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][6]  ( .D(\xmem_inst/mem[97][6] ), .CK(clk), .Q(\xmem_data[97][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][6]  ( .D(\xmem_inst/mem[63][6] ), .CK(clk), .Q(\xmem_data[63][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][6]  ( .D(\xmem_inst/mem[43][6] ), .CK(clk), .Q(\xmem_data[43][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][6]  ( .D(\xmem_inst/mem[41][6] ), .CK(clk), .Q(\xmem_data[41][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[29][7]  ( .D(\xmem_inst/mem[29][7] ), .CK(clk), .Q(\xmem_data[29][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][6]  ( .D(\xmem_inst/mem[125][6] ), .CK(
        clk), .Q(\xmem_data[125][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][5]  ( .D(\xmem_inst/mem[37][5] ), .CK(clk), .Q(\xmem_data[37][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][5]  ( .D(\xmem_inst/mem[75][5] ), .CK(clk), .Q(\xmem_data[75][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][6]  ( .D(\xmem_inst/mem[75][6] ), .CK(clk), .Q(\xmem_data[75][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][6]  ( .D(\xmem_inst/mem[69][6] ), .CK(clk), .Q(\xmem_data[69][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][7]  ( .D(\xmem_inst/mem[62][7] ), .CK(clk), .Q(\xmem_data[62][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][6]  ( .D(\xmem_inst/mem[2][6] ), .CK(clk), 
        .Q(\xmem_data[2][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][7]  ( .D(\xmem_inst/mem[38][7] ), .CK(clk), .Q(\xmem_data[38][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][6]  ( .D(\xmem_inst/mem[90][6] ), .CK(clk), .Q(\xmem_data[90][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][6]  ( .D(\xmem_inst/mem[84][6] ), .CK(clk), .Q(\xmem_data[84][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][6]  ( .D(\xmem_inst/mem[14][6] ), .CK(clk), .Q(\xmem_data[14][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][6]  ( .D(\xmem_inst/mem[78][6] ), .CK(clk), .Q(\xmem_data[78][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][6]  ( .D(\xmem_inst/mem[26][6] ), .CK(clk), .Q(\xmem_data[26][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][6]  ( .D(\xmem_inst/mem[52][6] ), .CK(clk), .Q(\xmem_data[52][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][6]  ( .D(\xmem_inst/mem[28][6] ), .CK(clk), .Q(\xmem_data[28][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][7]  ( .D(\xmem_inst/mem[58][7] ), .CK(clk), .Q(\xmem_data[58][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][0]  ( .D(\xmem_inst/mem[8][0] ), .CK(clk), 
        .Q(\xmem_data[8][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][5]  ( .D(\xmem_inst/mem[48][5] ), .CK(clk), .Q(\xmem_data[48][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][6]  ( .D(\xmem_inst/mem[24][6] ), .CK(clk), .Q(\xmem_data[24][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][7]  ( .D(\xmem_inst/mem[42][7] ), .CK(clk), .Q(\xmem_data[42][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][7]  ( .D(\xmem_inst/mem[36][7] ), .CK(clk), .Q(\xmem_data[36][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][6]  ( .D(\xmem_inst/mem[76][6] ), .CK(clk), .Q(\xmem_data[76][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][6]  ( .D(\xmem_inst/mem[106][6] ), .CK(
        clk), .Q(\xmem_data[106][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][5]  ( .D(\xmem_inst/mem[46][5] ), .CK(clk), .Q(\xmem_data[46][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][5]  ( .D(\xmem_inst/mem[38][5] ), .CK(clk), .Q(\xmem_data[38][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][5]  ( .D(\xmem_inst/mem[44][5] ), .CK(clk), .Q(\xmem_data[44][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][5]  ( .D(\xmem_inst/mem[58][5] ), .CK(clk), .Q(\xmem_data[58][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][5]  ( .D(\xmem_inst/mem[56][5] ), .CK(clk), .Q(\xmem_data[56][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][5]  ( .D(\xmem_inst/mem[52][5] ), .CK(clk), .Q(\xmem_data[52][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][7]  ( .D(\xmem_inst/mem[60][7] ), .CK(clk), .Q(\xmem_data[60][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][7]  ( .D(\xmem_inst/mem[56][7] ), .CK(clk), .Q(\xmem_data[56][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][7]  ( .D(\xmem_inst/mem[48][7] ), .CK(clk), .Q(\xmem_data[48][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][7]  ( .D(\xmem_inst/mem[46][7] ), .CK(clk), .Q(\xmem_data[46][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][4]  ( .D(\xmem_inst/mem[0][4] ), .CK(clk), 
        .Q(\xmem_data[0][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][6]  ( .D(\xmem_inst/mem[88][6] ), .CK(clk), .Q(\xmem_data[88][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][6]  ( .D(\xmem_inst/mem[70][6] ), .CK(clk), .Q(\xmem_data[70][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][6]  ( .D(\xmem_inst/mem[112][6] ), .CK(
        clk), .Q(\xmem_data[112][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][6]  ( .D(\xmem_inst/mem[56][6] ), .CK(clk), .Q(\xmem_data[56][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[48][6]  ( .D(\xmem_inst/mem[48][6] ), .CK(clk), .Q(\xmem_data[48][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][6]  ( .D(\xmem_inst/mem[46][6] ), .CK(clk), .Q(\xmem_data[46][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][6]  ( .D(\xmem_inst/mem[44][6] ), .CK(clk), .Q(\xmem_data[44][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[38][6]  ( .D(\xmem_inst/mem[38][6] ), .CK(clk), .Q(\xmem_data[38][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][5]  ( .D(\xmem_inst/mem[51][5] ), .CK(clk), .Q(\xmem_data[51][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][6]  ( .D(\xmem_inst/mem[37][6] ), .CK(clk), .Q(\xmem_data[37][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][6]  ( .D(\xmem_inst/mem[58][6] ), .CK(clk), .Q(\xmem_data[58][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][6]  ( .D(\xmem_inst/mem[104][6] ), .CK(
        clk), .Q(\xmem_data[104][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][1]  ( .D(\xmem_inst/mem[109][1] ), .CK(
        clk), .Q(\xmem_data[109][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][4]  ( .D(\xmem_inst/mem[103][4] ), .CK(
        clk), .Q(\xmem_data[103][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][2]  ( .D(\xmem_inst/mem[23][2] ), .CK(clk), .Q(\xmem_data[23][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][7]  ( .D(\xmem_inst/mem[10][7] ), .CK(clk), .Q(\xmem_data[10][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][1]  ( .D(\xmem_inst/mem[121][1] ), .CK(
        clk), .Q(\xmem_data[121][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][1]  ( .D(\xmem_inst/mem[119][1] ), .CK(
        clk), .Q(\xmem_data[119][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][1]  ( .D(\xmem_inst/mem[115][1] ), .CK(
        clk), .Q(\xmem_data[115][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][1]  ( .D(\xmem_inst/mem[87][1] ), .CK(clk), .Q(\xmem_data[87][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][1]  ( .D(\xmem_inst/mem[11][1] ), .CK(clk), .Q(\xmem_data[11][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][1]  ( .D(\xmem_inst/mem[35][1] ), .CK(clk), .Q(\xmem_data[35][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][3]  ( .D(\xmem_inst/mem[83][3] ), .CK(clk), .Q(\xmem_data[83][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][3]  ( .D(\xmem_inst/mem[115][3] ), .CK(
        clk), .Q(\xmem_data[115][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[57][3]  ( .D(\xmem_inst/mem[57][3] ), .CK(clk), .Q(\xmem_data[57][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][3]  ( .D(\xmem_inst/mem[55][3] ), .CK(clk), .Q(\xmem_data[55][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][3]  ( .D(\xmem_inst/mem[43][3] ), .CK(clk), .Q(\xmem_data[43][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][4]  ( .D(\xmem_inst/mem[55][4] ), .CK(clk), .Q(\xmem_data[55][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][4]  ( .D(\xmem_inst/mem[51][4] ), .CK(clk), .Q(\xmem_data[51][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][4]  ( .D(\xmem_inst/mem[119][4] ), .CK(
        clk), .Q(\xmem_data[119][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][4]  ( .D(\xmem_inst/mem[115][4] ), .CK(
        clk), .Q(\xmem_data[115][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][1]  ( .D(\xmem_inst/mem[89][1] ), .CK(clk), .Q(\xmem_data[89][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][1]  ( .D(\xmem_inst/mem[1][1] ), .CK(clk), 
        .Q(\xmem_data[1][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][1]  ( .D(\xmem_inst/mem[5][1] ), .CK(clk), 
        .Q(\xmem_data[5][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][2]  ( .D(\xmem_inst/mem[5][2] ), .CK(clk), 
        .Q(\xmem_data[5][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][3]  ( .D(\xmem_inst/mem[87][3] ), .CK(clk), .Q(\xmem_data[87][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[101][1]  ( .D(\xmem_inst/mem[101][1] ), .CK(
        clk), .Q(\xmem_data[101][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][4]  ( .D(\xmem_inst/mem[43][4] ), .CK(clk), .Q(\xmem_data[43][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][1]  ( .D(\xmem_inst/mem[23][1] ), .CK(clk), .Q(\xmem_data[23][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][3]  ( .D(\xmem_inst/mem[23][3] ), .CK(clk), .Q(\xmem_data[23][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][4]  ( .D(\xmem_inst/mem[60][4] ), .CK(clk), .Q(\xmem_data[60][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][1]  ( .D(\xmem_inst/mem[60][1] ), .CK(clk), .Q(\xmem_data[60][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][1]  ( .D(\xmem_inst/mem[20][1] ), .CK(clk), .Q(\xmem_data[20][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][1]  ( .D(\xmem_inst/mem[18][1] ), .CK(clk), .Q(\xmem_data[18][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][1]  ( .D(\xmem_inst/mem[16][1] ), .CK(clk), .Q(\xmem_data[16][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][1]  ( .D(\xmem_inst/mem[62][1] ), .CK(clk), .Q(\xmem_data[62][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[22][0]  ( .D(\xmem_inst/mem[22][0] ), .CK(clk), .Q(\xmem_data[22][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][3]  ( .D(\xmem_inst/mem[118][3] ), .CK(
        clk), .Q(\xmem_data[118][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][5]  ( .D(\xmem_inst/mem[18][5] ), .CK(clk), .Q(\xmem_data[18][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][1]  ( .D(\xmem_inst/mem[78][1] ), .CK(clk), .Q(\xmem_data[78][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][1]  ( .D(\xmem_inst/mem[28][1] ), .CK(clk), .Q(\xmem_data[28][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][1]  ( .D(\xmem_inst/mem[12][1] ), .CK(clk), .Q(\xmem_data[12][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][1]  ( .D(\xmem_inst/mem[42][1] ), .CK(clk), .Q(\xmem_data[42][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][4]  ( .D(\xmem_inst/mem[44][4] ), .CK(clk), .Q(\xmem_data[44][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][1]  ( .D(\xmem_inst/mem[122][1] ), .CK(
        clk), .Q(\xmem_data[122][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][1]  ( .D(\xmem_inst/mem[96][1] ), .CK(clk), .Q(\xmem_data[96][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][1]  ( .D(\xmem_inst/mem[90][1] ), .CK(clk), .Q(\xmem_data[90][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][1]  ( .D(\xmem_inst/mem[72][1] ), .CK(clk), .Q(\xmem_data[72][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][1]  ( .D(\xmem_inst/mem[74][1] ), .CK(clk), .Q(\xmem_data[74][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][1]  ( .D(\xmem_inst/mem[76][1] ), .CK(clk), .Q(\xmem_data[76][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][1]  ( .D(\xmem_inst/mem[64][1] ), .CK(clk), .Q(\xmem_data[64][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][1]  ( .D(\xmem_inst/mem[2][1] ), .CK(clk), 
        .Q(\xmem_data[2][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][1]  ( .D(\xmem_inst/mem[54][1] ), .CK(clk), .Q(\xmem_data[54][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][1]  ( .D(\xmem_inst/mem[50][1] ), .CK(clk), .Q(\xmem_data[50][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][1]  ( .D(\xmem_inst/mem[44][1] ), .CK(clk), .Q(\xmem_data[44][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][0]  ( .D(\xmem_inst/mem[24][0] ), .CK(clk), .Q(\xmem_data[24][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][7]  ( .D(\xmem_inst/mem[12][7] ), .CK(clk), .Q(\xmem_data[12][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][3]  ( .D(\xmem_inst/mem[64][3] ), .CK(clk), .Q(\xmem_data[64][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][3]  ( .D(\xmem_inst/mem[96][3] ), .CK(clk), .Q(\xmem_data[96][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][3]  ( .D(\xmem_inst/mem[62][3] ), .CK(clk), .Q(\xmem_data[62][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][3]  ( .D(\xmem_inst/mem[60][3] ), .CK(clk), .Q(\xmem_data[60][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][4]  ( .D(\xmem_inst/mem[36][4] ), .CK(clk), .Q(\xmem_data[36][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][4]  ( .D(\xmem_inst/mem[62][4] ), .CK(clk), .Q(\xmem_data[62][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][4]  ( .D(\xmem_inst/mem[40][4] ), .CK(clk), .Q(\xmem_data[40][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][4]  ( .D(\xmem_inst/mem[96][4] ), .CK(clk), .Q(\xmem_data[96][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][4]  ( .D(\xmem_inst/mem[122][4] ), .CK(
        clk), .Q(\xmem_data[122][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][4]  ( .D(\xmem_inst/mem[110][4] ), .CK(
        clk), .Q(\xmem_data[110][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][4]  ( .D(\xmem_inst/mem[108][4] ), .CK(
        clk), .Q(\xmem_data[108][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[112][4]  ( .D(\xmem_inst/mem[112][4] ), .CK(
        clk), .Q(\xmem_data[112][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[53][1]  ( .D(\xmem_inst/mem[53][1] ), .CK(clk), .Q(\xmem_data[53][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[49][1]  ( .D(\xmem_inst/mem[49][1] ), .CK(clk), .Q(\xmem_data[49][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][1]  ( .D(\xmem_inst/mem[116][1] ), .CK(
        clk), .Q(\xmem_data[116][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][5]  ( .D(\xmem_inst/mem[5][5] ), .CK(clk), 
        .Q(\xmem_data[5][5] ), .QN(n39026) );
  DFF_X2 \xmem_inst/data_out_reg[7][3]  ( .D(\xmem_inst/mem[7][3] ), .CK(clk), 
        .Q(\xmem_data[7][3] ), .QN(n39017) );
  DFF_X2 \xmem_inst/data_out_reg[7][1]  ( .D(\xmem_inst/mem[7][1] ), .CK(clk), 
        .Q(\xmem_data[7][1] ), .QN(n39020) );
  DFF_X2 \xmem_inst/data_out_reg[15][1]  ( .D(\xmem_inst/mem[15][1] ), .CK(clk), .Q(\xmem_data[15][1] ), .QN(n39016) );
  DFF_X2 \xmem_inst/data_out_reg[14][3]  ( .D(\xmem_inst/mem[14][3] ), .CK(clk), .Q(\xmem_data[14][3] ), .QN(n39022) );
  DFF_X2 \xmem_inst/data_out_reg[119][7]  ( .D(\xmem_inst/mem[119][7] ), .CK(
        clk), .Q(\xmem_data[119][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][7]  ( .D(\xmem_inst/mem[5][7] ), .CK(clk), 
        .Q(\xmem_data[5][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][0]  ( .D(\xmem_inst/mem[119][0] ), .CK(
        clk), .Q(\xmem_data[119][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][3]  ( .D(\xmem_inst/mem[111][3] ), .CK(
        clk), .Q(\xmem_data[111][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][6]  ( .D(\xmem_inst/mem[50][6] ), .CK(clk), .Q(\xmem_data[50][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][3]  ( .D(\xmem_inst/mem[12][3] ), .CK(clk), .Q(\xmem_data[12][3] ), .QN(n39011) );
  DFF_X2 \xmem_inst/data_out_reg[115][0]  ( .D(\xmem_inst/mem[115][0] ), .CK(
        clk), .Q(\xmem_data[115][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][0]  ( .D(\xmem_inst/mem[111][0] ), .CK(
        clk), .Q(\xmem_data[111][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][0]  ( .D(\xmem_inst/mem[121][0] ), .CK(
        clk), .Q(\xmem_data[121][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][0]  ( .D(\xmem_inst/mem[83][0] ), .CK(clk), .Q(\xmem_data[83][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][0]  ( .D(\xmem_inst/mem[79][0] ), .CK(clk), .Q(\xmem_data[79][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][0]  ( .D(\xmem_inst/mem[89][0] ), .CK(clk), .Q(\xmem_data[89][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][7]  ( .D(\xmem_inst/mem[111][7] ), .CK(
        clk), .Q(\xmem_data[111][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][7]  ( .D(\xmem_inst/mem[115][7] ), .CK(
        clk), .Q(\xmem_data[115][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][7]  ( .D(\xmem_inst/mem[121][7] ), .CK(
        clk), .Q(\xmem_data[121][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][3]  ( .D(\xmem_inst/mem[79][3] ), .CK(clk), .Q(\xmem_data[79][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[41][0]  ( .D(\xmem_inst/mem[41][0] ), .CK(clk), .Q(\xmem_data[41][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][6]  ( .D(\xmem_inst/mem[11][6] ), .CK(clk), .Q(\xmem_data[11][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][3]  ( .D(\xmem_inst/mem[5][3] ), .CK(clk), 
        .Q(\xmem_data[5][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][0]  ( .D(\xmem_inst/mem[1][0] ), .CK(clk), 
        .Q(\xmem_data[1][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][3]  ( .D(\xmem_inst/mem[10][3] ), .CK(clk), .Q(\xmem_data[10][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][4]  ( .D(\xmem_inst/mem[12][4] ), .CK(clk), .Q(\xmem_data[12][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][0]  ( .D(\xmem_inst/mem[62][0] ), .CK(clk), .Q(\xmem_data[62][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][0]  ( .D(\xmem_inst/mem[60][0] ), .CK(clk), .Q(\xmem_data[60][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[15][5]  ( .D(\xmem_inst/mem[15][5] ), .CK(clk), .Q(\xmem_data[15][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][4]  ( .D(\xmem_inst/mem[87][4] ), .CK(clk), .Q(\xmem_data[87][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][6]  ( .D(\xmem_inst/mem[8][6] ), .CK(clk), 
        .Q(\xmem_data[8][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][4]  ( .D(\xmem_inst/mem[10][4] ), .CK(clk), .Q(\xmem_data[10][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][5]  ( .D(\xmem_inst/mem[10][5] ), .CK(clk), .Q(\xmem_data[10][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][7]  ( .D(\xmem_inst/mem[108][7] ), .CK(
        clk), .Q(\xmem_data[108][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][7]  ( .D(\xmem_inst/mem[100][7] ), .CK(
        clk), .Q(\xmem_data[100][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][7]  ( .D(\xmem_inst/mem[98][7] ), .CK(clk), .Q(\xmem_data[98][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][7]  ( .D(\xmem_inst/mem[96][7] ), .CK(clk), .Q(\xmem_data[96][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][7]  ( .D(\xmem_inst/mem[122][7] ), .CK(
        clk), .Q(\xmem_data[122][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][0]  ( .D(\xmem_inst/mem[44][0] ), .CK(clk), .Q(\xmem_data[44][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][0]  ( .D(\xmem_inst/mem[42][0] ), .CK(clk), .Q(\xmem_data[42][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][0]  ( .D(\xmem_inst/mem[36][0] ), .CK(clk), .Q(\xmem_data[36][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][0]  ( .D(\xmem_inst/mem[34][0] ), .CK(clk), .Q(\xmem_data[34][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][0]  ( .D(\xmem_inst/mem[50][0] ), .CK(clk), .Q(\xmem_data[50][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[58][0]  ( .D(\xmem_inst/mem[58][0] ), .CK(clk), .Q(\xmem_data[58][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][4]  ( .D(\xmem_inst/mem[120][4] ), .CK(
        clk), .Q(\xmem_data[120][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][4]  ( .D(\xmem_inst/mem[82][4] ), .CK(clk), .Q(\xmem_data[82][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][4]  ( .D(\xmem_inst/mem[88][4] ), .CK(clk), .Q(\xmem_data[88][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][4]  ( .D(\xmem_inst/mem[74][4] ), .CK(clk), .Q(\xmem_data[74][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][3]  ( .D(\xmem_inst/mem[108][3] ), .CK(
        clk), .Q(\xmem_data[108][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][3]  ( .D(\xmem_inst/mem[76][3] ), .CK(clk), .Q(\xmem_data[76][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[106][3]  ( .D(\xmem_inst/mem[106][3] ), .CK(
        clk), .Q(\xmem_data[106][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][5]  ( .D(\xmem_inst/mem[119][5] ), .CK(
        clk), .Q(\xmem_data[119][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][3]  ( .D(\xmem_inst/mem[89][3] ), .CK(clk), .Q(\xmem_data[89][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][5]  ( .D(\xmem_inst/mem[23][5] ), .CK(clk), .Q(\xmem_data[23][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][0]  ( .D(\xmem_inst/mem[11][0] ), .CK(clk), .Q(\xmem_data[11][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][7]  ( .D(\xmem_inst/mem[83][7] ), .CK(clk), .Q(\xmem_data[83][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][7]  ( .D(\xmem_inst/mem[73][7] ), .CK(clk), .Q(\xmem_data[73][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][7]  ( .D(\xmem_inst/mem[67][7] ), .CK(clk), .Q(\xmem_data[67][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][5]  ( .D(\xmem_inst/mem[115][5] ), .CK(
        clk), .Q(\xmem_data[115][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][4]  ( .D(\xmem_inst/mem[69][4] ), .CK(clk), .Q(\xmem_data[69][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[95][4]  ( .D(\xmem_inst/mem[95][4] ), .CK(clk), .Q(\xmem_data[95][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][4]  ( .D(\xmem_inst/mem[77][4] ), .CK(clk), .Q(\xmem_data[77][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[73][4]  ( .D(\xmem_inst/mem[73][4] ), .CK(clk), .Q(\xmem_data[73][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[125][3]  ( .D(\xmem_inst/mem[125][3] ), .CK(
        clk), .Q(\xmem_data[125][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][3]  ( .D(\xmem_inst/mem[121][3] ), .CK(
        clk), .Q(\xmem_data[121][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][0]  ( .D(\xmem_inst/mem[27][0] ), .CK(clk), .Q(\xmem_data[27][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][2]  ( .D(\xmem_inst/mem[21][2] ), .CK(clk), .Q(\xmem_data[21][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][5]  ( .D(\xmem_inst/mem[93][5] ), .CK(clk), .Q(\xmem_data[93][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][5]  ( .D(\xmem_inst/mem[83][5] ), .CK(clk), .Q(\xmem_data[83][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][4]  ( .D(\xmem_inst/mem[67][4] ), .CK(clk), .Q(\xmem_data[67][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][5]  ( .D(\xmem_inst/mem[13][5] ), .CK(clk), .Q(\xmem_data[13][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[93][4]  ( .D(\xmem_inst/mem[93][4] ), .CK(clk), .Q(\xmem_data[93][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][0]  ( .D(\xmem_inst/mem[19][0] ), .CK(clk), .Q(\xmem_data[19][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[8][3]  ( .D(\xmem_inst/mem[8][3] ), .CK(clk), 
        .Q(\xmem_data[8][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[28][4]  ( .D(\xmem_inst/mem[28][4] ), .CK(clk), .Q(\xmem_data[28][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][2]  ( .D(\xmem_inst/mem[11][2] ), .CK(clk), .Q(\xmem_data[11][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][5]  ( .D(\xmem_inst/mem[0][5] ), .CK(clk), 
        .Q(\xmem_data[0][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][7]  ( .D(\xmem_inst/mem[86][7] ), .CK(clk), .Q(\xmem_data[86][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][0]  ( .D(\xmem_inst/mem[12][0] ), .CK(clk), .Q(\xmem_data[12][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[14][4]  ( .D(\xmem_inst/mem[14][4] ), .CK(clk), .Q(\xmem_data[14][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[2][5]  ( .D(\xmem_inst/mem[2][5] ), .CK(clk), 
        .Q(\xmem_data[2][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][3]  ( .D(\xmem_inst/mem[68][3] ), .CK(clk), .Q(\xmem_data[68][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][3]  ( .D(\xmem_inst/mem[36][3] ), .CK(clk), .Q(\xmem_data[36][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][0]  ( .D(\xmem_inst/mem[90][0] ), .CK(clk), .Q(\xmem_data[90][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][0]  ( .D(\xmem_inst/mem[100][0] ), .CK(
        clk), .Q(\xmem_data[100][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][0]  ( .D(\xmem_inst/mem[98][0] ), .CK(clk), .Q(\xmem_data[98][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][0]  ( .D(\xmem_inst/mem[96][0] ), .CK(clk), .Q(\xmem_data[96][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][0]  ( .D(\xmem_inst/mem[108][0] ), .CK(
        clk), .Q(\xmem_data[108][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][0]  ( .D(\xmem_inst/mem[124][0] ), .CK(
        clk), .Q(\xmem_data[124][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][0]  ( .D(\xmem_inst/mem[122][0] ), .CK(
        clk), .Q(\xmem_data[122][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][0]  ( .D(\xmem_inst/mem[68][0] ), .CK(clk), .Q(\xmem_data[68][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][0]  ( .D(\xmem_inst/mem[66][0] ), .CK(clk), .Q(\xmem_data[66][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][0]  ( .D(\xmem_inst/mem[64][0] ), .CK(clk), .Q(\xmem_data[64][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][0]  ( .D(\xmem_inst/mem[76][0] ), .CK(clk), .Q(\xmem_data[76][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][3]  ( .D(\xmem_inst/mem[18][3] ), .CK(clk), .Q(\xmem_data[18][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][7]  ( .D(\xmem_inst/mem[94][7] ), .CK(clk), .Q(\xmem_data[94][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][7]  ( .D(\xmem_inst/mem[92][7] ), .CK(clk), .Q(\xmem_data[92][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[90][7]  ( .D(\xmem_inst/mem[90][7] ), .CK(clk), .Q(\xmem_data[90][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][7]  ( .D(\xmem_inst/mem[88][7] ), .CK(clk), .Q(\xmem_data[88][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[76][7]  ( .D(\xmem_inst/mem[76][7] ), .CK(clk), .Q(\xmem_data[76][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][7]  ( .D(\xmem_inst/mem[74][7] ), .CK(clk), .Q(\xmem_data[74][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][7]  ( .D(\xmem_inst/mem[68][7] ), .CK(clk), .Q(\xmem_data[68][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][4]  ( .D(\xmem_inst/mem[34][4] ), .CK(clk), .Q(\xmem_data[34][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][3]  ( .D(\xmem_inst/mem[66][3] ), .CK(clk), .Q(\xmem_data[66][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][3]  ( .D(\xmem_inst/mem[122][3] ), .CK(
        clk), .Q(\xmem_data[122][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][3]  ( .D(\xmem_inst/mem[98][3] ), .CK(clk), .Q(\xmem_data[98][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[24][4]  ( .D(\xmem_inst/mem[24][4] ), .CK(clk), .Q(\xmem_data[24][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][2]  ( .D(\xmem_inst/mem[88][2] ), .CK(clk), .Q(\xmem_data[88][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][2]  ( .D(\xmem_inst/mem[120][2] ), .CK(
        clk), .Q(\xmem_data[120][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][2]  ( .D(\xmem_inst/mem[70][2] ), .CK(clk), .Q(\xmem_data[70][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][2]  ( .D(\xmem_inst/mem[34][2] ), .CK(clk), .Q(\xmem_data[34][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][2]  ( .D(\xmem_inst/mem[82][2] ), .CK(clk), .Q(\xmem_data[82][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][2]  ( .D(\xmem_inst/mem[114][2] ), .CK(
        clk), .Q(\xmem_data[114][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][0]  ( .D(\xmem_inst/mem[31][0] ), .CK(clk), .Q(\xmem_data[31][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][4]  ( .D(\xmem_inst/mem[27][4] ), .CK(clk), .Q(\xmem_data[27][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][5]  ( .D(\xmem_inst/mem[121][5] ), .CK(
        clk), .Q(\xmem_data[121][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][3]  ( .D(\xmem_inst/mem[20][3] ), .CK(clk), .Q(\xmem_data[20][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][5]  ( .D(\xmem_inst/mem[20][5] ), .CK(clk), .Q(\xmem_data[20][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][3]  ( .D(\xmem_inst/mem[50][3] ), .CK(clk), .Q(\xmem_data[50][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[25][3]  ( .D(\xmem_inst/mem[25][3] ), .CK(clk), .Q(\xmem_data[25][3] ), .QN(n39027) );
  DFF_X2 \xmem_inst/data_out_reg[20][0]  ( .D(\xmem_inst/mem[20][0] ), .CK(clk), .Q(\xmem_data[20][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[12][2]  ( .D(\xmem_inst/mem[12][2] ), .CK(clk), .Q(\xmem_data[12][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][5]  ( .D(\xmem_inst/mem[110][5] ), .CK(
        clk), .Q(\xmem_data[110][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][5]  ( .D(\xmem_inst/mem[94][5] ), .CK(clk), .Q(\xmem_data[94][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[79][2]  ( .D(\xmem_inst/mem[79][2] ), .CK(clk), .Q(\xmem_data[79][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[77][2]  ( .D(\xmem_inst/mem[77][2] ), .CK(clk), .Q(\xmem_data[77][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[61][2]  ( .D(\xmem_inst/mem[61][2] ), .CK(clk), .Q(\xmem_data[61][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[63][2]  ( .D(\xmem_inst/mem[63][2] ), .CK(clk), .Q(\xmem_data[63][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][2]  ( .D(\xmem_inst/mem[51][2] ), .CK(clk), .Q(\xmem_data[51][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][2]  ( .D(\xmem_inst/mem[45][2] ), .CK(clk), .Q(\xmem_data[45][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[37][2]  ( .D(\xmem_inst/mem[37][2] ), .CK(clk), .Q(\xmem_data[37][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][2]  ( .D(\xmem_inst/mem[111][2] ), .CK(
        clk), .Q(\xmem_data[111][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][2]  ( .D(\xmem_inst/mem[109][2] ), .CK(
        clk), .Q(\xmem_data[109][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][2]  ( .D(\xmem_inst/mem[97][2] ), .CK(clk), .Q(\xmem_data[97][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[91][2]  ( .D(\xmem_inst/mem[91][2] ), .CK(clk), .Q(\xmem_data[91][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][2]  ( .D(\xmem_inst/mem[65][2] ), .CK(clk), .Q(\xmem_data[65][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][4]  ( .D(\xmem_inst/mem[31][4] ), .CK(clk), .Q(\xmem_data[31][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][5]  ( .D(\xmem_inst/mem[66][5] ), .CK(clk), .Q(\xmem_data[66][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[7][6]  ( .D(\xmem_inst/mem[7][6] ), .CK(clk), 
        .Q(\xmem_data[7][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[19][4]  ( .D(\xmem_inst/mem[19][4] ), .CK(clk), .Q(\xmem_data[19][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[1][6]  ( .D(\xmem_inst/mem[1][6] ), .CK(clk), 
        .Q(\xmem_data[1][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[43][7]  ( .D(\xmem_inst/mem[43][7] ), .CK(clk), .Q(\xmem_data[43][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][6]  ( .D(\xmem_inst/mem[111][6] ), .CK(
        clk), .Q(\xmem_data[111][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[3][7]  ( .D(\xmem_inst/mem[3][7] ), .CK(clk), 
        .Q(\xmem_data[3][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][6]  ( .D(\xmem_inst/mem[54][6] ), .CK(clk), .Q(\xmem_data[54][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][6]  ( .D(\xmem_inst/mem[5][6] ), .CK(clk), 
        .Q(\xmem_data[5][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[21][4]  ( .D(\xmem_inst/mem[21][4] ), .CK(clk), .Q(\xmem_data[21][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][7]  ( .D(\xmem_inst/mem[55][7] ), .CK(clk), .Q(\xmem_data[55][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[45][7]  ( .D(\xmem_inst/mem[45][7] ), .CK(clk), .Q(\xmem_data[45][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][5]  ( .D(\xmem_inst/mem[55][5] ), .CK(clk), .Q(\xmem_data[55][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[69][5]  ( .D(\xmem_inst/mem[69][5] ), .CK(clk), .Q(\xmem_data[69][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[97][5]  ( .D(\xmem_inst/mem[97][5] ), .CK(clk), .Q(\xmem_data[97][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[109][5]  ( .D(\xmem_inst/mem[109][5] ), .CK(
        clk), .Q(\xmem_data[109][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][6]  ( .D(\xmem_inst/mem[115][6] ), .CK(
        clk), .Q(\xmem_data[115][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][4]  ( .D(\xmem_inst/mem[5][4] ), .CK(clk), 
        .Q(\xmem_data[5][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][6]  ( .D(\xmem_inst/mem[13][6] ), .CK(clk), .Q(\xmem_data[13][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[23][4]  ( .D(\xmem_inst/mem[23][4] ), .CK(clk), .Q(\xmem_data[23][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[17][4]  ( .D(\xmem_inst/mem[17][4] ), .CK(clk), .Q(\xmem_data[17][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][6]  ( .D(\xmem_inst/mem[16][6] ), .CK(clk), .Q(\xmem_data[16][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][5]  ( .D(\xmem_inst/mem[42][5] ), .CK(clk), .Q(\xmem_data[42][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][5]  ( .D(\xmem_inst/mem[36][5] ), .CK(clk), .Q(\xmem_data[36][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[74][6]  ( .D(\xmem_inst/mem[74][6] ), .CK(clk), .Q(\xmem_data[74][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[68][6]  ( .D(\xmem_inst/mem[68][6] ), .CK(clk), .Q(\xmem_data[68][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][6]  ( .D(\xmem_inst/mem[87][6] ), .CK(clk), .Q(\xmem_data[87][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[18][6]  ( .D(\xmem_inst/mem[18][6] ), .CK(clk), .Q(\xmem_data[18][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][6]  ( .D(\xmem_inst/mem[124][6] ), .CK(
        clk), .Q(\xmem_data[124][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[94][6]  ( .D(\xmem_inst/mem[94][6] ), .CK(clk), .Q(\xmem_data[94][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][5]  ( .D(\xmem_inst/mem[62][5] ), .CK(clk), .Q(\xmem_data[62][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][5]  ( .D(\xmem_inst/mem[60][5] ), .CK(clk), .Q(\xmem_data[60][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[52][7]  ( .D(\xmem_inst/mem[52][7] ), .CK(clk), .Q(\xmem_data[52][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][7]  ( .D(\xmem_inst/mem[50][7] ), .CK(clk), .Q(\xmem_data[50][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][7]  ( .D(\xmem_inst/mem[0][7] ), .CK(clk), 
        .Q(\xmem_data[0][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][6]  ( .D(\xmem_inst/mem[92][6] ), .CK(clk), .Q(\xmem_data[92][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][6]  ( .D(\xmem_inst/mem[82][6] ), .CK(clk), .Q(\xmem_data[82][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[80][6]  ( .D(\xmem_inst/mem[80][6] ), .CK(clk), .Q(\xmem_data[80][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][6]  ( .D(\xmem_inst/mem[72][6] ), .CK(clk), .Q(\xmem_data[72][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][6]  ( .D(\xmem_inst/mem[108][6] ), .CK(
        clk), .Q(\xmem_data[108][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][6]  ( .D(\xmem_inst/mem[102][6] ), .CK(
        clk), .Q(\xmem_data[102][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[100][6]  ( .D(\xmem_inst/mem[100][6] ), .CK(
        clk), .Q(\xmem_data[100][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[98][6]  ( .D(\xmem_inst/mem[98][6] ), .CK(clk), .Q(\xmem_data[98][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[96][6]  ( .D(\xmem_inst/mem[96][6] ), .CK(clk), .Q(\xmem_data[96][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[62][6]  ( .D(\xmem_inst/mem[62][6] ), .CK(clk), .Q(\xmem_data[62][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[60][6]  ( .D(\xmem_inst/mem[60][6] ), .CK(clk), .Q(\xmem_data[60][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][6]  ( .D(\xmem_inst/mem[42][6] ), .CK(clk), .Q(\xmem_data[42][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][5]  ( .D(\xmem_inst/mem[40][5] ), .CK(clk), .Q(\xmem_data[40][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[36][6]  ( .D(\xmem_inst/mem[36][6] ), .CK(clk), .Q(\xmem_data[36][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][5]  ( .D(\xmem_inst/mem[50][5] ), .CK(clk), .Q(\xmem_data[50][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][1]  ( .D(\xmem_inst/mem[82][1] ), .CK(clk), .Q(\xmem_data[82][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[105][1]  ( .D(\xmem_inst/mem[105][1] ), .CK(
        clk), .Q(\xmem_data[105][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][1]  ( .D(\xmem_inst/mem[31][1] ), .CK(clk), .Q(\xmem_data[31][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][1]  ( .D(\xmem_inst/mem[33][1] ), .CK(clk), .Q(\xmem_data[33][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][3]  ( .D(\xmem_inst/mem[103][3] ), .CK(
        clk), .Q(\xmem_data[103][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][3]  ( .D(\xmem_inst/mem[33][3] ), .CK(clk), .Q(\xmem_data[33][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[31][3]  ( .D(\xmem_inst/mem[31][3] ), .CK(clk), .Q(\xmem_data[31][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][4]  ( .D(\xmem_inst/mem[33][4] ), .CK(clk), .Q(\xmem_data[33][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[85][1]  ( .D(\xmem_inst/mem[85][1] ), .CK(clk), .Q(\xmem_data[85][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][1]  ( .D(\xmem_inst/mem[4][1] ), .CK(clk), 
        .Q(\xmem_data[4][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][2]  ( .D(\xmem_inst/mem[4][2] ), .CK(clk), 
        .Q(\xmem_data[4][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][3]  ( .D(\xmem_inst/mem[86][3] ), .CK(clk), .Q(\xmem_data[86][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][3]  ( .D(\xmem_inst/mem[70][3] ), .CK(clk), .Q(\xmem_data[70][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][4]  ( .D(\xmem_inst/mem[102][4] ), .CK(
        clk), .Q(\xmem_data[102][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][1]  ( .D(\xmem_inst/mem[120][1] ), .CK(
        clk), .Q(\xmem_data[120][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][1]  ( .D(\xmem_inst/mem[102][1] ), .CK(
        clk), .Q(\xmem_data[102][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][1]  ( .D(\xmem_inst/mem[110][1] ), .CK(
        clk), .Q(\xmem_data[110][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][1]  ( .D(\xmem_inst/mem[86][1] ), .CK(clk), .Q(\xmem_data[86][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][1]  ( .D(\xmem_inst/mem[10][1] ), .CK(clk), .Q(\xmem_data[10][1] ), .QN(n39033) );
  DFF_X2 \xmem_inst/data_out_reg[18][2]  ( .D(\xmem_inst/mem[18][2] ), .CK(clk), .Q(\xmem_data[18][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][3]  ( .D(\xmem_inst/mem[84][3] ), .CK(clk), .Q(\xmem_data[84][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][3]  ( .D(\xmem_inst/mem[82][3] ), .CK(clk), .Q(\xmem_data[82][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][3]  ( .D(\xmem_inst/mem[116][3] ), .CK(
        clk), .Q(\xmem_data[116][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][3]  ( .D(\xmem_inst/mem[114][3] ), .CK(
        clk), .Q(\xmem_data[114][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[56][3]  ( .D(\xmem_inst/mem[56][3] ), .CK(clk), .Q(\xmem_data[56][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][3]  ( .D(\xmem_inst/mem[54][3] ), .CK(clk), .Q(\xmem_data[54][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][3]  ( .D(\xmem_inst/mem[44][3] ), .CK(clk), .Q(\xmem_data[44][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[42][3]  ( .D(\xmem_inst/mem[42][3] ), .CK(clk), .Q(\xmem_data[42][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][3]  ( .D(\xmem_inst/mem[26][3] ), .CK(clk), .Q(\xmem_data[26][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][4]  ( .D(\xmem_inst/mem[54][4] ), .CK(clk), .Q(\xmem_data[54][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][4]  ( .D(\xmem_inst/mem[116][4] ), .CK(
        clk), .Q(\xmem_data[116][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][4]  ( .D(\xmem_inst/mem[114][4] ), .CK(
        clk), .Q(\xmem_data[114][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][1]  ( .D(\xmem_inst/mem[55][1] ), .CK(clk), .Q(\xmem_data[55][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][0]  ( .D(\xmem_inst/mem[4][0] ), .CK(clk), 
        .Q(\xmem_data[4][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][1]  ( .D(\xmem_inst/mem[118][1] ), .CK(
        clk), .Q(\xmem_data[118][1] ) );
  DFF_X2 \ctrl_conv_output_inst/load_xaddr_val_reg[5]  ( .D(n1814), .CK(clk), 
        .Q(load_xaddr_val[5]), .QN(n39041) );
  DFF_X2 \xmem_inst/data_out_reg[34][1]  ( .D(\xmem_inst/mem[34][1] ), .CK(clk), .Q(\xmem_data[34][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][7]  ( .D(\xmem_inst/mem[13][7] ), .CK(clk), .Q(\xmem_data[13][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][7]  ( .D(\xmem_inst/mem[6][7] ), .CK(clk), 
        .Q(\xmem_data[6][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][0]  ( .D(\xmem_inst/mem[103][0] ), .CK(
        clk), .Q(\xmem_data[103][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[87][0]  ( .D(\xmem_inst/mem[87][0] ), .CK(clk), .Q(\xmem_data[87][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[117][7]  ( .D(\xmem_inst/mem[117][7] ), .CK(
        clk), .Q(\xmem_data[117][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][7]  ( .D(\xmem_inst/mem[4][7] ), .CK(clk), 
        .Q(\xmem_data[4][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][0]  ( .D(\xmem_inst/mem[33][0] ), .CK(clk), .Q(\xmem_data[33][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][7]  ( .D(\xmem_inst/mem[118][7] ), .CK(
        clk), .Q(\xmem_data[118][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][6]  ( .D(\xmem_inst/mem[10][6] ), .CK(clk), .Q(\xmem_data[10][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][3]  ( .D(\xmem_inst/mem[4][3] ), .CK(clk), 
        .Q(\xmem_data[4][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[4][5]  ( .D(\xmem_inst/mem[4][5] ), .CK(clk), 
        .Q(\xmem_data[4][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][4]  ( .D(\xmem_inst/mem[64][4] ), .CK(clk), .Q(\xmem_data[64][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[0][3]  ( .D(\xmem_inst/mem[0][3] ), .CK(clk), 
        .Q(\xmem_data[0][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][7]  ( .D(\xmem_inst/mem[102][7] ), .CK(
        clk), .Q(\xmem_data[102][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][7]  ( .D(\xmem_inst/mem[120][7] ), .CK(
        clk), .Q(\xmem_data[120][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][3]  ( .D(\xmem_inst/mem[110][3] ), .CK(
        clk), .Q(\xmem_data[110][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][0]  ( .D(\xmem_inst/mem[40][0] ), .CK(clk), .Q(\xmem_data[40][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][3]  ( .D(\xmem_inst/mem[78][3] ), .CK(clk), .Q(\xmem_data[78][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][3]  ( .D(\xmem_inst/mem[11][3] ), .CK(clk), .Q(\xmem_data[11][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][3]  ( .D(\xmem_inst/mem[35][3] ), .CK(clk), .Q(\xmem_data[35][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][7]  ( .D(\xmem_inst/mem[65][7] ), .CK(clk), .Q(\xmem_data[65][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][4]  ( .D(\xmem_inst/mem[121][4] ), .CK(
        clk), .Q(\xmem_data[121][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[75][4]  ( .D(\xmem_inst/mem[75][4] ), .CK(clk), .Q(\xmem_data[75][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][4]  ( .D(\xmem_inst/mem[89][4] ), .CK(clk), .Q(\xmem_data[89][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[119][3]  ( .D(\xmem_inst/mem[119][3] ), .CK(
        clk), .Q(\xmem_data[119][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[11][5]  ( .D(\xmem_inst/mem[11][5] ), .CK(clk), .Q(\xmem_data[11][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][0]  ( .D(\xmem_inst/mem[116][0] ), .CK(
        clk), .Q(\xmem_data[116][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][0]  ( .D(\xmem_inst/mem[118][0] ), .CK(
        clk), .Q(\xmem_data[118][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[78][0]  ( .D(\xmem_inst/mem[78][0] ), .CK(clk), .Q(\xmem_data[78][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][0]  ( .D(\xmem_inst/mem[114][0] ), .CK(
        clk), .Q(\xmem_data[114][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][0]  ( .D(\xmem_inst/mem[110][0] ), .CK(
        clk), .Q(\xmem_data[110][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][0]  ( .D(\xmem_inst/mem[120][0] ), .CK(
        clk), .Q(\xmem_data[120][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][0]  ( .D(\xmem_inst/mem[70][0] ), .CK(clk), .Q(\xmem_data[70][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][0]  ( .D(\xmem_inst/mem[84][0] ), .CK(clk), .Q(\xmem_data[84][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][0]  ( .D(\xmem_inst/mem[82][0] ), .CK(clk), .Q(\xmem_data[82][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][0]  ( .D(\xmem_inst/mem[88][0] ), .CK(clk), .Q(\xmem_data[88][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[26][0]  ( .D(\xmem_inst/mem[26][0] ), .CK(clk), .Q(\xmem_data[26][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[72][7]  ( .D(\xmem_inst/mem[72][7] ), .CK(clk), .Q(\xmem_data[72][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][3]  ( .D(\xmem_inst/mem[120][3] ), .CK(
        clk), .Q(\xmem_data[120][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[20][2]  ( .D(\xmem_inst/mem[20][2] ), .CK(clk), .Q(\xmem_data[20][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[124][3]  ( .D(\xmem_inst/mem[124][3] ), .CK(
        clk), .Q(\xmem_data[124][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[27][5]  ( .D(\xmem_inst/mem[27][5] ), .CK(clk), .Q(\xmem_data[27][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[10][0]  ( .D(\xmem_inst/mem[10][0] ), .CK(clk), .Q(\xmem_data[10][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[71][2]  ( .D(\xmem_inst/mem[71][2] ), .CK(clk), .Q(\xmem_data[71][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[123][2]  ( .D(\xmem_inst/mem[123][2] ), .CK(
        clk), .Q(\xmem_data[123][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[115][2]  ( .D(\xmem_inst/mem[115][2] ), .CK(
        clk), .Q(\xmem_data[115][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][2]  ( .D(\xmem_inst/mem[33][2] ), .CK(clk), .Q(\xmem_data[33][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][2]  ( .D(\xmem_inst/mem[83][2] ), .CK(clk), .Q(\xmem_data[83][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[103][2]  ( .D(\xmem_inst/mem[103][2] ), .CK(
        clk), .Q(\xmem_data[103][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[89][2]  ( .D(\xmem_inst/mem[89][2] ), .CK(clk), .Q(\xmem_data[89][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][2]  ( .D(\xmem_inst/mem[121][2] ), .CK(
        clk), .Q(\xmem_data[121][2] ) );
  DFF_X2 \xmem_inst/data_out_reg[92][5]  ( .D(\xmem_inst/mem[92][5] ), .CK(clk), .Q(\xmem_data[92][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][5]  ( .D(\xmem_inst/mem[120][5] ), .CK(
        clk), .Q(\xmem_data[120][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][5]  ( .D(\xmem_inst/mem[116][5] ), .CK(
        clk), .Q(\xmem_data[116][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[30][0]  ( .D(\xmem_inst/mem[30][0] ), .CK(clk), .Q(\xmem_data[30][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[6][0]  ( .D(\xmem_inst/mem[6][0] ), .CK(clk), 
        .Q(\xmem_data[6][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][5]  ( .D(\xmem_inst/mem[35][5] ), .CK(clk), .Q(\xmem_data[35][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][7]  ( .D(\xmem_inst/mem[35][7] ), .CK(clk), .Q(\xmem_data[35][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[33][7]  ( .D(\xmem_inst/mem[33][7] ), .CK(clk), .Q(\xmem_data[33][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][5]  ( .D(\xmem_inst/mem[65][5] ), .CK(clk), .Q(\xmem_data[65][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[111][5]  ( .D(\xmem_inst/mem[111][5] ), .CK(
        clk), .Q(\xmem_data[111][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[121][6]  ( .D(\xmem_inst/mem[121][6] ), .CK(
        clk), .Q(\xmem_data[121][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[55][6]  ( .D(\xmem_inst/mem[55][6] ), .CK(clk), .Q(\xmem_data[55][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[22][6]  ( .D(\xmem_inst/mem[22][6] ), .CK(clk), .Q(\xmem_data[22][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][6]  ( .D(\xmem_inst/mem[116][6] ), .CK(
        clk), .Q(\xmem_data[116][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[122][6]  ( .D(\xmem_inst/mem[122][6] ), .CK(
        clk), .Q(\xmem_data[122][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[126][6]  ( .D(\xmem_inst/mem[126][6] ), .CK(
        clk), .Q(\xmem_data[126][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][5]  ( .D(\xmem_inst/mem[32][5] ), .CK(clk), .Q(\xmem_data[32][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][5]  ( .D(\xmem_inst/mem[54][5] ), .CK(clk), .Q(\xmem_data[54][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[44][7]  ( .D(\xmem_inst/mem[44][7] ), .CK(clk), .Q(\xmem_data[44][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][7]  ( .D(\xmem_inst/mem[40][7] ), .CK(clk), .Q(\xmem_data[40][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][6]  ( .D(\xmem_inst/mem[64][6] ), .CK(clk), .Q(\xmem_data[64][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][6]  ( .D(\xmem_inst/mem[118][6] ), .CK(
        clk), .Q(\xmem_data[118][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][6]  ( .D(\xmem_inst/mem[114][6] ), .CK(
        clk), .Q(\xmem_data[114][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[40][6]  ( .D(\xmem_inst/mem[40][6] ), .CK(clk), .Q(\xmem_data[40][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][6]  ( .D(\xmem_inst/mem[32][6] ), .CK(clk), .Q(\xmem_data[32][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][6]  ( .D(\xmem_inst/mem[86][6] ), .CK(clk), .Q(\xmem_data[86][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[16][0]  ( .D(\xmem_inst/mem[16][0] ), .CK(clk), .Q(\xmem_data[16][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][1]  ( .D(\xmem_inst/mem[88][1] ), .CK(clk), .Q(\xmem_data[88][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[84][1]  ( .D(\xmem_inst/mem[84][1] ), .CK(clk), .Q(\xmem_data[84][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[108][1]  ( .D(\xmem_inst/mem[108][1] ), .CK(
        clk), .Q(\xmem_data[108][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[104][1]  ( .D(\xmem_inst/mem[104][1] ), .CK(
        clk), .Q(\xmem_data[104][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[70][1]  ( .D(\xmem_inst/mem[70][1] ), .CK(clk), .Q(\xmem_data[70][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[46][1]  ( .D(\xmem_inst/mem[46][1] ), .CK(clk), .Q(\xmem_data[46][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][3]  ( .D(\xmem_inst/mem[102][3] ), .CK(
        clk), .Q(\xmem_data[102][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][3]  ( .D(\xmem_inst/mem[32][3] ), .CK(clk), .Q(\xmem_data[32][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][4]  ( .D(\xmem_inst/mem[32][4] ), .CK(clk), .Q(\xmem_data[32][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[50][4]  ( .D(\xmem_inst/mem[50][4] ), .CK(clk), .Q(\xmem_data[50][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[118][4]  ( .D(\xmem_inst/mem[118][4] ), .CK(
        clk), .Q(\xmem_data[118][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[102][5]  ( .D(\xmem_inst/mem[102][5] ), .CK(
        clk), .Q(\xmem_data[102][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][1]  ( .D(\xmem_inst/mem[114][1] ), .CK(
        clk), .Q(\xmem_data[114][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[5][0]  ( .D(\xmem_inst/mem[5][0] ), .CK(clk), 
        .Q(\xmem_data[5][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][1]  ( .D(\xmem_inst/mem[32][1] ), .CK(clk), .Q(\xmem_data[32][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][1]  ( .D(\xmem_inst/mem[83][1] ), .CK(clk), .Q(\xmem_data[83][1] ) );
  DFF_X2 \xmem_inst/data_out_reg[116][7]  ( .D(\xmem_inst/mem[116][7] ), .CK(
        clk), .Q(\xmem_data[116][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[110][7]  ( .D(\xmem_inst/mem[110][7] ), .CK(
        clk), .Q(\xmem_data[110][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][7]  ( .D(\xmem_inst/mem[114][7] ), .CK(
        clk), .Q(\xmem_data[114][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][0]  ( .D(\xmem_inst/mem[32][0] ), .CK(clk), .Q(\xmem_data[32][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[83][4]  ( .D(\xmem_inst/mem[83][4] ), .CK(clk), .Q(\xmem_data[83][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[65][4]  ( .D(\xmem_inst/mem[65][4] ), .CK(clk), .Q(\xmem_data[65][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[88][3]  ( .D(\xmem_inst/mem[88][3] ), .CK(clk), .Q(\xmem_data[88][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][3]  ( .D(\xmem_inst/mem[34][3] ), .CK(clk), .Q(\xmem_data[34][3] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][7]  ( .D(\xmem_inst/mem[82][7] ), .CK(clk), .Q(\xmem_data[82][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[66][7]  ( .D(\xmem_inst/mem[66][7] ), .CK(clk), .Q(\xmem_data[66][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[64][7]  ( .D(\xmem_inst/mem[64][7] ), .CK(clk), .Q(\xmem_data[64][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[82][5]  ( .D(\xmem_inst/mem[82][5] ), .CK(clk), .Q(\xmem_data[82][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[114][5]  ( .D(\xmem_inst/mem[114][5] ), .CK(
        clk), .Q(\xmem_data[114][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[13][4]  ( .D(\xmem_inst/mem[13][4] ), .CK(clk), .Q(\xmem_data[13][4] ) );
  DFF_X2 \xmem_inst/data_out_reg[51][6]  ( .D(\xmem_inst/mem[51][6] ), .CK(clk), .Q(\xmem_data[51][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[35][6]  ( .D(\xmem_inst/mem[35][6] ), .CK(clk), .Q(\xmem_data[35][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][5]  ( .D(\xmem_inst/mem[34][5] ), .CK(clk), .Q(\xmem_data[34][5] ) );
  DFF_X2 \xmem_inst/data_out_reg[54][7]  ( .D(\xmem_inst/mem[54][7] ), .CK(clk), .Q(\xmem_data[54][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][7]  ( .D(\xmem_inst/mem[34][7] ), .CK(clk), .Q(\xmem_data[34][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[32][7]  ( .D(\xmem_inst/mem[32][7] ), .CK(clk), .Q(\xmem_data[32][7] ) );
  DFF_X2 \xmem_inst/data_out_reg[120][6]  ( .D(\xmem_inst/mem[120][6] ), .CK(
        clk), .Q(\xmem_data[120][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[86][0]  ( .D(\xmem_inst/mem[86][0] ), .CK(clk), .Q(\xmem_data[86][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[7][0]  ( .D(\xmem_inst/mem[7][0] ), .CK(clk), 
        .Q(\xmem_data[7][0] ) );
  DFF_X2 \xmem_inst/data_out_reg[67][6]  ( .D(\xmem_inst/mem[67][6] ), .CK(clk), .Q(\xmem_data[67][6] ) );
  DFF_X2 \xmem_inst/data_out_reg[34][6]  ( .D(\xmem_inst/mem[34][6] ), .CK(clk), .Q(\xmem_data[34][6] ) );
  NAND3_X1 U3236 ( .A1(n11143), .A2(n11142), .A3(n11141), .ZN(n31996) );
  OR4_X1 U3237 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n8043) );
  OR4_X1 U3238 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n8098) );
  OR4_X1 U3239 ( .A1(n8019), .A2(n8018), .A3(n8017), .A4(n8016), .ZN(n8044) );
  NAND4_X1 U3240 ( .A1(n18239), .A2(n18238), .A3(n18237), .A4(n18236), .ZN(
        n33939) );
  NAND4_X1 U3241 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n33720)
         );
  OR4_X1 U3242 ( .A1(n8638), .A2(n8637), .A3(n8636), .A4(n8635), .ZN(n8639) );
  BUF_X1 U3243 ( .A(n8558), .Z(n3195) );
  BUF_X1 U3244 ( .A(n6234), .Z(n30219) );
  BUF_X1 U3245 ( .A(n8558), .Z(n3196) );
  BUF_X1 U3246 ( .A(n11850), .Z(n27814) );
  BUF_X1 U3247 ( .A(n8075), .Z(n28681) );
  BUF_X1 U3248 ( .A(n6281), .Z(n30251) );
  BUF_X1 U3249 ( .A(n8515), .Z(n3235) );
  BUF_X1 U3250 ( .A(n8513), .Z(n3243) );
  BUF_X1 U3251 ( .A(n8517), .Z(n3236) );
  BUF_X1 U3252 ( .A(n8519), .Z(n3237) );
  BUF_X1 U3253 ( .A(n6245), .Z(n30200) );
  BUF_X1 U3254 ( .A(n8503), .Z(n29865) );
  BUF_X1 U3255 ( .A(n8558), .Z(n3194) );
  BUF_X1 U3256 ( .A(n28111), .Z(n28165) );
  INV_X1 U3257 ( .A(n3123), .ZN(n3124) );
  BUF_X1 U3258 ( .A(n11454), .Z(n29583) );
  BUF_X1 U3259 ( .A(n11456), .Z(n29584) );
  BUF_X2 U3260 ( .A(n24625), .Z(n3203) );
  INV_X1 U3261 ( .A(n3118), .ZN(n3121) );
  INV_X1 U3262 ( .A(n27976), .ZN(n3327) );
  NAND4_X2 U3263 ( .A1(n27101), .A2(n27100), .A3(n27099), .A4(n27098), .ZN(
        n32937) );
  BUF_X1 U3264 ( .A(n32417), .Z(n3430) );
  BUF_X2 U3265 ( .A(n6247), .Z(n30256) );
  BUF_X2 U3266 ( .A(n36523), .Z(n3116) );
  BUF_X1 U3267 ( .A(n29389), .Z(n3117) );
  NAND4_X1 U3268 ( .A1(n30788), .A2(n30787), .A3(n30786), .A4(n30785), .ZN(
        n36523) );
  OR4_X2 U3269 ( .A1(n7492), .A2(n7491), .A3(n7490), .A4(n7489), .ZN(n7493) );
  BUF_X2 U3270 ( .A(n39053), .Z(n6586) );
  OR4_X2 U3271 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n8729) );
  NAND2_X2 U3272 ( .A1(n22150), .A2(n22149), .ZN(n32419) );
  INV_X2 U3273 ( .A(n28300), .ZN(n3118) );
  INV_X1 U3274 ( .A(n3118), .ZN(n3119) );
  INV_X2 U3275 ( .A(n3118), .ZN(n3120) );
  AOI21_X1 U3276 ( .B1(n7216), .B2(n6621), .A(n6816), .ZN(n6612) );
  BUF_X1 U3277 ( .A(n36442), .Z(n3122) );
  OR4_X2 U3278 ( .A1(n29561), .A2(n29563), .A3(n29562), .A4(n29564), .ZN(
        n29601) );
  INV_X1 U3279 ( .A(n8089), .ZN(n3123) );
  INV_X1 U3280 ( .A(n28741), .ZN(n3125) );
  INV_X2 U3281 ( .A(n3125), .ZN(n3126) );
  INV_X1 U3282 ( .A(n30942), .ZN(n3127) );
  INV_X1 U3283 ( .A(n3127), .ZN(n3128) );
  INV_X1 U3284 ( .A(n3127), .ZN(n3129) );
  INV_X1 U3285 ( .A(n30218), .ZN(n3130) );
  INV_X1 U3286 ( .A(n3130), .ZN(n3131) );
  INV_X1 U3287 ( .A(n3130), .ZN(n3132) );
  INV_X1 U3288 ( .A(n29401), .ZN(n3133) );
  INV_X1 U3289 ( .A(n3133), .ZN(n3134) );
  INV_X1 U3290 ( .A(n3133), .ZN(n3135) );
  INV_X1 U3291 ( .A(n30281), .ZN(n3136) );
  INV_X1 U3292 ( .A(n3136), .ZN(n3137) );
  INV_X1 U3293 ( .A(n3136), .ZN(n3138) );
  INV_X1 U3294 ( .A(n27762), .ZN(n3139) );
  INV_X2 U3295 ( .A(n3139), .ZN(n3140) );
  INV_X1 U3296 ( .A(n29620), .ZN(n3141) );
  INV_X2 U3297 ( .A(n3141), .ZN(n3142) );
  INV_X1 U3298 ( .A(n30758), .ZN(n3143) );
  INV_X2 U3299 ( .A(n3143), .ZN(n3144) );
  INV_X1 U3300 ( .A(n27817), .ZN(n3145) );
  INV_X1 U3301 ( .A(n3145), .ZN(n3146) );
  INV_X1 U3302 ( .A(n3145), .ZN(n3147) );
  INV_X1 U3303 ( .A(n27724), .ZN(n3148) );
  INV_X2 U3304 ( .A(n3148), .ZN(n3149) );
  INV_X1 U3305 ( .A(n29460), .ZN(n3150) );
  INV_X2 U3306 ( .A(n3150), .ZN(n3151) );
  INV_X1 U3307 ( .A(n30319), .ZN(n3152) );
  INV_X2 U3308 ( .A(n3152), .ZN(n3153) );
  INV_X1 U3309 ( .A(n11357), .ZN(n11350) );
  BUF_X2 U3310 ( .A(n4236), .Z(n13476) );
  INV_X2 U3311 ( .A(n4536), .ZN(n14933) );
  INV_X2 U3312 ( .A(n4254), .ZN(n13474) );
  BUF_X1 U3313 ( .A(n31276), .Z(n25707) );
  BUF_X2 U3314 ( .A(n30525), .Z(n3172) );
  BUF_X2 U3315 ( .A(n30525), .Z(n3171) );
  INV_X2 U3316 ( .A(n3331), .ZN(n3333) );
  BUF_X4 U3317 ( .A(n13474), .Z(n25514) );
  BUF_X2 U3318 ( .A(n29011), .Z(n3213) );
  BUF_X4 U3319 ( .A(n13188), .Z(n27516) );
  BUF_X1 U3320 ( .A(n15000), .Z(n29011) );
  BUF_X2 U3321 ( .A(n23794), .Z(n3207) );
  BUF_X1 U3322 ( .A(n14976), .Z(n30525) );
  BUF_X2 U3323 ( .A(n14912), .Z(n28492) );
  INV_X2 U3324 ( .A(n4237), .ZN(n14912) );
  INV_X2 U3325 ( .A(n4237), .ZN(n14970) );
  BUF_X2 U3326 ( .A(n10999), .Z(n20546) );
  BUF_X2 U3327 ( .A(n14991), .Z(n30295) );
  BUF_X4 U3328 ( .A(n14882), .Z(n25581) );
  INV_X2 U3329 ( .A(n4456), .ZN(n13487) );
  BUF_X2 U3330 ( .A(n13481), .Z(n29318) );
  BUF_X2 U3331 ( .A(n13481), .Z(n25435) );
  BUF_X2 U3332 ( .A(n13476), .Z(n25425) );
  AND3_X1 U3333 ( .A1(n3502), .A2(n3782), .A3(n8948), .ZN(n3154) );
  NAND4_X2 U3334 ( .A1(n16351), .A2(n16350), .A3(n16349), .A4(n16348), .ZN(
        n32787) );
  NAND4_X2 U3335 ( .A1(n17742), .A2(n17741), .A3(n17740), .A4(n17739), .ZN(
        n34626) );
  BUF_X4 U3336 ( .A(n11451), .Z(n29628) );
  AND2_X1 U3337 ( .A1(n8352), .A2(n8353), .ZN(n3155) );
  BUF_X2 U3338 ( .A(n11426), .Z(n3190) );
  BUF_X2 U3339 ( .A(n11426), .Z(n3191) );
  BUF_X2 U3340 ( .A(n11426), .Z(n3189) );
  BUF_X2 U3341 ( .A(n3181), .Z(n3188) );
  BUF_X2 U3342 ( .A(n3181), .Z(n3186) );
  AND4_X1 U3343 ( .A1(n28785), .A2(n28784), .A3(n28783), .A4(n28782), .ZN(
        n3156) );
  BUF_X2 U3344 ( .A(n3159), .Z(n3162) );
  BUF_X2 U3345 ( .A(n3159), .Z(n3163) );
  BUF_X2 U3346 ( .A(n3159), .Z(n3161) );
  BUF_X1 U3347 ( .A(n29770), .Z(n3157) );
  BUF_X4 U3348 ( .A(n29770), .Z(n3158) );
  OR4_X2 U3349 ( .A1(n15581), .A2(n15580), .A3(n15579), .A4(n15578), .ZN(
        n15582) );
  BUF_X4 U3350 ( .A(n14998), .Z(n24212) );
  BUF_X2 U3351 ( .A(n4177), .Z(n14998) );
  NOR2_X1 U3352 ( .A1(n8000), .A2(n11358), .ZN(n3159) );
  NOR2_X1 U3353 ( .A1(n8000), .A2(n11358), .ZN(n3160) );
  BUF_X4 U3354 ( .A(n3159), .Z(n3164) );
  BUF_X4 U3355 ( .A(n3160), .Z(n3165) );
  BUF_X4 U3356 ( .A(n11444), .Z(n3166) );
  BUF_X4 U3357 ( .A(n11444), .Z(n3167) );
  BUF_X4 U3358 ( .A(n11444), .Z(n3168) );
  NOR2_X1 U3359 ( .A1(n8000), .A2(n11358), .ZN(n11444) );
  CLKBUF_X1 U3360 ( .A(n30709), .Z(n3169) );
  BUF_X2 U3361 ( .A(n30709), .Z(n3170) );
  AOI22_X2 U3362 ( .A1(n12125), .A2(n28177), .B1(n12124), .B2(n28215), .ZN(
        n12126) );
  BUF_X2 U3363 ( .A(n14991), .Z(n30698) );
  BUF_X1 U3364 ( .A(n29474), .Z(n3173) );
  BUF_X2 U3365 ( .A(n29474), .Z(n3174) );
  BUF_X2 U3366 ( .A(n29475), .Z(n29438) );
  BUF_X4 U3367 ( .A(n10977), .Z(n28980) );
  BUF_X2 U3368 ( .A(n4526), .Z(n14981) );
  BUF_X2 U3369 ( .A(n27913), .Z(n3175) );
  BUF_X4 U3370 ( .A(n27913), .Z(n3176) );
  BUF_X1 U3371 ( .A(n24461), .Z(n3177) );
  BUF_X4 U3372 ( .A(n24461), .Z(n3178) );
  OAI21_X2 U3373 ( .B1(n35458), .B2(n35459), .A(n35457), .ZN(n35484) );
  BUF_X4 U3374 ( .A(n24523), .Z(n3179) );
  NOR2_X1 U3375 ( .A1(n11359), .A2(n8000), .ZN(n3180) );
  NOR2_X1 U3376 ( .A1(n11359), .A2(n8000), .ZN(n3181) );
  BUF_X4 U3377 ( .A(n3180), .Z(n3182) );
  BUF_X4 U3378 ( .A(n3180), .Z(n3183) );
  BUF_X4 U3379 ( .A(n3180), .Z(n3184) );
  BUF_X4 U3380 ( .A(n3180), .Z(n3185) );
  BUF_X4 U3381 ( .A(n3181), .Z(n3187) );
  NOR2_X1 U3382 ( .A1(n11359), .A2(n8000), .ZN(n11426) );
  CLKBUF_X1 U3383 ( .A(n30316), .Z(n3192) );
  BUF_X2 U3384 ( .A(n30316), .Z(n3193) );
  NAND2_X2 U3385 ( .A1(n6176), .A2(n11343), .ZN(n3378) );
  BUF_X4 U3386 ( .A(n14875), .Z(n28501) );
  BUF_X2 U3387 ( .A(n4247), .Z(n14875) );
  BUF_X1 U3388 ( .A(n27770), .Z(n3197) );
  BUF_X2 U3389 ( .A(n27770), .Z(n3198) );
  BUF_X2 U3390 ( .A(n6675), .Z(n3199) );
  BUF_X2 U3391 ( .A(n6675), .Z(n3200) );
  BUF_X2 U3392 ( .A(n6675), .Z(n3201) );
  AND2_X4 U3393 ( .A1(n4062), .A2(n4064), .ZN(n31263) );
  NOR2_X1 U3394 ( .A1(n6614), .A2(n6613), .ZN(n3202) );
  BUF_X2 U3395 ( .A(n8267), .Z(n28162) );
  INV_X2 U3396 ( .A(n3268), .ZN(n3269) );
  INV_X4 U3397 ( .A(n3373), .ZN(n3375) );
  INV_X2 U3398 ( .A(n3339), .ZN(n3342) );
  CLKBUF_X1 U3399 ( .A(n29189), .Z(n3204) );
  BUF_X2 U3400 ( .A(n29189), .Z(n3205) );
  BUF_X2 U3401 ( .A(n29189), .Z(n3206) );
  BUF_X4 U3402 ( .A(n23794), .Z(n3208) );
  BUF_X4 U3403 ( .A(n24523), .Z(n3209) );
  OR3_X2 U3404 ( .A1(n30122), .A2(n30121), .A3(n30120), .ZN(n36339) );
  BUF_X2 U3405 ( .A(n6246), .Z(n3210) );
  BUF_X2 U3406 ( .A(n6246), .Z(n3211) );
  BUF_X2 U3407 ( .A(n30259), .Z(n3420) );
  BUF_X2 U3408 ( .A(n29011), .Z(n3212) );
  BUF_X1 U3409 ( .A(n30171), .Z(n3214) );
  NOR2_X2 U3410 ( .A1(n3378), .A2(n6191), .ZN(n30171) );
  INV_X2 U3411 ( .A(n4489), .ZN(n14883) );
  BUF_X2 U3412 ( .A(n4404), .Z(n14999) );
  INV_X2 U3413 ( .A(n4516), .ZN(n14882) );
  BUF_X2 U3414 ( .A(n4248), .Z(n3215) );
  BUF_X2 U3415 ( .A(n4248), .Z(n3216) );
  BUF_X8 U3416 ( .A(n3215), .Z(n3217) );
  BUF_X8 U3417 ( .A(n3215), .Z(n3218) );
  BUF_X8 U3418 ( .A(n3215), .Z(n3219) );
  BUF_X8 U3419 ( .A(n3216), .Z(n3220) );
  BUF_X8 U3420 ( .A(n3216), .Z(n3221) );
  BUF_X8 U3421 ( .A(n3216), .Z(n3222) );
  BUF_X4 U3422 ( .A(n14933), .Z(n3358) );
  INV_X4 U3423 ( .A(n4037), .ZN(n14997) );
  BUF_X4 U3424 ( .A(n4478), .Z(n31276) );
  NAND4_X2 U3425 ( .A1(n19705), .A2(n19704), .A3(n19703), .A4(n19702), .ZN(
        n34624) );
  BUF_X1 U3426 ( .A(n15844), .Z(n29641) );
  CLKBUF_X1 U3427 ( .A(n6245), .Z(n30261) );
  BUF_X1 U3428 ( .A(n7903), .Z(n30654) );
  BUF_X1 U3429 ( .A(n11780), .Z(n27770) );
  BUF_X2 U3430 ( .A(n26878), .Z(n3223) );
  BUF_X2 U3431 ( .A(n26491), .Z(n3224) );
  BUF_X2 U3432 ( .A(n8518), .Z(n3225) );
  BUF_X1 U3433 ( .A(n8072), .Z(n28702) );
  BUF_X2 U3434 ( .A(n7640), .Z(n3226) );
  BUF_X2 U3435 ( .A(n8090), .Z(n3227) );
  INV_X1 U3436 ( .A(n3254), .ZN(n3256) );
  INV_X1 U3437 ( .A(n3268), .ZN(n3271) );
  INV_X1 U3438 ( .A(n3279), .ZN(n3281) );
  INV_X1 U3439 ( .A(n14890), .ZN(n3254) );
  INV_X2 U3440 ( .A(n3448), .ZN(n3228) );
  INV_X1 U3441 ( .A(n3423), .ZN(n3245) );
  INV_X2 U3442 ( .A(n3347), .ZN(n3229) );
  BUF_X1 U3443 ( .A(n14996), .Z(n20982) );
  BUF_X2 U3444 ( .A(n4078), .Z(n14926) );
  INV_X2 U3445 ( .A(n4242), .ZN(n13481) );
  INV_X1 U3446 ( .A(n8429), .ZN(n3230) );
  BUF_X1 U3447 ( .A(n13188), .Z(n25574) );
  INV_X2 U3448 ( .A(n4242), .ZN(n13452) );
  BUF_X4 U3449 ( .A(n14983), .Z(n3247) );
  BUF_X2 U3450 ( .A(n14928), .Z(n3231) );
  NAND2_X1 U3451 ( .A1(n4040), .A2(n4039), .ZN(n6179) );
  XNOR2_X1 U3452 ( .A(\fmem_data[24][3] ), .B(\fmem_data[24][4] ), .ZN(n34039)
         );
  AND2_X1 U3453 ( .A1(n37216), .A2(n37218), .ZN(n37214) );
  AND2_X1 U3454 ( .A1(n37216), .A2(n36012), .ZN(n37154) );
  OR2_X1 U3455 ( .A1(n37150), .A2(n37149), .ZN(n37216) );
  NOR2_X1 U3456 ( .A1(n37139), .A2(n37138), .ZN(n37264) );
  CLKBUF_X1 U3457 ( .A(n35471), .Z(n3355) );
  XNOR2_X1 U3458 ( .A(n36619), .B(n36618), .ZN(n36747) );
  CLKBUF_X1 U3459 ( .A(n34562), .Z(n3391) );
  OAI22_X1 U3460 ( .A1(n34359), .A2(n3662), .B1(n36242), .B2(n36241), .ZN(
        n36260) );
  NAND3_X1 U3461 ( .A1(n26147), .A2(n26146), .A3(n26145), .ZN(n33483) );
  XNOR2_X1 U3462 ( .A(n33321), .B(n34838), .ZN(n34826) );
  XNOR2_X1 U3463 ( .A(n33330), .B(n34832), .ZN(n34825) );
  OAI22_X1 U3464 ( .A1(n31014), .A2(n35493), .B1(n30447), .B2(n35494), .ZN(
        n26375) );
  OAI21_X1 U3465 ( .B1(n36339), .B2(n32292), .A(n32291), .ZN(n32327) );
  OAI22_X1 U3466 ( .A1(n33790), .A2(n34435), .B1(n34436), .B2(n34437), .ZN(
        n33910) );
  OAI22_X1 U3467 ( .A1(n3568), .A2(n33929), .B1(n32212), .B2(n36223), .ZN(
        n31877) );
  AND4_X1 U3468 ( .A1(n26687), .A2(n26686), .A3(n26685), .A4(n26684), .ZN(
        n34361) );
  OR3_X1 U3469 ( .A1(n6392), .A2(n6391), .A3(n6390), .ZN(n32597) );
  AND4_X2 U3470 ( .A1(n28264), .A2(n28263), .A3(n28262), .A4(n28261), .ZN(
        n36314) );
  OAI22_X1 U3471 ( .A1(n33778), .A2(n3577), .B1(n33777), .B2(n36196), .ZN(
        n33807) );
  OAI22_X1 U3472 ( .A1(n34042), .A2(n34039), .B1(n27582), .B2(n34041), .ZN(
        n31127) );
  NAND4_X1 U3473 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n35112) );
  NAND3_X1 U3474 ( .A1(n15403), .A2(n15402), .A3(n15401), .ZN(n32319) );
  AND2_X1 U3475 ( .A1(n30457), .A2(n30456), .ZN(n30476) );
  OAI22_X1 U3476 ( .A1(n32234), .A2(n34429), .B1(n32260), .B2(n34533), .ZN(
        n31392) );
  AOI21_X1 U3477 ( .B1(n36226), .B2(n3633), .A(n32152), .ZN(n26799) );
  OAI22_X1 U3478 ( .A1(n33040), .A2(n33643), .B1(n33183), .B2(n33642), .ZN(
        n17749) );
  NAND2_X1 U3479 ( .A1(n23477), .A2(n23476), .ZN(n33677) );
  OAI22_X1 U3480 ( .A1(n32536), .A2(n34535), .B1(n32714), .B2(n34537), .ZN(
        n31913) );
  NAND3_X1 U3481 ( .A1(n3723), .A2(n15015), .A3(n15014), .ZN(n31592) );
  NAND3_X1 U3482 ( .A1(n25245), .A2(n25244), .A3(n25243), .ZN(n35072) );
  OR2_X1 U3483 ( .A1(n16468), .A2(n16467), .ZN(n32612) );
  OAI22_X1 U3484 ( .A1(n33964), .A2(n33963), .B1(n33962), .B2(n33961), .ZN(
        n34000) );
  NAND4_X2 U3485 ( .A1(n29516), .A2(n29515), .A3(n29514), .A4(n29513), .ZN(
        n36315) );
  OAI22_X1 U3486 ( .A1(n25146), .A2(n35712), .B1(n32022), .B2(n35711), .ZN(
        n31646) );
  OR2_X1 U3487 ( .A1(n3267), .A2(n32752), .ZN(n32753) );
  NAND3_X1 U3488 ( .A1(n27972), .A2(n27971), .A3(n27970), .ZN(n34630) );
  OR2_X1 U3489 ( .A1(n35038), .A2(n3946), .ZN(n35283) );
  OAI21_X1 U3490 ( .B1(n29473), .B2(n29472), .A(n29471), .ZN(n29514) );
  NAND2_X1 U3491 ( .A1(n30012), .A2(n30011), .ZN(n36338) );
  NAND3_X1 U3492 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n31704) );
  NAND3_X1 U3493 ( .A1(n12714), .A2(n12713), .A3(n12712), .ZN(n32228) );
  NAND2_X1 U3494 ( .A1(n18631), .A2(n18630), .ZN(n31638) );
  NAND2_X1 U3495 ( .A1(n15115), .A2(n15114), .ZN(n32242) );
  NAND3_X1 U3496 ( .A1(n4268), .A2(n4267), .A3(n4266), .ZN(n32317) );
  NAND3_X1 U3497 ( .A1(n5867), .A2(n5866), .A3(n5865), .ZN(n32025) );
  AOI22_X1 U3498 ( .A1(n7882), .A2(n29471), .B1(n7881), .B2(n29511), .ZN(
        n32557) );
  NAND4_X1 U3499 ( .A1(n6074), .A2(n3721), .A3(n6073), .A4(n6072), .ZN(n31668)
         );
  NAND4_X1 U3500 ( .A1(n19415), .A2(n19414), .A3(n19413), .A4(n19412), .ZN(
        n33551) );
  NAND3_X1 U3501 ( .A1(n26369), .A2(n26368), .A3(n26367), .ZN(n33594) );
  NAND2_X1 U3502 ( .A1(n16565), .A2(n16564), .ZN(n31655) );
  OR2_X1 U3503 ( .A1(n33271), .A2(n3396), .ZN(n33272) );
  NAND3_X1 U3504 ( .A1(n3731), .A2(n13521), .A3(n13520), .ZN(n31511) );
  NAND4_X1 U3505 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n31489)
         );
  OR3_X1 U3506 ( .A1(n7704), .A2(n7703), .A3(n7702), .ZN(n31817) );
  OR3_X1 U3507 ( .A1(n4771), .A2(n4770), .A3(n4769), .ZN(n31957) );
  OAI211_X1 U3508 ( .C1(n13911), .C2(n25647), .A(n13910), .B(n13909), .ZN(
        n30451) );
  NAND3_X1 U3509 ( .A1(n5060), .A2(n5059), .A3(n5058), .ZN(n32543) );
  NAND4_X1 U3510 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n31798)
         );
  NAND3_X1 U3511 ( .A1(n3719), .A2(n28892), .A3(n28891), .ZN(n34531) );
  OR2_X1 U3512 ( .A1(n24589), .A2(n24588), .ZN(n34980) );
  NAND2_X1 U3513 ( .A1(n23572), .A2(n23571), .ZN(n33789) );
  NAND4_X1 U3514 ( .A1(n20487), .A2(n20486), .A3(n20485), .A4(n20484), .ZN(
        n33555) );
  OR4_X1 U3515 ( .A1(n30328), .A2(n30327), .A3(n30326), .A4(n30325), .ZN(
        n30330) );
  NOR2_X1 U3516 ( .A1(n28109), .A2(n3916), .ZN(n34588) );
  NAND4_X1 U3517 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n35340) );
  OR4_X1 U3518 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n8401) );
  OR3_X1 U3519 ( .A1(n6481), .A2(n6480), .A3(n6479), .ZN(n35122) );
  OR4_X1 U3520 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .ZN(n8231) );
  OR4_X1 U3521 ( .A1(n23913), .A2(n23912), .A3(n23911), .A4(n23910), .ZN(
        n23914) );
  NAND4_X1 U3522 ( .A1(n28635), .A2(n28634), .A3(n28633), .A4(n28632), .ZN(
        n32554) );
  NAND4_X1 U3523 ( .A1(n13110), .A2(n13109), .A3(n13108), .A4(n13107), .ZN(
        n33055) );
  NAND2_X1 U3524 ( .A1(n20706), .A2(n20705), .ZN(n34929) );
  NAND3_X1 U3525 ( .A1(n20005), .A2(n20004), .A3(n20003), .ZN(n33039) );
  NAND2_X1 U3526 ( .A1(n33465), .A2(n33466), .ZN(n34599) );
  NAND4_X2 U3527 ( .A1(n29843), .A2(n29842), .A3(n29841), .A4(n29840), .ZN(
        n36337) );
  NAND2_X1 U3528 ( .A1(n15496), .A2(n15495), .ZN(n31800) );
  NAND4_X1 U3529 ( .A1(n20285), .A2(n20284), .A3(n20283), .A4(n20282), .ZN(
        n33573) );
  NAND4_X1 U3530 ( .A1(n14572), .A2(n14571), .A3(n14570), .A4(n14569), .ZN(
        n35397) );
  NAND3_X1 U3531 ( .A1(n9685), .A2(n9684), .A3(n9683), .ZN(n31656) );
  OR4_X1 U3532 ( .A1(n12123), .A2(n12121), .A3(n12122), .A4(n12120), .ZN(
        n12124) );
  OR4_X1 U3533 ( .A1(n23645), .A2(n23644), .A3(n23643), .A4(n23642), .ZN(
        n23646) );
  OR3_X1 U3534 ( .A1(n9971), .A2(n9970), .A3(n9969), .ZN(n31799) );
  OR4_X1 U3535 ( .A1(n12081), .A2(n12079), .A3(n12080), .A4(n12078), .ZN(
        n12082) );
  NAND3_X1 U3536 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n31658) );
  OR4_X1 U3537 ( .A1(n23870), .A2(n23869), .A3(n23868), .A4(n23867), .ZN(
        n23871) );
  OR2_X1 U3538 ( .A1(n35005), .A2(n3937), .ZN(n35273) );
  NAND2_X1 U3539 ( .A1(n22977), .A2(n22976), .ZN(n32131) );
  NAND3_X1 U3540 ( .A1(n18917), .A2(n18916), .A3(n18915), .ZN(n32882) );
  NAND2_X1 U3541 ( .A1(n25475), .A2(n25474), .ZN(n35076) );
  OAI22_X1 U3542 ( .A1(n33799), .A2(n34039), .B1(n34041), .B2(n3651), .ZN(
        n33982) );
  NAND2_X1 U3543 ( .A1(n30631), .A2(n30630), .ZN(n32953) );
  NAND2_X1 U3544 ( .A1(n19904), .A2(n19903), .ZN(n32057) );
  NAND4_X1 U3545 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n31125) );
  AND2_X1 U3546 ( .A1(n34624), .A2(n32119), .ZN(n32687) );
  NAND3_X1 U3547 ( .A1(n29346), .A2(n3718), .A3(n29345), .ZN(n32899) );
  NAND3_X1 U3548 ( .A1(n25597), .A2(n25596), .A3(n25595), .ZN(n35074) );
  NAND4_X1 U3549 ( .A1(n28531), .A2(n28530), .A3(n28529), .A4(n28528), .ZN(
        n36245) );
  OR2_X1 U3550 ( .A1(n18069), .A2(n24151), .ZN(n18141) );
  OR4_X1 U3551 ( .A1(n13952), .A2(n13951), .A3(n13950), .A4(n13949), .ZN(
        n13953) );
  OR4_X1 U3552 ( .A1(n30006), .A2(n30005), .A3(n30004), .A4(n30003), .ZN(
        n30008) );
  OR4_X1 U3553 ( .A1(n3927), .A2(n13714), .A3(n13713), .A4(n13712), .ZN(n31492) );
  NAND4_X1 U3554 ( .A1(n23827), .A2(n23826), .A3(n23825), .A4(n23824), .ZN(
        n35324) );
  OR3_X1 U3555 ( .A1(n22641), .A2(n22640), .A3(n22639), .ZN(n33967) );
  OAI211_X1 U3556 ( .C1(n22548), .C2(n29341), .A(n22547), .B(n22546), .ZN(
        n32427) );
  NAND3_X1 U3557 ( .A1(n17554), .A2(n17553), .A3(n17552), .ZN(n36299) );
  NAND3_X1 U3558 ( .A1(n4576), .A2(n4575), .A3(n4574), .ZN(n31161) );
  NAND4_X1 U3559 ( .A1(n27303), .A2(n27302), .A3(n27301), .A4(n27300), .ZN(
        n32596) );
  NAND3_X1 U3560 ( .A1(n16752), .A2(n16751), .A3(n16750), .ZN(n35357) );
  OAI211_X1 U3561 ( .C1(n17850), .C2(n22298), .A(n17849), .B(n17848), .ZN(
        n33556) );
  NAND2_X1 U3562 ( .A1(n21672), .A2(n21671), .ZN(n36200) );
  OR4_X1 U3563 ( .A1(n24915), .A2(n24914), .A3(n24913), .A4(n24912), .ZN(
        n24916) );
  OR3_X1 U3564 ( .A1(n4965), .A2(n4964), .A3(n4963), .ZN(n32321) );
  OR3_X1 U3565 ( .A1(n13014), .A2(n13013), .A3(n13012), .ZN(n31895) );
  OAI21_X1 U3566 ( .B1(n29839), .B2(n29838), .A(n29837), .ZN(n29840) );
  NAND4_X1 U3567 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n32014)
         );
  OR4_X1 U3568 ( .A1(n26018), .A2(n26016), .A3(n26017), .A4(n26015), .ZN(
        n26019) );
  OR4_X1 U3569 ( .A1(n7067), .A2(n7066), .A3(n7065), .A4(n7064), .ZN(n7093) );
  OR4_X1 U3570 ( .A1(n25976), .A2(n25975), .A3(n25974), .A4(n25973), .ZN(
        n25977) );
  AND2_X1 U3571 ( .A1(n36101), .A2(n21284), .ZN(n33943) );
  OR4_X1 U3572 ( .A1(n26247), .A2(n26246), .A3(n26245), .A4(n26244), .ZN(
        n26248) );
  OAI21_X1 U3573 ( .B1(n29797), .B2(n29796), .A(n29795), .ZN(n29841) );
  OAI21_X1 U3574 ( .B1(n29760), .B2(n29759), .A(n29758), .ZN(n29842) );
  NAND4_X1 U3575 ( .A1(n20094), .A2(n20093), .A3(n20092), .A4(n20091), .ZN(
        n33214) );
  OR2_X1 U3576 ( .A1(n9660), .A2(n20188), .ZN(n9684) );
  NAND2_X1 U3577 ( .A1(n30978), .A2(n30977), .ZN(n36312) );
  NAND3_X1 U3578 ( .A1(n6584), .A2(n6583), .A3(n6582), .ZN(n35102) );
  OR4_X1 U3579 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7040) );
  NAND4_X1 U3580 ( .A1(n4469), .A2(n4468), .A3(n4467), .A4(n4466), .ZN(n35405)
         );
  NAND3_X1 U3581 ( .A1(n11048), .A2(n11047), .A3(n11046), .ZN(n31995) );
  NAND4_X1 U3582 ( .A1(n9297), .A2(n9296), .A3(n9295), .A4(n9294), .ZN(n35336)
         );
  NAND4_X1 U3583 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n33743) );
  NAND4_X1 U3584 ( .A1(n5454), .A2(n5453), .A3(n5452), .A4(n5451), .ZN(n32617)
         );
  OR4_X1 U3585 ( .A1(n18403), .A2(n18402), .A3(n18401), .A4(n18400), .ZN(
        n18426) );
  NAND4_X1 U3586 ( .A1(n20839), .A2(n20838), .A3(n20837), .A4(n20836), .ZN(
        n30156) );
  NAND3_X1 U3587 ( .A1(n25837), .A2(n25836), .A3(n25835), .ZN(n35328) );
  NAND4_X1 U3588 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n31657)
         );
  OR4_X1 U3589 ( .A1(n7261), .A2(n7262), .A3(n7263), .A4(n7260), .ZN(n7265) );
  OR4_X1 U3590 ( .A1(n18450), .A2(n18449), .A3(n18448), .A4(n18447), .ZN(
        n18451) );
  OR4_X1 U3591 ( .A1(n15538), .A2(n15537), .A3(n15536), .A4(n15535), .ZN(
        n15539) );
  OAI21_X1 U3592 ( .B1(n17694), .B2(n17693), .A(n29343), .ZN(n17741) );
  NAND4_X2 U3593 ( .A1(n20612), .A2(n20611), .A3(n20610), .A4(n20609), .ZN(
        n34615) );
  OR4_X1 U3594 ( .A1(n18423), .A2(n18424), .A3(n18422), .A4(n18421), .ZN(
        n18425) );
  NAND3_X1 U3595 ( .A1(n31381), .A2(n31380), .A3(n31379), .ZN(n36112) );
  OR4_X1 U3596 ( .A1(n14790), .A2(n14789), .A3(n14787), .A4(n14788), .ZN(
        n14791) );
  OR4_X1 U3597 ( .A1(n7420), .A2(n7419), .A3(n7418), .A4(n7417), .ZN(n7445) );
  OR3_X1 U3598 ( .A1(n29828), .A2(n29827), .A3(n29826), .ZN(n29839) );
  OR4_X1 U3599 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n8144) );
  NAND4_X1 U3600 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n33451) );
  OR2_X1 U3601 ( .A1(n5959), .A2(n5958), .ZN(n32586) );
  OR3_X1 U3602 ( .A1(n29752), .A2(n29751), .A3(n29750), .ZN(n29760) );
  OR3_X1 U3603 ( .A1(n29784), .A2(n29783), .A3(n29782), .ZN(n29797) );
  NAND4_X2 U3604 ( .A1(n21283), .A2(n21282), .A3(n21281), .A4(n21280), .ZN(
        n36101) );
  OR4_X1 U3605 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11840) );
  NAND4_X2 U3606 ( .A1(n17274), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n36228) );
  OR4_X1 U3607 ( .A1(n23020), .A2(n23019), .A3(n23018), .A4(n23017), .ZN(
        n23021) );
  OR4_X1 U3608 ( .A1(n12860), .A2(n12859), .A3(n12858), .A4(n12857), .ZN(
        n12861) );
  NAND4_X1 U3609 ( .A1(n15308), .A2(n15307), .A3(n15306), .A4(n15305), .ZN(
        n32582) );
  OR4_X1 U3610 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10854) );
  OR4_X1 U3611 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11797) );
  OR4_X1 U3612 ( .A1(n22405), .A2(n22404), .A3(n22403), .A4(n22402), .ZN(
        n22406) );
  OR4_X1 U3613 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n7837) );
  NAND4_X2 U3614 ( .A1(n22773), .A2(n22772), .A3(n22771), .A4(n22770), .ZN(
        n34623) );
  NAND4_X1 U3615 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n35326) );
  OR4_X1 U3616 ( .A1(n10903), .A2(n10901), .A3(n10902), .A4(n10900), .ZN(
        n10904) );
  OR4_X1 U3617 ( .A1(n14287), .A2(n14286), .A3(n14285), .A4(n14284), .ZN(
        n35338) );
  OR4_X1 U3618 ( .A1(n7442), .A2(n7441), .A3(n7443), .A4(n7440), .ZN(n7444) );
  OR4_X1 U3619 ( .A1(n18365), .A2(n18363), .A3(n18364), .A4(n18362), .ZN(
        n18383) );
  OR4_X1 U3620 ( .A1(n24009), .A2(n24008), .A3(n24007), .A4(n24006), .ZN(
        n24010) );
  OR4_X1 U3621 ( .A1(n7290), .A2(n7288), .A3(n7289), .A4(n7287), .ZN(n7293) );
  OR4_X1 U3622 ( .A1(n23043), .A2(n23042), .A3(n23041), .A4(n23040), .ZN(
        n23044) );
  OR3_X1 U3623 ( .A1(n22021), .A2(n22020), .A3(n22019), .ZN(n22024) );
  BUF_X1 U3624 ( .A(n30171), .Z(n30300) );
  BUF_X1 U3625 ( .A(n30171), .Z(n30192) );
  OR4_X1 U3626 ( .A1(n8879), .A2(n8878), .A3(n8877), .A4(n8876), .ZN(n8880) );
  BUF_X1 U3627 ( .A(n30259), .Z(n30317) );
  OR4_X1 U3628 ( .A1(n21626), .A2(n21625), .A3(n21624), .A4(n3972), .ZN(n21627) );
  AND4_X1 U3629 ( .A1(n26659), .A2(n26658), .A3(n26657), .A4(n26656), .ZN(
        n26660) );
  OR4_X1 U3630 ( .A1(n22178), .A2(n22177), .A3(n22176), .A4(n22175), .ZN(
        n22181) );
  OAI21_X1 U3631 ( .B1(n22737), .B2(n22736), .A(n22735), .ZN(n22771) );
  OR4_X1 U3632 ( .A1(n20385), .A2(n20384), .A3(n20383), .A4(n20382), .ZN(
        n20387) );
  OAI21_X1 U3633 ( .B1(n17435), .B2(n17434), .A(n24204), .ZN(n17460) );
  AND2_X1 U3634 ( .A1(n5160), .A2(n5159), .ZN(n20606) );
  OAI21_X1 U3635 ( .B1(n22700), .B2(n22699), .A(n22698), .ZN(n22772) );
  OR3_X1 U3636 ( .A1(n22726), .A2(n22725), .A3(n22724), .ZN(n22737) );
  OR4_X1 U3637 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12388) );
  OR4_X1 U3638 ( .A1(n18716), .A2(n18715), .A3(n18714), .A4(n18713), .ZN(
        n18717) );
  OR3_X1 U3639 ( .A1(n18749), .A2(n18748), .A3(n18747), .ZN(n18750) );
  OR3_X1 U3640 ( .A1(n28283), .A2(n28282), .A3(n28281), .ZN(n28290) );
  BUF_X1 U3641 ( .A(n8267), .Z(n28243) );
  BUF_X1 U3642 ( .A(n8266), .Z(n28244) );
  OR2_X1 U3643 ( .A1(n17433), .A2(n17432), .ZN(n17434) );
  OR2_X1 U3644 ( .A1(n17456), .A2(n17455), .ZN(n17457) );
  OAI21_X1 U3645 ( .B1(n28326), .B2(n28325), .A(n28324), .ZN(n28399) );
  BUF_X1 U3646 ( .A(n8266), .Z(n28163) );
  OAI21_X1 U3647 ( .B1(n28363), .B2(n28362), .A(n28361), .ZN(n28398) );
  BUF_X1 U3648 ( .A(n28111), .Z(n28196) );
  BUF_X1 U3649 ( .A(n8267), .Z(n28194) );
  BUF_X2 U3650 ( .A(n8464), .Z(n29976) );
  BUF_X1 U3651 ( .A(n11700), .Z(n29854) );
  BUF_X1 U3652 ( .A(n8489), .Z(n29855) );
  BUF_X1 U3653 ( .A(n8497), .Z(n29982) );
  BUF_X1 U3654 ( .A(n8496), .Z(n29980) );
  OR4_X1 U3655 ( .A1(n6531), .A2(n6530), .A3(n6529), .A4(n6528), .ZN(n6532) );
  BUF_X1 U3656 ( .A(n6247), .Z(n30316) );
  OR4_X1 U3657 ( .A1(n15302), .A2(n15301), .A3(n15300), .A4(n15299), .ZN(
        n15303) );
  INV_X1 U3658 ( .A(n20515), .ZN(n3232) );
  BUF_X1 U3659 ( .A(n7903), .Z(n27832) );
  AND2_X1 U3660 ( .A1(n4437), .A2(n4463), .ZN(n22735) );
  BUF_X1 U3661 ( .A(n8507), .Z(n29991) );
  BUF_X1 U3662 ( .A(n8518), .Z(n29880) );
  BUF_X1 U3663 ( .A(n8507), .Z(n29869) );
  BUF_X1 U3664 ( .A(n8506), .Z(n29919) );
  BUF_X1 U3665 ( .A(n8537), .Z(n29920) );
  OR4_X1 U3666 ( .A1(n18136), .A2(n18135), .A3(n18134), .A4(n18133), .ZN(
        n18137) );
  OR4_X1 U3667 ( .A1(n21419), .A2(n21418), .A3(n21417), .A4(n21416), .ZN(
        n21420) );
  OR4_X1 U3668 ( .A1(n13304), .A2(n13303), .A3(n13302), .A4(n13301), .ZN(
        n13305) );
  BUF_X1 U3669 ( .A(n11455), .Z(n29659) );
  AND2_X1 U3670 ( .A1(n5760), .A2(n5759), .ZN(n20765) );
  BUF_X2 U3671 ( .A(n8253), .Z(n3233) );
  OR3_X1 U3672 ( .A1(n28353), .A2(n28352), .A3(n28351), .ZN(n28363) );
  OR3_X1 U3673 ( .A1(n28316), .A2(n28315), .A3(n28314), .ZN(n28326) );
  BUF_X1 U3674 ( .A(n11476), .Z(n29617) );
  NOR2_X1 U3675 ( .A1(n8067), .A2(n8045), .ZN(n28662) );
  AND2_X1 U3676 ( .A1(n8302), .A2(n8303), .ZN(n28177) );
  BUF_X1 U3677 ( .A(n8293), .Z(n28206) );
  CLKBUF_X1 U3678 ( .A(n11453), .Z(n29655) );
  BUF_X1 U3679 ( .A(n7903), .Z(n30707) );
  BUF_X1 U3680 ( .A(n11561), .Z(n29568) );
  NOR2_X1 U3681 ( .A1(n5759), .A2(n5760), .ZN(n20833) );
  BUF_X2 U3682 ( .A(n8520), .Z(n3234) );
  BUF_X2 U3683 ( .A(n6680), .Z(n16979) );
  AND2_X1 U3684 ( .A1(n5862), .A2(n5838), .ZN(n31376) );
  BUF_X2 U3685 ( .A(n8516), .Z(n3238) );
  BUF_X2 U3686 ( .A(n11438), .Z(n3239) );
  AND2_X1 U3687 ( .A1(n7090), .A2(n7091), .ZN(n30782) );
  NOR2_X1 U3688 ( .A1(n8924), .A2(n8902), .ZN(n30628) );
  BUF_X1 U3689 ( .A(n7452), .Z(n29497) );
  BUF_X2 U3690 ( .A(n8259), .Z(n3240) );
  BUF_X2 U3691 ( .A(n8258), .Z(n3241) );
  BUF_X1 U3692 ( .A(n8074), .Z(n29462) );
  INV_X1 U3693 ( .A(n3339), .ZN(n3341) );
  BUF_X2 U3694 ( .A(n8514), .Z(n3242) );
  OR2_X1 U3695 ( .A1(n8448), .A2(n3230), .ZN(n8430) );
  NOR2_X1 U3696 ( .A1(n6067), .A2(n6066), .ZN(n24204) );
  NOR2_X1 U3697 ( .A1(n5360), .A2(n5336), .ZN(n29041) );
  BUF_X2 U3698 ( .A(n8080), .Z(n3244) );
  BUF_X1 U3699 ( .A(n8074), .Z(n27805) );
  BUF_X2 U3700 ( .A(n11439), .Z(n27754) );
  BUF_X1 U3701 ( .A(n7691), .Z(n29785) );
  NOR2_X1 U3702 ( .A1(n7091), .A2(n7090), .ZN(n30704) );
  BUF_X1 U3703 ( .A(n29475), .Z(n29397) );
  INV_X1 U3704 ( .A(n3448), .ZN(n3449) );
  INV_X1 U3705 ( .A(n3336), .ZN(n3338) );
  INV_X1 U3706 ( .A(n3327), .ZN(n3329) );
  INV_X1 U3707 ( .A(n3411), .ZN(n3414) );
  INV_X1 U3708 ( .A(n3347), .ZN(n3348) );
  INV_X1 U3709 ( .A(n3279), .ZN(n3282) );
  INV_X1 U3710 ( .A(n3268), .ZN(n3270) );
  INV_X1 U3711 ( .A(n3432), .ZN(n3384) );
  NOR2_X1 U3712 ( .A1(n6695), .A2(n6669), .ZN(n16966) );
  INV_X2 U3713 ( .A(n3432), .ZN(n3434) );
  INV_X1 U3714 ( .A(n3304), .ZN(n3306) );
  INV_X1 U3715 ( .A(n3304), .ZN(n3318) );
  INV_X1 U3716 ( .A(n3331), .ZN(n3334) );
  INV_X1 U3717 ( .A(n3268), .ZN(n3308) );
  INV_X1 U3718 ( .A(n3373), .ZN(n3374) );
  OR2_X1 U3719 ( .A1(n11368), .A2(n7005), .ZN(n11344) );
  BUF_X2 U3720 ( .A(n10802), .Z(n30766) );
  NAND2_X1 U3721 ( .A1(n11368), .A2(n11357), .ZN(n11363) );
  NOR2_X1 U3722 ( .A1(n8005), .A2(n7010), .ZN(n7446) );
  OR2_X1 U3723 ( .A1(n15009), .A2(n14967), .ZN(n15043) );
  INV_X1 U3724 ( .A(n3349), .ZN(n3352) );
  INV_X1 U3725 ( .A(n3385), .ZN(n3387) );
  NAND2_X1 U3726 ( .A1(n3230), .A2(n8448), .ZN(n8435) );
  INV_X1 U3727 ( .A(n14990), .ZN(n3339) );
  INV_X1 U3728 ( .A(n14991), .ZN(n3373) );
  CLKBUF_X1 U3729 ( .A(n11362), .Z(n3457) );
  CLKBUF_X1 U3730 ( .A(n6189), .Z(n3443) );
  INV_X1 U3731 ( .A(n14974), .ZN(n3268) );
  INV_X1 U3732 ( .A(n24466), .ZN(n3336) );
  BUF_X2 U3733 ( .A(n10977), .Z(n30891) );
  BUF_X1 U3734 ( .A(n14989), .Z(n25491) );
  OAI211_X1 U3735 ( .C1(n8415), .C2(n8414), .A(n8413), .B(n8412), .ZN(n8448)
         );
  INV_X1 U3736 ( .A(n14991), .ZN(n3279) );
  BUF_X2 U3737 ( .A(n13436), .Z(n30614) );
  INV_X1 U3738 ( .A(n17032), .ZN(n3385) );
  INV_X1 U3739 ( .A(n28077), .ZN(n3432) );
  NAND2_X1 U3740 ( .A1(n29180), .A2(\xmem_data[20][0] ), .ZN(n27340) );
  BUF_X1 U3741 ( .A(n4253), .Z(n13469) );
  BUF_X1 U3742 ( .A(n4177), .Z(n14934) );
  INV_X1 U3743 ( .A(n4516), .ZN(n14973) );
  BUF_X1 U3744 ( .A(n4158), .Z(n14972) );
  BUF_X1 U3745 ( .A(n4158), .Z(n14881) );
  CLKBUF_X1 U3746 ( .A(n7599), .Z(n7601) );
  BUF_X2 U3747 ( .A(n4253), .Z(n14989) );
  BUF_X1 U3748 ( .A(n4253), .Z(n14925) );
  BUF_X2 U3749 ( .A(n13420), .Z(n30901) );
  BUF_X1 U3750 ( .A(n31276), .Z(n30551) );
  BUF_X2 U3751 ( .A(n11362), .Z(n3246) );
  BUF_X2 U3752 ( .A(n4527), .Z(n13420) );
  INV_X1 U3753 ( .A(n4536), .ZN(n14996) );
  BUF_X4 U3754 ( .A(n4478), .Z(n27447) );
  BUF_X1 U3755 ( .A(n4526), .Z(n11008) );
  INV_X2 U3756 ( .A(n6179), .ZN(n29187) );
  INV_X1 U3757 ( .A(n4254), .ZN(n14928) );
  BUF_X4 U3758 ( .A(n4478), .Z(n25604) );
  INV_X1 U3759 ( .A(n4444), .ZN(n15000) );
  INV_X2 U3760 ( .A(n6179), .ZN(n3464) );
  BUF_X4 U3761 ( .A(n4478), .Z(n25422) );
  AND2_X2 U3762 ( .A1(n4040), .A2(n4062), .ZN(n4158) );
  AND2_X1 U3763 ( .A1(n6178), .A2(n6173), .ZN(n6177) );
  NAND2_X1 U3764 ( .A1(n4025), .A2(n4038), .ZN(n13132) );
  AND2_X1 U3765 ( .A1(n4024), .A2(n8409), .ZN(n4062) );
  OR2_X1 U3766 ( .A1(n10288), .A2(n4080), .ZN(n4444) );
  OR2_X1 U3767 ( .A1(n4065), .A2(n4058), .ZN(n4399) );
  INV_X1 U3768 ( .A(n6173), .ZN(n3248) );
  INV_X1 U3769 ( .A(n4391), .ZN(n37199) );
  XNOR2_X1 U3770 ( .A(\fmem_data[5][1] ), .B(\fmem_data[5][2] ), .ZN(n33850)
         );
  XNOR2_X1 U3771 ( .A(\fmem_data[9][6] ), .B(\fmem_data[9][5] ), .ZN(n35726)
         );
  XNOR2_X1 U3772 ( .A(\fmem_data[22][3] ), .B(\fmem_data[22][4] ), .ZN(n33963)
         );
  XNOR2_X1 U3773 ( .A(\fmem_data[31][6] ), .B(\fmem_data[31][5] ), .ZN(n35663)
         );
  XNOR2_X1 U3774 ( .A(\fmem_data[1][6] ), .B(\fmem_data[1][5] ), .ZN(n35701)
         );
  XNOR2_X1 U3775 ( .A(\fmem_data[21][6] ), .B(\fmem_data[21][5] ), .ZN(n35508)
         );
  XNOR2_X1 U3776 ( .A(\fmem_data[2][2] ), .B(\fmem_data[2][1] ), .ZN(n33797)
         );
  BUF_X1 U3777 ( .A(N345), .Z(n3402) );
  XNOR2_X1 U3778 ( .A(\fmem_data[0][4] ), .B(\fmem_data[0][3] ), .ZN(n33643)
         );
  XNOR2_X1 U3779 ( .A(\fmem_data[26][2] ), .B(\fmem_data[26][1] ), .ZN(n32780)
         );
  XNOR2_X1 U3780 ( .A(\fmem_data[8][6] ), .B(\fmem_data[8][5] ), .ZN(n35730)
         );
  XNOR2_X1 U3781 ( .A(\fmem_data[30][2] ), .B(\fmem_data[30][1] ), .ZN(n34435)
         );
  XNOR2_X1 U3782 ( .A(\fmem_data[14][1] ), .B(\fmem_data[14][2] ), .ZN(n33741)
         );
  XNOR2_X1 U3783 ( .A(\fmem_data[13][3] ), .B(\fmem_data[13][4] ), .ZN(n35182)
         );
  XNOR2_X1 U3784 ( .A(\fmem_data[28][2] ), .B(\fmem_data[28][1] ), .ZN(n33855)
         );
  XNOR2_X1 U3785 ( .A(\fmem_data[9][4] ), .B(\fmem_data[9][3] ), .ZN(n35041)
         );
  XNOR2_X1 U3786 ( .A(\fmem_data[26][6] ), .B(\fmem_data[26][5] ), .ZN(n35712)
         );
  XNOR2_X1 U3787 ( .A(\fmem_data[1][4] ), .B(\fmem_data[1][3] ), .ZN(n34942)
         );
  BUF_X1 U3788 ( .A(n11436), .Z(n3249) );
  NAND4_X1 U3789 ( .A1(n3250), .A2(n3251), .A3(n3252), .A4(n3253), .ZN(n8304)
         );
  AND4_X1 U3790 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), .ZN(n3250)
         );
  AND4_X1 U3791 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n3251)
         );
  AND4_X1 U3792 ( .A1(n8297), .A2(n8296), .A3(n8295), .A4(n8294), .ZN(n3252)
         );
  AND4_X1 U3793 ( .A1(n8301), .A2(n8300), .A3(n8299), .A4(n8298), .ZN(n3253)
         );
  NAND4_X1 U3794 ( .A1(n25047), .A2(n25046), .A3(n25045), .A4(n25044), .ZN(
        n32174) );
  INV_X1 U3795 ( .A(n3254), .ZN(n3255) );
  BUF_X2 U3796 ( .A(n7282), .Z(n29404) );
  NAND2_X1 U3797 ( .A1(n15585), .A2(n15584), .ZN(n3257) );
  AOI22_X1 U3798 ( .A1(n11798), .A2(n27801), .B1(n27839), .B2(n11797), .ZN(
        n3258) );
  XNOR2_X1 U3799 ( .A(n14874), .B(n34869), .ZN(n3259) );
  OAI22_X2 U3800 ( .A1(n23925), .A2(n35634), .B1(n24835), .B2(n35633), .ZN(
        n34869) );
  NAND3_X2 U3801 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n35110) );
  NAND4_X1 U3802 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n3260) );
  NAND2_X1 U3803 ( .A1(n3395), .A2(n3443), .ZN(n3261) );
  NAND4_X1 U3804 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), .ZN(n3262)
         );
  NAND4_X1 U3805 ( .A1(n3263), .A2(n3264), .A3(n3265), .A4(n3266), .ZN(n12083)
         );
  AND4_X1 U3806 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n3263) );
  AND4_X1 U3807 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n3264) );
  AND4_X1 U3808 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n3265) );
  AND4_X1 U3809 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n3266) );
  AND2_X1 U3810 ( .A1(n33725), .A2(n3678), .ZN(n3267) );
  BUF_X2 U3811 ( .A(n7659), .Z(n29709) );
  NAND3_X1 U3812 ( .A1(n12044), .A2(n12043), .A3(n12042), .ZN(n3272) );
  NAND3_X1 U3813 ( .A1(n12044), .A2(n12043), .A3(n12042), .ZN(n31386) );
  NOR2_X1 U3814 ( .A1(n37232), .A2(n3370), .ZN(n3273) );
  BUF_X4 U3815 ( .A(n7658), .Z(n29707) );
  BUF_X2 U3816 ( .A(n7275), .Z(n29419) );
  OR2_X1 U3817 ( .A1(n32189), .A2(n22359), .ZN(n29521) );
  AOI22_X1 U3818 ( .A1(n7838), .A2(n29428), .B1(n7837), .B2(n29376), .ZN(n3274) );
  AOI22_X1 U3819 ( .A1(n7838), .A2(n29428), .B1(n7837), .B2(n29376), .ZN(n3275) );
  AOI22_X1 U3820 ( .A1(n7838), .A2(n29428), .B1(n7837), .B2(n29376), .ZN(
        n32560) );
  NAND4_X1 U3821 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n3276)
         );
  NAND4_X1 U3822 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n31220)
         );
  BUF_X2 U3823 ( .A(n14926), .Z(n24697) );
  XNOR2_X1 U3824 ( .A(n31854), .B(n35433), .ZN(n3277) );
  NAND4_X1 U3825 ( .A1(n24014), .A2(n24013), .A3(n24012), .A4(n24011), .ZN(
        n3278) );
  NAND4_X1 U3826 ( .A1(n24014), .A2(n24013), .A3(n24012), .A4(n24011), .ZN(
        n31893) );
  NAND4_X2 U3827 ( .A1(n15695), .A2(n15694), .A3(n15693), .A4(n15692), .ZN(
        n32936) );
  INV_X1 U3828 ( .A(n3279), .ZN(n3280) );
  AND2_X1 U3829 ( .A1(n36433), .A2(n36432), .ZN(n3283) );
  AND2_X1 U3830 ( .A1(n4391), .A2(\add_x_2/A[0] ), .ZN(n6172) );
  BUF_X4 U3831 ( .A(n11489), .Z(n28136) );
  FA_X1 U3832 ( .A(n35468), .B(n35467), .CI(n35466), .S(n3284) );
  BUF_X4 U3833 ( .A(n7282), .Z(n29500) );
  BUF_X4 U3834 ( .A(n11489), .Z(n29788) );
  NAND2_X1 U3835 ( .A1(n29231), .A2(\xmem_data[96][6] ), .ZN(n3285) );
  NAND2_X1 U3836 ( .A1(n25450), .A2(\xmem_data[97][6] ), .ZN(n3286) );
  AND2_X1 U3837 ( .A1(n3285), .A2(n3286), .ZN(n11082) );
  XOR2_X1 U3838 ( .A(n33534), .B(n33536), .Z(n3287) );
  XOR2_X1 U3839 ( .A(n33535), .B(n3287), .Z(n36395) );
  NAND2_X1 U3840 ( .A1(n33535), .A2(n33534), .ZN(n3288) );
  NAND2_X1 U3841 ( .A1(n33535), .A2(n33536), .ZN(n3289) );
  NAND2_X1 U3842 ( .A1(n33534), .A2(n33536), .ZN(n3290) );
  NAND3_X1 U3843 ( .A1(n3288), .A2(n3289), .A3(n3290), .ZN(n33478) );
  BUF_X4 U3844 ( .A(n14928), .Z(n25450) );
  BUF_X4 U3845 ( .A(n13476), .Z(n28298) );
  AOI21_X1 U3846 ( .B1(n10976), .B2(n25790), .A(n10975), .ZN(n11048) );
  NAND2_X1 U3847 ( .A1(n13405), .A2(n13404), .ZN(n31664) );
  NAND2_X1 U3848 ( .A1(n14087), .A2(n14086), .ZN(n31892) );
  OAI211_X1 U3849 ( .C1(n3715), .C2(n11669), .A(n11668), .B(n11667), .ZN(
        n32938) );
  NAND2_X1 U3850 ( .A1(n11754), .A2(n11753), .ZN(n32442) );
  XNOR2_X1 U3851 ( .A(\fmem_data[5][4] ), .B(\fmem_data[5][3] ), .ZN(n33859)
         );
  OAI22_X1 U3852 ( .A1(n30381), .A2(n35508), .B1(n32756), .B2(n35507), .ZN(
        n30452) );
  XNOR2_X1 U3853 ( .A(\fmem_data[26][4] ), .B(\fmem_data[26][3] ), .ZN(n35034)
         );
  NAND2_X1 U3854 ( .A1(n9026), .A2(n35034), .ZN(n35033) );
  XOR2_X1 U3855 ( .A(\fmem_data[26][4] ), .B(\fmem_data[26][5] ), .Z(n9026) );
  NAND3_X1 U3856 ( .A1(n4671), .A2(n4670), .A3(n4669), .ZN(n31992) );
  AOI21_X1 U3857 ( .B1(n4647), .B2(n25287), .A(n4646), .ZN(n4670) );
  XNOR2_X1 U3858 ( .A(\fmem_data[17][1] ), .B(\fmem_data[17][2] ), .ZN(n33250)
         );
  NAND2_X1 U3859 ( .A1(n17556), .A2(n33250), .ZN(n33249) );
  XOR2_X1 U3860 ( .A(\fmem_data[17][3] ), .B(\fmem_data[17][2] ), .Z(n17556)
         );
  XNOR2_X1 U3861 ( .A(\fmem_data[10][4] ), .B(\fmem_data[10][3] ), .ZN(n35089)
         );
  XNOR2_X1 U3862 ( .A(\fmem_data[25][2] ), .B(\fmem_data[25][1] ), .ZN(n33059)
         );
  XNOR2_X1 U3863 ( .A(\fmem_data[31][4] ), .B(\fmem_data[31][3] ), .ZN(n34944)
         );
  XNOR2_X1 U3864 ( .A(\fmem_data[9][2] ), .B(\fmem_data[9][1] ), .ZN(n33873)
         );
  XNOR2_X1 U3865 ( .A(\fmem_data[8][4] ), .B(\fmem_data[8][3] ), .ZN(n35003)
         );
  XNOR2_X1 U3866 ( .A(\fmem_data[27][4] ), .B(\fmem_data[27][3] ), .ZN(n34903)
         );
  XNOR2_X1 U3867 ( .A(\fmem_data[19][4] ), .B(\fmem_data[19][3] ), .ZN(n34923)
         );
  XNOR2_X1 U3868 ( .A(\fmem_data[18][4] ), .B(\fmem_data[18][3] ), .ZN(n35006)
         );
  XNOR2_X1 U3869 ( .A(\fmem_data[22][1] ), .B(\fmem_data[22][2] ), .ZN(n34414)
         );
  XNOR2_X1 U3870 ( .A(\fmem_data[29][2] ), .B(\fmem_data[29][1] ), .ZN(n34422)
         );
  XNOR2_X1 U3871 ( .A(\fmem_data[30][3] ), .B(\fmem_data[30][4] ), .ZN(n33105)
         );
  XNOR2_X1 U3872 ( .A(\fmem_data[29][4] ), .B(\fmem_data[29][3] ), .ZN(n35083)
         );
  XNOR2_X1 U3873 ( .A(\fmem_data[15][4] ), .B(\fmem_data[15][3] ), .ZN(n34990)
         );
  NAND2_X1 U3874 ( .A1(n8643), .A2(n34942), .ZN(n34941) );
  OAI22_X1 U3875 ( .A1(n34034), .A2(n35711), .B1(n34033), .B2(n35712), .ZN(
        n34245) );
  XNOR2_X1 U3876 ( .A(\fmem_data[0][6] ), .B(\fmem_data[0][5] ), .ZN(n35494)
         );
  XNOR2_X1 U3877 ( .A(\fmem_data[16][2] ), .B(\fmem_data[16][1] ), .ZN(n34501)
         );
  XNOR2_X1 U3878 ( .A(\fmem_data[15][2] ), .B(\fmem_data[15][1] ), .ZN(n34364)
         );
  XNOR2_X1 U3879 ( .A(\fmem_data[31][2] ), .B(\fmem_data[31][1] ), .ZN(n34470)
         );
  XNOR2_X1 U3880 ( .A(\fmem_data[23][2] ), .B(\fmem_data[23][1] ), .ZN(n34412)
         );
  OAI22_X1 U3881 ( .A1(n30423), .A2(n34535), .B1(n30414), .B2(n34537), .ZN(
        n30466) );
  AND2_X1 U3882 ( .A1(n32223), .A2(n32222), .ZN(n30994) );
  OAI22_X1 U3883 ( .A1(n30398), .A2(n35508), .B1(n35507), .B2(n3600), .ZN(
        n30995) );
  OAI22_X1 U3884 ( .A1(n30397), .A2(n35712), .B1(n35711), .B2(n3655), .ZN(
        n30996) );
  NAND2_X1 U3885 ( .A1(n8553), .A2(n8552), .ZN(n31250) );
  NAND3_X1 U3886 ( .A1(n10675), .A2(n10674), .A3(n10673), .ZN(n31642) );
  NAND2_X1 U3887 ( .A1(n21189), .A2(n21188), .ZN(n28539) );
  NAND2_X1 U3888 ( .A1(n12715), .A2(n33859), .ZN(n33857) );
  OAI22_X1 U3889 ( .A1(n32022), .A2(n35712), .B1(n34033), .B2(n35711), .ZN(
        n33047) );
  OAI22_X1 U3890 ( .A1(n32017), .A2(n33328), .B1(n32016), .B2(n33326), .ZN(
        n33021) );
  OAI22_X1 U3891 ( .A1(n30460), .A2(n35089), .B1(n31999), .B2(n35088), .ZN(
        n30474) );
  NAND2_X1 U3892 ( .A1(n30168), .A2(n30167), .ZN(n30833) );
  NAND2_X1 U3893 ( .A1(n30479), .A2(n30478), .ZN(n30168) );
  OAI22_X1 U3894 ( .A1(n30159), .A2(n33850), .B1(n33180), .B2(n33851), .ZN(
        n30344) );
  OAI22_X1 U3895 ( .A1(n30460), .A2(n35088), .B1(n31666), .B2(n35089), .ZN(
        n11335) );
  AND2_X1 U3896 ( .A1(n33320), .A2(n33319), .ZN(n34838) );
  OAI22_X1 U3897 ( .A1(n33215), .A2(n34041), .B1(n33370), .B2(n34039), .ZN(
        n33302) );
  OAI22_X1 U3898 ( .A1(n33388), .A2(n35611), .B1(n33387), .B2(n35610), .ZN(
        n34911) );
  OAI22_X1 U3899 ( .A1(n33384), .A2(n35730), .B1(n33383), .B2(n35729), .ZN(
        n34913) );
  OAI22_X1 U3900 ( .A1(n33386), .A2(n33642), .B1(n33385), .B2(n33643), .ZN(
        n34912) );
  NAND2_X1 U3901 ( .A1(n8401), .A2(n28258), .ZN(n8402) );
  NAND2_X1 U3902 ( .A1(n23691), .A2(n23690), .ZN(n35030) );
  AOI22_X1 U3903 ( .A1(n23647), .A2(n30188), .B1(n23646), .B2(n30287), .ZN(
        n23691) );
  OAI22_X1 U3904 ( .A1(n35039), .A2(n35041), .B1(n34861), .B2(n35040), .ZN(
        n35143) );
  NAND2_X1 U3905 ( .A1(n23917), .A2(n23916), .ZN(n35316) );
  AOI22_X1 U3906 ( .A1(n23915), .A2(n30188), .B1(n23914), .B2(n30287), .ZN(
        n23916) );
  NAND2_X1 U3907 ( .A1(n27580), .A2(n27579), .ZN(n35178) );
  OAI22_X1 U3908 ( .A1(n31816), .A2(n35489), .B1(n35396), .B2(n35490), .ZN(
        n35166) );
  OR2_X1 U3909 ( .A1(n35008), .A2(n3948), .ZN(n35274) );
  OAI22_X1 U3910 ( .A1(n33316), .A2(n35515), .B1(n35123), .B2(n35516), .ZN(
        n35287) );
  OAI22_X1 U3911 ( .A1(n31661), .A2(n35507), .B1(n35404), .B2(n35508), .ZN(
        n35288) );
  OAI22_X1 U3912 ( .A1(n33325), .A2(n35721), .B1(n35337), .B2(n35722), .ZN(
        n35289) );
  OAI22_X1 U3913 ( .A1(n33314), .A2(n35580), .B1(n35075), .B2(n35581), .ZN(
        n35319) );
  OAI22_X1 U3914 ( .A1(n33384), .A2(n35729), .B1(n35329), .B2(n35730), .ZN(
        n35320) );
  INV_X1 U3915 ( .A(n31706), .ZN(n35318) );
  NAND2_X1 U3916 ( .A1(n29085), .A2(n29084), .ZN(n32616) );
  NAND2_X1 U3917 ( .A1(n16943), .A2(n16942), .ZN(n33592) );
  NAND4_X1 U3918 ( .A1(n8832), .A2(n8831), .A3(n8830), .A4(n8829), .ZN(n33484)
         );
  AND2_X1 U3919 ( .A1(n36339), .A2(n33813), .ZN(n33840) );
  NAND2_X1 U3920 ( .A1(n18820), .A2(n18819), .ZN(n31452) );
  INV_X1 U3921 ( .A(n24664), .ZN(n24724) );
  AND2_X1 U3922 ( .A1(n36111), .A2(n32077), .ZN(n32415) );
  XNOR2_X1 U3923 ( .A(n33750), .B(\fmem_data[17][5] ), .ZN(n32531) );
  OAI22_X1 U3924 ( .A1(n33224), .A2(n33963), .B1(n31993), .B2(n33961), .ZN(
        n19512) );
  XNOR2_X1 U3925 ( .A(\fmem_data[10][2] ), .B(\fmem_data[10][1] ), .ZN(n34736)
         );
  NAND2_X1 U3926 ( .A1(n12128), .A2(n34944), .ZN(n34945) );
  NAND3_X1 U3927 ( .A1(n25745), .A2(n25744), .A3(n25743), .ZN(n32117) );
  XNOR2_X1 U3928 ( .A(\fmem_data[23][4] ), .B(\fmem_data[23][3] ), .ZN(n34909)
         );
  NAND2_X1 U3929 ( .A1(n11049), .A2(n35003), .ZN(n35004) );
  OAI22_X1 U3930 ( .A1(n36228), .A2(n27325), .B1(n35740), .B2(n3484), .ZN(
        n30797) );
  XNOR2_X1 U3931 ( .A(\fmem_data[7][4] ), .B(\fmem_data[7][3] ), .ZN(n34835)
         );
  NAND2_X1 U3932 ( .A1(n25048), .A2(n34903), .ZN(n34904) );
  OAI22_X1 U3933 ( .A1(n30388), .A2(n35512), .B1(n35511), .B2(n3630), .ZN(
        n30991) );
  AND2_X1 U3934 ( .A1(n36312), .A2(n33572), .ZN(n33588) );
  OAI22_X1 U3935 ( .A1(n33574), .A2(n33853), .B1(n33854), .B2(n33855), .ZN(
        n33587) );
  NAND2_X1 U3936 ( .A1(n25333), .A2(n34414), .ZN(n34416) );
  NAND2_X1 U3937 ( .A1(n16753), .A2(n34422), .ZN(n34424) );
  OAI22_X1 U3938 ( .A1(n17555), .A2(n35753), .B1(n35752), .B2(n3621), .ZN(
        n26384) );
  OAI22_X1 U3939 ( .A1(n31994), .A2(n35730), .B1(n17744), .B2(n35729), .ZN(
        n26382) );
  OAI22_X1 U3940 ( .A1(n32067), .A2(n34199), .B1(n34200), .B2(n34201), .ZN(
        n31508) );
  XNOR2_X1 U3941 ( .A(\fmem_data[28][3] ), .B(\fmem_data[28][4] ), .ZN(n33828)
         );
  XNOR2_X1 U3942 ( .A(\fmem_data[20][3] ), .B(\fmem_data[20][4] ), .ZN(n35036)
         );
  NAND2_X1 U3943 ( .A1(n9492), .A2(n33105), .ZN(n33103) );
  XNOR2_X1 U3944 ( .A(\fmem_data[4][1] ), .B(\fmem_data[4][2] ), .ZN(n33174)
         );
  NAND2_X1 U3945 ( .A1(n23605), .A2(n34990), .ZN(n34989) );
  OAI22_X1 U3946 ( .A1(n33188), .A2(n33956), .B1(n33187), .B2(n33954), .ZN(
        n33231) );
  XNOR2_X1 U3947 ( .A(\fmem_data[11][4] ), .B(\fmem_data[11][3] ), .ZN(n34932)
         );
  OAI22_X1 U3948 ( .A1(n32255), .A2(n35638), .B1(n35637), .B2(n3656), .ZN(
        n32362) );
  OR2_X1 U3949 ( .A1(n36315), .A2(n3656), .ZN(n32255) );
  OAI22_X1 U3950 ( .A1(n35022), .A2(n35725), .B1(n35339), .B2(n35726), .ZN(
        n35261) );
  XNOR2_X1 U3951 ( .A(\fmem_data[15][6] ), .B(\fmem_data[15][5] ), .ZN(n35697)
         );
  XNOR2_X1 U3952 ( .A(\fmem_data[23][6] ), .B(\fmem_data[23][5] ), .ZN(n35652)
         );
  XNOR2_X1 U3953 ( .A(\fmem_data[10][6] ), .B(\fmem_data[10][5] ), .ZN(n35611)
         );
  NAND2_X1 U3954 ( .A1(n12811), .A2(n35494), .ZN(n35493) );
  XNOR2_X1 U3955 ( .A(\fmem_data[24][6] ), .B(\fmem_data[24][5] ), .ZN(n35490)
         );
  XNOR2_X1 U3956 ( .A(\fmem_data[5][6] ), .B(\fmem_data[5][5] ), .ZN(n35498)
         );
  XNOR2_X1 U3957 ( .A(\fmem_data[16][6] ), .B(\fmem_data[16][5] ), .ZN(n35753)
         );
  XNOR2_X1 U3958 ( .A(\fmem_data[28][6] ), .B(\fmem_data[28][5] ), .ZN(n35761)
         );
  XNOR2_X1 U3959 ( .A(\fmem_data[4][6] ), .B(\fmem_data[4][5] ), .ZN(n35749)
         );
  NAND4_X1 U3960 ( .A1(n22886), .A2(n22885), .A3(n22884), .A4(n22883), .ZN(
        n32979) );
  NAND3_X1 U3961 ( .A1(n17649), .A2(n17648), .A3(n17647), .ZN(n32898) );
  OAI22_X1 U3962 ( .A1(n32608), .A2(n34497), .B1(n34495), .B2(n3593), .ZN(
        n34539) );
  OAI22_X1 U3963 ( .A1(n32605), .A2(n33797), .B1(n33796), .B2(n3652), .ZN(
        n34541) );
  XNOR2_X1 U3964 ( .A(\fmem_data[0][1] ), .B(\fmem_data[0][2] ), .ZN(n34537)
         );
  XNOR2_X1 U3965 ( .A(\fmem_data[19][2] ), .B(\fmem_data[19][1] ), .ZN(n34472)
         );
  NAND2_X1 U3966 ( .A1(n14472), .A2(n34501), .ZN(n34499) );
  XNOR2_X1 U3967 ( .A(\fmem_data[20][1] ), .B(\fmem_data[20][2] ), .ZN(n34497)
         );
  NAND2_X1 U3968 ( .A1(n24113), .A2(n34364), .ZN(n34363) );
  XNOR2_X1 U3969 ( .A(\fmem_data[1][2] ), .B(\fmem_data[1][1] ), .ZN(n34779)
         );
  NAND2_X1 U3970 ( .A1(n8405), .A2(n34470), .ZN(n34468) );
  XNOR2_X1 U3971 ( .A(\fmem_data[8][2] ), .B(\fmem_data[8][1] ), .ZN(n34206)
         );
  OAI22_X1 U3972 ( .A1(n34438), .A2(n34435), .B1(n33678), .B2(n34437), .ZN(
        n33763) );
  OAI22_X1 U3973 ( .A1(n34434), .A2(n34431), .B1(n33684), .B2(n34433), .ZN(
        n33761) );
  XNOR2_X1 U3974 ( .A(\fmem_data[6][2] ), .B(\fmem_data[6][1] ), .ZN(n33596)
         );
  OAI22_X1 U3975 ( .A1(n32237), .A2(n35083), .B1(n35084), .B2(n3588), .ZN(
        n32446) );
  OAI22_X1 U3976 ( .A1(n32236), .A2(n34340), .B1(n33581), .B2(n33582), .ZN(
        n32447) );
  OAI22_X1 U3977 ( .A1(n34790), .A2(n3560), .B1(n34789), .B2(n34788), .ZN(
        n36234) );
  XNOR2_X1 U3978 ( .A(\fmem_data[3][2] ), .B(\fmem_data[3][1] ), .ZN(n34420)
         );
  OAI22_X1 U3979 ( .A1(n32238), .A2(n34739), .B1(n33969), .B2(n3563), .ZN(
        n31215) );
  OAI22_X1 U3980 ( .A1(n32236), .A2(n33582), .B1(n27583), .B2(n34340), .ZN(
        n31217) );
  XNOR2_X1 U3981 ( .A(\fmem_data[12][2] ), .B(\fmem_data[12][1] ), .ZN(n34340)
         );
  XNOR2_X1 U3982 ( .A(\fmem_data[12][6] ), .B(\fmem_data[12][5] ), .ZN(n35516)
         );
  XNOR2_X1 U3983 ( .A(\fmem_data[17][6] ), .B(\fmem_data[17][5] ), .ZN(n35581)
         );
  OAI22_X1 U3984 ( .A1(n32725), .A2(n34942), .B1(n31243), .B2(n34941), .ZN(
        n33637) );
  OAI22_X1 U3985 ( .A1(n31165), .A2(n35007), .B1(n27326), .B2(n35006), .ZN(
        n33635) );
  AND2_X1 U3986 ( .A1(n36339), .A2(n32891), .ZN(n36256) );
  AND2_X1 U3987 ( .A1(n36101), .A2(n31529), .ZN(n32960) );
  AND2_X1 U3988 ( .A1(n36105), .A2(n31581), .ZN(n32958) );
  AND2_X1 U3989 ( .A1(n34624), .A2(n31580), .ZN(n32959) );
  XNOR2_X1 U3990 ( .A(n32545), .B(n32566), .ZN(n34726) );
  XNOR2_X1 U3991 ( .A(n36967), .B(n36966), .ZN(n37025) );
  XNOR2_X1 U3992 ( .A(n36674), .B(n36673), .ZN(n36890) );
  XNOR2_X1 U3993 ( .A(n36672), .B(n36671), .ZN(n36674) );
  AND4_X1 U3994 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10147) );
  NOR2_X1 U3995 ( .A1(n25484), .A2(n25483), .ZN(n25500) );
  NAND2_X1 U3996 ( .A1(n7160), .A2(n30782), .ZN(n7161) );
  OAI21_X1 U3997 ( .B1(n20744), .B2(n20743), .A(n20742), .ZN(n20839) );
  OAI21_X1 U3998 ( .B1(n20835), .B2(n20834), .A(n20833), .ZN(n20836) );
  OAI21_X1 U3999 ( .B1(n20767), .B2(n20766), .A(n20765), .ZN(n20838) );
  AOI21_X1 U4000 ( .B1(n34736), .B2(n33690), .A(n33031), .ZN(n33032) );
  NAND2_X1 U4001 ( .A1(n30341), .A2(n30340), .ZN(n31758) );
  NAND2_X1 U4002 ( .A1(n30339), .A2(n30338), .ZN(n30340) );
  XNOR2_X1 U4003 ( .A(n31674), .B(\fmem_data[10][5] ), .ZN(n31666) );
  XNOR2_X1 U4004 ( .A(n32615), .B(\fmem_data[24][7] ), .ZN(n31639) );
  XNOR2_X1 U4005 ( .A(n35074), .B(\fmem_data[17][5] ), .ZN(n33127) );
  XNOR2_X1 U4006 ( .A(n35122), .B(\fmem_data[12][5] ), .ZN(n33373) );
  XNOR2_X1 U4007 ( .A(n35328), .B(\fmem_data[8][5] ), .ZN(n35005) );
  AOI21_X1 U4008 ( .B1(n33328), .B2(n33326), .A(n33329), .ZN(n31675) );
  XNOR2_X1 U4009 ( .A(n31673), .B(\fmem_data[10][7] ), .ZN(n33388) );
  AOI21_X1 U4010 ( .B1(n34039), .B2(n34041), .A(n33371), .ZN(n31803) );
  AOI21_X1 U4011 ( .B1(n33975), .B2(n33973), .A(n33373), .ZN(n31804) );
  NAND2_X1 U4012 ( .A1(n4573), .A2(n28107), .ZN(n4574) );
  OAI21_X1 U4013 ( .B1(n4503), .B2(n4502), .A(n25287), .ZN(n4576) );
  XNOR2_X1 U4014 ( .A(n36200), .B(\fmem_data[30][7] ), .ZN(n32667) );
  XNOR2_X1 U4015 ( .A(n35357), .B(\fmem_data[29][3] ), .ZN(n33017) );
  NAND2_X1 U4016 ( .A1(n9795), .A2(n27937), .ZN(n9874) );
  NAND2_X1 U4017 ( .A1(n9816), .A2(n27968), .ZN(n9873) );
  OAI21_X1 U4018 ( .B1(n9870), .B2(n9869), .A(n9896), .ZN(n9871) );
  NAND3_X1 U4019 ( .A1(n5364), .A2(n5363), .A3(n5362), .ZN(n32225) );
  NAND3_X1 U4020 ( .A1(n21491), .A2(n21490), .A3(n21489), .ZN(n33227) );
  NAND2_X1 U4021 ( .A1(n23163), .A2(n23162), .ZN(n33246) );
  NAND3_X1 U4022 ( .A1(n11237), .A2(n3716), .A3(n11236), .ZN(n31899) );
  NAND2_X1 U4023 ( .A1(n10467), .A2(n10466), .ZN(n31640) );
  NAND2_X1 U4024 ( .A1(n10465), .A2(n20980), .ZN(n10466) );
  AND2_X1 U4025 ( .A1(n10429), .A2(n20311), .ZN(n10430) );
  AND2_X1 U4026 ( .A1(n36111), .A2(n34052), .ZN(n34211) );
  NAND3_X1 U4027 ( .A1(n16849), .A2(n16848), .A3(n16847), .ZN(n32600) );
  XNOR2_X1 U4028 ( .A(n35102), .B(\fmem_data[14][1] ), .ZN(n33970) );
  OR2_X1 U4029 ( .A1(n36200), .A2(n3585), .ZN(n21674) );
  OR2_X1 U4030 ( .A1(n36244), .A2(n3598), .ZN(n21583) );
  XNOR2_X1 U4031 ( .A(n32612), .B(\fmem_data[30][7] ), .ZN(n31985) );
  NAND2_X1 U4032 ( .A1(n30402), .A2(n30401), .ZN(n32348) );
  OAI22_X1 U4033 ( .A1(n30471), .A2(n34431), .B1(n30983), .B2(n34433), .ZN(
        n31654) );
  OAI22_X1 U4034 ( .A1(n30473), .A2(n34045), .B1(n32322), .B2(n34043), .ZN(
        n31652) );
  NAND2_X1 U4035 ( .A1(n30390), .A2(n30389), .ZN(n30811) );
  NAND2_X1 U4036 ( .A1(n30824), .A2(n30823), .ZN(n30432) );
  NAND2_X1 U4037 ( .A1(n32044), .A2(n32043), .ZN(n32045) );
  OAI21_X1 U4038 ( .B1(n32044), .B2(n32043), .A(n32042), .ZN(n32046) );
  XNOR2_X1 U4039 ( .A(n33362), .B(n33054), .ZN(n33390) );
  XNOR2_X1 U4040 ( .A(n33364), .B(n33363), .ZN(n33054) );
  OAI22_X1 U4041 ( .A1(n33257), .A2(n35729), .B1(n33383), .B2(n35730), .ZN(
        n33123) );
  OAI22_X1 U4042 ( .A1(n35180), .A2(n35182), .B1(n33102), .B2(n35181), .ZN(
        n34993) );
  INV_X1 U4043 ( .A(n35012), .ZN(n35272) );
  AOI21_X1 U4044 ( .B1(n35011), .B2(n35010), .A(n35009), .ZN(n35012) );
  OAI22_X1 U4045 ( .A1(n35179), .A2(n35739), .B1(n31643), .B2(n35740), .ZN(
        n31712) );
  OAI22_X1 U4046 ( .A1(n31813), .A2(n35701), .B1(n33217), .B2(n35700), .ZN(
        n31797) );
  NAND3_X1 U4047 ( .A1(n17944), .A2(n17943), .A3(n17942), .ZN(n31660) );
  NAND4_X1 U4048 ( .A1(n13309), .A2(n13308), .A3(n13307), .A4(n13306), .ZN(
        n35023) );
  OR4_X1 U4049 ( .A1(n15733), .A2(n15735), .A3(n15734), .A4(n15736), .ZN(
        n15737) );
  NAND2_X1 U4050 ( .A1(n10067), .A2(n10066), .ZN(n35403) );
  NAND2_X1 U4051 ( .A1(n4394), .A2(n22768), .ZN(n4469) );
  OAI21_X1 U4052 ( .B1(n4439), .B2(n4438), .A(n22735), .ZN(n4467) );
  OAI21_X1 U4053 ( .B1(n4465), .B2(n4464), .A(n22698), .ZN(n4466) );
  INV_X1 U4054 ( .A(n31814), .ZN(n35162) );
  OAI22_X1 U4055 ( .A1(n31813), .A2(n35700), .B1(n35281), .B2(n35701), .ZN(
        n35163) );
  OAI22_X1 U4056 ( .A1(n35177), .A2(n35584), .B1(n35176), .B2(n35585), .ZN(
        n35394) );
  OAI22_X1 U4057 ( .A1(n35115), .A2(n35651), .B1(n35259), .B2(n35652), .ZN(
        n35137) );
  OAI22_X1 U4058 ( .A1(n35113), .A2(n35633), .B1(n35239), .B2(n35634), .ZN(
        n35138) );
  NAND4_X1 U4059 ( .A1(n20391), .A2(n20390), .A3(n20389), .A4(n20388), .ZN(
        n32065) );
  OAI21_X1 U4060 ( .B1(n20313), .B2(n20312), .A(n20311), .ZN(n20391) );
  NAND3_X1 U4061 ( .A1(n19303), .A2(n19302), .A3(n19301), .ZN(n32528) );
  AOI22_X1 U4062 ( .A1(n15540), .A2(n29837), .B1(n15539), .B2(n29758), .ZN(
        n15585) );
  NAND2_X1 U4063 ( .A1(n21953), .A2(n32780), .ZN(n32779) );
  XOR2_X1 U4064 ( .A(\fmem_data[26][2] ), .B(\fmem_data[26][3] ), .Z(n21953)
         );
  XNOR2_X1 U4065 ( .A(n32899), .B(\fmem_data[8][3] ), .ZN(n33831) );
  XNOR2_X1 U4066 ( .A(n31642), .B(\fmem_data[20][1] ), .ZN(n33878) );
  XNOR2_X1 U4067 ( .A(n34531), .B(\fmem_data[10][5] ), .ZN(n31123) );
  AND2_X1 U4068 ( .A1(n36200), .A2(n32252), .ZN(n32658) );
  AND2_X1 U4069 ( .A1(n36299), .A2(n32253), .ZN(n32657) );
  XNOR2_X1 U4070 ( .A(n32127), .B(\fmem_data[20][3] ), .ZN(n32418) );
  XNOR2_X1 U4071 ( .A(n32898), .B(\fmem_data[8][5] ), .ZN(n32130) );
  OR2_X1 U4072 ( .A1(n36299), .A2(n3596), .ZN(n32244) );
  OR2_X1 U4073 ( .A1(n36200), .A2(n3597), .ZN(n32245) );
  XNOR2_X1 U4074 ( .A(n31992), .B(\fmem_data[22][3] ), .ZN(n32125) );
  AND2_X1 U4075 ( .A1(n36105), .A2(n32120), .ZN(n32686) );
  INV_X1 U4076 ( .A(n35006), .ZN(n32120) );
  XNOR2_X1 U4077 ( .A(\fmem_data[12][3] ), .B(\fmem_data[12][4] ), .ZN(n33975)
         );
  XNOR2_X1 U4078 ( .A(n31656), .B(\fmem_data[28][1] ), .ZN(n32525) );
  NAND2_X1 U4079 ( .A1(n10167), .A2(n35089), .ZN(n35088) );
  XNOR2_X1 U4080 ( .A(n31663), .B(\fmem_data[12][1] ), .ZN(n30816) );
  NAND2_X1 U4081 ( .A1(n13111), .A2(n33059), .ZN(n33057) );
  XNOR2_X1 U4082 ( .A(n35270), .B(\fmem_data[19][1] ), .ZN(n32152) );
  NAND4_X1 U4083 ( .A1(n25936), .A2(n25935), .A3(n25934), .A4(n25933), .ZN(
        n31940) );
  XNOR2_X1 U4084 ( .A(n31799), .B(\fmem_data[14][1] ), .ZN(n33969) );
  OR2_X1 U4085 ( .A1(n36105), .A2(n3639), .ZN(n28401) );
  AND2_X1 U4086 ( .A1(n36338), .A2(n30013), .ZN(n31390) );
  AND2_X1 U4087 ( .A1(n36339), .A2(n30123), .ZN(n31391) );
  XNOR2_X1 U4088 ( .A(\fmem_data[3][4] ), .B(\fmem_data[3][3] ), .ZN(n34919)
         );
  OAI211_X1 U4089 ( .C1(n6166), .C2(n24151), .A(n6165), .B(n6164), .ZN(n31669)
         );
  NAND2_X1 U4090 ( .A1(n24334), .A2(n24333), .ZN(n32235) );
  AOI22_X1 U4091 ( .A1(n24332), .A2(n31342), .B1(n24331), .B2(n31376), .ZN(
        n24333) );
  NAND2_X1 U4092 ( .A1(n25598), .A2(n34909), .ZN(n34908) );
  NAND2_X1 U4093 ( .A1(n12343), .A2(n33873), .ZN(n33875) );
  OAI22_X1 U4094 ( .A1(n30493), .A2(n35726), .B1(n35725), .B2(n3625), .ZN(
        n30987) );
  NAND2_X1 U4095 ( .A1(n27323), .A2(n34835), .ZN(n34836) );
  OAI22_X1 U4096 ( .A1(n33951), .A2(n35615), .B1(n35614), .B2(n3602), .ZN(
        n34080) );
  OAI22_X1 U4097 ( .A1(n33948), .A2(n3567), .B1(n33947), .B2(n34777), .ZN(
        n34082) );
  OAI22_X1 U4098 ( .A1(n33649), .A2(n34598), .B1(n33648), .B2(n3569), .ZN(
        n34350) );
  AND2_X1 U4099 ( .A1(n36338), .A2(n33647), .ZN(n34352) );
  OAI22_X1 U4100 ( .A1(n33601), .A2(n36114), .B1(n33600), .B2(n3561), .ZN(
        n33651) );
  OAI22_X1 U4101 ( .A1(n33604), .A2(n33603), .B1(n33602), .B2(n33741), .ZN(
        n33650) );
  OAI22_X1 U4102 ( .A1(n33599), .A2(n33598), .B1(n33597), .B2(n33596), .ZN(
        n33652) );
  NAND2_X1 U4103 ( .A1(n18429), .A2(n34923), .ZN(n34922) );
  NAND2_X1 U4104 ( .A1(n6896), .A2(n35006), .ZN(n35007) );
  XNOR2_X1 U4105 ( .A(n32528), .B(\fmem_data[29][3] ), .ZN(n34423) );
  XNOR2_X1 U4106 ( .A(n33789), .B(\fmem_data[30][3] ), .ZN(n34436) );
  XNOR2_X1 U4107 ( .A(\fmem_data[16][3] ), .B(\fmem_data[16][4] ), .ZN(n33328)
         );
  OAI22_X1 U4108 ( .A1(n33200), .A2(n35592), .B1(n17464), .B2(n35591), .ZN(
        n23583) );
  OAI22_X1 U4109 ( .A1(n33186), .A2(n35083), .B1(n26370), .B2(n35084), .ZN(
        n23575) );
  NAND2_X1 U4110 ( .A1(n9686), .A2(n33828), .ZN(n33827) );
  NAND2_X1 U4111 ( .A1(n10767), .A2(n35036), .ZN(n35037) );
  XNOR2_X1 U4112 ( .A(n31640), .B(\fmem_data[0][1] ), .ZN(n31126) );
  OAI22_X1 U4113 ( .A1(n33843), .A2(n35019), .B1(n35018), .B2(n3620), .ZN(
        n33898) );
  XNOR2_X1 U4114 ( .A(n31492), .B(\fmem_data[25][5] ), .ZN(n32514) );
  XNOR2_X1 U4115 ( .A(\fmem_data[25][4] ), .B(\fmem_data[25][3] ), .ZN(n34986)
         );
  NAND2_X1 U4116 ( .A1(n25049), .A2(n34986), .ZN(n34985) );
  XOR2_X1 U4117 ( .A(\fmem_data[25][4] ), .B(\fmem_data[25][5] ), .Z(n25049)
         );
  OAI22_X1 U4118 ( .A1(n33860), .A2(n33859), .B1(n33858), .B2(n33857), .ZN(
        n34213) );
  OAI22_X1 U4119 ( .A1(n33856), .A2(n33855), .B1(n33854), .B2(n33853), .ZN(
        n34214) );
  XNOR2_X1 U4120 ( .A(\fmem_data[17][3] ), .B(\fmem_data[17][4] ), .ZN(n34045)
         );
  NAND2_X1 U4121 ( .A1(n14670), .A2(n34045), .ZN(n34043) );
  XOR2_X1 U4122 ( .A(\fmem_data[17][5] ), .B(\fmem_data[17][4] ), .Z(n14670)
         );
  XNOR2_X1 U4123 ( .A(\fmem_data[21][2] ), .B(\fmem_data[21][1] ), .ZN(n34201)
         );
  XNOR2_X1 U4124 ( .A(\fmem_data[14][3] ), .B(\fmem_data[14][4] ), .ZN(n33100)
         );
  NAND2_X1 U4125 ( .A1(n33166), .A2(n33165), .ZN(n33245) );
  OAI22_X1 U4126 ( .A1(n33168), .A2(n34903), .B1(n33167), .B2(n34904), .ZN(
        n33244) );
  OAI22_X1 U4127 ( .A1(n33170), .A2(n34364), .B1(n33169), .B2(n34363), .ZN(
        n33243) );
  OAI22_X1 U4128 ( .A1(n33257), .A2(n35730), .B1(n33256), .B2(n35729), .ZN(
        n33339) );
  OAI22_X1 U4129 ( .A1(n34242), .A2(n35726), .B1(n34241), .B2(n35725), .ZN(
        n34666) );
  OAI22_X1 U4130 ( .A1(n34240), .A2(n35652), .B1(n34239), .B2(n35651), .ZN(
        n34667) );
  OAI21_X1 U4131 ( .B1(n32769), .B2(n32768), .A(n32770), .ZN(n32674) );
  OAI22_X1 U4132 ( .A1(n32259), .A2(n35662), .B1(n35663), .B2(n32258), .ZN(
        n32366) );
  OAI22_X1 U4133 ( .A1(n32261), .A2(n34533), .B1(n32260), .B2(n34429), .ZN(
        n32365) );
  OAI22_X1 U4134 ( .A1(n24112), .A2(n35083), .B1(n33185), .B2(n35084), .ZN(
        n26041) );
  OAI22_X1 U4135 ( .A1(n24016), .A2(n35003), .B1(n24015), .B2(n35004), .ZN(
        n26043) );
  OAI22_X1 U4136 ( .A1(n31947), .A2(n35584), .B1(n35585), .B2(n24111), .ZN(
        n26042) );
  OAI21_X1 U4137 ( .B1(n33089), .B2(n33090), .A(n33088), .ZN(n33092) );
  NAND2_X1 U4138 ( .A1(n32471), .A2(n32469), .ZN(n31923) );
  INV_X1 U4139 ( .A(n34943), .ZN(n35368) );
  OAI22_X1 U4140 ( .A1(n35086), .A2(n35083), .B1(n33131), .B2(n35084), .ZN(
        n35046) );
  AOI21_X1 U4141 ( .B1(n13999), .B2(n30007), .A(n13998), .ZN(n14000) );
  NAND2_X1 U4142 ( .A1(n6393), .A2(n35697), .ZN(n35696) );
  OAI22_X1 U4143 ( .A1(n31819), .A2(n35704), .B1(n35109), .B2(n35705), .ZN(
        n35118) );
  XNOR2_X1 U4144 ( .A(\fmem_data[11][6] ), .B(\fmem_data[11][5] ), .ZN(n35634)
         );
  XNOR2_X1 U4145 ( .A(\fmem_data[3][6] ), .B(\fmem_data[3][5] ), .ZN(n35638)
         );
  XNOR2_X1 U4146 ( .A(\fmem_data[27][6] ), .B(\fmem_data[27][5] ), .ZN(n35642)
         );
  XNOR2_X1 U4147 ( .A(\fmem_data[29][6] ), .B(\fmem_data[29][5] ), .ZN(n35615)
         );
  NAND2_X1 U4148 ( .A1(n15217), .A2(n35611), .ZN(n35610) );
  NAND2_X1 U4149 ( .A1(n5266), .A2(n35508), .ZN(n35507) );
  XNOR2_X1 U4150 ( .A(n35403), .B(\fmem_data[21][7] ), .ZN(n35506) );
  NAND3_X1 U4151 ( .A1(n24240), .A2(n24239), .A3(n24238), .ZN(n35104) );
  XNOR2_X1 U4152 ( .A(\fmem_data[14][6] ), .B(\fmem_data[14][5] ), .ZN(n35577)
         );
  XNOR2_X1 U4153 ( .A(\fmem_data[22][6] ), .B(\fmem_data[22][5] ), .ZN(n35585)
         );
  XNOR2_X1 U4154 ( .A(n35401), .B(\fmem_data[0][7] ), .ZN(n35492) );
  NAND2_X1 U4155 ( .A1(n24725), .A2(n35490), .ZN(n35489) );
  XNOR2_X1 U4156 ( .A(n35395), .B(\fmem_data[24][7] ), .ZN(n35488) );
  NAND2_X1 U4157 ( .A1(n5667), .A2(n35498), .ZN(n35497) );
  XNOR2_X1 U4158 ( .A(n35405), .B(\fmem_data[5][7] ), .ZN(n35496) );
  NAND2_X1 U4159 ( .A1(n13615), .A2(n35753), .ZN(n35752) );
  NAND2_X1 U4160 ( .A1(n19609), .A2(n35761), .ZN(n35760) );
  XNOR2_X1 U4161 ( .A(\fmem_data[25][6] ), .B(\fmem_data[25][5] ), .ZN(n35745)
         );
  NAND2_X1 U4162 ( .A1(n4269), .A2(n35749), .ZN(n35748) );
  XNOR2_X1 U4163 ( .A(\fmem_data[20][6] ), .B(\fmem_data[20][5] ), .ZN(n35739)
         );
  NAND2_X1 U4164 ( .A1(n35071), .A2(n35070), .ZN(n35734) );
  NAND2_X1 U4165 ( .A1(n35069), .A2(n35068), .ZN(n35070) );
  OAI21_X1 U4166 ( .B1(n35069), .B2(n35068), .A(n35067), .ZN(n35071) );
  INV_X1 U4167 ( .A(n3385), .ZN(n3388) );
  NOR2_X1 U4168 ( .A1(n6890), .A2(n6889), .ZN(n28395) );
  NAND3_X1 U4169 ( .A1(n31110), .A2(n31109), .A3(n31108), .ZN(n34610) );
  NAND3_X1 U4170 ( .A1(n19209), .A2(n19208), .A3(n19207), .ZN(n33750) );
  NAND2_X1 U4171 ( .A1(n11239), .A2(n34537), .ZN(n34535) );
  XNOR2_X1 U4172 ( .A(n32057), .B(\fmem_data[21][1] ), .ZN(n34485) );
  NAND2_X1 U4173 ( .A1(n7705), .A2(n34472), .ZN(n34474) );
  NAND2_X1 U4174 ( .A1(n14188), .A2(n34497), .ZN(n34495) );
  XNOR2_X1 U4175 ( .A(\fmem_data[11][2] ), .B(\fmem_data[11][1] ), .ZN(n34533)
         );
  AND2_X1 U4176 ( .A1(n36244), .A2(n33742), .ZN(n34609) );
  OR2_X1 U4177 ( .A1(n36339), .A2(n3609), .ZN(n34365) );
  XNOR2_X1 U4178 ( .A(n36338), .B(\fmem_data[1][3] ), .ZN(n34467) );
  XNOR2_X1 U4179 ( .A(\fmem_data[27][2] ), .B(\fmem_data[27][1] ), .ZN(n34463)
         );
  NAND2_X1 U4180 ( .A1(n25148), .A2(n34779), .ZN(n34466) );
  AND2_X1 U4181 ( .A1(n36299), .A2(n34339), .ZN(n34621) );
  AND2_X1 U4182 ( .A1(n36112), .A2(n34341), .ZN(n34620) );
  OAI22_X1 U4183 ( .A1(n32551), .A2(n33855), .B1(n33853), .B2(n3604), .ZN(
        n32887) );
  NAND2_X1 U4184 ( .A1(n25838), .A2(n34206), .ZN(n34208) );
  OAI22_X1 U4185 ( .A1(n33691), .A2(n34736), .B1(n33690), .B2(n3611), .ZN(
        n33765) );
  OAI22_X1 U4186 ( .A1(n33689), .A2(n36221), .B1(n33688), .B2(n3558), .ZN(
        n33766) );
  XNOR2_X1 U4187 ( .A(n33806), .B(n33805), .ZN(n33808) );
  NAND2_X1 U4188 ( .A1(n31507), .A2(n31506), .ZN(n33564) );
  NAND2_X1 U4189 ( .A1(n33490), .A2(n33491), .ZN(n31506) );
  OAI21_X1 U4190 ( .B1(n33490), .B2(n33491), .A(n33489), .ZN(n31507) );
  XNOR2_X1 U4191 ( .A(n33576), .B(n33575), .ZN(n33566) );
  OAI22_X1 U4192 ( .A1(n31251), .A2(n34990), .B1(n34989), .B2(n3619), .ZN(
        n31555) );
  OAI22_X1 U4193 ( .A1(n31543), .A2(n33603), .B1(n33604), .B2(n33741), .ZN(
        n33548) );
  OAI22_X1 U4194 ( .A1(n31544), .A2(n33741), .B1(n33603), .B2(n3617), .ZN(
        n33547) );
  OR2_X1 U4195 ( .A1(n36244), .A2(n3617), .ZN(n31544) );
  OAI22_X1 U4196 ( .A1(n31218), .A2(n34942), .B1(n34941), .B2(n3583), .ZN(
        n31575) );
  OR2_X1 U4197 ( .A1(n36338), .A2(n3583), .ZN(n31218) );
  NAND2_X1 U4198 ( .A1(n33487), .A2(n33486), .ZN(n31593) );
  OAI22_X1 U4199 ( .A1(n31173), .A2(n35083), .B1(n31172), .B2(n35084), .ZN(
        n32492) );
  OAI22_X1 U4200 ( .A1(n31169), .A2(n33105), .B1(n31168), .B2(n33103), .ZN(
        n32490) );
  OAI22_X1 U4201 ( .A1(n31170), .A2(n34932), .B1(n34933), .B2(n3697), .ZN(
        n32489) );
  XNOR2_X1 U4202 ( .A(n32612), .B(\fmem_data[30][3] ), .ZN(n33790) );
  XNOR2_X1 U4203 ( .A(\fmem_data[24][2] ), .B(\fmem_data[24][1] ), .ZN(n34431)
         );
  NAND2_X1 U4204 ( .A1(n18142), .A2(n34435), .ZN(n34437) );
  OAI22_X1 U4205 ( .A1(n32203), .A2(n33098), .B1(n32202), .B2(n33100), .ZN(
        n32411) );
  XNOR2_X1 U4206 ( .A(n36244), .B(\fmem_data[14][5] ), .ZN(n32203) );
  OAI22_X1 U4207 ( .A1(n32204), .A2(n33100), .B1(n33098), .B2(n3584), .ZN(
        n32410) );
  OR2_X1 U4208 ( .A1(n36244), .A2(n3584), .ZN(n32204) );
  OAI22_X1 U4209 ( .A1(n34471), .A2(n34468), .B1(n32621), .B2(n34470), .ZN(
        n34773) );
  OAI22_X1 U4210 ( .A1(n32187), .A2(n35663), .B1(n35662), .B2(n3487), .ZN(
        n32635) );
  OAI22_X1 U4211 ( .A1(n32162), .A2(n35701), .B1(n35700), .B2(n3601), .ZN(
        n32198) );
  OR2_X1 U4212 ( .A1(n36338), .A2(n3601), .ZN(n32162) );
  OAI22_X1 U4213 ( .A1(n31014), .A2(n35494), .B1(n31013), .B2(n35493), .ZN(
        n31114) );
  OAI22_X1 U4214 ( .A1(n32132), .A2(n33176), .B1(n28265), .B2(n33174), .ZN(
        n31212) );
  XNOR2_X1 U4215 ( .A(\fmem_data[6][6] ), .B(\fmem_data[6][5] ), .ZN(n35512)
         );
  NAND2_X1 U4216 ( .A1(n6482), .A2(n34340), .ZN(n33582) );
  XNOR2_X1 U4217 ( .A(\fmem_data[7][2] ), .B(\fmem_data[7][1] ), .ZN(n34505)
         );
  XNOR2_X1 U4218 ( .A(\fmem_data[7][6] ), .B(\fmem_data[7][5] ), .ZN(n35619)
         );
  XNOR2_X1 U4219 ( .A(\fmem_data[13][1] ), .B(\fmem_data[13][2] ), .ZN(n33568)
         );
  NAND2_X1 U4220 ( .A1(n21190), .A2(n33568), .ZN(n33570) );
  XOR2_X1 U4221 ( .A(\fmem_data[13][3] ), .B(\fmem_data[13][2] ), .Z(n21190)
         );
  NAND2_X1 U4222 ( .A1(n5868), .A2(n35516), .ZN(n35515) );
  NAND2_X1 U4223 ( .A1(n4966), .A2(n35581), .ZN(n35580) );
  XNOR2_X1 U4224 ( .A(n31193), .B(n31192), .ZN(n31606) );
  OAI22_X1 U4225 ( .A1(n34417), .A2(n34416), .B1(n34415), .B2(n34414), .ZN(
        n34490) );
  OAI22_X1 U4226 ( .A1(n34413), .A2(n34412), .B1(n34411), .B2(n34410), .ZN(
        n34491) );
  OAI22_X1 U4227 ( .A1(n32751), .A2(n34364), .B1(n34363), .B2(n26805), .ZN(
        n33629) );
  OAI22_X1 U4228 ( .A1(n35661), .A2(n35663), .B1(n35257), .B2(n35662), .ZN(
        n35520) );
  OAI22_X1 U4229 ( .A1(n35650), .A2(n35652), .B1(n35259), .B2(n35651), .ZN(
        n35519) );
  XNOR2_X1 U4230 ( .A(\fmem_data[19][6] ), .B(\fmem_data[19][5] ), .ZN(n35656)
         );
  XNOR2_X1 U4231 ( .A(\fmem_data[2][6] ), .B(\fmem_data[2][5] ), .ZN(n35722)
         );
  XNOR2_X1 U4232 ( .A(\fmem_data[13][6] ), .B(\fmem_data[13][5] ), .ZN(n35592)
         );
  NAND2_X1 U4233 ( .A1(n21279), .A2(n21278), .ZN(n21280) );
  XNOR2_X1 U4234 ( .A(n34610), .B(\fmem_data[12][1] ), .ZN(n34735) );
  XNOR2_X1 U4235 ( .A(n33750), .B(\fmem_data[17][1] ), .ZN(n34530) );
  OR2_X1 U4236 ( .A1(n36200), .A2(n3672), .ZN(n34628) );
  NAND2_X1 U4237 ( .A1(\fmem_data[12][1] ), .A2(n3572), .ZN(n34734) );
  NAND4_X1 U4238 ( .A1(n22054), .A2(n22053), .A3(n22052), .A4(n22051), .ZN(
        n33553) );
  NAND2_X1 U4239 ( .A1(n36789), .A2(n36787), .ZN(n36212) );
  OAI22_X1 U4240 ( .A1(n34772), .A2(n3565), .B1(n34771), .B2(n36100), .ZN(
        n36140) );
  NAND2_X1 U4241 ( .A1(n36472), .A2(n36473), .ZN(n33558) );
  NAND2_X1 U4242 ( .A1(n36696), .A2(n36695), .ZN(n36250) );
  NAND2_X1 U4243 ( .A1(n36351), .A2(n36350), .ZN(n32964) );
  OAI22_X1 U4244 ( .A1(n33601), .A2(n3561), .B1(n34532), .B2(n36114), .ZN(
        n32987) );
  OAI22_X1 U4245 ( .A1(n33599), .A2(n33596), .B1(n31450), .B2(n33598), .ZN(
        n32988) );
  NAND2_X1 U4246 ( .A1(n36175), .A2(n36176), .ZN(n32902) );
  NAND2_X1 U4247 ( .A1(n32831), .A2(n32829), .ZN(n32628) );
  NAND2_X1 U4248 ( .A1(n35388), .A2(n35387), .ZN(n35540) );
  NAND2_X1 U4249 ( .A1(n35386), .A2(n35385), .ZN(n35387) );
  OAI21_X1 U4250 ( .B1(n35385), .B2(n35386), .A(n35384), .ZN(n35388) );
  XNOR2_X1 U4251 ( .A(\fmem_data[30][6] ), .B(\fmem_data[30][5] ), .ZN(n35709)
         );
  XNOR2_X1 U4252 ( .A(\fmem_data[18][6] ), .B(\fmem_data[18][5] ), .ZN(n35705)
         );
  AND2_X1 U4253 ( .A1(n34615), .A2(\fmem_data[21][0] ), .ZN(n36201) );
  INV_X1 U4254 ( .A(n28437), .ZN(n28531) );
  NAND3_X1 U4255 ( .A1(n28737), .A2(n28736), .A3(n28735), .ZN(n28764) );
  AND2_X1 U4256 ( .A1(n29435), .A2(n29434), .ZN(n29445) );
  NAND4_X2 U4257 ( .A1(n17462), .A2(n17461), .A3(n17460), .A4(n17459), .ZN(
        n33800) );
  OAI21_X1 U4258 ( .B1(n17412), .B2(n17411), .A(n24236), .ZN(n17461) );
  OAI21_X1 U4259 ( .B1(n17458), .B2(n17457), .A(n24205), .ZN(n17459) );
  NAND2_X1 U4260 ( .A1(n17390), .A2(n17389), .ZN(n17462) );
  NAND2_X1 U4261 ( .A1(\fmem_data[10][1] ), .A2(n3561), .ZN(n36114) );
  OR2_X1 U4262 ( .A1(n36338), .A2(n3661), .ZN(n36220) );
  OR2_X1 U4263 ( .A1(n36299), .A2(n3680), .ZN(n34622) );
  OAI22_X1 U4264 ( .A1(n34596), .A2(n3560), .B1(n36200), .B2(n34788), .ZN(
        n36571) );
  OAI22_X1 U4265 ( .A1(n34746), .A2(n3562), .B1(n34624), .B2(n34745), .ZN(
        n36531) );
  XNOR2_X1 U4266 ( .A(n36307), .B(n36306), .ZN(n36710) );
  NAND2_X1 U4267 ( .A1(n36924), .A2(n36923), .ZN(n36587) );
  NAND2_X1 U4268 ( .A1(n37086), .A2(n37084), .ZN(n37027) );
  XNOR2_X1 U4269 ( .A(n36737), .B(n36736), .ZN(n36939) );
  XNOR2_X1 U4270 ( .A(n36735), .B(n36734), .ZN(n36736) );
  XNOR2_X1 U4271 ( .A(n36678), .B(n36677), .ZN(n36938) );
  NAND2_X1 U4272 ( .A1(n36884), .A2(n36883), .ZN(n36822) );
  XNOR2_X1 U4273 ( .A(n36666), .B(n36665), .ZN(n36825) );
  NOR2_X1 U4274 ( .A1(n37152), .A2(n37151), .ZN(n37228) );
  NAND2_X1 U4275 ( .A1(n37145), .A2(n3436), .ZN(n37234) );
  NAND3_X1 U4276 ( .A1(n19926), .A2(n19925), .A3(n19924), .ZN(n19929) );
  INV_X1 U4277 ( .A(n3339), .ZN(n3340) );
  INV_X1 U4278 ( .A(n24795), .ZN(n24796) );
  INV_X1 U4279 ( .A(n24794), .ZN(n24797) );
  AND4_X1 U4280 ( .A1(n26194), .A2(n26193), .A3(n26192), .A4(n26191), .ZN(
        n26197) );
  INV_X1 U4281 ( .A(n3339), .ZN(n3322) );
  INV_X1 U4282 ( .A(n23518), .ZN(n23519) );
  INV_X1 U4283 ( .A(n14357), .ZN(n14358) );
  OR2_X1 U4284 ( .A1(n18595), .A2(n18594), .ZN(n18596) );
  AND2_X1 U4285 ( .A1(n16986), .A2(\xmem_data[22][5] ), .ZN(n18594) );
  NOR2_X1 U4286 ( .A1(n16308), .A2(n16307), .ZN(n16319) );
  AND2_X1 U4287 ( .A1(n16302), .A2(n16301), .ZN(n16320) );
  NAND3_X1 U4288 ( .A1(n24989), .A2(n24988), .A3(n24987), .ZN(n24990) );
  NAND3_X1 U4289 ( .A1(n24962), .A2(n24961), .A3(n24960), .ZN(n24963) );
  AOI22_X1 U4290 ( .A1(n27754), .A2(\xmem_data[104][6] ), .B1(n30237), .B2(
        \xmem_data[105][6] ), .ZN(n12277) );
  INV_X1 U4291 ( .A(n4781), .ZN(n4786) );
  NOR2_X1 U4292 ( .A1(n13840), .A2(n13839), .ZN(n13841) );
  INV_X1 U4293 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U4294 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  INV_X1 U4295 ( .A(n10457), .ZN(n10461) );
  INV_X1 U4296 ( .A(n10452), .ZN(n10453) );
  NOR2_X1 U4297 ( .A1(n10447), .A2(n10446), .ZN(n10464) );
  NAND2_X1 U4298 ( .A1(n10433), .A2(n10432), .ZN(n10447) );
  NAND2_X1 U4299 ( .A1(n21010), .A2(\xmem_data[6][5] ), .ZN(n10432) );
  NOR2_X1 U4300 ( .A1(n11983), .A2(n11982), .ZN(n11984) );
  NAND2_X1 U4301 ( .A1(n11981), .A2(n11980), .ZN(n11982) );
  NAND2_X1 U4302 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  AND4_X1 U4303 ( .A1(n18033), .A2(n18032), .A3(n18031), .A4(n18030), .ZN(
        n18036) );
  AOI22_X1 U4304 ( .A1(n27710), .A2(\xmem_data[28][4] ), .B1(n30707), .B2(
        \xmem_data[29][4] ), .ZN(n8173) );
  NOR2_X1 U4305 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  INV_X1 U4306 ( .A(n24482), .ZN(n24485) );
  AND2_X1 U4307 ( .A1(n24443), .A2(\xmem_data[2][7] ), .ZN(n14474) );
  AND2_X1 U4308 ( .A1(n24470), .A2(\xmem_data[31][7] ), .ZN(n14473) );
  INV_X1 U4309 ( .A(n23444), .ZN(n23445) );
  INV_X1 U4310 ( .A(n3343), .ZN(n3344) );
  NAND3_X1 U4311 ( .A1(n18828), .A2(n18827), .A3(n18826), .ZN(n18829) );
  AND4_X1 U4312 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11898) );
  NAND2_X1 U4313 ( .A1(n29272), .A2(\xmem_data[6][3] ), .ZN(n22478) );
  AND4_X1 U4314 ( .A1(n15611), .A2(n15610), .A3(n15609), .A4(n15608), .ZN(
        n15628) );
  NAND3_X1 U4315 ( .A1(n8746), .A2(n8745), .A3(n8744), .ZN(n8747) );
  INV_X1 U4316 ( .A(n4634), .ZN(n4635) );
  OR2_X1 U4317 ( .A1(n16405), .A2(n16404), .ZN(n16406) );
  OR2_X1 U4318 ( .A1(n24619), .A2(n24618), .ZN(n24621) );
  NAND2_X1 U4319 ( .A1(n24617), .A2(n24616), .ZN(n24618) );
  NAND2_X1 U4320 ( .A1(n24615), .A2(\xmem_data[30][3] ), .ZN(n24616) );
  OAI21_X1 U4321 ( .B1(n5954), .B2(n5953), .A(n31284), .ZN(n5955) );
  OR4_X1 U4322 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n5953) );
  NAND2_X1 U4323 ( .A1(n9843), .A2(n27935), .ZN(n9872) );
  OR4_X1 U4324 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n9843) );
  NAND3_X1 U4325 ( .A1(n15798), .A2(n15797), .A3(n15796), .ZN(n15799) );
  OR4_X1 U4326 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n5429) );
  OR3_X1 U4327 ( .A1(n5379), .A2(n5378), .A3(n5377), .ZN(n5385) );
  NAND2_X1 U4328 ( .A1(n5407), .A2(n29041), .ZN(n5453) );
  OR4_X1 U4329 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(n5407) );
  XNOR2_X1 U4330 ( .A(n35178), .B(\fmem_data[20][3] ), .ZN(n32012) );
  XNOR2_X1 U4331 ( .A(n31489), .B(\fmem_data[21][5] ), .ZN(n33269) );
  NAND2_X1 U4332 ( .A1(n34688), .A2(n34687), .ZN(n34689) );
  XNOR2_X1 U4333 ( .A(n33227), .B(\fmem_data[14][7] ), .ZN(n33311) );
  XNOR2_X1 U4334 ( .A(n32543), .B(\fmem_data[17][7] ), .ZN(n33313) );
  NAND2_X1 U4335 ( .A1(n30476), .A2(n30475), .ZN(n30461) );
  XNOR2_X1 U4336 ( .A(n32528), .B(\fmem_data[29][7] ), .ZN(n30449) );
  NOR2_X1 U4337 ( .A1(n31867), .A2(n31866), .ZN(n30372) );
  NAND2_X1 U4338 ( .A1(n31867), .A2(n31866), .ZN(n30371) );
  INV_X1 U4339 ( .A(n30351), .ZN(n31695) );
  AOI21_X1 U4340 ( .B1(n34472), .B2(n34474), .A(n30350), .ZN(n30351) );
  XNOR2_X1 U4341 ( .A(n33039), .B(\fmem_data[0][5] ), .ZN(n33386) );
  AOI21_X1 U4342 ( .B1(n33059), .B2(n33057), .A(n33060), .ZN(n13213) );
  XNOR2_X1 U4343 ( .A(n35023), .B(\fmem_data[5][5] ), .ZN(n33309) );
  XNOR2_X1 U4344 ( .A(n30156), .B(\fmem_data[28][7] ), .ZN(n33317) );
  XNOR2_X1 U4345 ( .A(n31817), .B(\fmem_data[19][5] ), .ZN(n33219) );
  XNOR2_X1 U4346 ( .A(n35072), .B(\fmem_data[22][5] ), .ZN(n33130) );
  AND2_X1 U4347 ( .A1(n25492), .A2(\xmem_data[6][7] ), .ZN(n24146) );
  XNOR2_X1 U4348 ( .A(n31638), .B(\fmem_data[24][7] ), .ZN(n31816) );
  XNOR2_X1 U4349 ( .A(n31664), .B(\fmem_data[22][7] ), .ZN(n35177) );
  XNOR2_X1 U4350 ( .A(n31640), .B(\fmem_data[0][7] ), .ZN(n31824) );
  XNOR2_X1 U4351 ( .A(n34929), .B(\fmem_data[6][5] ), .ZN(n33369) );
  AOI21_X1 U4352 ( .B1(n35089), .B2(n35088), .A(n35087), .ZN(n35090) );
  AOI21_X1 U4353 ( .B1(n33828), .B2(n33827), .A(n33323), .ZN(n31676) );
  XNOR2_X1 U4354 ( .A(n31656), .B(\fmem_data[28][7] ), .ZN(n33318) );
  XNOR2_X1 U4355 ( .A(n31704), .B(\fmem_data[17][7] ), .ZN(n33314) );
  INV_X1 U4356 ( .A(n3327), .ZN(n3302) );
  NAND4_X1 U4357 ( .A1(n31025), .A2(n31024), .A3(n31023), .A4(n31022), .ZN(
        n31040) );
  NAND4_X1 U4358 ( .A1(n17309), .A2(n17308), .A3(n17307), .A4(n17306), .ZN(
        n17315) );
  NAND2_X1 U4359 ( .A1(n22858), .A2(n22857), .ZN(n22864) );
  NOR2_X1 U4360 ( .A1(n22856), .A2(n22855), .ZN(n22857) );
  NAND2_X1 U4361 ( .A1(n13475), .A2(\xmem_data[31][1] ), .ZN(n22852) );
  INV_X1 U4362 ( .A(n3432), .ZN(n3433) );
  NAND3_X1 U4363 ( .A1(n29129), .A2(n29128), .A3(n29127), .ZN(n29134) );
  NAND3_X1 U4364 ( .A1(n29132), .A2(n29131), .A3(n29130), .ZN(n29133) );
  NAND2_X1 U4365 ( .A1(n9113), .A2(n9112), .ZN(n32163) );
  XNOR2_X1 U4366 ( .A(n36101), .B(\fmem_data[24][7] ), .ZN(n32665) );
  XNOR2_X1 U4367 ( .A(n33677), .B(\fmem_data[30][7] ), .ZN(n32668) );
  AOI21_X1 U4368 ( .B1(n36295), .B2(n3564), .A(n31966), .ZN(n31967) );
  AOI21_X1 U4369 ( .B1(n34745), .B2(n3562), .A(n31959), .ZN(n31960) );
  XNOR2_X1 U4370 ( .A(n33214), .B(\fmem_data[24][3] ), .ZN(n30983) );
  OAI21_X1 U4371 ( .B1(n30423), .B2(n34537), .A(n30422), .ZN(n30824) );
  INV_X1 U4372 ( .A(n34535), .ZN(n30421) );
  OAI21_X1 U4373 ( .B1(n14352), .B2(n14351), .A(n31342), .ZN(n14380) );
  OAI21_X1 U4374 ( .B1(n14331), .B2(n14330), .A(n31376), .ZN(n14381) );
  XNOR2_X1 U4375 ( .A(n32131), .B(\fmem_data[4][7] ), .ZN(n30408) );
  XNOR2_X1 U4376 ( .A(n32065), .B(\fmem_data[0][7] ), .ZN(n30447) );
  XNOR2_X1 U4377 ( .A(n31664), .B(\fmem_data[22][5] ), .ZN(n33224) );
  XNOR2_X1 U4378 ( .A(n32600), .B(\fmem_data[14][7] ), .ZN(n33228) );
  OAI21_X1 U4379 ( .B1(n15304), .B2(n15303), .A(n10213), .ZN(n15305) );
  NAND4_X1 U4380 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n31233)
         );
  NAND2_X1 U4381 ( .A1(n7179), .A2(n30704), .ZN(n7186) );
  NAND2_X1 U4382 ( .A1(n7174), .A2(n30782), .ZN(n7187) );
  NAND2_X1 U4383 ( .A1(n7112), .A2(n30704), .ZN(n7130) );
  NAND2_X1 U4384 ( .A1(n7127), .A2(n30659), .ZN(n7128) );
  NAND2_X1 U4385 ( .A1(n7100), .A2(n30782), .ZN(n7107) );
  NAND4_X1 U4386 ( .A1(n7164), .A2(n7163), .A3(n7162), .A4(n7161), .ZN(n7190)
         );
  AOI22_X1 U4387 ( .A1(n30782), .A2(n7155), .B1(n7154), .B2(n30659), .ZN(n7162) );
  NAND2_X1 U4388 ( .A1(n7135), .A2(n30659), .ZN(n7164) );
  NAND4_X1 U4389 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n31670)
         );
  NAND3_X1 U4390 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n31673) );
  OR2_X1 U4391 ( .A1(n4363), .A2(n22877), .ZN(n4364) );
  NAND3_X1 U4392 ( .A1(n4866), .A2(n4865), .A3(n4864), .ZN(n31958) );
  XNOR2_X1 U4393 ( .A(n33451), .B(\fmem_data[9][5] ), .ZN(n33846) );
  OAI21_X1 U4394 ( .B1(n7564), .B2(n7563), .A(n27801), .ZN(n7591) );
  NAND3_X1 U4395 ( .A1(n18042), .A2(n18041), .A3(n18040), .ZN(n30846) );
  OR2_X1 U4396 ( .A1(n18039), .A2(n24151), .ZN(n18040) );
  XNOR2_X1 U4397 ( .A(n32584), .B(\fmem_data[4][1] ), .ZN(n33648) );
  XNOR2_X1 U4398 ( .A(n31958), .B(\fmem_data[6][5] ), .ZN(n33187) );
  XNOR2_X1 U4399 ( .A(n31250), .B(\fmem_data[1][5] ), .ZN(n31973) );
  XNOR2_X1 U4400 ( .A(n31957), .B(\fmem_data[6][5] ), .ZN(n33957) );
  XNOR2_X1 U4401 ( .A(n31995), .B(\fmem_data[8][3] ), .ZN(n33968) );
  OR2_X1 U4402 ( .A1(n36112), .A2(n3615), .ZN(n33926) );
  XNOR2_X1 U4403 ( .A(n31669), .B(\fmem_data[13][1] ), .ZN(n33927) );
  XNOR2_X1 U4404 ( .A(n35104), .B(\fmem_data[13][1] ), .ZN(n33928) );
  NAND2_X1 U4405 ( .A1(n33901), .A2(n33900), .ZN(n33902) );
  XNOR2_X1 U4406 ( .A(n33789), .B(\fmem_data[30][7] ), .ZN(n31984) );
  XNOR2_X1 U4407 ( .A(n33551), .B(\fmem_data[20][5] ), .ZN(n32523) );
  XNOR2_X1 U4408 ( .A(n30406), .B(n30405), .ZN(n32347) );
  XNOR2_X1 U4409 ( .A(n30404), .B(n30403), .ZN(n30406) );
  XNOR2_X1 U4410 ( .A(n32025), .B(\fmem_data[12][5] ), .ZN(n33976) );
  XNOR2_X1 U4411 ( .A(n31800), .B(\fmem_data[29][3] ), .ZN(n32320) );
  INV_X1 U4412 ( .A(n32327), .ZN(n32293) );
  AOI21_X1 U4413 ( .B1(n34739), .B2(n3563), .A(n33970), .ZN(n30827) );
  NAND2_X1 U4414 ( .A1(n32348), .A2(n32347), .ZN(n30411) );
  XNOR2_X1 U4415 ( .A(n31592), .B(\fmem_data[29][7] ), .ZN(n30450) );
  XNOR2_X1 U4416 ( .A(n32582), .B(\fmem_data[10][7] ), .ZN(n33387) );
  AOI21_X1 U4417 ( .B1(n33741), .B2(n33603), .A(n25602), .ZN(n6585) );
  OAI22_X1 U4418 ( .A1(n33325), .A2(n35722), .B1(n33324), .B2(n35721), .ZN(
        n34830) );
  OAI22_X1 U4419 ( .A1(n33318), .A2(n35761), .B1(n33317), .B2(n35760), .ZN(
        n34840) );
  OAI22_X1 U4420 ( .A1(n33316), .A2(n35516), .B1(n33315), .B2(n35515), .ZN(
        n34839) );
  XNOR2_X1 U4421 ( .A(n32597), .B(\fmem_data[15][7] ), .ZN(n33235) );
  OAI22_X1 U4422 ( .A1(n33253), .A2(n35037), .B1(n33252), .B2(n35036), .ZN(
        n33377) );
  XNOR2_X1 U4423 ( .A(n31655), .B(\fmem_data[30][7] ), .ZN(n33307) );
  XNOR2_X1 U4424 ( .A(n31658), .B(\fmem_data[30][7] ), .ZN(n33308) );
  NAND2_X1 U4425 ( .A1(n31756), .A2(n31757), .ZN(n30342) );
  AOI21_X1 U4426 ( .B1(n34909), .B2(n34908), .A(n34907), .ZN(n34910) );
  XNOR2_X1 U4427 ( .A(n31668), .B(\fmem_data[13][7] ), .ZN(n33133) );
  XNOR2_X1 U4428 ( .A(n35316), .B(\fmem_data[15][5] ), .ZN(n34988) );
  OAI22_X1 U4429 ( .A1(n30459), .A2(n35740), .B1(n31643), .B2(n35739), .ZN(
        n34876) );
  OAI22_X1 U4430 ( .A1(n24016), .A2(n35004), .B1(n31826), .B2(n35003), .ZN(
        n34877) );
  OAI22_X1 U4431 ( .A1(n34984), .A2(n34986), .B1(n31825), .B2(n34985), .ZN(
        n34882) );
  OAI22_X1 U4432 ( .A1(n31826), .A2(n35004), .B1(n35005), .B2(n35003), .ZN(
        n34881) );
  OR2_X1 U4433 ( .A1(n32021), .A2(n3956), .ZN(n26032) );
  XNOR2_X1 U4434 ( .A(n31892), .B(\fmem_data[1][5] ), .ZN(n31972) );
  OR2_X1 U4435 ( .A1(n33127), .A2(n3943), .ZN(n35125) );
  AOI21_X1 U4436 ( .B1(n13997), .B2(n13996), .A(n13995), .ZN(n13998) );
  INV_X1 U4437 ( .A(n30009), .ZN(n13995) );
  NOR2_X1 U4438 ( .A1(n13984), .A2(n13983), .ZN(n13997) );
  NOR2_X1 U4439 ( .A1(n13994), .A2(n13993), .ZN(n13996) );
  NAND2_X1 U4440 ( .A1(n10260), .A2(n10259), .ZN(n31674) );
  NAND3_X1 U4441 ( .A1(n14768), .A2(n14767), .A3(n14766), .ZN(n31705) );
  NAND2_X1 U4442 ( .A1(n14734), .A2(n25593), .ZN(n14767) );
  NAND3_X1 U4443 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n31659) );
  NAND4_X1 U4444 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n35238) );
  NAND2_X1 U4445 ( .A1(n16749), .A2(n28490), .ZN(n16750) );
  INV_X1 U4446 ( .A(n16728), .ZN(n16751) );
  NAND2_X1 U4447 ( .A1(n16661), .A2(n16660), .ZN(n35355) );
  NAND3_X1 U4448 ( .A1(n4155), .A2(n4154), .A3(n4153), .ZN(n35120) );
  OAI21_X1 U4449 ( .B1(n25507), .B2(n25506), .A(n19110), .ZN(n25597) );
  OAI22_X1 U4450 ( .A1(n31824), .A2(n35493), .B1(n35402), .B2(n35494), .ZN(
        n35133) );
  INV_X1 U4451 ( .A(n35124), .ZN(n35129) );
  NOR2_X1 U4452 ( .A1(n35126), .A2(n35125), .ZN(n35128) );
  NAND2_X1 U4453 ( .A1(n35126), .A2(n35125), .ZN(n35127) );
  XNOR2_X1 U4454 ( .A(n31817), .B(\fmem_data[19][7] ), .ZN(n35271) );
  OAI21_X1 U4455 ( .B1(n35274), .B2(n35273), .A(n35272), .ZN(n35276) );
  OAI22_X1 U4456 ( .A1(n34983), .A2(n35744), .B1(n35327), .B2(n35745), .ZN(
        n35268) );
  OAI22_X1 U4457 ( .A1(n34981), .A2(n35752), .B1(n35398), .B2(n35753), .ZN(
        n35269) );
  AND2_X1 U4458 ( .A1(n37199), .A2(n6586), .ZN(n6485) );
  AND2_X1 U4459 ( .A1(n4062), .A2(n4049), .ZN(n4078) );
  OR2_X1 U4460 ( .A1(n27203), .A2(n27202), .ZN(n27204) );
  AOI22_X1 U4461 ( .A1(n29647), .A2(\xmem_data[48][1] ), .B1(n29589), .B2(
        \xmem_data[49][1] ), .ZN(n26670) );
  OR2_X1 U4462 ( .A1(n19329), .A2(n19328), .ZN(n19331) );
  NAND2_X1 U4463 ( .A1(n24457), .A2(\xmem_data[17][1] ), .ZN(n17780) );
  NAND3_X1 U4464 ( .A1(n3711), .A2(n29200), .A3(n29199), .ZN(n29202) );
  NAND4_X1 U4465 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n32978) );
  OR2_X1 U4466 ( .A1(n36111), .A2(n3658), .ZN(n32781) );
  XNOR2_X1 U4467 ( .A(n32225), .B(\fmem_data[9][1] ), .ZN(n34198) );
  XNOR2_X1 U4468 ( .A(n32115), .B(\fmem_data[21][3] ), .ZN(n34202) );
  NAND2_X1 U4469 ( .A1(n34355), .A2(n34354), .ZN(n34356) );
  XNOR2_X1 U4470 ( .A(n34531), .B(\fmem_data[10][3] ), .ZN(n33590) );
  AND2_X1 U4471 ( .A1(n28534), .A2(n26485), .ZN(n31470) );
  XNOR2_X1 U4472 ( .A(n31899), .B(\fmem_data[20][1] ), .ZN(n32059) );
  XNOR2_X1 U4473 ( .A(n32115), .B(\fmem_data[21][1] ), .ZN(n32058) );
  XNOR2_X1 U4474 ( .A(n33451), .B(\fmem_data[9][3] ), .ZN(n32783) );
  XNOR2_X1 U4475 ( .A(n33743), .B(\fmem_data[9][3] ), .ZN(n31394) );
  OR2_X1 U4476 ( .A1(n36315), .A2(n3688), .ZN(n31245) );
  XNOR2_X1 U4477 ( .A(n31900), .B(\fmem_data[20][1] ), .ZN(n31446) );
  XNOR2_X1 U4478 ( .A(n33594), .B(\fmem_data[29][5] ), .ZN(n31173) );
  OR2_X1 U4479 ( .A1(n36312), .A2(n3595), .ZN(n31912) );
  XNOR2_X1 U4480 ( .A(n31638), .B(\fmem_data[24][1] ), .ZN(n31911) );
  XNOR2_X1 U4481 ( .A(n34615), .B(\fmem_data[21][3] ), .ZN(n32066) );
  NAND2_X1 U4482 ( .A1(n16466), .A2(n3955), .ZN(n16467) );
  NAND3_X1 U4483 ( .A1(n18721), .A2(n18720), .A3(n18719), .ZN(n32615) );
  OAI22_X1 U4484 ( .A1(n34346), .A2(n36226), .B1(n32426), .B2(n3633), .ZN(
        n32867) );
  XNOR2_X1 U4485 ( .A(n33967), .B(\fmem_data[8][1] ), .ZN(n32428) );
  XNOR2_X1 U4486 ( .A(n31995), .B(\fmem_data[8][1] ), .ZN(n32126) );
  XNOR2_X1 U4487 ( .A(n31899), .B(\fmem_data[20][3] ), .ZN(n32128) );
  XNOR2_X1 U4488 ( .A(n36112), .B(\fmem_data[12][5] ), .ZN(n32136) );
  XNOR2_X1 U4489 ( .A(n32582), .B(\fmem_data[10][1] ), .ZN(n33600) );
  XNOR2_X1 U4490 ( .A(n32612), .B(\fmem_data[30][1] ), .ZN(n34790) );
  OAI22_X1 U4491 ( .A1(n32424), .A2(n33850), .B1(n32423), .B2(n33851), .ZN(
        n34791) );
  OAI22_X1 U4492 ( .A1(n32420), .A2(n3576), .B1(n34482), .B2(n34483), .ZN(
        n34793) );
  OAI21_X1 U4493 ( .B1(n32687), .B2(n32686), .A(n32685), .ZN(n32123) );
  NAND2_X1 U4494 ( .A1(n32687), .A2(n32686), .ZN(n32122) );
  AND2_X1 U4495 ( .A1(n36101), .A2(n32578), .ZN(n32692) );
  XNOR2_X1 U4496 ( .A(n32979), .B(\fmem_data[4][3] ), .ZN(n32690) );
  OR2_X1 U4497 ( .A1(n36112), .A2(n3589), .ZN(n32239) );
  NAND2_X1 U4498 ( .A1(n14383), .A2(n33975), .ZN(n33973) );
  AND2_X1 U4499 ( .A1(n36112), .A2(n32285), .ZN(n32663) );
  NAND2_X1 U4500 ( .A1(n32568), .A2(n32567), .ZN(n32569) );
  XNOR2_X1 U4501 ( .A(n33594), .B(\fmem_data[29][7] ), .ZN(n32651) );
  OAI22_X1 U4502 ( .A1(n32177), .A2(n34779), .B1(n33994), .B2(n34466), .ZN(
        n32332) );
  OAI22_X1 U4503 ( .A1(n32180), .A2(n35700), .B1(n32179), .B2(n35701), .ZN(
        n32336) );
  XNOR2_X1 U4504 ( .A(\fmem_data[18][2] ), .B(\fmem_data[18][1] ), .ZN(n33681)
         );
  NAND2_X1 U4505 ( .A1(n25145), .A2(n33681), .ZN(n33679) );
  XOR2_X1 U4506 ( .A(\fmem_data[18][2] ), .B(\fmem_data[18][3] ), .Z(n25145)
         );
  XNOR2_X1 U4507 ( .A(n31704), .B(\fmem_data[17][1] ), .ZN(n32544) );
  XNOR2_X1 U4508 ( .A(n31738), .B(n31737), .ZN(n30832) );
  OAI22_X1 U4509 ( .A1(n32516), .A2(n35748), .B1(n30408), .B2(n35749), .ZN(
        n31007) );
  XNOR2_X1 U4510 ( .A(n3390), .B(\fmem_data[10][3] ), .ZN(n32572) );
  XNOR2_X1 U4511 ( .A(n32065), .B(\fmem_data[0][5] ), .ZN(n32562) );
  XNOR2_X1 U4512 ( .A(n34615), .B(\fmem_data[21][7] ), .ZN(n20613) );
  XNOR2_X1 U4513 ( .A(n34929), .B(\fmem_data[6][1] ), .ZN(n34016) );
  INV_X1 U4514 ( .A(n36240), .ZN(n17753) );
  XNOR2_X1 U4515 ( .A(n33556), .B(\fmem_data[16][7] ), .ZN(n31888) );
  NAND2_X1 U4516 ( .A1(n3586), .A2(n16566), .ZN(n16567) );
  INV_X1 U4517 ( .A(n26799), .ZN(n16566) );
  XNOR2_X1 U4518 ( .A(\fmem_data[21][3] ), .B(\fmem_data[21][4] ), .ZN(n34195)
         );
  NAND2_X1 U4519 ( .A1(n19905), .A2(n34195), .ZN(n34194) );
  XOR2_X1 U4520 ( .A(\fmem_data[21][5] ), .B(\fmem_data[21][4] ), .Z(n19905)
         );
  XNOR2_X1 U4521 ( .A(n32582), .B(\fmem_data[10][3] ), .ZN(n30817) );
  NAND2_X1 U4522 ( .A1(n16662), .A2(n34736), .ZN(n33690) );
  NAND2_X1 U4523 ( .A1(n23919), .A2(n35041), .ZN(n35040) );
  XNOR2_X1 U4524 ( .A(n31233), .B(\fmem_data[5][3] ), .ZN(n32229) );
  XNOR2_X1 U4525 ( .A(n34862), .B(\fmem_data[16][3] ), .ZN(n34038) );
  XNOR2_X1 U4526 ( .A(n33484), .B(\fmem_data[31][7] ), .ZN(n26148) );
  XNOR2_X1 U4527 ( .A(n32614), .B(\fmem_data[24][5] ), .ZN(n34042) );
  OR2_X1 U4528 ( .A1(n36101), .A2(n3599), .ZN(n27581) );
  XNOR2_X1 U4529 ( .A(\fmem_data[2][4] ), .B(\fmem_data[2][3] ), .ZN(n35019)
         );
  XNOR2_X1 U4530 ( .A(n32317), .B(\fmem_data[4][3] ), .ZN(n32132) );
  NAND2_X1 U4531 ( .A1(n13406), .A2(n33963), .ZN(n33961) );
  NAND2_X1 U4532 ( .A1(n6555), .A2(n27935), .ZN(n6583) );
  OAI21_X1 U4533 ( .B1(n6581), .B2(n6580), .A(n9896), .ZN(n6582) );
  AOI22_X1 U4534 ( .A1(n27968), .A2(n6533), .B1(n6532), .B2(n27937), .ZN(n6584) );
  INV_X1 U4535 ( .A(n6457), .ZN(n6480) );
  INV_X1 U4536 ( .A(n9899), .ZN(n9971) );
  NAND2_X1 U4537 ( .A1(n14471), .A2(n14470), .ZN(n31663) );
  XNOR2_X1 U4538 ( .A(n32882), .B(\fmem_data[6][5] ), .ZN(n32576) );
  XNOR2_X1 U4539 ( .A(\fmem_data[6][3] ), .B(\fmem_data[6][4] ), .ZN(n33956)
         );
  NAND2_X1 U4540 ( .A1(n28541), .A2(n33956), .ZN(n33954) );
  XOR2_X1 U4541 ( .A(\fmem_data[6][5] ), .B(\fmem_data[6][4] ), .Z(n28541) );
  NAND2_X1 U4542 ( .A1(n7399), .A2(n34919), .ZN(n34918) );
  XNOR2_X1 U4543 ( .A(n30451), .B(\fmem_data[6][3] ), .ZN(n31881) );
  XNOR2_X1 U4544 ( .A(n32427), .B(\fmem_data[8][5] ), .ZN(n30819) );
  XNOR2_X1 U4545 ( .A(n33967), .B(\fmem_data[8][5] ), .ZN(n24015) );
  OAI22_X1 U4546 ( .A1(n32125), .A2(n34416), .B1(n32003), .B2(n34414), .ZN(
        n31387) );
  AND2_X1 U4547 ( .A1(n36315), .A2(n29517), .ZN(n31388) );
  OAI22_X1 U4548 ( .A1(n27433), .A2(n35745), .B1(n35744), .B2(n3622), .ZN(
        n30492) );
  XNOR2_X1 U4549 ( .A(n32176), .B(\fmem_data[1][5] ), .ZN(n30169) );
  XNOR2_X1 U4550 ( .A(n35073), .B(\fmem_data[22][3] ), .ZN(n30370) );
  XNOR2_X1 U4551 ( .A(n33227), .B(\fmem_data[14][5] ), .ZN(n30415) );
  XNOR2_X1 U4552 ( .A(n33225), .B(\fmem_data[16][5] ), .ZN(n32016) );
  XNOR2_X1 U4553 ( .A(n32939), .B(\fmem_data[1][5] ), .ZN(n31243) );
  NAND2_X1 U4554 ( .A1(n36057), .A2(n36056), .ZN(n34369) );
  XNOR2_X1 U4555 ( .A(n31492), .B(\fmem_data[25][1] ), .ZN(n34441) );
  XNOR2_X1 U4556 ( .A(n33677), .B(\fmem_data[30][3] ), .ZN(n34438) );
  AND2_X1 U4557 ( .A1(n36315), .A2(n33705), .ZN(n33822) );
  OAI22_X1 U4558 ( .A1(n22778), .A2(n33859), .B1(n31884), .B2(n33857), .ZN(
        n29533) );
  OAI22_X1 U4559 ( .A1(n22775), .A2(n35498), .B1(n22774), .B2(n35497), .ZN(
        n29535) );
  OAI22_X1 U4560 ( .A1(n22777), .A2(n35722), .B1(n22776), .B2(n35721), .ZN(
        n29534) );
  OAI22_X1 U4561 ( .A1(n33878), .A2(n36227), .B1(n33877), .B2(n3647), .ZN(
        n34014) );
  XNOR2_X1 U4562 ( .A(n31958), .B(\fmem_data[6][1] ), .ZN(n33811) );
  NAND2_X1 U4563 ( .A1(n24437), .A2(n33328), .ZN(n33326) );
  XNOR2_X1 U4564 ( .A(n33789), .B(\fmem_data[30][5] ), .ZN(n30997) );
  NAND2_X1 U4565 ( .A1(n18722), .A2(n34039), .ZN(n34041) );
  OAI21_X1 U4566 ( .B1(n33891), .B2(n33890), .A(n33889), .ZN(n33893) );
  OAI22_X1 U4567 ( .A1(n33794), .A2(n34986), .B1(n34985), .B2(n3644), .ZN(
        n33869) );
  OAI22_X1 U4568 ( .A1(n33795), .A2(n35036), .B1(n35037), .B2(n3628), .ZN(
        n33868) );
  XNOR2_X1 U4569 ( .A(\fmem_data[4][4] ), .B(\fmem_data[4][3] ), .ZN(n35011)
         );
  NAND2_X1 U4570 ( .A1(n13015), .A2(n35011), .ZN(n35010) );
  XOR2_X1 U4571 ( .A(\fmem_data[4][4] ), .B(\fmem_data[4][5] ), .Z(n13015) );
  XNOR2_X1 U4572 ( .A(n31592), .B(\fmem_data[29][5] ), .ZN(n33186) );
  XNOR2_X1 U4573 ( .A(n31125), .B(\fmem_data[0][5] ), .ZN(n33183) );
  XNOR2_X1 U4574 ( .A(n32242), .B(\fmem_data[29][5] ), .ZN(n33185) );
  NAND2_X1 U4575 ( .A1(n10562), .A2(n33643), .ZN(n33642) );
  NAND2_X1 U4576 ( .A1(n15404), .A2(n35083), .ZN(n35084) );
  XNOR2_X1 U4577 ( .A(n35023), .B(\fmem_data[5][3] ), .ZN(n33180) );
  XNOR2_X1 U4578 ( .A(n34211), .B(n34210), .ZN(n34212) );
  XNOR2_X1 U4579 ( .A(n33967), .B(\fmem_data[8][3] ), .ZN(n34207) );
  NAND2_X1 U4580 ( .A1(n6075), .A2(n35182), .ZN(n35181) );
  NAND2_X1 U4581 ( .A1(n9972), .A2(n34201), .ZN(n34199) );
  XNOR2_X1 U4582 ( .A(n32600), .B(\fmem_data[14][5] ), .ZN(n32734) );
  XNOR2_X1 U4583 ( .A(n33592), .B(\fmem_data[14][5] ), .ZN(n32733) );
  NAND2_X1 U4584 ( .A1(n9875), .A2(n33100), .ZN(n33098) );
  OAI22_X1 U4585 ( .A1(n31954), .A2(n35490), .B1(n31953), .B2(n35489), .ZN(
        n33081) );
  OAI22_X1 U4586 ( .A1(n29208), .A2(n33057), .B1(n33058), .B2(n33059), .ZN(
        n34077) );
  NAND2_X1 U4587 ( .A1(n8197), .A2(n34932), .ZN(n34933) );
  OAI22_X1 U4588 ( .A1(n34042), .A2(n34041), .B1(n34040), .B2(n34039), .ZN(
        n34263) );
  OAI22_X1 U4589 ( .A1(n34233), .A2(n34835), .B1(n34232), .B2(n34836), .ZN(
        n34664) );
  OAI22_X1 U4590 ( .A1(n34235), .A2(n34909), .B1(n34234), .B2(n34908), .ZN(
        n34663) );
  NAND2_X1 U4591 ( .A1(n21397), .A2(n21396), .ZN(n34004) );
  XNOR2_X1 U4592 ( .A(n32211), .B(\fmem_data[15][3] ), .ZN(n32751) );
  OAI22_X1 U4593 ( .A1(n32755), .A2(n33827), .B1(n32754), .B2(n33828), .ZN(
        n33255) );
  OAI22_X1 U4594 ( .A1(n32757), .A2(n35507), .B1(n32756), .B2(n35508), .ZN(
        n33254) );
  XNOR2_X1 U4595 ( .A(n35030), .B(\fmem_data[15][3] ), .ZN(n33169) );
  OAI22_X1 U4596 ( .A1(n32525), .A2(n3562), .B1(n32524), .B2(n34745), .ZN(
        n32777) );
  OAI22_X1 U4597 ( .A1(n32523), .A2(n35037), .B1(n32522), .B2(n35036), .ZN(
        n32791) );
  NAND2_X1 U4598 ( .A1(n30470), .A2(n30469), .ZN(n31732) );
  XNOR2_X1 U4599 ( .A(n30809), .B(n30808), .ZN(n30810) );
  XNOR2_X1 U4600 ( .A(n30836), .B(n30835), .ZN(n31932) );
  AND2_X1 U4601 ( .A1(n34363), .A2(n34364), .ZN(n24114) );
  NAND2_X1 U4602 ( .A1(n34977), .A2(n34976), .ZN(n34978) );
  INV_X1 U4603 ( .A(n31714), .ZN(n31719) );
  XNOR2_X1 U4604 ( .A(n35013), .B(n35272), .ZN(n35279) );
  XNOR2_X1 U4605 ( .A(n35273), .B(n35274), .ZN(n35013) );
  NAND4_X1 U4606 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n35270)
         );
  NAND2_X1 U4607 ( .A1(n26023), .A2(n35652), .ZN(n35651) );
  XNOR2_X1 U4608 ( .A(n31674), .B(\fmem_data[10][7] ), .ZN(n35356) );
  XNOR2_X1 U4609 ( .A(n31705), .B(\fmem_data[17][7] ), .ZN(n35075) );
  XNOR2_X1 U4610 ( .A(n31659), .B(\fmem_data[30][7] ), .ZN(n35077) );
  XNOR2_X1 U4611 ( .A(n31799), .B(\fmem_data[14][7] ), .ZN(n35103) );
  NAND2_X1 U4612 ( .A1(n14873), .A2(n35634), .ZN(n35633) );
  NAND2_X1 U4613 ( .A1(n7991), .A2(n35638), .ZN(n35637) );
  NAND2_X1 U4614 ( .A1(n11955), .A2(n35642), .ZN(n35641) );
  XNOR2_X1 U4615 ( .A(n35357), .B(\fmem_data[29][7] ), .ZN(n35613) );
  NAND2_X1 U4616 ( .A1(n15016), .A2(n35615), .ZN(n35614) );
  XNOR2_X1 U4617 ( .A(n35120), .B(\fmem_data[6][7] ), .ZN(n35510) );
  XNOR2_X1 U4618 ( .A(n35122), .B(\fmem_data[12][7] ), .ZN(n35514) );
  NAND2_X1 U4619 ( .A1(n16944), .A2(n35577), .ZN(n35576) );
  XNOR2_X1 U4620 ( .A(n35102), .B(\fmem_data[14][7] ), .ZN(n35575) );
  NAND2_X1 U4621 ( .A1(n4577), .A2(n35585), .ZN(n35584) );
  OAI22_X1 U4622 ( .A1(n35699), .A2(n35701), .B1(n35281), .B2(n35700), .ZN(
        n35523) );
  NAND2_X1 U4623 ( .A1(n35286), .A2(n35285), .ZN(n35522) );
  NAND2_X1 U4624 ( .A1(n35284), .A2(n35283), .ZN(n35285) );
  OAI22_X1 U4625 ( .A1(n35695), .A2(n35697), .B1(n35317), .B2(n35696), .ZN(
        n35573) );
  INV_X1 U4626 ( .A(n3423), .ZN(n3335) );
  NAND2_X1 U4627 ( .A1(n6487), .A2(n6488), .ZN(n6489) );
  INV_X1 U4628 ( .A(n13429), .ZN(n6487) );
  BUF_X2 U4629 ( .A(n7446), .Z(n27804) );
  INV_X1 U4630 ( .A(n21310), .ZN(n21317) );
  NAND2_X1 U4631 ( .A1(n21314), .A2(n21313), .ZN(n21315) );
  AND4_X1 U4632 ( .A1(n21325), .A2(n21324), .A3(n21323), .A4(n21322), .ZN(
        n21326) );
  BUF_X2 U4633 ( .A(n8700), .Z(n26884) );
  OR4_X1 U4634 ( .A1(n22998), .A2(n22997), .A3(n22996), .A4(n22995), .ZN(
        n22999) );
  NAND4_X1 U4635 ( .A1(n17368), .A2(n17367), .A3(n17366), .A4(n17365), .ZN(
        n33749) );
  NAND2_X1 U4636 ( .A1(n17296), .A2(n24236), .ZN(n17368) );
  NAND4_X1 U4637 ( .A1(n19506), .A2(n19505), .A3(n19504), .A4(n19503), .ZN(
        n32127) );
  NAND3_X1 U4638 ( .A1(n19608), .A2(n19607), .A3(n19606), .ZN(n33756) );
  XNOR2_X1 U4639 ( .A(n32065), .B(\fmem_data[0][1] ), .ZN(n33755) );
  OAI22_X1 U4640 ( .A1(n34530), .A2(n34529), .B1(n34528), .B2(n3566), .ZN(
        n36118) );
  XNOR2_X1 U4641 ( .A(n33733), .B(\fmem_data[11][3] ), .ZN(n34430) );
  NAND2_X1 U4642 ( .A1(n12342), .A2(n34533), .ZN(n34429) );
  XNOR2_X1 U4643 ( .A(n32427), .B(\fmem_data[8][1] ), .ZN(n33748) );
  XNOR2_X1 U4644 ( .A(n32939), .B(\fmem_data[1][3] ), .ZN(n34465) );
  NAND2_X1 U4645 ( .A1(n7594), .A2(n34463), .ZN(n34462) );
  XNOR2_X1 U4646 ( .A(n32936), .B(\fmem_data[19][1] ), .ZN(n34345) );
  OAI22_X1 U4647 ( .A1(n32435), .A2(n33250), .B1(n33249), .B2(n3654), .ZN(
        n32894) );
  OAI22_X1 U4648 ( .A1(n32431), .A2(n33873), .B1(n33875), .B2(n3607), .ZN(
        n32897) );
  NAND2_X1 U4649 ( .A1(n16945), .A2(n33174), .ZN(n33176) );
  XNOR2_X1 U4650 ( .A(n32614), .B(\fmem_data[24][1] ), .ZN(n34772) );
  XNOR2_X1 U4651 ( .A(n34624), .B(\fmem_data[28][3] ), .ZN(n32072) );
  NAND2_X1 U4652 ( .A1(n5668), .A2(n33855), .ZN(n33853) );
  XNOR2_X1 U4653 ( .A(n33573), .B(\fmem_data[28][1] ), .ZN(n34744) );
  INV_X1 U4654 ( .A(n31540), .ZN(n31541) );
  OAI22_X1 U4655 ( .A1(n34615), .A2(n31539), .B1(n34199), .B2(n3684), .ZN(
        n31540) );
  OR2_X1 U4656 ( .A1(n34201), .A2(n3684), .ZN(n31539) );
  XNOR2_X1 U4657 ( .A(n31511), .B(\fmem_data[16][1] ), .ZN(n32599) );
  INV_X1 U4658 ( .A(n36480), .ZN(n33759) );
  NAND2_X1 U4659 ( .A1(n33738), .A2(n33737), .ZN(n33703) );
  OAI22_X1 U4660 ( .A1(n33583), .A2(n33582), .B1(n33581), .B2(n34340), .ZN(
        n33695) );
  XNOR2_X1 U4661 ( .A(n32597), .B(\fmem_data[15][1] ), .ZN(n34402) );
  OAI22_X1 U4662 ( .A1(n33832), .A2(n34208), .B1(n33831), .B2(n34206), .ZN(
        n34508) );
  OAI22_X1 U4663 ( .A1(n34485), .A2(n34613), .B1(n32058), .B2(n3570), .ZN(
        n32966) );
  NAND2_X1 U4664 ( .A1(n4366), .A2(n33850), .ZN(n33851) );
  XOR2_X1 U4665 ( .A(\fmem_data[5][3] ), .B(\fmem_data[5][2] ), .Z(n4366) );
  NAND2_X1 U4666 ( .A1(n4156), .A2(n33596), .ZN(n33598) );
  OAI22_X1 U4667 ( .A1(n34790), .A2(n34788), .B1(n32573), .B2(n3560), .ZN(
        n32992) );
  OAI22_X1 U4668 ( .A1(n33867), .A2(n3558), .B1(n32443), .B2(n36221), .ZN(
        n31562) );
  OAI22_X1 U4669 ( .A1(n33907), .A2(n34470), .B1(n32621), .B2(n34468), .ZN(
        n31561) );
  OAI22_X1 U4670 ( .A1(n33992), .A2(n34505), .B1(n32604), .B2(n34503), .ZN(
        n31607) );
  OAI22_X1 U4671 ( .A1(n31225), .A2(n34923), .B1(n34922), .B2(n3606), .ZN(
        n31609) );
  OAI22_X1 U4672 ( .A1(n34502), .A2(n34499), .B1(n31453), .B2(n34501), .ZN(
        n32974) );
  OAI22_X1 U4673 ( .A1(n31126), .A2(n3564), .B1(n33577), .B2(n36295), .ZN(
        n31459) );
  OAI22_X1 U4674 ( .A1(n31122), .A2(n33741), .B1(n33602), .B2(n33603), .ZN(
        n31461) );
  OAI22_X1 U4675 ( .A1(n31124), .A2(n35088), .B1(n31123), .B2(n35089), .ZN(
        n31460) );
  OAI22_X1 U4676 ( .A1(n31595), .A2(n34435), .B1(n34437), .B2(n3592), .ZN(
        n33445) );
  OAI22_X1 U4677 ( .A1(n31596), .A2(n34414), .B1(n34416), .B2(n3603), .ZN(
        n33444) );
  OAI22_X1 U4678 ( .A1(n33812), .A2(n3559), .B1(n32883), .B2(n34017), .ZN(
        n33443) );
  OAI22_X1 U4679 ( .A1(n31162), .A2(n3567), .B1(n33809), .B2(n34777), .ZN(
        n32084) );
  OAI22_X1 U4680 ( .A1(n33731), .A2(n34363), .B1(n32602), .B2(n34364), .ZN(
        n32872) );
  XNOR2_X1 U4681 ( .A(n32614), .B(\fmem_data[24][3] ), .ZN(n33804) );
  NAND2_X1 U4682 ( .A1(n10363), .A2(n34431), .ZN(n34433) );
  OAI22_X1 U4683 ( .A1(n32443), .A2(n3558), .B1(n33688), .B2(n36221), .ZN(
        n32843) );
  OAI22_X1 U4684 ( .A1(n32536), .A2(n34537), .B1(n32535), .B2(n34535), .ZN(
        n32546) );
  NAND2_X1 U4685 ( .A1(n36139), .A2(n36137), .ZN(n34750) );
  XNOR2_X1 U4686 ( .A(n36177), .B(n36176), .ZN(n36774) );
  XNOR2_X1 U4687 ( .A(n36175), .B(n36174), .ZN(n36177) );
  OAI21_X1 U4688 ( .B1(n32831), .B2(n32829), .A(n32830), .ZN(n32629) );
  NAND2_X1 U4689 ( .A1(n32272), .A2(n32274), .ZN(n32213) );
  OAI22_X1 U4690 ( .A1(n31122), .A2(n33603), .B1(n26271), .B2(n33741), .ZN(
        n28895) );
  OAI22_X1 U4691 ( .A1(n31162), .A2(n34777), .B1(n33947), .B2(n3567), .ZN(
        n28897) );
  INV_X1 U4692 ( .A(n23175), .ZN(n20288) );
  OAI22_X1 U4693 ( .A1(n31443), .A2(n33057), .B1(n29209), .B2(n33059), .ZN(
        n28536) );
  OAI22_X1 U4694 ( .A1(n31445), .A2(n35010), .B1(n34099), .B2(n35011), .ZN(
        n28535) );
  OAI22_X1 U4695 ( .A1(n32177), .A2(n34466), .B1(n33189), .B2(n34779), .ZN(
        n28942) );
  NAND2_X1 U4696 ( .A1(n7193), .A2(n34412), .ZN(n34410) );
  NAND2_X1 U4697 ( .A1(n10943), .A2(n34420), .ZN(n34418) );
  NAND2_X1 U4698 ( .A1(n4772), .A2(n35512), .ZN(n35511) );
  OAI22_X1 U4699 ( .A1(n29518), .A2(n35722), .B1(n35721), .B2(n3624), .ZN(
        n29687) );
  NAND2_X1 U4700 ( .A1(n11585), .A2(n35619), .ZN(n35618) );
  OAI22_X1 U4701 ( .A1(n31990), .A2(n3573), .B1(n32167), .B2(n36298), .ZN(
        n29530) );
  OAI22_X1 U4702 ( .A1(n26252), .A2(n33873), .B1(n33874), .B2(n33875), .ZN(
        n29532) );
  OAI22_X1 U4703 ( .A1(n30795), .A2(n35739), .B1(n30794), .B2(n35740), .ZN(
        n31891) );
  XNOR2_X1 U4704 ( .A(n36228), .B(\fmem_data[20][7] ), .ZN(n30794) );
  OAI22_X1 U4705 ( .A1(n32107), .A2(n34836), .B1(n34232), .B2(n34835), .ZN(
        n30803) );
  XNOR2_X1 U4706 ( .A(n31484), .B(n31483), .ZN(n33630) );
  XNOR2_X1 U4707 ( .A(n31482), .B(n31481), .ZN(n31484) );
  NAND2_X1 U4708 ( .A1(n34520), .A2(n34519), .ZN(n34442) );
  XNOR2_X1 U4709 ( .A(n33543), .B(n33542), .ZN(n36490) );
  XNOR2_X1 U4710 ( .A(n33541), .B(n33540), .ZN(n33543) );
  NAND2_X1 U4711 ( .A1(n33911), .A2(n33910), .ZN(n33912) );
  OAI22_X1 U4712 ( .A1(n32518), .A2(n34497), .B1(n32517), .B2(n34495), .ZN(
        n33171) );
  OAI22_X1 U4713 ( .A1(n34046), .A2(n34045), .B1(n34044), .B2(n34043), .ZN(
        n34205) );
  OAI22_X1 U4714 ( .A1(n32726), .A2(n35611), .B1(n35610), .B2(n3631), .ZN(
        n32759) );
  NAND2_X1 U4715 ( .A1(n34458), .A2(n34459), .ZN(n34444) );
  NAND2_X1 U4716 ( .A1(n32674), .A2(n32673), .ZN(n32814) );
  XNOR2_X1 U4717 ( .A(n34817), .B(n34816), .ZN(n35469) );
  NAND2_X1 U4718 ( .A1(n33396), .A2(n33395), .ZN(n34956) );
  NAND2_X1 U4719 ( .A1(n33394), .A2(n33393), .ZN(n33395) );
  OAI21_X1 U4720 ( .B1(n33394), .B2(n33393), .A(n33392), .ZN(n33396) );
  OAI21_X1 U4721 ( .B1(n35375), .B2(n35374), .A(n35373), .ZN(n35377) );
  NAND2_X1 U4722 ( .A1(n35375), .A2(n35374), .ZN(n35376) );
  OAI21_X1 U4723 ( .B1(n34829), .B2(n34828), .A(n34827), .ZN(n35371) );
  INV_X1 U4724 ( .A(n34824), .ZN(n34829) );
  NAND2_X1 U4725 ( .A1(n34826), .A2(n34825), .ZN(n34827) );
  OAI21_X1 U4726 ( .B1(n35366), .B2(n35365), .A(n35364), .ZN(n35764) );
  INV_X1 U4727 ( .A(n35361), .ZN(n35366) );
  NAND2_X1 U4728 ( .A1(n35363), .A2(n35362), .ZN(n35364) );
  OAI22_X1 U4729 ( .A1(n35031), .A2(n35696), .B1(n35317), .B2(n35697), .ZN(
        n35265) );
  XNOR2_X1 U4730 ( .A(n35043), .B(n35284), .ZN(n35264) );
  XNOR2_X1 U4731 ( .A(n35282), .B(n35283), .ZN(n35043) );
  NAND2_X1 U4732 ( .A1(n35567), .A2(n35566), .ZN(n35571) );
  OR2_X1 U4733 ( .A1(n35569), .A2(n35568), .ZN(n35566) );
  NAND2_X1 U4734 ( .A1(n35569), .A2(n35568), .ZN(n35570) );
  OAI21_X1 U4735 ( .B1(n35563), .B2(n35562), .A(n35561), .ZN(n35565) );
  XNOR2_X1 U4736 ( .A(n35270), .B(\fmem_data[19][7] ), .ZN(n35654) );
  NAND2_X1 U4737 ( .A1(n15696), .A2(n35656), .ZN(n35655) );
  OAI22_X1 U4738 ( .A1(n35506), .A2(n35508), .B1(n35404), .B2(n35507), .ZN(
        n35659) );
  OAI22_X1 U4739 ( .A1(n35402), .A2(n35493), .B1(n35492), .B2(n35494), .ZN(
        n35660) );
  AOI21_X1 U4740 ( .B1(n35652), .B2(n35651), .A(n35650), .ZN(n35653) );
  OAI22_X1 U4741 ( .A1(n35488), .A2(n35490), .B1(n35396), .B2(n35489), .ZN(
        n35667) );
  OAI22_X1 U4742 ( .A1(n35751), .A2(n35753), .B1(n35398), .B2(n35752), .ZN(
        n35666) );
  NAND2_X1 U4743 ( .A1(n8833), .A2(n35663), .ZN(n35662) );
  NAND2_X1 U4744 ( .A1(n9114), .A2(n35712), .ZN(n35711) );
  AOI21_X1 U4745 ( .B1(n35512), .B2(n35511), .A(n35510), .ZN(n35513) );
  AOI21_X1 U4746 ( .B1(n35508), .B2(n35507), .A(n35506), .ZN(n35509) );
  AOI21_X1 U4747 ( .B1(n35516), .B2(n35515), .A(n35514), .ZN(n35517) );
  NAND2_X1 U4748 ( .A1(n17463), .A2(n35592), .ZN(n35591) );
  OAI22_X1 U4749 ( .A1(n35743), .A2(n35745), .B1(n35327), .B2(n35744), .ZN(
        n35595) );
  OAI22_X1 U4750 ( .A1(n35329), .A2(n35729), .B1(n35728), .B2(n35730), .ZN(
        n35594) );
  OAI22_X1 U4751 ( .A1(n35747), .A2(n35749), .B1(n35325), .B2(n35748), .ZN(
        n35596) );
  OAI22_X1 U4752 ( .A1(n35724), .A2(n35726), .B1(n35339), .B2(n35725), .ZN(
        n35588) );
  OAI22_X1 U4753 ( .A1(n35738), .A2(n35739), .B1(n35341), .B2(n35740), .ZN(
        n35587) );
  OAI22_X1 U4754 ( .A1(n35720), .A2(n35722), .B1(n35337), .B2(n35721), .ZN(
        n35589) );
  AOI21_X1 U4755 ( .B1(n35494), .B2(n35493), .A(n35492), .ZN(n35495) );
  AOI21_X1 U4756 ( .B1(n35490), .B2(n35489), .A(n35488), .ZN(n35491) );
  AOI21_X1 U4757 ( .B1(n35498), .B2(n35497), .A(n35496), .ZN(n35499) );
  OR2_X1 U4758 ( .A1(n17680), .A2(n17679), .ZN(n17681) );
  BUF_X2 U4759 ( .A(n14928), .Z(n28007) );
  AND2_X1 U4760 ( .A1(n28207), .A2(\xmem_data[62][0] ), .ZN(n28708) );
  NAND2_X1 U4761 ( .A1(n28683), .A2(n28682), .ZN(n28695) );
  NOR2_X1 U4762 ( .A1(n27824), .A2(n27823), .ZN(n27829) );
  NAND3_X1 U4763 ( .A1(n27822), .A2(n27821), .A3(n27820), .ZN(n27823) );
  BUF_X2 U4764 ( .A(n10861), .Z(n30100) );
  NAND2_X1 U4765 ( .A1(n27212), .A2(n27211), .ZN(n32940) );
  NAND2_X1 U4766 ( .A1(n23288), .A2(n23287), .ZN(n33683) );
  NAND3_X1 U4767 ( .A1(n30333), .A2(n30332), .A3(n30331), .ZN(n33479) );
  NAND2_X1 U4768 ( .A1(n21090), .A2(n21089), .ZN(n33754) );
  OR2_X1 U4769 ( .A1(n36112), .A2(n3673), .ZN(n34629) );
  XNOR2_X1 U4770 ( .A(n33677), .B(\fmem_data[30][1] ), .ZN(n34596) );
  NAND2_X1 U4771 ( .A1(\fmem_data[30][1] ), .A2(n3560), .ZN(n34788) );
  NAND2_X1 U4772 ( .A1(\fmem_data[14][1] ), .A2(n3563), .ZN(n34739) );
  OR3_X1 U4773 ( .A1(n20605), .A2(n20604), .A3(n20603), .ZN(n20607) );
  NAND2_X1 U4774 ( .A1(n22769), .A2(n22768), .ZN(n22770) );
  NAND2_X1 U4775 ( .A1(\fmem_data[9][1] ), .A2(n3579), .ZN(n34476) );
  XNOR2_X1 U4776 ( .A(n32882), .B(\fmem_data[6][1] ), .ZN(n33757) );
  NAND2_X1 U4777 ( .A1(\fmem_data[28][1] ), .A2(n3562), .ZN(n34745) );
  NAND2_X1 U4778 ( .A1(n36534), .A2(n36533), .ZN(n33752) );
  OAI22_X1 U4779 ( .A1(n36297), .A2(n36295), .B1(n33755), .B2(n3564), .ZN(
        n36478) );
  XNOR2_X1 U4780 ( .A(n32898), .B(\fmem_data[8][1] ), .ZN(n34627) );
  OAI22_X1 U4781 ( .A1(n34486), .A2(n34613), .B1(n34485), .B2(n3570), .ZN(
        n34585) );
  OAI22_X1 U4782 ( .A1(n34478), .A2(n3579), .B1(n34477), .B2(n34476), .ZN(
        n34578) );
  OAI22_X1 U4783 ( .A1(n34502), .A2(n34501), .B1(n34500), .B2(n34499), .ZN(
        n34583) );
  OAI22_X1 U4784 ( .A1(n34506), .A2(n34505), .B1(n34504), .B2(n34503), .ZN(
        n34582) );
  OAI22_X1 U4785 ( .A1(n34596), .A2(n34788), .B1(n34789), .B2(n3560), .ZN(
        n36350) );
  OAI22_X1 U4786 ( .A1(n31526), .A2(n34340), .B1(n33582), .B2(n3616), .ZN(
        n33498) );
  OAI22_X1 U4787 ( .A1(n33781), .A2(n3572), .B1(n34733), .B2(n34734), .ZN(
        n33496) );
  OR2_X1 U4788 ( .A1(n36112), .A2(n3616), .ZN(n31526) );
  OAI22_X1 U4789 ( .A1(n33810), .A2(n3567), .B1(n34776), .B2(n34777), .ZN(
        n33499) );
  XNOR2_X1 U4790 ( .A(n33473), .B(n33472), .ZN(n36354) );
  XNOR2_X1 U4791 ( .A(n33471), .B(n33470), .ZN(n33472) );
  NAND2_X1 U4792 ( .A1(n36507), .A2(n36509), .ZN(n33729) );
  XNOR2_X1 U4793 ( .A(n36490), .B(n36489), .ZN(n36491) );
  NAND2_X1 U4794 ( .A1(n36504), .A2(n36503), .ZN(n33770) );
  NAND2_X1 U4795 ( .A1(n33561), .A2(n33560), .ZN(n36467) );
  NAND2_X1 U4796 ( .A1(n36484), .A2(n36482), .ZN(n33560) );
  OAI21_X1 U4797 ( .B1(n36484), .B2(n36482), .A(n36483), .ZN(n33561) );
  XNOR2_X1 U4798 ( .A(n32993), .B(n32992), .ZN(n32994) );
  NAND2_X1 U4799 ( .A1(n34753), .A2(n34752), .ZN(n32697) );
  XNOR2_X1 U4800 ( .A(n32826), .B(n32825), .ZN(n32828) );
  XNOR2_X1 U4801 ( .A(n26801), .B(n3586), .ZN(n34153) );
  XNOR2_X1 U4802 ( .A(n26800), .B(n26799), .ZN(n26801) );
  INV_X1 U4803 ( .A(n26798), .ZN(n26800) );
  OAI22_X1 U4804 ( .A1(n24335), .A2(n35516), .B1(n33182), .B2(n35515), .ZN(
        n29537) );
  OAI22_X1 U4805 ( .A1(n33052), .A2(n33568), .B1(n31964), .B2(n33570), .ZN(
        n29538) );
  NAND2_X1 U4806 ( .A1(n32088), .A2(n32089), .ZN(n31920) );
  NAND2_X1 U4807 ( .A1(n36419), .A2(n36420), .ZN(n33607) );
  XNOR2_X1 U4808 ( .A(n34449), .B(n34448), .ZN(n36049) );
  NAND2_X1 U4809 ( .A1(n35625), .A2(n35624), .ZN(n35787) );
  NAND2_X1 U4810 ( .A1(n35623), .A2(n35622), .ZN(n35624) );
  OAI21_X1 U4811 ( .B1(n35623), .B2(n35622), .A(n35621), .ZN(n35625) );
  AOI21_X1 U4812 ( .B1(n35701), .B2(n35700), .A(n35699), .ZN(n35702) );
  NAND2_X1 U4813 ( .A1(n21673), .A2(n35709), .ZN(n35708) );
  XNOR2_X1 U4814 ( .A(n35076), .B(\fmem_data[30][7] ), .ZN(n35707) );
  NAND2_X1 U4815 ( .A1(n24435), .A2(n35705), .ZN(n35704) );
  AOI21_X1 U4816 ( .B1(n35712), .B2(n35711), .A(n35710), .ZN(n35713) );
  OAI21_X1 U4817 ( .B1(n17040), .B2(n17039), .A(n17038), .ZN(n17076) );
  OR3_X1 U4818 ( .A1(n27422), .A2(n27421), .A3(n27420), .ZN(n27428) );
  NAND4_X2 U4819 ( .A1(n19023), .A2(n19022), .A3(n19021), .A4(n19020), .ZN(
        n34612) );
  OAI21_X1 U4820 ( .B1(n28290), .B2(n28289), .A(n28288), .ZN(n28400) );
  XNOR2_X1 U4821 ( .A(n32940), .B(\fmem_data[18][1] ), .ZN(n36106) );
  NAND2_X1 U4822 ( .A1(\fmem_data[18][1] ), .A2(n3580), .ZN(n36104) );
  NAND2_X1 U4823 ( .A1(\fmem_data[23][1] ), .A2(n3662), .ZN(n36241) );
  NAND2_X1 U4824 ( .A1(\fmem_data[19][1] ), .A2(n3633), .ZN(n36226) );
  OR2_X1 U4825 ( .A1(n33454), .A2(n3945), .ZN(n33458) );
  NAND2_X1 U4826 ( .A1(\fmem_data[7][1] ), .A2(n3581), .ZN(n36218) );
  NAND2_X1 U4827 ( .A1(\fmem_data[15][1] ), .A2(n3568), .ZN(n36223) );
  NAND2_X1 U4828 ( .A1(\fmem_data[31][1] ), .A2(n3931), .ZN(n36216) );
  XNOR2_X1 U4829 ( .A(n32939), .B(\fmem_data[1][1] ), .ZN(n36209) );
  NAND2_X1 U4830 ( .A1(\fmem_data[27][1] ), .A2(n3482), .ZN(n36240) );
  NAND2_X1 U4831 ( .A1(\fmem_data[1][1] ), .A2(n3558), .ZN(n36221) );
  XNOR2_X1 U4832 ( .A(n33754), .B(\fmem_data[0][1] ), .ZN(n36297) );
  XNOR2_X1 U4833 ( .A(n33556), .B(\fmem_data[16][1] ), .ZN(n36300) );
  NAND2_X1 U4834 ( .A1(\fmem_data[16][1] ), .A2(n3573), .ZN(n36298) );
  NAND2_X1 U4835 ( .A1(\fmem_data[0][1] ), .A2(n3564), .ZN(n36295) );
  INV_X1 U4836 ( .A(n34616), .ZN(n34617) );
  NAND2_X1 U4837 ( .A1(\fmem_data[8][1] ), .A2(n3574), .ZN(n34625) );
  NAND2_X1 U4838 ( .A1(\fmem_data[20][1] ), .A2(n3647), .ZN(n36227) );
  NAND2_X1 U4839 ( .A1(\fmem_data[26][1] ), .A2(n3678), .ZN(n33725) );
  NAND2_X1 U4840 ( .A1(\fmem_data[13][1] ), .A2(n3571), .ZN(n34742) );
  NAND2_X1 U4841 ( .A1(\fmem_data[17][1] ), .A2(n3566), .ZN(n34529) );
  NAND2_X1 U4842 ( .A1(\fmem_data[24][1] ), .A2(n3565), .ZN(n36100) );
  NAND2_X1 U4843 ( .A1(\fmem_data[5][1] ), .A2(n3576), .ZN(n34483) );
  XNOR2_X1 U4844 ( .A(n36510), .B(n36509), .ZN(n36903) );
  XNOR2_X1 U4845 ( .A(n36506), .B(n36505), .ZN(n36904) );
  XNOR2_X1 U4846 ( .A(n36508), .B(n36507), .ZN(n36510) );
  XNOR2_X1 U4847 ( .A(n36291), .B(n36290), .ZN(n36704) );
  XNOR2_X1 U4848 ( .A(n36189), .B(n36188), .ZN(n36809) );
  NAND2_X1 U4849 ( .A1(n36388), .A2(n36389), .ZN(n33521) );
  XNOR2_X1 U4850 ( .A(n36049), .B(n36048), .ZN(n36051) );
  NAND2_X1 U4851 ( .A1(n3431), .A2(n35778), .ZN(n35780) );
  BUF_X1 U4852 ( .A(n35779), .Z(n3431) );
  XNOR2_X1 U4853 ( .A(n35909), .B(n35910), .ZN(n35539) );
  AOI21_X1 U4854 ( .B1(n35709), .B2(n35708), .A(n35707), .ZN(n35869) );
  NAND4_X1 U4855 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n3353) );
  OAI21_X1 U4856 ( .B1(n3722), .B2(n17154), .A(n21088), .ZN(n17177) );
  AOI22_X1 U4857 ( .A1(n21628), .A2(n25396), .B1(n21627), .B2(n16443), .ZN(
        n21672) );
  NAND2_X1 U4858 ( .A1(n17527), .A2(n24508), .ZN(n17553) );
  OAI21_X1 U4859 ( .B1(n17551), .B2(n17550), .A(n22180), .ZN(n17552) );
  NAND2_X1 U4860 ( .A1(n21579), .A2(n27968), .ZN(n21580) );
  OAI21_X1 U4861 ( .B1(n21558), .B2(n21557), .A(n9896), .ZN(n21581) );
  NAND2_X1 U4862 ( .A1(n28459), .A2(n28458), .ZN(n28530) );
  NAND2_X1 U4863 ( .A1(n28491), .A2(n28490), .ZN(n28529) );
  NAND2_X1 U4864 ( .A1(n21737), .A2(n28107), .ZN(n21764) );
  OAI21_X1 U4865 ( .B1(n27639), .B2(n27638), .A(n29598), .ZN(n27696) );
  OAI21_X1 U4866 ( .B1(n27693), .B2(n27692), .A(n29600), .ZN(n27694) );
  OAI21_X1 U4867 ( .B1(n28217), .B2(n28216), .A(n28215), .ZN(n28262) );
  OAI21_X1 U4868 ( .B1(n28135), .B2(n28134), .A(n28133), .ZN(n28264) );
  AND2_X1 U4869 ( .A1(n36101), .A2(\fmem_data[24][0] ), .ZN(n36525) );
  AOI22_X1 U4870 ( .A1(n30010), .A2(n30009), .B1(n30008), .B2(n30007), .ZN(
        n30011) );
  OR2_X1 U4871 ( .A1(n36312), .A2(n3681), .ZN(n36113) );
  OR2_X1 U4872 ( .A1(n36315), .A2(n3695), .ZN(n36198) );
  XNOR2_X1 U4873 ( .A(n36948), .B(n36947), .ZN(n37000) );
  XNOR2_X1 U4874 ( .A(n36743), .B(n36742), .ZN(n36933) );
  NAND2_X1 U4875 ( .A1(n36938), .A2(n36941), .ZN(n36738) );
  INV_X1 U4876 ( .A(n37128), .ZN(n36650) );
  CLKBUF_X1 U4877 ( .A(n36448), .Z(n36449) );
  INV_X1 U4878 ( .A(n35962), .ZN(n35952) );
  XNOR2_X1 U4879 ( .A(n36730), .B(n36729), .ZN(n37011) );
  NAND2_X1 U4880 ( .A1(n37110), .A2(n37109), .ZN(n37111) );
  NAND2_X1 U4881 ( .A1(n37108), .A2(n37107), .ZN(n37109) );
  OAI21_X1 U4882 ( .B1(n37108), .B2(n37107), .A(n37106), .ZN(n37110) );
  INV_X1 U4883 ( .A(n36008), .ZN(n37166) );
  AOI22_X1 U4884 ( .A1(n36007), .A2(n36006), .B1(n36005), .B2(n36004), .ZN(
        n36008) );
  NAND2_X1 U4885 ( .A1(n36003), .A2(n36002), .ZN(n36006) );
  INV_X1 U4886 ( .A(n37182), .ZN(n37178) );
  NOR2_X1 U4887 ( .A1(n37079), .A2(n37078), .ZN(n37303) );
  NAND2_X1 U4888 ( .A1(n37079), .A2(n37078), .ZN(n37304) );
  AND2_X1 U4889 ( .A1(n37099), .A2(n37098), .ZN(n37285) );
  OR2_X1 U4890 ( .A1(n37112), .A2(n37111), .ZN(n37276) );
  XNOR2_X1 U4891 ( .A(n36662), .B(n36661), .ZN(n37127) );
  INV_X1 U4892 ( .A(n37187), .ZN(n37252) );
  INV_X1 U4893 ( .A(n37208), .ZN(n37209) );
  INV_X1 U4894 ( .A(n37202), .ZN(n37243) );
  NOR2_X1 U4895 ( .A1(n37181), .A2(n37180), .ZN(n37202) );
  NOR2_X1 U4896 ( .A1(n37183), .A2(n37182), .ZN(n37246) );
  NAND2_X1 U4897 ( .A1(n37183), .A2(n37182), .ZN(n37247) );
  OR2_X1 U4898 ( .A1(n37244), .A2(n37164), .ZN(n37204) );
  NAND2_X1 U4899 ( .A1(n10440), .A2(n10439), .ZN(n10441) );
  AND2_X1 U4900 ( .A1(n19736), .A2(n19735), .ZN(n19739) );
  INV_X1 U4901 ( .A(n13372), .ZN(n13373) );
  NOR4_X1 U4902 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10445) );
  INV_X1 U4903 ( .A(n10436), .ZN(n10443) );
  INV_X1 U4904 ( .A(n10435), .ZN(n10444) );
  NAND2_X1 U4905 ( .A1(n10438), .A2(n10437), .ZN(n10442) );
  AND2_X1 U4906 ( .A1(n31255), .A2(\xmem_data[55][5] ), .ZN(n18464) );
  INV_X1 U4907 ( .A(n7994), .ZN(n7995) );
  INV_X1 U4908 ( .A(n7992), .ZN(n7996) );
  NAND3_X1 U4909 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10206) );
  NAND3_X1 U4910 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(n9497) );
  NAND3_X1 U4911 ( .A1(n16637), .A2(n16636), .A3(n16635), .ZN(n16638) );
  NAND2_X1 U4912 ( .A1(n10977), .A2(\xmem_data[22][7] ), .ZN(n10264) );
  NAND2_X1 U4913 ( .A1(n24597), .A2(\xmem_data[23][7] ), .ZN(n10265) );
  NAND3_X1 U4914 ( .A1(n14487), .A2(n14486), .A3(n14485), .ZN(n14491) );
  INV_X1 U4915 ( .A(n14100), .ZN(n14107) );
  NAND3_X1 U4916 ( .A1(n7887), .A2(n7886), .A3(n7885), .ZN(n7888) );
  NAND3_X1 U4917 ( .A1(n7917), .A2(n7916), .A3(n7915), .ZN(n7918) );
  NOR2_X1 U4918 ( .A1(n24789), .A2(n24788), .ZN(n24790) );
  INV_X1 U4919 ( .A(n24787), .ZN(n24788) );
  INV_X1 U4920 ( .A(n24786), .ZN(n24789) );
  NOR2_X1 U4921 ( .A1(n24743), .A2(n24742), .ZN(n24744) );
  INV_X1 U4922 ( .A(n24741), .ZN(n24742) );
  INV_X1 U4923 ( .A(n24740), .ZN(n24743) );
  INV_X1 U4924 ( .A(n3268), .ZN(n3307) );
  AOI22_X1 U4925 ( .A1(n30261), .A2(\xmem_data[126][2] ), .B1(n3434), .B2(
        \xmem_data[127][2] ), .ZN(n18195) );
  AND2_X1 U4926 ( .A1(n18176), .A2(n18175), .ZN(n18178) );
  NAND3_X1 U4927 ( .A1(n3726), .A2(n13443), .A3(n13442), .ZN(n13448) );
  NAND2_X1 U4928 ( .A1(n24443), .A2(\xmem_data[2][3] ), .ZN(n13451) );
  NAND3_X1 U4929 ( .A1(n15139), .A2(n15138), .A3(n15137), .ZN(n15140) );
  NAND3_X1 U4930 ( .A1(n16472), .A2(n16471), .A3(n16470), .ZN(n16475) );
  INV_X1 U4931 ( .A(n16473), .ZN(n16474) );
  NAND3_X1 U4932 ( .A1(n14834), .A2(n14833), .A3(n14832), .ZN(n14835) );
  NAND3_X1 U4933 ( .A1(n19789), .A2(n19788), .A3(n19787), .ZN(n19790) );
  AND2_X1 U4934 ( .A1(n19730), .A2(n19729), .ZN(n19753) );
  NAND3_X1 U4935 ( .A1(n5166), .A2(n5168), .A3(n5167), .ZN(n5179) );
  AOI21_X1 U4936 ( .B1(n30503), .B2(\xmem_data[76][6] ), .A(n8943), .ZN(n8948)
         );
  NAND3_X1 U4937 ( .A1(n8957), .A2(n8956), .A3(n8955), .ZN(n8963) );
  AOI22_X1 U4938 ( .A1(n28516), .A2(\xmem_data[58][6] ), .B1(n30542), .B2(
        \xmem_data[59][6] ), .ZN(n8967) );
  NOR2_X1 U4939 ( .A1(n25627), .A2(n25626), .ZN(n25645) );
  INV_X1 U4940 ( .A(n25625), .ZN(n25626) );
  INV_X1 U4941 ( .A(n25623), .ZN(n25627) );
  NOR2_X1 U4942 ( .A1(n15847), .A2(n15846), .ZN(n15848) );
  NOR2_X1 U4943 ( .A1(n9412), .A2(n9411), .ZN(n9413) );
  INV_X1 U4944 ( .A(n9410), .ZN(n9411) );
  NAND2_X1 U4945 ( .A1(n25486), .A2(\xmem_data[8][3] ), .ZN(n4936) );
  NAND2_X1 U4946 ( .A1(n25481), .A2(\xmem_data[12][3] ), .ZN(n4937) );
  NAND3_X1 U4947 ( .A1(n25010), .A2(n25009), .A3(n25008), .ZN(n25011) );
  NAND3_X1 U4948 ( .A1(n25031), .A2(n25030), .A3(n25029), .ZN(n25032) );
  INV_X1 U4949 ( .A(n21415), .ZN(n21416) );
  AOI22_X1 U4950 ( .A1(n27761), .A2(\xmem_data[37][6] ), .B1(n30743), .B2(
        \xmem_data[36][6] ), .ZN(n12240) );
  NAND3_X1 U4951 ( .A1(n12318), .A2(n12317), .A3(n12316), .ZN(n12319) );
  AND2_X1 U4952 ( .A1(n27741), .A2(\xmem_data[28][6] ), .ZN(n12331) );
  NAND3_X1 U4953 ( .A1(n12258), .A2(n12257), .A3(n12256), .ZN(n12269) );
  INV_X1 U4954 ( .A(n11198), .ZN(n11204) );
  NOR2_X1 U4955 ( .A1(n11193), .A2(n11192), .ZN(n11196) );
  INV_X1 U4956 ( .A(n11191), .ZN(n11192) );
  NAND3_X1 U4957 ( .A1(n13727), .A2(n13726), .A3(n13725), .ZN(n13728) );
  NAND3_X1 U4958 ( .A1(n5462), .A2(n5461), .A3(n5460), .ZN(n5463) );
  NAND3_X1 U4959 ( .A1(n5530), .A2(n5529), .A3(n5528), .ZN(n5531) );
  AND2_X1 U4960 ( .A1(n27563), .A2(\xmem_data[19][5] ), .ZN(n13000) );
  INV_X1 U4961 ( .A(n12981), .ZN(n12987) );
  NAND3_X1 U4962 ( .A1(n7536), .A2(n7535), .A3(n7534), .ZN(n7537) );
  NAND3_X1 U4963 ( .A1(n5069), .A2(n5068), .A3(n5067), .ZN(n5070) );
  NAND2_X1 U4964 ( .A1(n30294), .A2(\xmem_data[40][5] ), .ZN(n18473) );
  NAND2_X1 U4965 ( .A1(n29589), .A2(\xmem_data[45][5] ), .ZN(n18475) );
  INV_X1 U4966 ( .A(n16816), .ZN(n16817) );
  OR3_X1 U4967 ( .A1(n20764), .A2(n20763), .A3(n20762), .ZN(n20766) );
  OR3_X1 U4968 ( .A1(n20825), .A2(n20824), .A3(n20823), .ZN(n20835) );
  OR3_X1 U4969 ( .A1(n20741), .A2(n20740), .A3(n20739), .ZN(n20743) );
  NAND3_X1 U4970 ( .A1(n19919), .A2(n19918), .A3(n19917), .ZN(n19936) );
  NAND3_X1 U4971 ( .A1(n19934), .A2(n19933), .A3(n19932), .ZN(n19935) );
  AND2_X1 U4972 ( .A1(n19931), .A2(n19930), .ZN(n19932) );
  NAND3_X1 U4973 ( .A1(n14759), .A2(n14758), .A3(n14757), .ZN(n14760) );
  NOR2_X1 U4974 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  INV_X1 U4975 ( .A(n12129), .ZN(n12132) );
  INV_X1 U4976 ( .A(n12130), .ZN(n12131) );
  NAND3_X1 U4977 ( .A1(n12181), .A2(n12180), .A3(n12179), .ZN(n12187) );
  OR3_X1 U4978 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(n10016) );
  NAND3_X1 U4979 ( .A1(n11254), .A2(n11253), .A3(n11252), .ZN(n11258) );
  NOR2_X1 U4980 ( .A1(n31021), .A2(n31020), .ZN(n31025) );
  INV_X1 U4981 ( .A(n31019), .ZN(n31020) );
  INV_X1 U4982 ( .A(n3385), .ZN(n3317) );
  AND2_X1 U4983 ( .A1(n27871), .A2(n27870), .ZN(n27872) );
  INV_X1 U4984 ( .A(n22854), .ZN(n22855) );
  AND2_X1 U4985 ( .A1(n23813), .A2(\xmem_data[30][1] ), .ZN(n22856) );
  INV_X1 U4986 ( .A(n19567), .ZN(n19573) );
  NAND3_X1 U4987 ( .A1(n20352), .A2(n20351), .A3(n20350), .ZN(n20355) );
  NAND3_X1 U4988 ( .A1(n20328), .A2(n20327), .A3(n20326), .ZN(n20331) );
  NOR2_X1 U4989 ( .A1(n24797), .A2(n24796), .ZN(n24798) );
  NAND3_X1 U4990 ( .A1(n24767), .A2(n24766), .A3(n24765), .ZN(n24768) );
  AND2_X1 U4991 ( .A1(n20568), .A2(\xmem_data[102][2] ), .ZN(n19858) );
  NOR2_X1 U4992 ( .A1(n29036), .A2(n29035), .ZN(n29037) );
  OR2_X1 U4993 ( .A1(n29034), .A2(n29033), .ZN(n29035) );
  NAND2_X1 U4994 ( .A1(n28990), .A2(n28989), .ZN(n28991) );
  NOR2_X1 U4995 ( .A1(n29073), .A2(n29072), .ZN(n29074) );
  OR2_X1 U4996 ( .A1(n29071), .A2(n29070), .ZN(n29072) );
  AND2_X1 U4997 ( .A1(n29390), .A2(\xmem_data[52][2] ), .ZN(n11940) );
  NAND3_X1 U4998 ( .A1(n26505), .A2(n26504), .A3(n26503), .ZN(n26506) );
  OR2_X1 U4999 ( .A1(n26199), .A2(n26198), .ZN(n26202) );
  NAND3_X1 U5000 ( .A1(n26197), .A2(n26196), .A3(n26195), .ZN(n26199) );
  AND3_X1 U5001 ( .A1(n15678), .A2(n15677), .A3(n15676), .ZN(n15679) );
  NAND3_X1 U5002 ( .A1(n15599), .A2(n15598), .A3(n15597), .ZN(n15602) );
  NAND3_X1 U5003 ( .A1(n15659), .A2(n15658), .A3(n15657), .ZN(n15660) );
  NAND2_X1 U5004 ( .A1(n23522), .A2(n23521), .ZN(n23523) );
  NOR2_X1 U5005 ( .A1(n23520), .A2(n23519), .ZN(n23521) );
  NAND3_X1 U5006 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(n8770) );
  NAND3_X1 U5007 ( .A1(n8793), .A2(n8792), .A3(n8791), .ZN(n8794) );
  INV_X1 U5008 ( .A(n20095), .ZN(n20101) );
  NOR2_X1 U5009 ( .A1(n24038), .A2(n24037), .ZN(n24039) );
  INV_X1 U5010 ( .A(n24036), .ZN(n24037) );
  INV_X1 U5011 ( .A(n18157), .ZN(n18162) );
  AND2_X1 U5012 ( .A1(n30318), .A2(\xmem_data[60][4] ), .ZN(n6338) );
  INV_X1 U5013 ( .A(n15116), .ZN(n15122) );
  OR2_X1 U5014 ( .A1(n4496), .A2(n4495), .ZN(n4502) );
  OR2_X1 U5015 ( .A1(n4494), .A2(n3966), .ZN(n4495) );
  OR2_X1 U5016 ( .A1(n18712), .A2(n18711), .ZN(n18713) );
  NOR2_X1 U5017 ( .A1(n30424), .A2(\fmem_data[13][0] ), .ZN(n30425) );
  INV_X1 U5018 ( .A(n34742), .ZN(n30424) );
  OR3_X1 U5019 ( .A1(n14329), .A2(n14328), .A3(n14327), .ZN(n14330) );
  OR3_X1 U5020 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n14351) );
  OAI21_X1 U5021 ( .B1(n14378), .B2(n14377), .A(n31284), .ZN(n14379) );
  NAND4_X1 U5022 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14378) );
  NOR2_X1 U5023 ( .A1(n18599), .A2(n18598), .ZN(n18600) );
  OR2_X1 U5024 ( .A1(n18597), .A2(n18596), .ZN(n18598) );
  AND2_X1 U5025 ( .A1(n3231), .A2(\xmem_data[3][4] ), .ZN(n15300) );
  NAND3_X1 U5026 ( .A1(n5619), .A2(n5618), .A3(n5617), .ZN(n5620) );
  NAND3_X1 U5027 ( .A1(n3712), .A2(n5626), .A3(n5625), .ZN(n5638) );
  AOI21_X1 U5028 ( .B1(n22181), .B2(n22180), .A(n3881), .ZN(n22251) );
  AOI22_X1 U5029 ( .A1(n28138), .A2(\xmem_data[86][6] ), .B1(n29431), .B2(
        \xmem_data[87][6] ), .ZN(n10866) );
  NAND3_X1 U5030 ( .A1(n25854), .A2(n25853), .A3(n25852), .ZN(n25855) );
  OAI21_X1 U5031 ( .B1(n5932), .B2(n5931), .A(n31342), .ZN(n5956) );
  OR3_X1 U5032 ( .A1(n5930), .A2(n5929), .A3(n5928), .ZN(n5931) );
  OAI21_X1 U5033 ( .B1(n5911), .B2(n5910), .A(n31376), .ZN(n5957) );
  OR4_X1 U5034 ( .A1(n9857), .A2(n9856), .A3(n3504), .A4(n3947), .ZN(n9870) );
  OR2_X1 U5035 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  OR4_X1 U5036 ( .A1(n9815), .A2(n9814), .A3(n9813), .A4(n9812), .ZN(n9816) );
  OR4_X1 U5037 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(n9795) );
  NAND4_X1 U5038 ( .A1(n16320), .A2(n16319), .A3(n3703), .A4(n16318), .ZN(
        n16321) );
  NAND3_X1 U5039 ( .A1(n16271), .A2(n16270), .A3(n16269), .ZN(n16272) );
  OR2_X1 U5040 ( .A1(n16331), .A2(n16330), .ZN(n16347) );
  AND2_X1 U5041 ( .A1(n8998), .A2(n8997), .ZN(n9020) );
  OR4_X1 U5042 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10163) );
  NAND2_X1 U5043 ( .A1(n10153), .A2(n3950), .ZN(n10158) );
  AND4_X1 U5044 ( .A1(n6438), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n6450)
         );
  NAND3_X1 U5045 ( .A1(n24928), .A2(n24927), .A3(n24926), .ZN(n24929) );
  NAND3_X1 U5046 ( .A1(n24271), .A2(n3706), .A3(n24270), .ZN(n24277) );
  AND4_X1 U5047 ( .A1(n24265), .A2(n24264), .A3(n24263), .A4(n24262), .ZN(
        n24271) );
  AOI21_X1 U5048 ( .B1(\xmem_data[24][3] ), .B2(n28036), .A(n5815), .ZN(n5822)
         );
  NAND2_X1 U5049 ( .A1(n31261), .A2(\xmem_data[25][3] ), .ZN(n5813) );
  NAND3_X1 U5050 ( .A1(n24994), .A2(n24993), .A3(n24992), .ZN(n24995) );
  AND4_X1 U5051 ( .A1(n24955), .A2(n24954), .A3(n24953), .A4(n24952), .ZN(
        n24967) );
  NAND3_X1 U5052 ( .A1(n3709), .A2(n12249), .A3(n12248), .ZN(n12250) );
  NAND3_X1 U5053 ( .A1(n12279), .A2(n12278), .A3(n12277), .ZN(n12285) );
  NOR2_X1 U5054 ( .A1(n4797), .A2(n4796), .ZN(n4798) );
  NAND2_X1 U5055 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  NAND4_X1 U5056 ( .A1(n10464), .A2(n10463), .A3(n3710), .A4(n10462), .ZN(
        n10465) );
  NOR2_X1 U5057 ( .A1(n3990), .A2(n10453), .ZN(n10463) );
  NOR2_X1 U5058 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  OR2_X1 U5059 ( .A1(n36111), .A2(n3655), .ZN(n30397) );
  OR2_X1 U5060 ( .A1(n34615), .A2(n3600), .ZN(n30398) );
  AND2_X1 U5061 ( .A1(n34615), .A2(n30400), .ZN(n32222) );
  NAND3_X1 U5062 ( .A1(n7392), .A2(n7391), .A3(n7390), .ZN(n7393) );
  NAND3_X1 U5063 ( .A1(n7377), .A2(n7376), .A3(n7375), .ZN(n7383) );
  OR3_X1 U5064 ( .A1(n11997), .A2(n11996), .A3(n11995), .ZN(n11998) );
  NOR3_X1 U5065 ( .A1(n10571), .A2(n10570), .A3(n10569), .ZN(n10588) );
  OAI21_X1 U5066 ( .B1(n12957), .B2(n12956), .A(n23713), .ZN(n12958) );
  OR3_X1 U5067 ( .A1(n12955), .A2(n12954), .A3(n12953), .ZN(n12956) );
  OR2_X1 U5068 ( .A1(n7556), .A2(n7555), .ZN(n7564) );
  OR3_X1 U5069 ( .A1(n7516), .A2(n7515), .A3(n7514), .ZN(n7517) );
  OAI21_X1 U5070 ( .B1(n22612), .B2(n22611), .A(n29343), .ZN(n22637) );
  OR2_X1 U5071 ( .A1(n22626), .A2(n22625), .ZN(n22627) );
  NAND3_X1 U5072 ( .A1(n18036), .A2(n18035), .A3(n18034), .ZN(n18037) );
  AND3_X1 U5073 ( .A1(n18063), .A2(n18062), .A3(n18061), .ZN(n18066) );
  NOR2_X1 U5074 ( .A1(n11619), .A2(n11618), .ZN(n11624) );
  NAND4_X1 U5075 ( .A1(n3471), .A2(n3727), .A3(n3497), .A4(n3473), .ZN(n11709)
         );
  OR4_X1 U5076 ( .A1(n8191), .A2(n8190), .A3(n8189), .A4(n8188), .ZN(n8192) );
  OR4_X1 U5077 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8118), .ZN(n8122) );
  NAND3_X1 U5078 ( .A1(n7841), .A2(n7840), .A3(n7839), .ZN(n7842) );
  AOI22_X1 U5079 ( .A1(n8044), .A2(n28762), .B1(n28662), .B2(n8043), .ZN(n8100) );
  NOR2_X1 U5080 ( .A1(n34614), .A2(\fmem_data[21][0] ), .ZN(n31942) );
  NAND2_X1 U5081 ( .A1(n34683), .A2(n34682), .ZN(n34684) );
  XNOR2_X1 U5082 ( .A(n31673), .B(\fmem_data[10][5] ), .ZN(n30460) );
  AOI21_X1 U5083 ( .B1(n33250), .B2(n33249), .A(n33248), .ZN(n33251) );
  AND2_X1 U5084 ( .A1(n34418), .A2(n34420), .ZN(n30441) );
  XNOR2_X1 U5085 ( .A(n35104), .B(\fmem_data[13][5] ), .ZN(n35180) );
  XNOR2_X1 U5086 ( .A(n35076), .B(\fmem_data[30][5] ), .ZN(n33106) );
  XNOR2_X1 U5087 ( .A(n33967), .B(\fmem_data[8][7] ), .ZN(n33383) );
  XNOR2_X1 U5088 ( .A(n35401), .B(\fmem_data[0][5] ), .ZN(n33385) );
  AND2_X1 U5089 ( .A1(n8365), .A2(n8364), .ZN(n8378) );
  AND4_X1 U5090 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n8379)
         );
  AOI21_X1 U5091 ( .B1(n33850), .B2(n33851), .A(n30159), .ZN(n4470) );
  XNOR2_X1 U5092 ( .A(n31996), .B(\fmem_data[8][5] ), .ZN(n31826) );
  XNOR2_X1 U5093 ( .A(n32115), .B(\fmem_data[21][7] ), .ZN(n30381) );
  INV_X1 U5094 ( .A(n3411), .ZN(n3413) );
  OR4_X1 U5095 ( .A1(n17893), .A2(n17892), .A3(n17891), .A4(n17890), .ZN(
        n17894) );
  OR2_X1 U5096 ( .A1(n24497), .A2(n24496), .ZN(n24507) );
  OR3_X1 U5097 ( .A1(n24580), .A2(n24579), .A3(n24578), .ZN(n24582) );
  NAND2_X1 U5098 ( .A1(n9707), .A2(n20795), .ZN(n9774) );
  NAND3_X1 U5099 ( .A1(n12209), .A2(n12208), .A3(n12207), .ZN(n12220) );
  NOR2_X1 U5100 ( .A1(n3720), .A2(n12153), .ZN(n12154) );
  AND4_X1 U5101 ( .A1(n10781), .A2(n10780), .A3(n10779), .A4(n10778), .ZN(
        n10787) );
  AOI21_X1 U5102 ( .B1(n27568), .B2(\xmem_data[85][7] ), .A(n14264), .ZN(
        n14268) );
  AND2_X1 U5103 ( .A1(n23725), .A2(\xmem_data[84][7] ), .ZN(n14264) );
  INV_X1 U5104 ( .A(n3336), .ZN(n3337) );
  NAND4_X1 U5105 ( .A1(n3738), .A2(n25500), .A3(n25499), .A4(n25498), .ZN(
        n25507) );
  NOR2_X1 U5106 ( .A1(n25497), .A2(n25496), .ZN(n25498) );
  OR2_X1 U5107 ( .A1(n25174), .A2(n25173), .ZN(n25175) );
  OR3_X1 U5108 ( .A1(n4455), .A2(n4454), .A3(n4453), .ZN(n4465) );
  OR3_X1 U5109 ( .A1(n4436), .A2(n4435), .A3(n4434), .ZN(n4438) );
  NAND2_X1 U5110 ( .A1(n28007), .A2(\xmem_data[30][7] ), .ZN(n4389) );
  OAI21_X1 U5111 ( .B1(n4417), .B2(n4416), .A(n22663), .ZN(n4468) );
  OR3_X1 U5112 ( .A1(n4415), .A2(n4414), .A3(n4413), .ZN(n4416) );
  NOR2_X1 U5113 ( .A1(n14474), .A2(n14473), .ZN(n14501) );
  OR3_X1 U5114 ( .A1(n14159), .A2(n14158), .A3(n14157), .ZN(n14160) );
  XNOR2_X1 U5115 ( .A(n31250), .B(\fmem_data[1][7] ), .ZN(n31813) );
  AOI21_X1 U5116 ( .B1(n35182), .B2(n35181), .A(n35180), .ZN(n35183) );
  XNOR2_X1 U5117 ( .A(n31642), .B(\fmem_data[20][7] ), .ZN(n35179) );
  AOI21_X1 U5118 ( .B1(n34986), .B2(n34985), .A(n34984), .ZN(n34987) );
  XNOR2_X1 U5119 ( .A(n34859), .B(\fmem_data[25][7] ), .ZN(n34983) );
  XNOR2_X1 U5120 ( .A(n31995), .B(\fmem_data[8][7] ), .ZN(n33384) );
  NAND3_X1 U5121 ( .A1(n27188), .A2(n27187), .A3(n27186), .ZN(n27189) );
  INV_X1 U5122 ( .A(n3331), .ZN(n3332) );
  AND2_X1 U5123 ( .A1(n26840), .A2(n26839), .ZN(n26841) );
  NOR2_X1 U5124 ( .A1(n19318), .A2(n19317), .ZN(n19322) );
  NAND2_X1 U5125 ( .A1(n19316), .A2(n19315), .ZN(n19317) );
  AND2_X1 U5126 ( .A1(n26722), .A2(n26721), .ZN(n26723) );
  OR2_X1 U5127 ( .A1(n20948), .A2(n3924), .ZN(n20977) );
  INV_X1 U5128 ( .A(n31026), .ZN(n31032) );
  NAND3_X1 U5129 ( .A1(n19156), .A2(n19155), .A3(n19154), .ZN(n19157) );
  NOR2_X1 U5130 ( .A1(n23446), .A2(n23445), .ZN(n23447) );
  INV_X1 U5131 ( .A(n3327), .ZN(n3330) );
  NAND3_X1 U5132 ( .A1(n29112), .A2(n29111), .A3(n29110), .ZN(n29113) );
  NAND3_X1 U5133 ( .A1(n29092), .A2(n29091), .A3(n29090), .ZN(n29093) );
  OR2_X1 U5134 ( .A1(n20366), .A2(n3928), .ZN(n20385) );
  AND2_X1 U5135 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  OR4_X1 U5136 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .ZN(n8686) );
  NAND3_X1 U5137 ( .A1(n11898), .A2(n11897), .A3(n11896), .ZN(n11899) );
  OR2_X1 U5138 ( .A1(n22481), .A2(n22480), .ZN(n22482) );
  NAND2_X1 U5139 ( .A1(n22479), .A2(n22478), .ZN(n22480) );
  NAND3_X1 U5140 ( .A1(n26513), .A2(n26512), .A3(n26511), .ZN(n26514) );
  OR3_X1 U5141 ( .A1(n26561), .A2(n26560), .A3(n26559), .ZN(n26567) );
  AND2_X1 U5142 ( .A1(n15625), .A2(n15624), .ZN(n15626) );
  OR2_X1 U5143 ( .A1(n8761), .A2(n8760), .ZN(n8780) );
  AND2_X1 U5144 ( .A1(n8738), .A2(n8737), .ZN(n8755) );
  NAND3_X1 U5145 ( .A1(n20216), .A2(n20215), .A3(n20214), .ZN(n20217) );
  NOR2_X1 U5146 ( .A1(n4629), .A2(n4628), .ZN(n4644) );
  NOR2_X1 U5147 ( .A1(n4636), .A2(n4635), .ZN(n4643) );
  AND4_X1 U5148 ( .A1(n18217), .A2(n18216), .A3(n18215), .A4(n18214), .ZN(
        n18229) );
  AND2_X1 U5149 ( .A1(n18298), .A2(n18297), .ZN(n18305) );
  NAND2_X1 U5150 ( .A1(n6387), .A2(n30228), .ZN(n6388) );
  AND2_X1 U5151 ( .A1(n36112), .A2(n31382), .ZN(n31522) );
  NOR2_X1 U5152 ( .A1(n16407), .A2(n16406), .ZN(n16408) );
  OAI21_X1 U5153 ( .B1(n24663), .B2(n24662), .A(n24661), .ZN(n24664) );
  AOI21_X1 U5154 ( .B1(n24660), .B2(n24659), .A(n24658), .ZN(n24661) );
  XNOR2_X1 U5155 ( .A(n33554), .B(\fmem_data[2][3] ), .ZN(n32422) );
  INV_X1 U5156 ( .A(n35641), .ZN(n32287) );
  XNOR2_X1 U5157 ( .A(n36338), .B(\fmem_data[1][7] ), .ZN(n32180) );
  XNOR2_X1 U5158 ( .A(n32442), .B(\fmem_data[1][7] ), .ZN(n33216) );
  XNOR2_X1 U5159 ( .A(n31161), .B(\fmem_data[22][5] ), .ZN(n31993) );
  XNOR2_X1 U5160 ( .A(n31492), .B(\fmem_data[25][7] ), .ZN(n33247) );
  AND4_X1 U5161 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n10881) );
  AND2_X1 U5162 ( .A1(n6577), .A2(n6576), .ZN(n6580) );
  OR2_X1 U5163 ( .A1(n6575), .A2(n25514), .ZN(n6577) );
  OR2_X1 U5164 ( .A1(n6575), .A2(\xmem_data[7][7] ), .ZN(n6576) );
  OR4_X1 U5165 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n6555) );
  OR4_X1 U5166 ( .A1(n25669), .A2(n25668), .A3(n25667), .A4(n25666), .ZN(
        n25705) );
  AND2_X1 U5167 ( .A1(n15839), .A2(n15838), .ZN(n15857) );
  NAND3_X1 U5168 ( .A1(n15804), .A2(n15803), .A3(n15802), .ZN(n15805) );
  NAND3_X1 U5169 ( .A1(n15830), .A2(n15829), .A3(n15828), .ZN(n15831) );
  OAI21_X1 U5170 ( .B1(n15880), .B2(n15879), .A(n29683), .ZN(n15881) );
  OR2_X1 U5171 ( .A1(n15867), .A2(n15866), .ZN(n15880) );
  OR2_X1 U5172 ( .A1(n15878), .A2(n15877), .ZN(n15879) );
  NAND3_X1 U5173 ( .A1(n24893), .A2(n24892), .A3(n24891), .ZN(n24894) );
  AND2_X1 U5174 ( .A1(n24882), .A2(n24881), .ZN(n24883) );
  AND4_X1 U5175 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11530) );
  NOR3_X1 U5176 ( .A1(n24374), .A2(n24373), .A3(n24372), .ZN(n24383) );
  OAI21_X1 U5177 ( .B1(n5450), .B2(n5449), .A(n29002), .ZN(n5451) );
  OAI21_X1 U5178 ( .B1(n5385), .B2(n5384), .A(n28968), .ZN(n5454) );
  NAND2_X1 U5179 ( .A1(n5429), .A2(n29078), .ZN(n5452) );
  NAND2_X1 U5180 ( .A1(n27324), .A2(\fmem_data[20][7] ), .ZN(n27325) );
  OAI22_X1 U5181 ( .A1(n32651), .A2(n35614), .B1(n30449), .B2(n35615), .ZN(
        n30486) );
  OR2_X1 U5182 ( .A1(n35749), .A2(n3614), .ZN(n30386) );
  AOI21_X1 U5183 ( .B1(n34788), .B2(n3560), .A(n33978), .ZN(n30468) );
  OR2_X1 U5184 ( .A1(n32012), .A2(n34497), .ZN(n30160) );
  XNOR2_X1 U5185 ( .A(n32176), .B(\fmem_data[1][3] ), .ZN(n33994) );
  OR2_X1 U5186 ( .A1(n36299), .A2(n3621), .ZN(n17555) );
  OR2_X1 U5187 ( .A1(n35011), .A2(n3632), .ZN(n28540) );
  OR2_X1 U5188 ( .A1(n33956), .A2(n3696), .ZN(n28542) );
  OR2_X1 U5189 ( .A1(n35006), .A2(n3649), .ZN(n33826) );
  XNOR2_X1 U5190 ( .A(n33573), .B(\fmem_data[28][3] ), .ZN(n33854) );
  XNOR2_X1 U5191 ( .A(n33553), .B(\fmem_data[5][5] ), .ZN(n33860) );
  XNOR2_X1 U5192 ( .A(n32614), .B(\fmem_data[24][7] ), .ZN(n31954) );
  XNOR2_X1 U5193 ( .A(n30451), .B(\fmem_data[6][5] ), .ZN(n33188) );
  XNOR2_X1 U5194 ( .A(n32427), .B(\fmem_data[8][7] ), .ZN(n33257) );
  XNOR2_X1 U5195 ( .A(n35076), .B(\fmem_data[30][1] ), .ZN(n33978) );
  XNOR2_X1 U5196 ( .A(n32235), .B(\fmem_data[12][5] ), .ZN(n33974) );
  XNOR2_X1 U5197 ( .A(n31992), .B(\fmem_data[22][5] ), .ZN(n33964) );
  AND2_X1 U5198 ( .A1(n36105), .A2(n33959), .ZN(n34069) );
  AND2_X1 U5199 ( .A1(n34624), .A2(n33958), .ZN(n34070) );
  XNOR2_X1 U5200 ( .A(n32616), .B(\fmem_data[9][7] ), .ZN(n34242) );
  OAI22_X1 U5201 ( .A1(n33274), .A2(n33582), .B1(n33273), .B2(n34340), .ZN(
        n34103) );
  OAI22_X1 U5202 ( .A1(n33270), .A2(n34194), .B1(n33269), .B2(n34195), .ZN(
        n34104) );
  OAI21_X1 U5203 ( .B1(n33943), .B2(n33941), .A(n33942), .ZN(n21397) );
  NAND2_X1 U5204 ( .A1(n33943), .A2(n33941), .ZN(n21396) );
  XNOR2_X1 U5205 ( .A(n30156), .B(\fmem_data[28][5] ), .ZN(n32754) );
  XNOR2_X1 U5206 ( .A(n32057), .B(\fmem_data[21][7] ), .ZN(n32756) );
  XNOR2_X1 U5207 ( .A(n36105), .B(\fmem_data[18][7] ), .ZN(n32007) );
  XNOR2_X1 U5208 ( .A(n31161), .B(\fmem_data[22][3] ), .ZN(n32003) );
  OAI22_X1 U5209 ( .A1(n30437), .A2(n35592), .B1(n33199), .B2(n35591), .ZN(
        n31961) );
  OAI22_X1 U5210 ( .A1(n30436), .A2(n34195), .B1(n33269), .B2(n34194), .ZN(
        n31962) );
  OAI22_X1 U5211 ( .A1(n30435), .A2(n33859), .B1(n30434), .B2(n33857), .ZN(
        n31963) );
  XNOR2_X1 U5212 ( .A(n32543), .B(\fmem_data[17][5] ), .ZN(n32322) );
  NAND2_X1 U5213 ( .A1(n30484), .A2(n30482), .ZN(n30469) );
  XNOR2_X1 U5214 ( .A(n32939), .B(\fmem_data[1][7] ), .ZN(n32179) );
  AOI21_X1 U5215 ( .B1(n33873), .B2(n33875), .A(n33044), .ZN(n14288) );
  XNOR2_X1 U5216 ( .A(n31995), .B(\fmem_data[8][5] ), .ZN(n24016) );
  NAND2_X1 U5217 ( .A1(n34856), .A2(n34855), .ZN(n34857) );
  NAND2_X1 U5218 ( .A1(n32036), .A2(n32035), .ZN(n34970) );
  OAI21_X1 U5219 ( .B1(n33086), .B2(n33085), .A(n33084), .ZN(n32036) );
  NAND2_X1 U5220 ( .A1(n33085), .A2(n33086), .ZN(n32035) );
  OAI22_X1 U5221 ( .A1(n24431), .A2(n35580), .B1(n33313), .B2(n35581), .ZN(
        n33341) );
  INV_X1 U5222 ( .A(n33032), .ZN(n33136) );
  OAI22_X1 U5223 ( .A1(n34233), .A2(n34836), .B1(n33028), .B2(n34835), .ZN(
        n33138) );
  OAI22_X1 U5224 ( .A1(n31973), .A2(n34941), .B1(n31972), .B2(n34942), .ZN(
        n33140) );
  OAI22_X1 U5225 ( .A1(n31975), .A2(n35662), .B1(n31974), .B2(n35663), .ZN(
        n33139) );
  AOI21_X1 U5226 ( .B1(n34422), .B2(n34424), .A(n33017), .ZN(n33018) );
  NAND2_X1 U5227 ( .A1(n10945), .A2(n10944), .ZN(n12721) );
  NAND2_X1 U5228 ( .A1(n17750), .A2(n17749), .ZN(n10944) );
  INV_X1 U5229 ( .A(n33053), .ZN(n33363) );
  AOI21_X1 U5230 ( .B1(n33568), .B2(n33570), .A(n33052), .ZN(n33053) );
  INV_X1 U5231 ( .A(n33051), .ZN(n33364) );
  OAI22_X1 U5232 ( .A1(n33040), .A2(n33642), .B1(n33386), .B2(n33643), .ZN(
        n33375) );
  OAI21_X1 U5233 ( .B1(n34839), .B2(n34840), .A(n34838), .ZN(n34842) );
  NAND2_X1 U5234 ( .A1(n34840), .A2(n34839), .ZN(n34841) );
  NAND2_X1 U5235 ( .A1(n34832), .A2(n34831), .ZN(n34833) );
  OAI22_X1 U5236 ( .A1(n33228), .A2(n35576), .B1(n33311), .B2(n35577), .ZN(
        n33380) );
  OAI22_X1 U5237 ( .A1(n33224), .A2(n33961), .B1(n33223), .B2(n33963), .ZN(
        n33382) );
  OAI22_X1 U5238 ( .A1(n33226), .A2(n35752), .B1(n34863), .B2(n35753), .ZN(
        n33381) );
  OAI22_X1 U5239 ( .A1(n33310), .A2(n33859), .B1(n33309), .B2(n33857), .ZN(
        n34950) );
  OAI22_X1 U5240 ( .A1(n33314), .A2(n35581), .B1(n33313), .B2(n35580), .ZN(
        n34948) );
  OAI22_X1 U5241 ( .A1(n33312), .A2(n35577), .B1(n33311), .B2(n35576), .ZN(
        n34949) );
  OAI22_X1 U5242 ( .A1(n24726), .A2(n35181), .B1(n33102), .B2(n35182), .ZN(
        n11339) );
  OR2_X1 U5243 ( .A1(n30464), .A2(n30463), .ZN(n31687) );
  AND2_X1 U5244 ( .A1(n34410), .A2(n34412), .ZN(n30463) );
  OAI22_X1 U5245 ( .A1(n30446), .A2(n33596), .B1(n30445), .B2(n33598), .ZN(
        n31735) );
  OAI22_X1 U5246 ( .A1(n30450), .A2(n35615), .B1(n30449), .B2(n35614), .ZN(
        n31733) );
  OAI22_X1 U5247 ( .A1(n33188), .A2(n33954), .B1(n33369), .B2(n33956), .ZN(
        n31681) );
  OAI21_X1 U5248 ( .B1(n30443), .B2(n31693), .A(n31692), .ZN(n31722) );
  NAND2_X1 U5249 ( .A1(n31691), .A2(n31690), .ZN(n31692) );
  NOR2_X1 U5250 ( .A1(n31691), .A2(n31690), .ZN(n31693) );
  NAND2_X1 U5251 ( .A1(n31696), .A2(n31695), .ZN(n31697) );
  OAI22_X1 U5252 ( .A1(n31985), .A2(n35708), .B1(n33307), .B2(n35709), .ZN(
        n31727) );
  XNOR2_X1 U5253 ( .A(n32225), .B(\fmem_data[9][7] ), .ZN(n35022) );
  OAI22_X1 U5254 ( .A1(n33130), .A2(n33963), .B1(n33223), .B2(n33961), .ZN(
        n35014) );
  OAI22_X1 U5255 ( .A1(n33127), .A2(n34045), .B1(n34043), .B2(n33126), .ZN(
        n35016) );
  OAI22_X1 U5256 ( .A1(n33129), .A2(n35615), .B1(n33128), .B2(n35614), .ZN(
        n35015) );
  OAI22_X1 U5257 ( .A1(n35177), .A2(n35585), .B1(n31665), .B2(n35584), .ZN(
        n31701) );
  OAI22_X1 U5258 ( .A1(n35087), .A2(n35089), .B1(n31666), .B2(n35088), .ZN(
        n31700) );
  AND2_X1 U5259 ( .A1(n34466), .A2(n34779), .ZN(n25149) );
  OAI22_X1 U5260 ( .A1(n30435), .A2(n33857), .B1(n33309), .B2(n33859), .ZN(
        n23921) );
  OAI22_X1 U5261 ( .A1(n30354), .A2(n35760), .B1(n33317), .B2(n35761), .ZN(
        n25599) );
  OAI22_X1 U5262 ( .A1(n31824), .A2(n35494), .B1(n31641), .B2(n35493), .ZN(
        n31708) );
  OAI22_X1 U5263 ( .A1(n31816), .A2(n35490), .B1(n31639), .B2(n35489), .ZN(
        n31709) );
  OAI22_X1 U5264 ( .A1(n34921), .A2(n34923), .B1(n33219), .B2(n34922), .ZN(
        n31782) );
  AND4_X1 U5265 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n7721)
         );
  OR4_X1 U5266 ( .A1(n24148), .A2(n24147), .A3(n24146), .A4(n24145), .ZN(
        n24149) );
  OAI22_X1 U5267 ( .A1(n34930), .A2(n35511), .B1(n35121), .B2(n35512), .ZN(
        n35069) );
  OAI22_X1 U5268 ( .A1(n33371), .A2(n34039), .B1(n33370), .B2(n34041), .ZN(
        n34937) );
  OAI22_X1 U5269 ( .A1(n33373), .A2(n33975), .B1(n33372), .B2(n33973), .ZN(
        n34936) );
  INV_X1 U5270 ( .A(n35090), .ZN(n35117) );
  XNOR2_X1 U5271 ( .A(n31892), .B(\fmem_data[1][7] ), .ZN(n35281) );
  OAI22_X1 U5272 ( .A1(n33388), .A2(n35610), .B1(n35356), .B2(n35611), .ZN(
        n35323) );
  INV_X1 U5273 ( .A(n31676), .ZN(n35321) );
  INV_X1 U5274 ( .A(n31675), .ZN(n35322) );
  OAI22_X1 U5275 ( .A1(n33129), .A2(n35614), .B1(n35358), .B2(n35615), .ZN(
        n35331) );
  OAI22_X1 U5276 ( .A1(n33312), .A2(n35576), .B1(n35103), .B2(n35577), .ZN(
        n35332) );
  OAI22_X1 U5277 ( .A1(n33133), .A2(n35591), .B1(n35105), .B2(n35592), .ZN(
        n35334) );
  INV_X1 U5278 ( .A(n31804), .ZN(n35342) );
  INV_X1 U5279 ( .A(n31803), .ZN(n35343) );
  OAI22_X1 U5280 ( .A1(n33308), .A2(n35708), .B1(n35077), .B2(n35709), .ZN(
        n35313) );
  OAI22_X1 U5281 ( .A1(n33306), .A2(n35748), .B1(n35325), .B2(n35749), .ZN(
        n35314) );
  OAI22_X1 U5282 ( .A1(n33318), .A2(n35760), .B1(n35400), .B2(n35761), .ZN(
        n35315) );
  BUF_X2 U5283 ( .A(n17042), .Z(n17019) );
  CLKBUF_X1 U5284 ( .A(n39053), .Z(n3346) );
  INV_X1 U5285 ( .A(n3304), .ZN(n3383) );
  AND2_X1 U5286 ( .A1(n4062), .A2(n7216), .ZN(n4236) );
  INV_X1 U5287 ( .A(n17032), .ZN(n3448) );
  INV_X1 U5288 ( .A(n30961), .ZN(n3331) );
  CLKBUF_X1 U5289 ( .A(n28973), .Z(n30961) );
  AND2_X1 U5290 ( .A1(n13432), .A2(n5691), .ZN(n5692) );
  INV_X1 U5291 ( .A(n5985), .ZN(n5691) );
  INV_X1 U5292 ( .A(n30961), .ZN(n3411) );
  XNOR2_X1 U5293 ( .A(n5289), .B(load_xaddr_val[6]), .ZN(n5359) );
  NAND2_X1 U5294 ( .A1(n5288), .A2(n37191), .ZN(n5289) );
  NOR2_X1 U5295 ( .A1(n7206), .A2(n8005), .ZN(n7640) );
  NAND2_X1 U5296 ( .A1(n6201), .A2(n11357), .ZN(n6202) );
  NAND3_X1 U5297 ( .A1(n11343), .A2(n11342), .A3(n6173), .ZN(n7010) );
  INV_X1 U5298 ( .A(n3230), .ZN(n8420) );
  AND3_X1 U5299 ( .A1(n23051), .A2(n23050), .A3(n23049), .ZN(n23069) );
  INV_X1 U5300 ( .A(n3304), .ZN(n3305) );
  AOI22_X1 U5301 ( .A1(n27031), .A2(\xmem_data[118][1] ), .B1(n25678), .B2(
        \xmem_data[119][1] ), .ZN(n27032) );
  NAND3_X1 U5302 ( .A1(n27089), .A2(n27088), .A3(n27087), .ZN(n27092) );
  NAND3_X1 U5303 ( .A1(n26995), .A2(n26994), .A3(n26993), .ZN(n26996) );
  AND2_X1 U5304 ( .A1(n17318), .A2(n17389), .ZN(n17320) );
  NOR2_X1 U5305 ( .A1(n22864), .A2(n22863), .ZN(n22876) );
  NAND2_X1 U5306 ( .A1(n22880), .A2(n3953), .ZN(n22881) );
  NAND2_X1 U5307 ( .A1(n22878), .A2(n28007), .ZN(n22880) );
  CLKBUF_X1 U5308 ( .A(n28973), .Z(n28077) );
  INV_X1 U5309 ( .A(n30907), .ZN(n3349) );
  CLKBUF_X1 U5310 ( .A(n28973), .Z(n30907) );
  NAND3_X1 U5311 ( .A1(n22032), .A2(n22031), .A3(n22030), .ZN(n22033) );
  OAI21_X1 U5312 ( .B1(n19502), .B2(n19501), .A(n19410), .ZN(n19503) );
  OR4_X1 U5313 ( .A1(n19500), .A2(n19499), .A3(n19498), .A4(n19497), .ZN(
        n19501) );
  AND2_X1 U5314 ( .A1(n18848), .A2(n18847), .ZN(n18849) );
  OR2_X1 U5315 ( .A1(n36228), .A2(n3593), .ZN(n32608) );
  OR2_X1 U5316 ( .A1(n34624), .A2(n3604), .ZN(n32551) );
  OR2_X1 U5317 ( .A1(n36105), .A2(n3664), .ZN(n32550) );
  XNOR2_X1 U5318 ( .A(n32317), .B(\fmem_data[4][1] ), .ZN(n33649) );
  OR2_X1 U5319 ( .A1(n36312), .A2(n3611), .ZN(n33691) );
  XNOR2_X1 U5320 ( .A(n31592), .B(\fmem_data[29][1] ), .ZN(n33580) );
  OAI22_X1 U5321 ( .A1(n33787), .A2(n35033), .B1(n33786), .B2(n35034), .ZN(
        n33899) );
  OR2_X1 U5322 ( .A1(n35003), .A2(n3594), .ZN(n33785) );
  OAI22_X1 U5323 ( .A1(n33781), .A2(n34734), .B1(n33780), .B2(n3572), .ZN(
        n33806) );
  XNOR2_X1 U5324 ( .A(n36105), .B(\fmem_data[18][3] ), .ZN(n33680) );
  XNOR2_X1 U5325 ( .A(n36101), .B(\fmem_data[24][3] ), .ZN(n33684) );
  XNOR2_X1 U5326 ( .A(n36200), .B(\fmem_data[30][3] ), .ZN(n33678) );
  OAI22_X1 U5327 ( .A1(n32563), .A2(n33643), .B1(n31469), .B2(n33642), .ZN(
        n33673) );
  OAI22_X1 U5328 ( .A1(n31505), .A2(n34422), .B1(n34424), .B2(n3587), .ZN(
        n33489) );
  NAND3_X1 U5329 ( .A1(n6796), .A2(n6795), .A3(n6794), .ZN(n31221) );
  NAND4_X1 U5330 ( .A1(n16155), .A2(n16154), .A3(n16153), .A4(n16152), .ZN(
        n31219) );
  NAND2_X1 U5331 ( .A1(n31523), .A2(n31522), .ZN(n31384) );
  OR2_X1 U5332 ( .A1(n36339), .A2(n3619), .ZN(n31251) );
  XNOR2_X1 U5333 ( .A(n33592), .B(\fmem_data[14][3] ), .ZN(n33602) );
  XNOR2_X1 U5334 ( .A(n31125), .B(\fmem_data[0][1] ), .ZN(n33577) );
  OR2_X1 U5335 ( .A1(n36200), .A2(n3592), .ZN(n31595) );
  XNOR2_X1 U5336 ( .A(n36200), .B(\fmem_data[30][5] ), .ZN(n31168) );
  XNOR2_X1 U5337 ( .A(n36105), .B(\fmem_data[18][5] ), .ZN(n31164) );
  NAND2_X1 U5338 ( .A1(n12810), .A2(n33797), .ZN(n33796) );
  XOR2_X1 U5339 ( .A(\fmem_data[2][2] ), .B(\fmem_data[2][3] ), .Z(n12810) );
  XNOR2_X1 U5340 ( .A(n32235), .B(\fmem_data[12][3] ), .ZN(n33581) );
  XNOR2_X1 U5341 ( .A(n32176), .B(\fmem_data[1][1] ), .ZN(n32443) );
  XNOR2_X1 U5342 ( .A(n32442), .B(\fmem_data[1][1] ), .ZN(n33688) );
  XNOR2_X1 U5343 ( .A(n33484), .B(\fmem_data[31][3] ), .ZN(n32621) );
  XNOR2_X1 U5344 ( .A(n32543), .B(\fmem_data[17][1] ), .ZN(n33833) );
  XNOR2_X1 U5345 ( .A(n32065), .B(\fmem_data[0][3] ), .ZN(n32535) );
  OR2_X1 U5346 ( .A1(n35697), .A2(n3486), .ZN(n32292) );
  NAND2_X1 U5347 ( .A1(n32290), .A2(\fmem_data[15][7] ), .ZN(n32291) );
  INV_X1 U5348 ( .A(n35696), .ZN(n32290) );
  OAI22_X1 U5349 ( .A1(n34198), .A2(n34476), .B1(n32226), .B2(n3579), .ZN(
        n32313) );
  OAI22_X1 U5350 ( .A1(n33846), .A2(n35040), .B1(n32227), .B2(n35041), .ZN(
        n32312) );
  OAI22_X1 U5351 ( .A1(n32229), .A2(n33850), .B1(n33851), .B2(n33849), .ZN(
        n32311) );
  OAI22_X1 U5352 ( .A1(n32668), .A2(n35709), .B1(n32667), .B2(n35708), .ZN(
        n32719) );
  OAI22_X1 U5353 ( .A1(n32666), .A2(n35490), .B1(n32665), .B2(n35489), .ZN(
        n32720) );
  AND2_X1 U5354 ( .A1(n36244), .A2(n32114), .ZN(n32231) );
  OAI22_X1 U5355 ( .A1(n34202), .A2(n34199), .B1(n32116), .B2(n34201), .ZN(
        n32230) );
  OAI22_X1 U5356 ( .A1(n31965), .A2(n33570), .B1(n31964), .B2(n33568), .ZN(
        n32173) );
  INV_X1 U5357 ( .A(n31969), .ZN(n32171) );
  OAI22_X1 U5358 ( .A1(n33957), .A2(n33954), .B1(n33187), .B2(n33956), .ZN(
        n32185) );
  NAND2_X1 U5359 ( .A1(n31914), .A2(n31913), .ZN(n31111) );
  XNOR2_X1 U5360 ( .A(n33754), .B(\fmem_data[0][7] ), .ZN(n31014) );
  OAI22_X1 U5361 ( .A1(n32717), .A2(n34433), .B1(n30983), .B2(n34431), .ZN(
        n31743) );
  XNOR2_X1 U5362 ( .A(n31640), .B(\fmem_data[0][5] ), .ZN(n33040) );
  XNOR2_X1 U5363 ( .A(n31638), .B(\fmem_data[24][5] ), .ZN(n33215) );
  XNOR2_X1 U5364 ( .A(n35073), .B(\fmem_data[22][1] ), .ZN(n33947) );
  XNOR2_X1 U5365 ( .A(n33227), .B(\fmem_data[14][3] ), .ZN(n26271) );
  XNOR2_X1 U5366 ( .A(n31664), .B(\fmem_data[22][1] ), .ZN(n31162) );
  NAND2_X1 U5367 ( .A1(n26376), .A2(n26375), .ZN(n21091) );
  OAI22_X1 U5368 ( .A1(n33017), .A2(n34422), .B1(n32320), .B2(n34424), .ZN(
        n23829) );
  XNOR2_X1 U5369 ( .A(n32617), .B(\fmem_data[9][5] ), .ZN(n30360) );
  NAND2_X1 U5370 ( .A1(n7107), .A2(n7106), .ZN(n7192) );
  NAND2_X1 U5371 ( .A1(n9386), .A2(n35019), .ZN(n35018) );
  XNOR2_X1 U5372 ( .A(n32117), .B(\fmem_data[6][5] ), .ZN(n33955) );
  XNOR2_X1 U5373 ( .A(n32617), .B(\fmem_data[9][3] ), .ZN(n33874) );
  XNOR2_X1 U5374 ( .A(n33551), .B(\fmem_data[20][7] ), .ZN(n30795) );
  OAI22_X1 U5375 ( .A1(n32529), .A2(n34424), .B1(n33965), .B2(n34422), .ZN(
        n31915) );
  OAI22_X1 U5376 ( .A1(n31123), .A2(n35088), .B1(n30800), .B2(n35089), .ZN(
        n31907) );
  AOI21_X1 U5377 ( .B1(n34529), .B2(n3566), .A(n33950), .ZN(n30163) );
  OAI22_X1 U5378 ( .A1(n32058), .A2(n34613), .B1(n34024), .B2(n3570), .ZN(
        n33576) );
  OAI22_X1 U5379 ( .A1(n33646), .A2(n33681), .B1(n33645), .B2(n33679), .ZN(
        n34065) );
  OAI22_X1 U5380 ( .A1(n32523), .A2(n35036), .B1(n31195), .B2(n35037), .ZN(
        n31495) );
  OAI22_X1 U5381 ( .A1(n34209), .A2(n34206), .B1(n33831), .B2(n34208), .ZN(
        n31497) );
  OAI22_X1 U5382 ( .A1(n34403), .A2(n36223), .B1(n32212), .B2(n3568), .ZN(
        n32271) );
  NAND2_X1 U5383 ( .A1(n32411), .A2(n32410), .ZN(n32206) );
  OAI22_X1 U5384 ( .A1(n32059), .A2(n36227), .B1(n31446), .B2(n3647), .ZN(
        n31486) );
  OAI22_X1 U5385 ( .A1(n31911), .A2(n36100), .B1(n26806), .B2(n3565), .ZN(
        n28900) );
  OAI22_X1 U5386 ( .A1(n30998), .A2(n33105), .B1(n30997), .B2(n33103), .ZN(
        n31155) );
  OAI22_X1 U5387 ( .A1(n32126), .A2(n34625), .B1(n29519), .B2(n3574), .ZN(
        n31228) );
  XNOR2_X1 U5388 ( .A(n31250), .B(\fmem_data[1][1] ), .ZN(n33867) );
  XNOR2_X1 U5389 ( .A(n31892), .B(\fmem_data[1][1] ), .ZN(n33866) );
  OAI22_X1 U5390 ( .A1(n34018), .A2(n34017), .B1(n34016), .B2(n3559), .ZN(
        n34316) );
  XNOR2_X1 U5391 ( .A(n28539), .B(\fmem_data[13][5] ), .ZN(n33163) );
  AOI21_X1 U5392 ( .B1(n34476), .B2(n3579), .A(n33197), .ZN(n33198) );
  OAI22_X1 U5393 ( .A1(n32576), .A2(n33956), .B1(n32575), .B2(n33954), .ZN(
        n32798) );
  OAI22_X1 U5394 ( .A1(n32585), .A2(n3569), .B1(n33648), .B2(n34598), .ZN(
        n32774) );
  OR2_X1 U5395 ( .A1(n36312), .A2(n3631), .ZN(n32726) );
  OAI22_X1 U5396 ( .A1(n31973), .A2(n34942), .B1(n30169), .B2(n34941), .ZN(
        n34272) );
  OAI22_X1 U5397 ( .A1(n33978), .A2(n3560), .B1(n34788), .B2(n33977), .ZN(
        n34007) );
  OAI22_X1 U5398 ( .A1(n33976), .A2(n33975), .B1(n33974), .B2(n33973), .ZN(
        n34006) );
  OAI22_X1 U5399 ( .A1(n33968), .A2(n34206), .B1(n34207), .B2(n34208), .ZN(
        n34060) );
  OAI22_X1 U5400 ( .A1(n33970), .A2(n3563), .B1(n33969), .B2(n34739), .ZN(
        n34059) );
  NAND2_X1 U5401 ( .A1(n33931), .A2(n33930), .ZN(n34228) );
  NAND2_X1 U5402 ( .A1(n36223), .A2(n3568), .ZN(n33930) );
  INV_X1 U5403 ( .A(n33929), .ZN(n33931) );
  OAI22_X1 U5404 ( .A1(n33928), .A2(n3571), .B1(n33927), .B2(n34742), .ZN(
        n33936) );
  OAI22_X1 U5405 ( .A1(n33926), .A2(n35516), .B1(n35515), .B2(n3615), .ZN(
        n33937) );
  OAI22_X1 U5406 ( .A1(n33925), .A2(n35515), .B1(n33924), .B2(n35516), .ZN(
        n33938) );
  INV_X1 U5407 ( .A(n34079), .ZN(n34247) );
  OAI22_X1 U5408 ( .A1(n21766), .A2(n35585), .B1(n35584), .B2(n3645), .ZN(
        n34010) );
  OAI22_X1 U5409 ( .A1(n21583), .A2(n35577), .B1(n35576), .B2(n3598), .ZN(
        n34012) );
  OAI22_X1 U5410 ( .A1(n21674), .A2(n35709), .B1(n35708), .B2(n3585), .ZN(
        n34011) );
  OAI22_X1 U5411 ( .A1(n27327), .A2(n35007), .B1(n33033), .B2(n35006), .ZN(
        n34238) );
  OAI22_X1 U5412 ( .A1(n31985), .A2(n35709), .B1(n31984), .B2(n35708), .ZN(
        n33026) );
  NAND2_X1 U5413 ( .A1(n32358), .A2(n32357), .ZN(n32033) );
  OAI22_X1 U5414 ( .A1(n32715), .A2(n35610), .B1(n33268), .B2(n35611), .ZN(
        n32743) );
  NAND2_X1 U5415 ( .A1(n32769), .A2(n32768), .ZN(n32673) );
  XNOR2_X1 U5416 ( .A(n33278), .B(n3360), .ZN(n32655) );
  CLKBUF_X1 U5417 ( .A(n33277), .Z(n3360) );
  NAND2_X1 U5418 ( .A1(n30809), .A2(n30808), .ZN(n30392) );
  OAI22_X1 U5419 ( .A1(n30417), .A2(n35610), .B1(n33387), .B2(n35611), .ZN(
        n34879) );
  OAI22_X1 U5420 ( .A1(n24112), .A2(n35084), .B1(n33131), .B2(n35083), .ZN(
        n34878) );
  NAND2_X1 U5421 ( .A1(n31857), .A2(n31856), .ZN(n31763) );
  NAND2_X1 U5422 ( .A1(n34971), .A2(n34970), .ZN(n34972) );
  NAND2_X1 U5423 ( .A1(n33348), .A2(n33347), .ZN(n34848) );
  NAND2_X1 U5424 ( .A1(n34693), .A2(n34691), .ZN(n33347) );
  OAI21_X1 U5425 ( .B1(n34693), .B2(n34691), .A(n34692), .ZN(n33348) );
  XNOR2_X1 U5426 ( .A(n33242), .B(n33241), .ZN(n33354) );
  XNOR2_X1 U5427 ( .A(n33240), .B(n33239), .ZN(n33242) );
  NAND2_X1 U5428 ( .A1(n35293), .A2(n35292), .ZN(n35294) );
  XNOR2_X1 U5429 ( .A(n34831), .B(n34830), .ZN(n33330) );
  XNOR2_X1 U5430 ( .A(n34839), .B(n34840), .ZN(n33321) );
  INV_X1 U5431 ( .A(n33233), .ZN(n33333) );
  NOR2_X1 U5432 ( .A1(n34826), .A2(n34825), .ZN(n34828) );
  OAI22_X1 U5433 ( .A1(n33304), .A2(n34195), .B1(n33303), .B2(n34194), .ZN(
        n34927) );
  OAI22_X1 U5434 ( .A1(n33306), .A2(n35749), .B1(n33305), .B2(n35748), .ZN(
        n34926) );
  OAI22_X1 U5435 ( .A1(n33308), .A2(n35709), .B1(n33307), .B2(n35708), .ZN(
        n34925) );
  NOR2_X1 U5436 ( .A1(n35363), .A2(n35362), .ZN(n35365) );
  NOR2_X1 U5437 ( .A1(n31715), .A2(n31716), .ZN(n31718) );
  NAND2_X1 U5438 ( .A1(n31716), .A2(n31715), .ZN(n31717) );
  INV_X1 U5439 ( .A(n34991), .ZN(n35248) );
  AOI21_X1 U5440 ( .B1(n34990), .B2(n34989), .A(n34988), .ZN(n34991) );
  NAND2_X1 U5441 ( .A1(n34906), .A2(n34905), .ZN(n35246) );
  NAND2_X1 U5442 ( .A1(n34904), .A2(n34903), .ZN(n34905) );
  AOI21_X1 U5443 ( .B1(n35041), .B2(n35040), .A(n35039), .ZN(n35042) );
  XNOR2_X1 U5444 ( .A(n32211), .B(\fmem_data[15][7] ), .ZN(n35031) );
  XNOR2_X1 U5445 ( .A(n35030), .B(\fmem_data[15][7] ), .ZN(n35317) );
  XNOR2_X1 U5446 ( .A(n31827), .B(n35132), .ZN(n35170) );
  XNOR2_X1 U5447 ( .A(n35134), .B(n35133), .ZN(n31827) );
  NAND2_X1 U5448 ( .A1(n35186), .A2(n35185), .ZN(n35187) );
  INV_X1 U5449 ( .A(n31836), .ZN(n31840) );
  OAI22_X1 U5450 ( .A1(n34930), .A2(n35512), .B1(n13912), .B2(n35511), .ZN(
        n31835) );
  OAI22_X1 U5451 ( .A1(n34940), .A2(n34942), .B1(n31972), .B2(n34941), .ZN(
        n31834) );
  XNOR2_X1 U5452 ( .A(n35124), .B(n31832), .ZN(n35410) );
  XNOR2_X1 U5453 ( .A(n35126), .B(n35125), .ZN(n31832) );
  XNOR2_X1 U5454 ( .A(n35316), .B(\fmem_data[15][7] ), .ZN(n35695) );
  XNOR2_X1 U5455 ( .A(n31660), .B(\fmem_data[21][7] ), .ZN(n35404) );
  XNOR2_X1 U5456 ( .A(n35023), .B(\fmem_data[5][7] ), .ZN(n35406) );
  XNOR2_X1 U5457 ( .A(n34980), .B(\fmem_data[16][7] ), .ZN(n35398) );
  XNOR2_X1 U5458 ( .A(n33055), .B(\fmem_data[4][7] ), .ZN(n35325) );
  XNOR2_X1 U5459 ( .A(n31996), .B(\fmem_data[8][7] ), .ZN(n35329) );
  XNOR2_X1 U5460 ( .A(n32014), .B(\fmem_data[2][7] ), .ZN(n35337) );
  XNOR2_X1 U5461 ( .A(n35178), .B(\fmem_data[20][7] ), .ZN(n35341) );
  XNOR2_X1 U5462 ( .A(n35021), .B(\fmem_data[9][7] ), .ZN(n35339) );
  NAND2_X1 U5463 ( .A1(n13814), .A2(n35745), .ZN(n35744) );
  XNOR2_X1 U5464 ( .A(n35324), .B(\fmem_data[4][7] ), .ZN(n35747) );
  NAND2_X1 U5465 ( .A1(n11238), .A2(n35739), .ZN(n35740) );
  OAI21_X1 U5466 ( .B1(n35129), .B2(n35128), .A(n35127), .ZN(n35645) );
  NAND2_X1 U5467 ( .A1(n35134), .A2(n35133), .ZN(n35135) );
  OAI22_X1 U5468 ( .A1(n35640), .A2(n35642), .B1(n35243), .B2(n35641), .ZN(
        n35500) );
  OAI22_X1 U5469 ( .A1(n35632), .A2(n35634), .B1(n35239), .B2(n35633), .ZN(
        n35502) );
  OAI22_X1 U5470 ( .A1(n35654), .A2(n35656), .B1(n35271), .B2(n35655), .ZN(
        n35504) );
  NAND2_X1 U5471 ( .A1(n35276), .A2(n35275), .ZN(n35503) );
  NAND2_X1 U5472 ( .A1(n35274), .A2(n35273), .ZN(n35275) );
  AND2_X1 U5473 ( .A1(n17144), .A2(n17143), .ZN(n17145) );
  INV_X1 U5474 ( .A(n28973), .ZN(n3423) );
  AND2_X1 U5475 ( .A1(n14989), .A2(\xmem_data[9][0] ), .ZN(n17194) );
  AND2_X1 U5476 ( .A1(n27339), .A2(n27338), .ZN(n27341) );
  INV_X1 U5477 ( .A(n3327), .ZN(n3301) );
  CLKBUF_X1 U5478 ( .A(n28973), .Z(n17032) );
  NAND2_X1 U5479 ( .A1(n5985), .A2(n10589), .ZN(n5767) );
  INV_X1 U5480 ( .A(n28365), .ZN(n3304) );
  CLKBUF_X1 U5481 ( .A(n28973), .Z(n28365) );
  INV_X1 U5482 ( .A(n30590), .ZN(n3347) );
  CLKBUF_X1 U5483 ( .A(n28973), .Z(n30590) );
  AOI22_X1 U5484 ( .A1(n25724), .A2(\xmem_data[52][0] ), .B1(n31262), .B2(
        \xmem_data[53][0] ), .ZN(n18974) );
  BUF_X2 U5485 ( .A(n14937), .Z(n25573) );
  NAND2_X1 U5486 ( .A1(n10589), .A2(load_xaddr_val[5]), .ZN(n13429) );
  INV_X1 U5487 ( .A(n29567), .ZN(n3343) );
  CLKBUF_X1 U5488 ( .A(n14991), .Z(n29567) );
  INV_X1 U5489 ( .A(n28745), .ZN(n28746) );
  INV_X1 U5490 ( .A(n28742), .ZN(n28747) );
  CLKBUF_X1 U5491 ( .A(n8020), .Z(n3444) );
  INV_X1 U5492 ( .A(n31263), .ZN(n3379) );
  AND3_X1 U5493 ( .A1(n27782), .A2(n27781), .A3(n27780), .ZN(n27783) );
  NAND3_X1 U5494 ( .A1(n21369), .A2(n21368), .A3(n21367), .ZN(n21370) );
  NOR2_X1 U5495 ( .A1(n5360), .A2(n5359), .ZN(n29002) );
  NAND2_X1 U5496 ( .A1(n21286), .A2(n21285), .ZN(n21292) );
  INV_X1 U5497 ( .A(n21295), .ZN(n21296) );
  INV_X1 U5498 ( .A(n3349), .ZN(n3351) );
  OR2_X1 U5499 ( .A1(n17431), .A2(n17430), .ZN(n17432) );
  OR2_X1 U5500 ( .A1(n27148), .A2(n27147), .ZN(n27149) );
  NOR2_X1 U5501 ( .A1(n27205), .A2(n27204), .ZN(n27207) );
  NOR2_X1 U5502 ( .A1(n27172), .A2(n27171), .ZN(n27182) );
  NOR2_X1 U5503 ( .A1(n27118), .A2(n27117), .ZN(n27128) );
  OR3_X1 U5504 ( .A1(n26613), .A2(n26612), .A3(n26611), .ZN(n26614) );
  OR3_X1 U5505 ( .A1(n26681), .A2(n26680), .A3(n26679), .ZN(n26682) );
  AND2_X1 U5506 ( .A1(n27084), .A2(n27083), .ZN(n27085) );
  AOI21_X1 U5507 ( .B1(n19354), .B2(n19410), .A(n19353), .ZN(n19415) );
  AND4_X1 U5508 ( .A1(n30255), .A2(n30254), .A3(n30253), .A4(n30252), .ZN(
        n30277) );
  OR2_X1 U5509 ( .A1(n17783), .A2(n17782), .ZN(n17784) );
  NAND2_X1 U5510 ( .A1(n17781), .A2(n17780), .ZN(n17782) );
  OR2_X1 U5511 ( .A1(n20417), .A2(n3232), .ZN(n20487) );
  NAND3_X1 U5512 ( .A1(n3713), .A2(n21986), .A3(n21985), .ZN(n21998) );
  NAND3_X1 U5513 ( .A1(n29206), .A2(n29205), .A3(n29204), .ZN(n32078) );
  NAND2_X1 U5514 ( .A1(n29172), .A2(n29171), .ZN(n29205) );
  OAI22_X1 U5515 ( .A1(n36106), .A2(n36104), .B1(n32941), .B2(n3580), .ZN(
        n36304) );
  XNOR2_X1 U5516 ( .A(n32528), .B(\fmem_data[29][1] ), .ZN(n32928) );
  XNOR2_X1 U5517 ( .A(n33556), .B(\fmem_data[16][3] ), .ZN(n34502) );
  XNOR2_X1 U5518 ( .A(n36299), .B(\fmem_data[16][3] ), .ZN(n34500) );
  XNOR2_X1 U5519 ( .A(n36228), .B(\fmem_data[20][3] ), .ZN(n34496) );
  OR2_X1 U5520 ( .A1(n33174), .A2(n3610), .ZN(n32552) );
  OAI22_X1 U5521 ( .A1(n32790), .A2(n33568), .B1(n33570), .B2(n3641), .ZN(
        n34768) );
  OAI22_X1 U5522 ( .A1(n32789), .A2(n34431), .B1(n34433), .B2(n3605), .ZN(
        n34769) );
  OAI22_X1 U5523 ( .A1(n32778), .A2(n33059), .B1(n33057), .B2(n3634), .ZN(
        n34767) );
  OAI22_X1 U5524 ( .A1(n32781), .A2(n32780), .B1(n32779), .B2(n3658), .ZN(
        n34766) );
  XNOR2_X1 U5525 ( .A(n32025), .B(\fmem_data[12][1] ), .ZN(n33781) );
  AND2_X1 U5526 ( .A1(n36111), .A2(n31498), .ZN(n33471) );
  OAI22_X1 U5527 ( .A1(n33649), .A2(n3569), .B1(n32980), .B2(n34598), .ZN(
        n33485) );
  AND2_X1 U5528 ( .A1(n36200), .A2(n33723), .ZN(n34606) );
  OAI22_X1 U5529 ( .A1(n32690), .A2(n33174), .B1(n31494), .B2(n33176), .ZN(
        n33717) );
  OAI22_X1 U5530 ( .A1(n34441), .A2(n3483), .B1(n34440), .B2(n31500), .ZN(
        n33719) );
  OAI22_X1 U5531 ( .A1(n33591), .A2(n33690), .B1(n33590), .B2(n34736), .ZN(
        n33716) );
  OAI22_X1 U5532 ( .A1(n34337), .A2(n34472), .B1(n34474), .B2(n3686), .ZN(
        n34631) );
  OAI22_X1 U5533 ( .A1(n34336), .A2(n34412), .B1(n34410), .B2(n3674), .ZN(
        n34632) );
  NAND2_X1 U5534 ( .A1(n33839), .A2(n33838), .ZN(n34640) );
  NAND2_X1 U5535 ( .A1(n33837), .A2(n33836), .ZN(n33838) );
  XNOR2_X1 U5536 ( .A(n3390), .B(\fmem_data[10][1] ), .ZN(n33601) );
  XNOR2_X1 U5537 ( .A(n32882), .B(\fmem_data[6][3] ), .ZN(n33599) );
  OAI22_X1 U5538 ( .A1(n31242), .A2(n34944), .B1(n34945), .B2(n3488), .ZN(
        n31566) );
  OAI22_X1 U5539 ( .A1(n31397), .A2(n34903), .B1(n34904), .B2(n3636), .ZN(
        n31572) );
  OAI22_X1 U5540 ( .A1(n31198), .A2(n34909), .B1(n34908), .B2(n3687), .ZN(
        n31516) );
  OAI22_X1 U5541 ( .A1(n33895), .A2(n34420), .B1(n34421), .B2(n34418), .ZN(
        n31517) );
  NAND2_X1 U5542 ( .A1(n36306), .A2(n36305), .ZN(n32942) );
  OAI22_X1 U5543 ( .A1(n32783), .A2(n33875), .B1(n31394), .B2(n33873), .ZN(
        n31531) );
  OAI22_X1 U5544 ( .A1(n31396), .A2(n34922), .B1(n31395), .B2(n34923), .ZN(
        n31576) );
  OAI22_X1 U5545 ( .A1(n31245), .A2(n34919), .B1(n34918), .B2(n3688), .ZN(
        n31612) );
  OAI22_X1 U5546 ( .A1(n33878), .A2(n3647), .B1(n31446), .B2(n36227), .ZN(
        n31917) );
  OAI22_X1 U5547 ( .A1(n31912), .A2(n35089), .B1(n35088), .B2(n3595), .ZN(
        n32487) );
  OAI22_X1 U5548 ( .A1(n32075), .A2(n33963), .B1(n33961), .B2(n3591), .ZN(
        n32210) );
  OAI22_X1 U5549 ( .A1(n32081), .A2(n33961), .B1(n32080), .B2(n33963), .ZN(
        n32208) );
  NAND2_X1 U5550 ( .A1(n32967), .A2(n32966), .ZN(n32062) );
  OAI22_X1 U5551 ( .A1(n32069), .A2(n33250), .B1(n32068), .B2(n33249), .ZN(
        n32933) );
  XNOR2_X1 U5552 ( .A(n32869), .B(n32868), .ZN(n36172) );
  XNOR2_X1 U5553 ( .A(n32867), .B(n32866), .ZN(n32868) );
  OAI22_X1 U5554 ( .A1(n33593), .A2(n34739), .B1(n32601), .B2(n3563), .ZN(
        n34525) );
  OAI22_X1 U5555 ( .A1(n32599), .A2(n36298), .B1(n34025), .B2(n3573), .ZN(
        n34526) );
  XNOR2_X1 U5556 ( .A(n32794), .B(n32793), .ZN(n34720) );
  XNOR2_X1 U5557 ( .A(n32792), .B(n32791), .ZN(n32794) );
  OAI22_X1 U5558 ( .A1(n32130), .A2(n35003), .B1(n32129), .B2(n35004), .ZN(
        n32795) );
  OAI22_X1 U5559 ( .A1(n32128), .A2(n34497), .B1(n32418), .B2(n34495), .ZN(
        n32796) );
  OAI22_X1 U5560 ( .A1(n32136), .A2(n33973), .B1(n32135), .B2(n33975), .ZN(
        n32801) );
  OAI22_X1 U5561 ( .A1(n32134), .A2(n33250), .B1(n32133), .B2(n33249), .ZN(
        n32802) );
  OAI22_X1 U5562 ( .A1(n32132), .A2(n33174), .B1(n32689), .B2(n33176), .ZN(
        n32803) );
  OAI22_X1 U5563 ( .A1(n32583), .A2(n3561), .B1(n33600), .B2(n36114), .ZN(
        n32622) );
  OAI22_X1 U5564 ( .A1(n32245), .A2(n33105), .B1(n33103), .B2(n3597), .ZN(
        n32625) );
  OAI22_X1 U5565 ( .A1(n32244), .A2(n33328), .B1(n33326), .B2(n3596), .ZN(
        n32626) );
  NAND2_X1 U5566 ( .A1(n36172), .A2(n36171), .ZN(n32876) );
  NAND2_X1 U5567 ( .A1(n36778), .A2(n36777), .ZN(n36230) );
  OAI22_X1 U5568 ( .A1(n32594), .A2(n34779), .B1(n34465), .B2(n34466), .ZN(
        n34732) );
  OAI22_X1 U5569 ( .A1(n33682), .A2(n33679), .B1(n33645), .B2(n33681), .ZN(
        n34730) );
  NAND2_X1 U5570 ( .A1(n32123), .A2(n32122), .ZN(n32683) );
  OAI22_X1 U5571 ( .A1(n32125), .A2(n34414), .B1(n34415), .B2(n34416), .ZN(
        n32682) );
  OAI22_X1 U5572 ( .A1(n32690), .A2(n33176), .B1(n32689), .B2(n33174), .ZN(
        n34728) );
  OAI22_X1 U5573 ( .A1(n32239), .A2(n33975), .B1(n33973), .B2(n3589), .ZN(
        n32695) );
  OAI22_X1 U5574 ( .A1(n32238), .A2(n3563), .B1(n32601), .B2(n34739), .ZN(
        n32696) );
  OAI22_X1 U5575 ( .A1(n32565), .A2(n33326), .B1(n32564), .B2(n33328), .ZN(
        n32746) );
  OAI22_X1 U5576 ( .A1(n32563), .A2(n33642), .B1(n32562), .B2(n33643), .ZN(
        n32747) );
  OAI22_X1 U5577 ( .A1(n32651), .A2(n35615), .B1(n32650), .B2(n35614), .ZN(
        n32750) );
  OAI21_X1 U5578 ( .B1(n32827), .B2(n32825), .A(n32826), .ZN(n32593) );
  NAND2_X1 U5579 ( .A1(n32827), .A2(n32825), .ZN(n32592) );
  OAI22_X1 U5580 ( .A1(n32106), .A2(n35656), .B1(n35655), .B2(n3640), .ZN(
        n32316) );
  OAI22_X1 U5581 ( .A1(n32140), .A2(n35642), .B1(n35641), .B2(n3698), .ZN(
        n32630) );
  OAI22_X1 U5582 ( .A1(n32139), .A2(n35041), .B1(n32227), .B2(n35040), .ZN(
        n32631) );
  OAI22_X1 U5583 ( .A1(n32155), .A2(n35652), .B1(n35651), .B2(n3668), .ZN(
        n32249) );
  OAI22_X1 U5584 ( .A1(n32152), .A2(n3633), .B1(n32151), .B2(n36226), .ZN(
        n32251) );
  OAI22_X1 U5585 ( .A1(n32527), .A2(n34343), .B1(n30982), .B2(n3578), .ZN(
        n31120) );
  OAI22_X1 U5586 ( .A1(n32525), .A2(n34745), .B1(n30981), .B2(n3562), .ZN(
        n31121) );
  AND2_X1 U5587 ( .A1(n36312), .A2(n30979), .ZN(n31138) );
  OAI22_X1 U5588 ( .A1(n32581), .A2(n33827), .B1(n30980), .B2(n33828), .ZN(
        n31137) );
  NAND2_X1 U5589 ( .A1(n32495), .A2(n32492), .ZN(n31176) );
  XNOR2_X1 U5590 ( .A(n30832), .B(n31736), .ZN(n30999) );
  XNOR2_X1 U5591 ( .A(n31009), .B(n31008), .ZN(n31871) );
  XNOR2_X1 U5592 ( .A(n31007), .B(n31006), .ZN(n31008) );
  OAI22_X1 U5593 ( .A1(n30819), .A2(n35003), .B1(n30818), .B2(n35004), .ZN(
        n31876) );
  OAI22_X1 U5594 ( .A1(n32572), .A2(n33690), .B1(n30817), .B2(n34736), .ZN(
        n31116) );
  OAI22_X1 U5595 ( .A1(n32587), .A2(n34734), .B1(n30816), .B2(n3572), .ZN(
        n31117) );
  OAI22_X1 U5596 ( .A1(n31888), .A2(n35753), .B1(n31887), .B2(n35752), .ZN(
        n32159) );
  OAI22_X1 U5597 ( .A1(n31881), .A2(n33596), .B1(n31880), .B2(n33598), .ZN(
        n32161) );
  XNOR2_X1 U5598 ( .A(n36299), .B(\fmem_data[16][7] ), .ZN(n31887) );
  OAI22_X1 U5599 ( .A1(n32757), .A2(n35508), .B1(n20613), .B2(n35507), .ZN(
        n26268) );
  OAI22_X1 U5600 ( .A1(n31888), .A2(n35752), .B1(n17851), .B2(n35753), .ZN(
        n23581) );
  NOR2_X1 U5601 ( .A1(n17753), .A2(\fmem_data[27][0] ), .ZN(n17754) );
  OAI22_X1 U5602 ( .A1(n32002), .A2(n35512), .B1(n19024), .B2(n35511), .ZN(
        n23589) );
  OAI22_X1 U5603 ( .A1(n31968), .A2(n3576), .B1(n31886), .B2(n34483), .ZN(
        n23591) );
  NAND2_X1 U5604 ( .A1(n23577), .A2(n23574), .ZN(n19304) );
  OAI22_X1 U5605 ( .A1(n31949), .A2(n34736), .B1(n30817), .B2(n33690), .ZN(
        n23166) );
  OAI22_X1 U5606 ( .A1(n30828), .A2(n3572), .B1(n30816), .B2(n34734), .ZN(
        n23168) );
  NOR2_X1 U5607 ( .A1(n16357), .A2(n3489), .ZN(n16358) );
  INV_X1 U5608 ( .A(n36216), .ZN(n16357) );
  AOI21_X1 U5609 ( .B1(n36241), .B2(n3662), .A(n32191), .ZN(n17745) );
  NOR2_X1 U5610 ( .A1(n22358), .A2(\fmem_data[3][0] ), .ZN(n22359) );
  INV_X1 U5611 ( .A(n36199), .ZN(n22358) );
  INV_X1 U5612 ( .A(n22360), .ZN(n29520) );
  OAI22_X1 U5613 ( .A1(n33181), .A2(n33850), .B1(n32229), .B2(n33851), .ZN(
        n29527) );
  XNOR2_X1 U5614 ( .A(n31391), .B(n31390), .ZN(n31393) );
  OAI22_X1 U5615 ( .A1(n27581), .A2(n35490), .B1(n35489), .B2(n3599), .ZN(
        n28936) );
  OAI22_X1 U5616 ( .A1(n32202), .A2(n33098), .B1(n32733), .B2(n33100), .ZN(
        n31140) );
  NAND2_X1 U5617 ( .A1(n6484), .A2(n33741), .ZN(n33603) );
  NAND2_X1 U5618 ( .A1(n15885), .A2(n34505), .ZN(n34503) );
  OAI22_X1 U5619 ( .A1(n28402), .A2(n35592), .B1(n35591), .B2(n3613), .ZN(
        n29845) );
  OAI22_X1 U5620 ( .A1(n28401), .A2(n35705), .B1(n35704), .B2(n3639), .ZN(
        n29846) );
  XNOR2_X1 U5621 ( .A(n31669), .B(\fmem_data[13][3] ), .ZN(n31964) );
  XNOR2_X1 U5622 ( .A(n35104), .B(\fmem_data[13][3] ), .ZN(n33052) );
  XNOR2_X1 U5623 ( .A(n32321), .B(\fmem_data[17][7] ), .ZN(n24431) );
  OAI22_X1 U5624 ( .A1(n32183), .A2(n34922), .B1(n22454), .B2(n34923), .ZN(
        n28908) );
  OAI22_X1 U5625 ( .A1(n30819), .A2(n35004), .B1(n24015), .B2(n35003), .ZN(
        n28912) );
  AOI21_X1 U5626 ( .B1(n36196), .B2(n3577), .A(n32112), .ZN(n22642) );
  OAI22_X1 U5627 ( .A1(n32734), .A2(n33098), .B1(n30415), .B2(n33100), .ZN(
        n30840) );
  OAI22_X1 U5628 ( .A1(n34425), .A2(n34424), .B1(n34423), .B2(n34422), .ZN(
        n34512) );
  OAI22_X1 U5629 ( .A1(n34438), .A2(n34437), .B1(n34436), .B2(n34435), .ZN(
        n34523) );
  OAI22_X1 U5630 ( .A1(n34434), .A2(n34433), .B1(n34432), .B2(n34431), .ZN(
        n34524) );
  NAND2_X1 U5631 ( .A1(n33822), .A2(n33821), .ZN(n33823) );
  NAND2_X1 U5632 ( .A1(n31440), .A2(n31439), .ZN(n31223) );
  NAND2_X1 U5633 ( .A1(n34332), .A2(n34330), .ZN(n33884) );
  NAND2_X1 U5634 ( .A1(n34568), .A2(n34569), .ZN(n33863) );
  OAI22_X1 U5635 ( .A1(n34018), .A2(n3559), .B1(n33811), .B2(n34017), .ZN(
        n33586) );
  OAI22_X1 U5636 ( .A1(n32565), .A2(n33328), .B1(n28409), .B2(n33326), .ZN(
        n33585) );
  XNOR2_X1 U5637 ( .A(n36299), .B(\fmem_data[16][5] ), .ZN(n28409) );
  XNOR2_X1 U5638 ( .A(n28536), .B(n28535), .ZN(n28538) );
  OAI22_X1 U5639 ( .A1(n31987), .A2(n35036), .B1(n32522), .B2(n35037), .ZN(
        n23187) );
  OAI22_X1 U5640 ( .A1(n31126), .A2(n36295), .B1(n23573), .B2(n3564), .ZN(
        n28901) );
  NAND2_X1 U5641 ( .A1(n33665), .A2(n33663), .ZN(n33653) );
  OAI21_X1 U5642 ( .B1(n33665), .B2(n33663), .A(n33664), .ZN(n33654) );
  NAND2_X1 U5643 ( .A1(n33632), .A2(n33631), .ZN(n33633) );
  NAND2_X1 U5644 ( .A1(n33893), .A2(n33892), .ZN(n34091) );
  OAI22_X1 U5645 ( .A1(n33186), .A2(n35084), .B1(n33185), .B2(n35083), .ZN(
        n33191) );
  OAI22_X1 U5646 ( .A1(n33181), .A2(n33851), .B1(n33180), .B2(n33850), .ZN(
        n33260) );
  OAI22_X1 U5647 ( .A1(n34209), .A2(n34208), .B1(n34207), .B2(n34206), .ZN(
        n34401) );
  OAI22_X1 U5648 ( .A1(n32734), .A2(n33100), .B1(n32733), .B2(n33098), .ZN(
        n33205) );
  NAND2_X1 U5649 ( .A1(n34264), .A2(n34263), .ZN(n34265) );
  OAI22_X1 U5650 ( .A1(n32751), .A2(n34363), .B1(n33169), .B2(n34364), .ZN(
        n33157) );
  NAND2_X1 U5651 ( .A1(n32792), .A2(n32791), .ZN(n32537) );
  XNOR2_X1 U5652 ( .A(n32358), .B(n32357), .ZN(n32359) );
  NAND2_X1 U5653 ( .A1(n32500), .A2(n32499), .ZN(n31199) );
  XNOR2_X1 U5654 ( .A(n30140), .B(n30139), .ZN(n30376) );
  XNOR2_X1 U5655 ( .A(n30138), .B(n3618), .ZN(n30140) );
  NAND2_X1 U5656 ( .A1(n33090), .A2(n33089), .ZN(n33091) );
  NAND2_X1 U5657 ( .A1(n35157), .A2(n35156), .ZN(n35204) );
  NAND2_X1 U5658 ( .A1(n11670), .A2(n35701), .ZN(n35700) );
  AOI21_X1 U5659 ( .B1(n35697), .B2(n35696), .A(n35695), .ZN(n35698) );
  OAI22_X1 U5660 ( .A1(n35609), .A2(n35611), .B1(n35356), .B2(n35610), .ZN(
        n35737) );
  OAI22_X1 U5661 ( .A1(n35613), .A2(n35615), .B1(n35358), .B2(n35614), .ZN(
        n35736) );
  OAI22_X1 U5662 ( .A1(n35583), .A2(n35585), .B1(n35176), .B2(n35584), .ZN(
        n35716) );
  OAI22_X1 U5663 ( .A1(n35579), .A2(n35581), .B1(n35075), .B2(n35580), .ZN(
        n35715) );
  OAI22_X1 U5664 ( .A1(n35590), .A2(n35592), .B1(n35105), .B2(n35591), .ZN(
        n35718) );
  OAI22_X1 U5665 ( .A1(n35575), .A2(n35577), .B1(n35103), .B2(n35576), .ZN(
        n35719) );
  AOI21_X1 U5666 ( .B1(n35634), .B2(n35633), .A(n35632), .ZN(n35635) );
  AOI21_X1 U5667 ( .B1(n35638), .B2(n35637), .A(n35636), .ZN(n35639) );
  AOI21_X1 U5668 ( .B1(n35642), .B2(n35641), .A(n35640), .ZN(n35643) );
  AOI21_X1 U5669 ( .B1(n35615), .B2(n35614), .A(n35613), .ZN(n35616) );
  AOI21_X1 U5670 ( .B1(n35611), .B2(n35610), .A(n35609), .ZN(n35612) );
  NAND2_X1 U5671 ( .A1(n6701), .A2(n35722), .ZN(n35721) );
  XNOR2_X1 U5672 ( .A(n35338), .B(\fmem_data[9][7] ), .ZN(n35724) );
  NAND2_X1 U5673 ( .A1(n5455), .A2(n35726), .ZN(n35725) );
  NAND2_X1 U5674 ( .A1(n17743), .A2(n35730), .ZN(n35729) );
  AOI21_X1 U5675 ( .B1(n35577), .B2(n35576), .A(n35575), .ZN(n35578) );
  AOI21_X1 U5676 ( .B1(n35581), .B2(n35580), .A(n35579), .ZN(n35582) );
  AOI21_X1 U5677 ( .B1(n35585), .B2(n35584), .A(n35583), .ZN(n35586) );
  AOI21_X1 U5678 ( .B1(n35753), .B2(n35752), .A(n35751), .ZN(n35754) );
  AOI21_X1 U5679 ( .B1(n35761), .B2(n35760), .A(n35759), .ZN(n35762) );
  NAND3_X1 U5680 ( .A1(n17007), .A2(n17006), .A3(n17005), .ZN(n17008) );
  INV_X1 U5681 ( .A(n3423), .ZN(n3424) );
  OR2_X1 U5682 ( .A1(n20896), .A2(n20895), .ZN(n20912) );
  OR3_X1 U5683 ( .A1(n20882), .A2(n20881), .A3(n20880), .ZN(n20883) );
  OR3_X1 U5684 ( .A1(n20860), .A2(n20859), .A3(n20858), .ZN(n20861) );
  NOR2_X1 U5685 ( .A1(n27348), .A2(n3739), .ZN(n27349) );
  AND2_X1 U5686 ( .A1(n8924), .A2(n8923), .ZN(n30626) );
  AND2_X1 U5687 ( .A1(n4129), .A2(n4130), .ZN(n25741) );
  NAND2_X1 U5688 ( .A1(n13431), .A2(n13430), .ZN(n13467) );
  NAND2_X1 U5689 ( .A1(n13429), .A2(load_xaddr_val[6]), .ZN(n13430) );
  NAND2_X1 U5690 ( .A1(n6488), .A2(n10589), .ZN(n6491) );
  INV_X1 U5691 ( .A(n27584), .ZN(n27589) );
  NOR2_X1 U5692 ( .A1(n11383), .A2(n3941), .ZN(n11467) );
  INV_X2 U5693 ( .A(n3343), .ZN(n3345) );
  NAND2_X1 U5694 ( .A1(n27650), .A2(n27649), .ZN(n27651) );
  INV_X1 U5695 ( .A(n27640), .ZN(n27645) );
  NAND3_X1 U5696 ( .A1(n28775), .A2(n28774), .A3(n28773), .ZN(n28776) );
  NAND3_X1 U5697 ( .A1(n28723), .A2(n28722), .A3(n28721), .ZN(n28731) );
  INV_X1 U5698 ( .A(n30848), .ZN(n30860) );
  AND2_X1 U5699 ( .A1(n10135), .A2(n10162), .ZN(n30918) );
  NOR2_X1 U5700 ( .A1(n3913), .A2(n27727), .ZN(n27735) );
  NOR2_X1 U5701 ( .A1(n19697), .A2(n3742), .ZN(n19698) );
  OR2_X1 U5702 ( .A1(n21362), .A2(n21361), .ZN(n21363) );
  OR2_X1 U5703 ( .A1(n21352), .A2(n21351), .ZN(n21364) );
  OR2_X1 U5704 ( .A1(n3961), .A2(n21335), .ZN(n21336) );
  OR2_X1 U5705 ( .A1(n17450), .A2(n17449), .ZN(n17456) );
  OR3_X1 U5706 ( .A1(n17410), .A2(n17409), .A3(n17408), .ZN(n17411) );
  NAND2_X1 U5707 ( .A1(n22999), .A2(n29376), .ZN(n23074) );
  NOR2_X1 U5708 ( .A1(n6890), .A2(n6867), .ZN(n28324) );
  OR2_X1 U5709 ( .A1(n34624), .A2(n3671), .ZN(n33469) );
  OAI21_X1 U5710 ( .B1(n34615), .B2(n3999), .A(n34613), .ZN(n34616) );
  AND2_X1 U5711 ( .A1(n36203), .A2(n36201), .ZN(n34618) );
  XNOR2_X1 U5712 ( .A(n32979), .B(\fmem_data[4][1] ), .ZN(n34600) );
  NAND2_X1 U5713 ( .A1(\fmem_data[4][1] ), .A2(n3569), .ZN(n34598) );
  NAND3_X1 U5714 ( .A1(n34588), .A2(n34589), .A3(n3693), .ZN(n34593) );
  OR2_X1 U5715 ( .A1(n36244), .A2(n3675), .ZN(n34594) );
  NAND2_X1 U5716 ( .A1(\fmem_data[22][1] ), .A2(n3567), .ZN(n34777) );
  OR3_X1 U5717 ( .A1(n20537), .A2(n20536), .A3(n20535), .ZN(n20539) );
  OR3_X1 U5718 ( .A1(n20566), .A2(n20565), .A3(n20564), .ZN(n20575) );
  OR3_X1 U5719 ( .A1(n20514), .A2(n20513), .A3(n20512), .ZN(n20516) );
  OR3_X1 U5720 ( .A1(n22692), .A2(n22691), .A3(n22690), .ZN(n22700) );
  OR2_X1 U5721 ( .A1(n36105), .A2(n3690), .ZN(n32955) );
  NAND2_X1 U5722 ( .A1(\fmem_data[6][1] ), .A2(n3559), .ZN(n34017) );
  AND2_X1 U5723 ( .A1(n36338), .A2(n34780), .ZN(n36247) );
  OAI22_X1 U5724 ( .A1(n34538), .A2(n34537), .B1(n34536), .B2(n34535), .ZN(
        n36108) );
  OAI22_X1 U5725 ( .A1(n33702), .A2(n3931), .B1(n33701), .B2(n36216), .ZN(
        n33739) );
  OAI22_X1 U5726 ( .A1(n33700), .A2(n3581), .B1(n33699), .B2(n36218), .ZN(
        n33738) );
  OAI22_X1 U5727 ( .A1(n33736), .A2(n3482), .B1(n33735), .B2(n36240), .ZN(
        n33814) );
  OAI22_X1 U5728 ( .A1(n33748), .A2(n3574), .B1(n33747), .B2(n34625), .ZN(
        n34347) );
  OAI22_X1 U5729 ( .A1(n33746), .A2(n34779), .B1(n34466), .B2(n3590), .ZN(
        n34348) );
  OR2_X1 U5730 ( .A1(n36338), .A2(n3590), .ZN(n33746) );
  OAI22_X1 U5731 ( .A1(n34365), .A2(n34364), .B1(n34363), .B2(n3609), .ZN(
        n36091) );
  OAI22_X1 U5732 ( .A1(n34464), .A2(n34463), .B1(n34462), .B2(n3643), .ZN(
        n36087) );
  OAI22_X1 U5733 ( .A1(n34471), .A2(n34470), .B1(n34469), .B2(n34468), .ZN(
        n36085) );
  OAI22_X1 U5734 ( .A1(n34467), .A2(n34466), .B1(n34465), .B2(n34779), .ZN(
        n36086) );
  OAI22_X1 U5735 ( .A1(n34338), .A2(n34470), .B1(n34468), .B2(n3485), .ZN(
        n36090) );
  OAI22_X1 U5736 ( .A1(n34346), .A2(n3633), .B1(n34345), .B2(n36226), .ZN(
        n36088) );
  OAI22_X1 U5737 ( .A1(n34743), .A2(n34742), .B1(n34741), .B2(n3571), .ZN(
        n36099) );
  AND2_X1 U5738 ( .A1(n36312), .A2(n34737), .ZN(n36095) );
  NAND2_X1 U5739 ( .A1(n36205), .A2(n36204), .ZN(n32885) );
  OAI22_X1 U5740 ( .A1(n32071), .A2(n3562), .B1(n34744), .B2(n34745), .ZN(
        n32985) );
  OAI22_X1 U5741 ( .A1(n32070), .A2(n33570), .B1(n33568), .B2(n33571), .ZN(
        n32986) );
  OAI22_X1 U5742 ( .A1(n33574), .A2(n33855), .B1(n32072), .B2(n33853), .ZN(
        n32984) );
  XNOR2_X1 U5743 ( .A(n31542), .B(n31541), .ZN(n33493) );
  AND2_X1 U5744 ( .A1(n34480), .A2(n34479), .ZN(n31542) );
  OAI22_X1 U5745 ( .A1(n33834), .A2(n3566), .B1(n34528), .B2(n34529), .ZN(
        n33545) );
  OAI22_X1 U5746 ( .A1(n32599), .A2(n3573), .B1(n33557), .B2(n36298), .ZN(
        n33546) );
  OAI22_X1 U5747 ( .A1(n36223), .A2(n33480), .B1(n32598), .B2(n3568), .ZN(
        n33544) );
  OAI21_X1 U5748 ( .B1(n33760), .B2(n33759), .A(n33758), .ZN(n36488) );
  NAND2_X1 U5749 ( .A1(n36479), .A2(n36478), .ZN(n33758) );
  NOR2_X1 U5750 ( .A1(n36479), .A2(n36478), .ZN(n33760) );
  OAI22_X1 U5751 ( .A1(n34403), .A2(n3568), .B1(n34402), .B2(n36223), .ZN(
        n34494) );
  NAND2_X1 U5752 ( .A1(n32995), .A2(n32992), .ZN(n31560) );
  NAND2_X1 U5753 ( .A1(n36289), .A2(n36288), .ZN(n32969) );
  NOR2_X1 U5754 ( .A1(n36403), .A2(n36402), .ZN(n33474) );
  AOI21_X1 U5755 ( .B1(n36402), .B2(n36403), .A(n36404), .ZN(n33475) );
  OAI22_X1 U5756 ( .A1(n33804), .A2(n34433), .B1(n32716), .B2(n34431), .ZN(
        n32670) );
  XNOR2_X1 U5757 ( .A(n32411), .B(n32410), .ZN(n32412) );
  NAND2_X1 U5758 ( .A1(n34762), .A2(n34761), .ZN(n32449) );
  NAND2_X1 U5759 ( .A1(n32705), .A2(n32703), .ZN(n32215) );
  XNOR2_X1 U5760 ( .A(n34375), .B(n34374), .ZN(n34554) );
  NAND2_X1 U5761 ( .A1(n27700), .A2(n27699), .ZN(n31208) );
  NAND2_X1 U5762 ( .A1(n31129), .A2(n31127), .ZN(n27699) );
  OAI21_X1 U5763 ( .B1(n31129), .B2(n31127), .A(n31128), .ZN(n27700) );
  NAND2_X1 U5764 ( .A1(n36071), .A2(n36070), .ZN(n34542) );
  NAND2_X1 U5765 ( .A1(n36734), .A2(n36737), .ZN(n36417) );
  NAND2_X1 U5766 ( .A1(n36490), .A2(n36492), .ZN(n33605) );
  NAND2_X1 U5767 ( .A1(n36456), .A2(n36455), .ZN(n33775) );
  NAND2_X1 U5768 ( .A1(n36393), .A2(n36392), .ZN(n33516) );
  NAND2_X1 U5769 ( .A1(n34808), .A2(n34806), .ZN(n32708) );
  NAND2_X1 U5770 ( .A1(n34896), .A2(n34895), .ZN(n34897) );
  NAND2_X1 U5771 ( .A1(n35377), .A2(n35376), .ZN(n35537) );
  NAND2_X1 U5772 ( .A1(n35565), .A2(n35564), .ZN(n35833) );
  NAND2_X1 U5773 ( .A1(n35571), .A2(n35570), .ZN(n35832) );
  NAND2_X1 U5774 ( .A1(n35563), .A2(n35562), .ZN(n35564) );
  AOI21_X1 U5775 ( .B1(n35656), .B2(n35655), .A(n35654), .ZN(n35657) );
  AOI21_X1 U5776 ( .B1(n35663), .B2(n35662), .A(n35661), .ZN(n35664) );
  AOI21_X1 U5777 ( .B1(n35726), .B2(n35725), .A(n35724), .ZN(n35727) );
  AOI21_X1 U5778 ( .B1(n35730), .B2(n35729), .A(n35728), .ZN(n35731) );
  INV_X1 U5779 ( .A(n35517), .ZN(n35822) );
  INV_X1 U5780 ( .A(n35509), .ZN(n35824) );
  INV_X1 U5781 ( .A(n35513), .ZN(n35823) );
  AOI21_X1 U5782 ( .B1(n35592), .B2(n35591), .A(n35590), .ZN(n35593) );
  INV_X1 U5783 ( .A(n35499), .ZN(n35810) );
  INV_X1 U5784 ( .A(n35491), .ZN(n35812) );
  INV_X1 U5785 ( .A(n35495), .ZN(n35811) );
  OR2_X1 U5786 ( .A1(n17115), .A2(n17114), .ZN(n3987) );
  NAND4_X1 U5787 ( .A1(n17113), .A2(n17112), .A3(n17111), .A4(n17110), .ZN(
        n17114) );
  NAND2_X1 U5788 ( .A1(n19111), .A2(n19110), .ZN(n19112) );
  OR2_X1 U5789 ( .A1(n17700), .A2(n17699), .ZN(n17717) );
  OR2_X1 U5790 ( .A1(n17682), .A2(n17681), .ZN(n17694) );
  AND4_X1 U5791 ( .A1(n26424), .A2(n26423), .A3(n26422), .A4(n26421), .ZN(
        n26426) );
  OR4_X1 U5792 ( .A1(n17504), .A2(n17503), .A3(n17502), .A4(n17501), .ZN(
        n17505) );
  OR2_X1 U5793 ( .A1(n17549), .A2(n3958), .ZN(n17550) );
  AND2_X1 U5794 ( .A1(n13496), .A2(n13497), .ZN(n24508) );
  OR2_X1 U5795 ( .A1(n21556), .A2(n3957), .ZN(n21557) );
  OR2_X1 U5796 ( .A1(n21760), .A2(n3960), .ZN(n21761) );
  AND2_X1 U5797 ( .A1(n4571), .A2(n4525), .ZN(n28071) );
  OR2_X1 U5798 ( .A1(n27687), .A2(n27686), .ZN(n27693) );
  AND3_X1 U5799 ( .A1(n28699), .A2(n28698), .A3(n28697), .ZN(n28710) );
  AND2_X1 U5800 ( .A1(n28637), .A2(n28636), .ZN(n28651) );
  NOR2_X1 U5801 ( .A1(n8067), .A2(n8066), .ZN(n28794) );
  AND2_X1 U5802 ( .A1(n27827), .A2(n27826), .ZN(n27828) );
  NOR2_X1 U5803 ( .A1(n7471), .A2(n7470), .ZN(n27839) );
  AND2_X1 U5804 ( .A1(n7470), .A2(n7471), .ZN(n27737) );
  NOR2_X1 U5805 ( .A1(n7471), .A2(n7469), .ZN(n27778) );
  AND4_X1 U5806 ( .A1(n29367), .A2(n29366), .A3(n29365), .A4(n29364), .ZN(
        n29368) );
  NOR2_X1 U5807 ( .A1(n7292), .A2(n7291), .ZN(n29511) );
  NOR2_X1 U5808 ( .A1(n28189), .A2(n28188), .ZN(n28205) );
  NOR2_X1 U5809 ( .A1(n7619), .A2(n7618), .ZN(n29758) );
  AND4_X1 U5810 ( .A1(n29713), .A2(n29712), .A3(n29711), .A4(n29710), .ZN(
        n29731) );
  NOR2_X1 U5811 ( .A1(n7619), .A2(n7612), .ZN(n29733) );
  AOI21_X1 U5812 ( .B1(n30042), .B2(n30228), .A(n30041), .ZN(n30056) );
  NAND2_X1 U5813 ( .A1(n30047), .A2(n30228), .ZN(n30055) );
  NAND2_X1 U5814 ( .A1(n30053), .A2(n30329), .ZN(n30054) );
  NAND2_X1 U5815 ( .A1(n30018), .A2(n30329), .ZN(n30057) );
  AOI22_X1 U5816 ( .A1(n30287), .A2(n30069), .B1(n30068), .B2(n30329), .ZN(
        n30099) );
  NAND2_X1 U5817 ( .A1(n30116), .A2(n30188), .ZN(n30117) );
  NAND2_X1 U5818 ( .A1(n30105), .A2(n30329), .ZN(n30119) );
  NAND2_X1 U5819 ( .A1(n30111), .A2(n30287), .ZN(n30118) );
  XNOR2_X1 U5820 ( .A(n33594), .B(\fmem_data[29][1] ), .ZN(n36121) );
  NAND2_X1 U5821 ( .A1(\fmem_data[29][1] ), .A2(n3575), .ZN(n36120) );
  OR2_X1 U5822 ( .A1(n36339), .A2(n3692), .ZN(n36217) );
  NAND2_X1 U5823 ( .A1(\fmem_data[3][1] ), .A2(n3582), .ZN(n36199) );
  NAND2_X1 U5824 ( .A1(\fmem_data[11][1] ), .A2(n3577), .ZN(n36196) );
  OAI22_X1 U5825 ( .A1(n36244), .A2(n34739), .B1(n34740), .B2(n3563), .ZN(
        n36527) );
  OR2_X1 U5826 ( .A1(n36101), .A2(n3670), .ZN(n32949) );
  OR2_X1 U5827 ( .A1(n36111), .A2(n3732), .ZN(n33450) );
  OAI22_X1 U5828 ( .A1(n36229), .A2(n36227), .B1(n33552), .B2(n3647), .ZN(
        n36472) );
  XNOR2_X1 U5829 ( .A(n36249), .B(n36248), .ZN(n36697) );
  XNOR2_X1 U5830 ( .A(n36247), .B(n36246), .ZN(n36249) );
  OAI22_X1 U5831 ( .A1(n34627), .A2(n34625), .B1(n33747), .B2(n3574), .ZN(
        n36238) );
  AND2_X1 U5832 ( .A1(n36315), .A2(n32900), .ZN(n36237) );
  XNOR2_X1 U5833 ( .A(n34581), .B(n34580), .ZN(n36605) );
  XNOR2_X1 U5834 ( .A(n34579), .B(n34578), .ZN(n34581) );
  XNOR2_X1 U5835 ( .A(n36351), .B(n36350), .ZN(n36353) );
  XNOR2_X1 U5836 ( .A(n36492), .B(n36491), .ZN(n36835) );
  XNOR2_X1 U5837 ( .A(n32977), .B(n32976), .ZN(n36321) );
  XNOR2_X1 U5838 ( .A(n32995), .B(n32994), .ZN(n36319) );
  OAI21_X1 U5839 ( .B1(n36363), .B2(n36362), .A(n36361), .ZN(n36681) );
  INV_X1 U5840 ( .A(n36707), .ZN(n36363) );
  NAND2_X1 U5841 ( .A1(n36706), .A2(n36705), .ZN(n36361) );
  NOR2_X1 U5842 ( .A1(n36706), .A2(n36705), .ZN(n36362) );
  NAND2_X1 U5843 ( .A1(n36186), .A2(n36187), .ZN(n34794) );
  XNOR2_X1 U5844 ( .A(n36741), .B(n36740), .ZN(n36742) );
  NAND2_X1 U5845 ( .A1(n36078), .A2(n36080), .ZN(n32848) );
  NAND2_X1 U5846 ( .A1(n36769), .A2(n36770), .ZN(n36263) );
  NAND2_X1 U5847 ( .A1(n34374), .A2(n34373), .ZN(n34177) );
  NAND2_X1 U5848 ( .A1(n36050), .A2(n36049), .ZN(n34546) );
  XNOR2_X1 U5849 ( .A(n30337), .B(n30338), .ZN(n29688) );
  XNOR2_X1 U5850 ( .A(n32502), .B(n32501), .ZN(n33419) );
  XNOR2_X1 U5851 ( .A(n32500), .B(n32499), .ZN(n32502) );
  XNOR2_X1 U5852 ( .A(n36613), .B(n36612), .ZN(n36896) );
  NAND2_X1 U5853 ( .A1(n36876), .A2(n36874), .ZN(n36543) );
  XNOR2_X1 U5854 ( .A(n36376), .B(n36375), .ZN(n36672) );
  NAND2_X1 U5855 ( .A1(n32908), .A2(n32907), .ZN(n36038) );
  NAND2_X1 U5856 ( .A1(n36153), .A2(n36154), .ZN(n32907) );
  OAI21_X1 U5857 ( .B1(n36154), .B2(n36153), .A(n36155), .ZN(n32908) );
  NAND2_X1 U5858 ( .A1(n36639), .A2(n36637), .ZN(n33922) );
  XNOR2_X1 U5859 ( .A(n36031), .B(n36030), .ZN(n36446) );
  AOI21_X1 U5860 ( .B1(n35705), .B2(n35704), .A(n35703), .ZN(n35706) );
  AND2_X1 U5861 ( .A1(n34624), .A2(\fmem_data[28][0] ), .ZN(n36520) );
  AND2_X1 U5862 ( .A1(n36105), .A2(\fmem_data[18][0] ), .ZN(n36522) );
  OAI22_X1 U5863 ( .A1(n36312), .A2(n36114), .B1(n36103), .B2(n3561), .ZN(
        n36582) );
  OAI22_X1 U5864 ( .A1(n36106), .A2(n3580), .B1(n36105), .B2(n36104), .ZN(
        n36581) );
  OAI22_X1 U5865 ( .A1(n36229), .A2(n3647), .B1(n36228), .B2(n36227), .ZN(
        n36692) );
  OAI22_X1 U5866 ( .A1(n36339), .A2(n36223), .B1(n36222), .B2(n3568), .ZN(
        n36791) );
  OAI22_X1 U5867 ( .A1(n36338), .A2(n36221), .B1(n36209), .B2(n3558), .ZN(
        n36795) );
  OAI22_X1 U5868 ( .A1(n36211), .A2(n3931), .B1(n36216), .B2(n36210), .ZN(
        n36794) );
  OAI22_X1 U5869 ( .A1(n36300), .A2(n3573), .B1(n36299), .B2(n36298), .ZN(
        n36716) );
  XNOR2_X1 U5870 ( .A(n36536), .B(n36535), .ZN(n36912) );
  XNOR2_X1 U5871 ( .A(n36534), .B(n36533), .ZN(n36536) );
  OAI22_X1 U5872 ( .A1(n34486), .A2(n3570), .B1(n34615), .B2(n34613), .ZN(
        n36328) );
  NAND2_X1 U5873 ( .A1(n36979), .A2(n36977), .ZN(n36869) );
  XNOR2_X1 U5874 ( .A(n36816), .B(n36815), .ZN(n36883) );
  XNOR2_X1 U5875 ( .A(n36814), .B(n36813), .ZN(n36816) );
  XNOR2_X1 U5876 ( .A(n36617), .B(n36616), .ZN(n36619) );
  XNOR2_X1 U5877 ( .A(n36051), .B(n36050), .ZN(n36764) );
  XNOR2_X1 U5878 ( .A(n36041), .B(n36040), .ZN(n36043) );
  NAND2_X1 U5879 ( .A1(n36664), .A2(n36663), .ZN(n36428) );
  INV_X1 U5880 ( .A(n36655), .ZN(n36438) );
  NAND2_X1 U5881 ( .A1(n35975), .A2(n35974), .ZN(n35976) );
  INV_X1 U5882 ( .A(n36005), .ZN(n36002) );
  INV_X1 U5883 ( .A(n36004), .ZN(n36003) );
  AND2_X1 U5884 ( .A1(n36111), .A2(\fmem_data[26][0] ), .ZN(n36564) );
  AND2_X1 U5885 ( .A1(n36112), .A2(\fmem_data[12][0] ), .ZN(n36563) );
  AND2_X1 U5886 ( .A1(n36200), .A2(\fmem_data[30][0] ), .ZN(n36723) );
  AND2_X1 U5887 ( .A1(n36299), .A2(\fmem_data[16][0] ), .ZN(n36722) );
  AND2_X1 U5888 ( .A1(n36244), .A2(\fmem_data[14][0] ), .ZN(n36719) );
  AND2_X1 U5889 ( .A1(n36312), .A2(\fmem_data[10][0] ), .ZN(n36725) );
  AND2_X1 U5890 ( .A1(n36315), .A2(\fmem_data[3][0] ), .ZN(n36861) );
  AND2_X1 U5891 ( .A1(n36339), .A2(\fmem_data[15][0] ), .ZN(n36857) );
  AND2_X1 U5892 ( .A1(n36338), .A2(\fmem_data[1][0] ), .ZN(n36858) );
  XNOR2_X1 U5893 ( .A(n36980), .B(n36979), .ZN(n37060) );
  XNOR2_X1 U5894 ( .A(n36978), .B(n36977), .ZN(n36980) );
  XNOR2_X1 U5895 ( .A(n37023), .B(n37022), .ZN(n37052) );
  XNOR2_X1 U5896 ( .A(n37021), .B(n37020), .ZN(n37023) );
  XNOR2_X1 U5897 ( .A(n36941), .B(n36940), .ZN(n37050) );
  XNOR2_X1 U5898 ( .A(n36939), .B(n36938), .ZN(n36940) );
  XNOR2_X1 U5899 ( .A(n36895), .B(n36894), .ZN(n37043) );
  XNOR2_X1 U5900 ( .A(n36893), .B(n36892), .ZN(n36895) );
  NAND2_X1 U5901 ( .A1(n36654), .A2(n36653), .ZN(n37160) );
  OAI21_X1 U5902 ( .B1(n35953), .B2(n35952), .A(n35951), .ZN(n35982) );
  OAI21_X1 U5903 ( .B1(n37218), .B2(n37228), .A(n37229), .ZN(n37153) );
  NOR2_X1 U5904 ( .A1(n37083), .A2(n37082), .ZN(n37298) );
  INV_X1 U5905 ( .A(n37081), .ZN(n37301) );
  OAI21_X1 U5906 ( .B1(n37303), .B2(n37080), .A(n37304), .ZN(n37081) );
  NAND2_X1 U5907 ( .A1(n37083), .A2(n37082), .ZN(n37299) );
  OAI21_X1 U5908 ( .B1(n37298), .B2(n37301), .A(n37299), .ZN(n37296) );
  OR2_X1 U5909 ( .A1(n37096), .A2(n37095), .ZN(n37291) );
  NAND2_X1 U5910 ( .A1(n37103), .A2(n37102), .ZN(n36887) );
  NAND2_X1 U5911 ( .A1(n37104), .A2(n36886), .ZN(n36888) );
  OR2_X1 U5912 ( .A1(n37103), .A2(n37102), .ZN(n36886) );
  NAND2_X1 U5913 ( .A1(n37152), .A2(n37151), .ZN(n37229) );
  AOI21_X1 U5914 ( .B1(n37222), .B2(n37221), .A(n37220), .ZN(n37223) );
  OAI21_X1 U5915 ( .B1(n37238), .B2(n37219), .A(n37218), .ZN(n37220) );
  NOR2_X1 U5916 ( .A1(n8406), .A2(n8414), .ZN(n8408) );
  NAND2_X1 U5917 ( .A1(n6172), .A2(n8415), .ZN(n8406) );
  INV_X1 U5918 ( .A(n37285), .ZN(n37286) );
  INV_X1 U5919 ( .A(n37275), .ZN(n37277) );
  INV_X1 U5920 ( .A(n37264), .ZN(n37266) );
  OAI21_X1 U5921 ( .B1(n37267), .B2(n37264), .A(n37265), .ZN(n37263) );
  INV_X1 U5922 ( .A(n37254), .ZN(n37256) );
  NOR2_X1 U5923 ( .A1(n37232), .A2(n37231), .ZN(n37237) );
  NAND2_X1 U5924 ( .A1(n37243), .A2(n37241), .ZN(n37203) );
  INV_X1 U5925 ( .A(n37246), .ZN(n37248) );
  NOR2_X1 U5926 ( .A1(n37202), .A2(n37246), .ZN(n37185) );
  OAI21_X1 U5927 ( .B1(n37241), .B2(n37246), .A(n37247), .ZN(n37184) );
  OAI22_X1 U5928 ( .A1(n36243), .A2(n34777), .B1(n34778), .B2(n3567), .ZN(
        n36568) );
  OR2_X1 U5929 ( .A1(n36243), .A2(n3693), .ZN(n34597) );
  XNOR2_X1 U5930 ( .A(n36243), .B(\fmem_data[22][5] ), .ZN(n32081) );
  XNOR2_X1 U5931 ( .A(n36243), .B(\fmem_data[22][3] ), .ZN(n31504) );
  OR2_X1 U5932 ( .A1(n36243), .A2(n3591), .ZN(n32075) );
  AND2_X1 U5933 ( .A1(n36243), .A2(n33745), .ZN(n34607) );
  AND2_X1 U5934 ( .A1(n36243), .A2(n31232), .ZN(n31532) );
  AND2_X1 U5935 ( .A1(n36243), .A2(\fmem_data[22][0] ), .ZN(n36720) );
  AND2_X1 U5936 ( .A1(n36243), .A2(n32113), .ZN(n32232) );
  OR2_X1 U5937 ( .A1(n36243), .A2(n3645), .ZN(n21766) );
  OR2_X1 U5938 ( .A1(n36243), .A2(n3603), .ZN(n31596) );
  NAND2_X1 U5939 ( .A1(n11333), .A2(n11332), .ZN(n35401) );
  INV_X1 U5940 ( .A(n29448), .ZN(n29456) );
  AOI21_X1 U5941 ( .B1(n36120), .B2(n3575), .A(n32732), .ZN(n27434) );
  XNOR2_X1 U5942 ( .A(n32225), .B(\fmem_data[9][5] ), .ZN(n30359) );
  OAI22_X1 U5943 ( .A1(n30360), .A2(n35040), .B1(n30359), .B2(n35041), .ZN(
        n30403) );
  OAI22_X1 U5944 ( .A1(n30359), .A2(n35040), .B1(n34861), .B2(n35041), .ZN(
        n25601) );
  XOR2_X1 U5945 ( .A(n30429), .B(n30428), .Z(n3291) );
  XOR2_X1 U5946 ( .A(n3291), .B(n30430), .Z(n31188) );
  NAND2_X1 U5947 ( .A1(n30430), .A2(n30429), .ZN(n3292) );
  NAND2_X1 U5948 ( .A1(n30430), .A2(n30428), .ZN(n3293) );
  NAND2_X1 U5949 ( .A1(n30429), .A2(n30428), .ZN(n3294) );
  NAND3_X1 U5950 ( .A1(n3292), .A2(n3293), .A3(n3294), .ZN(n30826) );
  OAI22_X1 U5951 ( .A1(n27973), .A2(n35498), .B1(n35497), .B2(n3623), .ZN(
        n30428) );
  NAND3_X1 U5952 ( .A1(n18141), .A2(n18140), .A3(n18139), .ZN(n3295) );
  NAND3_X1 U5953 ( .A1(n18141), .A2(n18140), .A3(n18139), .ZN(n32541) );
  BUF_X4 U5954 ( .A(n13476), .Z(n16986) );
  XNOR2_X1 U5955 ( .A(n32975), .B(n32974), .ZN(n32976) );
  NAND2_X1 U5956 ( .A1(n32975), .A2(n32974), .ZN(n31457) );
  OAI22_X1 U5957 ( .A1(n34538), .A2(n34535), .B1(n32535), .B2(n34537), .ZN(
        n32975) );
  BUF_X2 U5958 ( .A(n14928), .Z(n28045) );
  AND4_X1 U5959 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11918) );
  XOR2_X1 U5960 ( .A(n31520), .B(n31519), .Z(n3296) );
  XOR2_X1 U5961 ( .A(n31521), .B(n3296), .Z(n33439) );
  NAND2_X1 U5962 ( .A1(n31521), .A2(n31520), .ZN(n3297) );
  NAND2_X1 U5963 ( .A1(n31521), .A2(n31519), .ZN(n3298) );
  NAND2_X1 U5964 ( .A1(n31520), .A2(n31519), .ZN(n3299) );
  NAND3_X1 U5965 ( .A1(n3297), .A2(n3298), .A3(n3299), .ZN(n31570) );
  AND2_X1 U5966 ( .A1(n36299), .A2(n31400), .ZN(n31520) );
  AND2_X1 U5967 ( .A1(n36200), .A2(n31401), .ZN(n31519) );
  XNOR2_X1 U5968 ( .A(n32321), .B(\fmem_data[17][5] ), .ZN(n34046) );
  OAI22_X1 U5969 ( .A1(n34046), .A2(n34043), .B1(n32322), .B2(n34045), .ZN(
        n33066) );
  INV_X1 U5970 ( .A(n3336), .ZN(n3300) );
  AOI21_X1 U5971 ( .B1(n34435), .B2(n34437), .A(n33232), .ZN(n33233) );
  OAI22_X1 U5972 ( .A1(n33757), .A2(n3559), .B1(n34612), .B2(n34017), .ZN(
        n36530) );
  OAI22_X1 U5973 ( .A1(n34612), .A2(n28542), .B1(n33954), .B2(n3696), .ZN(
        n33987) );
  XNOR2_X1 U5974 ( .A(n34612), .B(\fmem_data[6][3] ), .ZN(n31450) );
  XNOR2_X1 U5975 ( .A(n34612), .B(\fmem_data[6][5] ), .ZN(n32575) );
  AND2_X1 U5976 ( .A1(n34612), .A2(n30399), .ZN(n32223) );
  AND2_X1 U5977 ( .A1(n34612), .A2(\fmem_data[6][0] ), .ZN(n36203) );
  XNOR2_X1 U5978 ( .A(n34612), .B(\fmem_data[6][7] ), .ZN(n19024) );
  AND2_X1 U5979 ( .A1(n34612), .A2(n26483), .ZN(n28534) );
  AND2_X1 U5980 ( .A1(n34612), .A2(n31537), .ZN(n34480) );
  OR2_X1 U5981 ( .A1(n34612), .A2(n3630), .ZN(n30388) );
  AOI21_X1 U5982 ( .B1(n34414), .B2(n34416), .A(n33050), .ZN(n33051) );
  NAND2_X1 U5983 ( .A1(n8732), .A2(n8731), .ZN(n3303) );
  NOR2_X1 U5984 ( .A1(n28988), .A2(n28987), .ZN(n28989) );
  XNOR2_X1 U5985 ( .A(n32615), .B(\fmem_data[24][3] ), .ZN(n32716) );
  AND2_X1 U5986 ( .A1(n3309), .A2(n3310), .ZN(n27879) );
  NOR2_X1 U5987 ( .A1(n27862), .A2(n27861), .ZN(n3309) );
  NOR3_X1 U5988 ( .A1(n27876), .A2(n27875), .A3(n27874), .ZN(n3310) );
  OR2_X1 U5989 ( .A1(n4061), .A2(n4063), .ZN(n4242) );
  NOR2_X1 U5990 ( .A1(n10288), .A2(n9417), .ZN(n9420) );
  XNOR2_X1 U5991 ( .A(n30846), .B(\fmem_data[13][7] ), .ZN(n30437) );
  AND2_X1 U5992 ( .A1(n16165), .A2(n16164), .ZN(n16166) );
  NAND2_X1 U5993 ( .A1(n16247), .A2(n16246), .ZN(n33554) );
  OAI22_X1 U5994 ( .A1(n31911), .A2(n3565), .B1(n31910), .B2(n36100), .ZN(
        n32488) );
  OAI22_X1 U5995 ( .A1(n34772), .A2(n36100), .B1(n31910), .B2(n3565), .ZN(
        n32993) );
  OAI22_X1 U5996 ( .A1(n31894), .A2(n34462), .B1(n22453), .B2(n34463), .ZN(
        n28909) );
  OAI22_X1 U5997 ( .A1(n32516), .A2(n35749), .B1(n32515), .B2(n35748), .ZN(
        n33172) );
  XNOR2_X1 U5998 ( .A(n32979), .B(\fmem_data[4][7] ), .ZN(n32516) );
  AOI21_X1 U5999 ( .B1(n22882), .B2(n23822), .A(n22881), .ZN(n22883) );
  XNOR2_X1 U6000 ( .A(n33592), .B(\fmem_data[14][7] ), .ZN(n31952) );
  OAI22_X1 U6001 ( .A1(n31955), .A2(n3559), .B1(n34016), .B2(n34017), .ZN(
        n26267) );
  AOI21_X1 U6002 ( .B1(n34017), .B2(n3559), .A(n31955), .ZN(n31956) );
  XNOR2_X1 U6003 ( .A(n3452), .B(\fmem_data[11][5] ), .ZN(n31979) );
  XNOR2_X1 U6004 ( .A(n32228), .B(\fmem_data[5][5] ), .ZN(n22778) );
  XNOR2_X1 U6005 ( .A(n32228), .B(\fmem_data[5][1] ), .ZN(n32420) );
  OAI22_X1 U6006 ( .A1(n35017), .A2(n35019), .B1(n12809), .B2(n35018), .ZN(
        n31828) );
  AOI21_X1 U6007 ( .B1(n35019), .B2(n35018), .A(n35017), .ZN(n35020) );
  AND2_X1 U6008 ( .A1(n5540), .A2(n3311), .ZN(n5543) );
  AND2_X1 U6009 ( .A1(n5542), .A2(n5541), .ZN(n3311) );
  XNOR2_X1 U6010 ( .A(n3312), .B(n3688), .ZN(n32154) );
  AND2_X1 U6011 ( .A1(n3274), .A2(n32557), .ZN(n3312) );
  INV_X1 U6012 ( .A(n31667), .ZN(n35335) );
  OAI22_X1 U6013 ( .A1(n33164), .A2(n35181), .B1(n33163), .B2(n35182), .ZN(
        n33203) );
  NAND4_X1 U6014 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n3313) );
  NAND4_X1 U6015 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n33459) );
  AND2_X1 U6016 ( .A1(n30223), .A2(\xmem_data[84][2] ), .ZN(n7907) );
  AND2_X1 U6017 ( .A1(n30223), .A2(\xmem_data[116][2] ), .ZN(n7959) );
  NAND2_X1 U6018 ( .A1(n12020), .A2(n28258), .ZN(n12043) );
  INV_X1 U6019 ( .A(n15313), .ZN(n3314) );
  NAND2_X1 U6020 ( .A1(n15309), .A2(n3315), .ZN(n15319) );
  NOR2_X1 U6021 ( .A1(n15312), .A2(n3314), .ZN(n3315) );
  NAND4_X1 U6022 ( .A1(n8196), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n3316)
         );
  NAND4_X1 U6023 ( .A1(n8196), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n31247)
         );
  XNOR2_X1 U6024 ( .A(n35256), .B(\fmem_data[31][7] ), .ZN(n35661) );
  OAI22_X1 U6025 ( .A1(n30368), .A2(n35701), .B1(n32179), .B2(n35700), .ZN(
        n30990) );
  OAI22_X1 U6026 ( .A1(n30368), .A2(n35700), .B1(n33216), .B2(n35701), .ZN(
        n20290) );
  OAI21_X1 U6027 ( .B1(n3724), .B2(n17105), .A(n20311), .ZN(n17179) );
  XNOR2_X1 U6028 ( .A(n31657), .B(\fmem_data[28][3] ), .ZN(n32643) );
  OAI22_X1 U6029 ( .A1(n33798), .A2(n33797), .B1(n3456), .B2(n33796), .ZN(
        n3319) );
  XNOR2_X1 U6030 ( .A(n23174), .B(n23173), .ZN(n23176) );
  NOR3_X1 U6031 ( .A1(n10486), .A2(n10485), .A3(n10484), .ZN(n10493) );
  AND2_X1 U6032 ( .A1(n29626), .A2(\xmem_data[124][7] ), .ZN(n12153) );
  NAND2_X1 U6033 ( .A1(n30143), .A2(n30142), .ZN(n30144) );
  OAI21_X1 U6034 ( .B1(n30143), .B2(n30142), .A(n30141), .ZN(n30145) );
  XNOR2_X1 U6035 ( .A(n35340), .B(\fmem_data[20][7] ), .ZN(n35738) );
  XNOR2_X1 U6036 ( .A(n35340), .B(\fmem_data[20][3] ), .ZN(n32013) );
  NAND2_X1 U6037 ( .A1(n12127), .A2(n12126), .ZN(n3320) );
  NAND2_X1 U6038 ( .A1(n28922), .A2(n28920), .ZN(n23578) );
  XNOR2_X1 U6039 ( .A(n33803), .B(\fmem_data[24][3] ), .ZN(n34432) );
  XNOR2_X1 U6040 ( .A(n33803), .B(\fmem_data[24][7] ), .ZN(n31953) );
  NAND4_X1 U6041 ( .A1(n22452), .A2(n22451), .A3(n22450), .A4(n22449), .ZN(
        n3321) );
  NAND4_X1 U6042 ( .A1(n22452), .A2(n22451), .A3(n22450), .A4(n22449), .ZN(
        n31980) );
  INV_X1 U6043 ( .A(n25480), .ZN(n25484) );
  NAND2_X1 U6044 ( .A1(n34050), .A2(n34049), .ZN(n3323) );
  BUF_X1 U6045 ( .A(n4158), .Z(n3324) );
  BUF_X1 U6046 ( .A(n3324), .Z(n3325) );
  BUF_X1 U6047 ( .A(n3324), .Z(n3326) );
  NAND2_X1 U6048 ( .A1(n10434), .A2(n10445), .ZN(n10446) );
  AND2_X1 U6049 ( .A1(n36228), .A2(n27324), .ZN(n26272) );
  AND2_X1 U6050 ( .A1(n36228), .A2(n31536), .ZN(n33462) );
  AND2_X1 U6051 ( .A1(n36228), .A2(\fmem_data[20][0] ), .ZN(n36557) );
  OR2_X1 U6052 ( .A1(n36228), .A2(n3628), .ZN(n33795) );
  AND2_X1 U6053 ( .A1(n36228), .A2(n32590), .ZN(n32784) );
  XNOR2_X1 U6054 ( .A(n31798), .B(\fmem_data[14][7] ), .ZN(n33312) );
  XNOR2_X1 U6055 ( .A(n31798), .B(\fmem_data[14][1] ), .ZN(n32238) );
  XNOR2_X1 U6056 ( .A(n31798), .B(\fmem_data[14][5] ), .ZN(n30416) );
  NAND3_X1 U6057 ( .A1(n9851), .A2(n9850), .A3(n9849), .ZN(n9857) );
  INV_X1 U6058 ( .A(n3327), .ZN(n3328) );
  BUF_X2 U6059 ( .A(n11453), .Z(n29579) );
  AND2_X1 U6060 ( .A1(n36110), .A2(\fmem_data[25][0] ), .ZN(n36565) );
  AND2_X1 U6061 ( .A1(n36110), .A2(n32076), .ZN(n32416) );
  OR2_X1 U6062 ( .A1(n36110), .A2(n3679), .ZN(n33481) );
  OR2_X1 U6063 ( .A1(n36110), .A2(n3634), .ZN(n32778) );
  AND2_X1 U6064 ( .A1(n36110), .A2(n31499), .ZN(n33470) );
  AND2_X1 U6065 ( .A1(n36110), .A2(n34051), .ZN(n34210) );
  OR2_X1 U6066 ( .A1(n36110), .A2(n3644), .ZN(n33794) );
  OR2_X1 U6067 ( .A1(n36110), .A2(n3622), .ZN(n27433) );
  NAND4_X2 U6068 ( .A1(n27432), .A2(n27431), .A3(n27430), .A4(n27429), .ZN(
        n36110) );
  OAI22_X1 U6069 ( .A1(n32056), .A2(n34742), .B1(n32240), .B2(n3571), .ZN(
        n31488) );
  OAI22_X1 U6070 ( .A1(n32241), .A2(n3571), .B1(n32240), .B2(n34742), .ZN(
        n32694) );
  XNOR2_X1 U6071 ( .A(n31662), .B(\fmem_data[12][3] ), .ZN(n33274) );
  XNOR2_X1 U6072 ( .A(n31662), .B(\fmem_data[12][7] ), .ZN(n33316) );
  XNOR2_X1 U6073 ( .A(n31662), .B(\fmem_data[12][5] ), .ZN(n30472) );
  NAND4_X1 U6074 ( .A1(n14382), .A2(n14381), .A3(n14380), .A4(n14379), .ZN(
        n31662) );
  OAI22_X1 U6075 ( .A1(n35024), .A2(n35497), .B1(n35406), .B2(n35498), .ZN(
        n35260) );
  OAI22_X1 U6076 ( .A1(n35024), .A2(n35498), .B1(n23920), .B2(n35497), .ZN(
        n35091) );
  NAND2_X1 U6077 ( .A1(n34685), .A2(n34684), .ZN(n34890) );
  NAND2_X1 U6078 ( .A1(n34300), .A2(n34301), .ZN(n34142) );
  OAI22_X1 U6079 ( .A1(n34600), .A2(n3569), .B1(n34599), .B2(n34598), .ZN(
        n36569) );
  XNOR2_X1 U6080 ( .A(n34599), .B(\fmem_data[4][3] ), .ZN(n31494) );
  XNOR2_X1 U6081 ( .A(n34599), .B(\fmem_data[4][5] ), .ZN(n31444) );
  OAI22_X1 U6082 ( .A1(n34599), .A2(n30386), .B1(n35748), .B2(n3614), .ZN(
        n30993) );
  OAI22_X1 U6083 ( .A1(n34599), .A2(n32552), .B1(n33176), .B2(n3610), .ZN(
        n34749) );
  OAI22_X1 U6084 ( .A1(n34599), .A2(n28540), .B1(n35010), .B2(n3632), .ZN(
        n33988) );
  XNOR2_X1 U6085 ( .A(n34599), .B(\fmem_data[4][7] ), .ZN(n32515) );
  AND2_X1 U6086 ( .A1(n34599), .A2(\fmem_data[4][0] ), .ZN(n36562) );
  AND2_X1 U6087 ( .A1(n34599), .A2(n31449), .ZN(n33446) );
  AND2_X1 U6088 ( .A1(n34599), .A2(n20937), .ZN(n34108) );
  NOR2_X1 U6089 ( .A1(n11359), .A2(n6202), .ZN(n6247) );
  XNOR2_X1 U6090 ( .A(n34610), .B(\fmem_data[12][3] ), .ZN(n33583) );
  OAI22_X1 U6091 ( .A1(n31533), .A2(n33582), .B1(n33583), .B2(n34340), .ZN(
        n33495) );
  NAND3_X1 U6092 ( .A1(n8351), .A2(n3828), .A3(n3155), .ZN(n8354) );
  XNOR2_X1 U6093 ( .A(n32938), .B(\fmem_data[1][3] ), .ZN(n32594) );
  XNOR2_X1 U6094 ( .A(n32938), .B(\fmem_data[1][7] ), .ZN(n30368) );
  INV_X1 U6095 ( .A(n3349), .ZN(n3350) );
  NAND4_X1 U6096 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n3354) );
  NAND4_X1 U6097 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n34611) );
  OAI22_X1 U6098 ( .A1(n36102), .A2(n3565), .B1(n36101), .B2(n36100), .ZN(
        n36583) );
  XNOR2_X1 U6099 ( .A(n33683), .B(\fmem_data[24][1] ), .ZN(n36102) );
  XNOR2_X1 U6100 ( .A(n35401), .B(\fmem_data[0][1] ), .ZN(n31966) );
  OR2_X2 U6101 ( .A1(n10972), .A2(n4059), .ZN(n4536) );
  OAI22_X1 U6102 ( .A1(n34425), .A2(n34422), .B1(n33595), .B2(n34424), .ZN(
        n33714) );
  XNOR2_X1 U6103 ( .A(n33594), .B(\fmem_data[29][3] ), .ZN(n34425) );
  XNOR2_X1 U6104 ( .A(n28919), .B(n28918), .ZN(n33622) );
  NAND2_X1 U6105 ( .A1(n28917), .A2(n28916), .ZN(n26373) );
  OAI22_X1 U6106 ( .A1(n31163), .A2(n34501), .B1(n31453), .B2(n34499), .ZN(
        n32083) );
  OAI22_X1 U6107 ( .A1(n31163), .A2(n34499), .B1(n26270), .B2(n34501), .ZN(
        n28896) );
  INV_X1 U6108 ( .A(n26377), .ZN(n21093) );
  XNOR2_X1 U6109 ( .A(n28905), .B(n28904), .ZN(n28907) );
  NAND2_X1 U6110 ( .A1(n28906), .A2(n28905), .ZN(n26255) );
  XNOR2_X1 U6111 ( .A(n28907), .B(n28906), .ZN(n30131) );
  OAI22_X1 U6112 ( .A1(n32150), .A2(n34908), .B1(n34234), .B2(n34909), .ZN(
        n28905) );
  XNOR2_X1 U6113 ( .A(n31704), .B(\fmem_data[17][5] ), .ZN(n30473) );
  OAI22_X1 U6114 ( .A1(n33200), .A2(n35591), .B1(n33199), .B2(n35592), .ZN(
        n33258) );
  XNOR2_X1 U6115 ( .A(n32541), .B(\fmem_data[13][7] ), .ZN(n33199) );
  NAND4_X1 U6116 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n3356)
         );
  BUF_X2 U6117 ( .A(n14933), .Z(n3357) );
  OAI22_X1 U6118 ( .A1(n33689), .A2(n3558), .B1(n36209), .B2(n36221), .ZN(
        n36305) );
  XNOR2_X1 U6119 ( .A(n34862), .B(\fmem_data[16][5] ), .ZN(n32017) );
  NAND3_X1 U6120 ( .A1(n14738), .A2(n14737), .A3(n14736), .ZN(n14743) );
  OAI22_X1 U6121 ( .A1(n34078), .A2(n3558), .B1(n33866), .B2(n36221), .ZN(
        n32158) );
  AOI21_X1 U6122 ( .B1(n36221), .B2(n3558), .A(n34078), .ZN(n34079) );
  NAND3_X1 U6123 ( .A1(n3361), .A2(n12808), .A3(n12807), .ZN(n3359) );
  OAI21_X1 U6124 ( .B1(n3362), .B2(n3363), .A(n17073), .ZN(n3361) );
  NAND2_X1 U6125 ( .A1(n12744), .A2(n12743), .ZN(n3362) );
  OR2_X1 U6126 ( .A1(n12751), .A2(n12750), .ZN(n3363) );
  OAI22_X1 U6127 ( .A1(n33994), .A2(n34779), .B1(n33993), .B2(n34466), .ZN(
        n34063) );
  OAI22_X1 U6128 ( .A1(n33578), .A2(n36295), .B1(n33577), .B2(n3564), .ZN(
        n33697) );
  NAND2_X1 U6129 ( .A1(n32945), .A2(n32944), .ZN(n32073) );
  BUF_X2 U6130 ( .A(n7452), .Z(n29418) );
  BUF_X2 U6131 ( .A(n8088), .Z(n28765) );
  AND2_X1 U6132 ( .A1(n17095), .A2(n17094), .ZN(n17096) );
  NAND2_X1 U6133 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  OR2_X1 U6134 ( .A1(n6589), .A2(n37199), .ZN(n3364) );
  NAND2_X1 U6135 ( .A1(n3364), .A2(n10069), .ZN(n6611) );
  BUF_X2 U6136 ( .A(n7452), .Z(n27743) );
  XNOR2_X1 U6137 ( .A(n31125), .B(\fmem_data[0][7] ), .ZN(n31641) );
  NAND4_X1 U6138 ( .A1(n21393), .A2(n21392), .A3(n21391), .A4(n21390), .ZN(
        n3365) );
  NAND4_X1 U6139 ( .A1(n21393), .A2(n21392), .A3(n21391), .A4(n21390), .ZN(
        n33844) );
  OAI22_X1 U6140 ( .A1(n32002), .A2(n35511), .B1(n35512), .B2(n32001), .ZN(
        n33072) );
  XNOR2_X1 U6141 ( .A(n32882), .B(\fmem_data[6][7] ), .ZN(n32002) );
  BUF_X2 U6142 ( .A(n8073), .Z(n28725) );
  NAND4_X1 U6143 ( .A1(n7297), .A2(n7296), .A3(n7295), .A4(n7294), .ZN(n3366)
         );
  NAND4_X1 U6144 ( .A1(n7297), .A2(n7296), .A3(n7295), .A4(n7294), .ZN(n3367)
         );
  BUF_X1 U6145 ( .A(n11437), .Z(n3368) );
  BUF_X1 U6146 ( .A(n11437), .Z(n3369) );
  NAND4_X1 U6147 ( .A1(n7297), .A2(n7296), .A3(n7295), .A4(n7294), .ZN(n31402)
         );
  NAND2_X1 U6148 ( .A1(n36179), .A2(n36178), .ZN(n36805) );
  NAND3_X1 U6149 ( .A1(n8893), .A2(n8892), .A3(n8891), .ZN(n8894) );
  XNOR2_X1 U6150 ( .A(n30826), .B(n30825), .ZN(n31000) );
  NAND2_X1 U6151 ( .A1(n37154), .A2(n37239), .ZN(n3370) );
  BUF_X2 U6152 ( .A(n7452), .Z(n27812) );
  XNOR2_X1 U6153 ( .A(n31393), .B(n31392), .ZN(n31462) );
  NAND2_X1 U6154 ( .A1(n31426), .A2(n31427), .ZN(n31410) );
  NAND4_X1 U6155 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n3371)
         );
  BUF_X1 U6156 ( .A(n14882), .Z(n3372) );
  OAI22_X1 U6157 ( .A1(n33106), .A2(n33105), .B1(n33104), .B2(n33103), .ZN(
        n34992) );
  XNOR2_X1 U6158 ( .A(n31658), .B(\fmem_data[30][5] ), .ZN(n30420) );
  XNOR2_X1 U6159 ( .A(n34032), .B(n34031), .ZN(n34188) );
  XNOR2_X1 U6160 ( .A(n34030), .B(n34029), .ZN(n34032) );
  NAND3_X1 U6161 ( .A1(n24834), .A2(n24833), .A3(n24832), .ZN(n3376) );
  NAND2_X1 U6162 ( .A1(n6176), .A2(n11343), .ZN(n3377) );
  NAND2_X1 U6163 ( .A1(n6176), .A2(n11343), .ZN(n11360) );
  NOR2_X2 U6164 ( .A1(n6183), .A2(n3248), .ZN(n6176) );
  INV_X1 U6165 ( .A(n3379), .ZN(n3380) );
  AND3_X1 U6166 ( .A1(n29182), .A2(n3381), .A3(n29183), .ZN(n29184) );
  NAND2_X1 U6167 ( .A1(n30885), .A2(\xmem_data[83][1] ), .ZN(n3381) );
  BUF_X2 U6168 ( .A(n11437), .Z(n29646) );
  INV_X1 U6169 ( .A(n3347), .ZN(n3382) );
  NAND3_X1 U6170 ( .A1(n20117), .A2(n20116), .A3(n20115), .ZN(n20121) );
  INV_X1 U6171 ( .A(n3385), .ZN(n3386) );
  XNOR2_X1 U6172 ( .A(n33555), .B(\fmem_data[21][1] ), .ZN(n34486) );
  XNOR2_X1 U6173 ( .A(n33555), .B(\fmem_data[21][7] ), .ZN(n32757) );
  XNOR2_X1 U6174 ( .A(n36664), .B(n36663), .ZN(n36665) );
  OR2_X1 U6175 ( .A1(n33800), .A2(n3683), .ZN(n32950) );
  XNOR2_X1 U6176 ( .A(n33800), .B(\fmem_data[13][3] ), .ZN(n32070) );
  XNOR2_X1 U6177 ( .A(n33800), .B(\fmem_data[13][7] ), .ZN(n17464) );
  AND2_X1 U6178 ( .A1(n33800), .A2(\fmem_data[13][0] ), .ZN(n36524) );
  OR2_X1 U6179 ( .A1(n33800), .A2(n3641), .ZN(n32790) );
  AND2_X1 U6180 ( .A1(n33800), .A2(n32579), .ZN(n32691) );
  OR2_X1 U6181 ( .A1(n33800), .A2(n3613), .ZN(n28402) );
  OR2_X1 U6182 ( .A1(n33800), .A2(n3612), .ZN(n33801) );
  AND2_X1 U6183 ( .A1(n33800), .A2(n21395), .ZN(n33942) );
  AND2_X1 U6184 ( .A1(n33800), .A2(n31528), .ZN(n32961) );
  XNOR2_X1 U6185 ( .A(n35403), .B(\fmem_data[21][1] ), .ZN(n31943) );
  XNOR2_X1 U6186 ( .A(n3257), .B(\fmem_data[19][1] ), .ZN(n34346) );
  AOI22_X1 U6187 ( .A1(n29683), .A2(n29682), .B1(n29681), .B2(n29680), .ZN(
        n3389) );
  NAND4_X1 U6188 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n3390) );
  NAND4_X1 U6189 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n31451) );
  OAI22_X1 U6190 ( .A1(n32134), .A2(n33249), .B1(n30791), .B2(n33250), .ZN(
        n31192) );
  OAI22_X1 U6191 ( .A1(n34242), .A2(n35725), .B1(n31977), .B2(n35726), .ZN(
        n33108) );
  OR3_X1 U6192 ( .A1(n5448), .A2(n5447), .A3(n5446), .ZN(n5449) );
  AND2_X1 U6193 ( .A1(n27741), .A2(\xmem_data[8][3] ), .ZN(n26198) );
  OAI22_X1 U6194 ( .A1(n31971), .A2(n34945), .B1(n31970), .B2(n34944), .ZN(
        n33141) );
  OAI22_X1 U6195 ( .A1(n34627), .A2(n3574), .B1(n34626), .B2(n34625), .ZN(
        n36517) );
  OR2_X1 U6196 ( .A1(n34626), .A2(n3666), .ZN(n32952) );
  XNOR2_X1 U6197 ( .A(n34626), .B(\fmem_data[8][5] ), .ZN(n32129) );
  AND2_X1 U6198 ( .A1(n34626), .A2(\fmem_data[8][0] ), .ZN(n36561) );
  AND2_X1 U6199 ( .A1(n34626), .A2(n32533), .ZN(n32619) );
  AND2_X1 U6200 ( .A1(n34626), .A2(n31448), .ZN(n33447) );
  AND2_X1 U6201 ( .A1(n34626), .A2(n20841), .ZN(n34109) );
  NAND3_X1 U6202 ( .A1(n17670), .A2(n17669), .A3(n3702), .ZN(n17671) );
  NAND3_X1 U6203 ( .A1(n17662), .A2(n17661), .A3(n17660), .ZN(n17663) );
  OAI22_X1 U6204 ( .A1(n32071), .A2(n34745), .B1(n32524), .B2(n3562), .ZN(
        n31487) );
  XNOR2_X1 U6205 ( .A(n30156), .B(\fmem_data[28][1] ), .ZN(n32524) );
  OAI22_X1 U6206 ( .A1(n34530), .A2(n3566), .B1(n33751), .B2(n34529), .ZN(
        n36533) );
  OR2_X1 U6207 ( .A1(n33751), .A2(n3669), .ZN(n32948) );
  XNOR2_X1 U6208 ( .A(n33751), .B(\fmem_data[17][3] ), .ZN(n32068) );
  AND2_X1 U6209 ( .A1(n33751), .A2(\fmem_data[17][0] ), .ZN(n36560) );
  AND2_X1 U6210 ( .A1(n33751), .A2(n32532), .ZN(n32620) );
  OR2_X1 U6211 ( .A1(n33751), .A2(n3654), .ZN(n32435) );
  OR2_X1 U6212 ( .A1(n33751), .A2(n3626), .ZN(n31473) );
  AND2_X1 U6213 ( .A1(n33751), .A2(n31447), .ZN(n33448) );
  AND2_X1 U6214 ( .A1(n33751), .A2(n20840), .ZN(n34110) );
  NAND4_X2 U6215 ( .A1(n19115), .A2(n19114), .A3(n19113), .A4(n19112), .ZN(
        n33751) );
  XNOR2_X1 U6216 ( .A(n33749), .B(\fmem_data[13][5] ), .ZN(n32539) );
  XNOR2_X1 U6217 ( .A(n33749), .B(\fmem_data[13][7] ), .ZN(n33200) );
  NAND4_X1 U6218 ( .A1(n17300), .A2(n17299), .A3(n17298), .A4(n17297), .ZN(
        n17317) );
  NAND3_X1 U6219 ( .A1(n29504), .A2(n29503), .A3(n29502), .ZN(n29505) );
  BUF_X4 U6220 ( .A(n18518), .Z(n30765) );
  NOR2_X1 U6221 ( .A1(n36314), .A2(n3931), .ZN(n36862) );
  NAND2_X1 U6222 ( .A1(n36314), .A2(\fmem_data[31][1] ), .ZN(n36215) );
  NAND2_X1 U6223 ( .A1(n36314), .A2(\fmem_data[31][3] ), .ZN(n34338) );
  XNOR2_X1 U6224 ( .A(n36314), .B(n3485), .ZN(n34469) );
  XNOR2_X1 U6225 ( .A(n36314), .B(n3487), .ZN(n32259) );
  NAND2_X1 U6226 ( .A1(n36314), .A2(\fmem_data[31][7] ), .ZN(n32187) );
  NOR2_X1 U6227 ( .A1(n36314), .A2(n34470), .ZN(n36257) );
  NOR2_X1 U6228 ( .A1(n36314), .A2(n35663), .ZN(n31213) );
  NAND2_X1 U6229 ( .A1(n36314), .A2(\fmem_data[31][5] ), .ZN(n31242) );
  NOR2_X1 U6230 ( .A1(n36314), .A2(n34944), .ZN(n34351) );
  NAND2_X1 U6231 ( .A1(n6486), .A2(n6485), .ZN(n6488) );
  NAND2_X1 U6232 ( .A1(n6486), .A2(n6586), .ZN(n5985) );
  NOR2_X1 U6233 ( .A1(n6486), .A2(n8416), .ZN(n8415) );
  BUF_X2 U6234 ( .A(n11451), .Z(n3392) );
  OAI22_X1 U6235 ( .A1(n32669), .A2(n35634), .B1(n35633), .B2(n3663), .ZN(
        n32718) );
  OAI21_X1 U6236 ( .B1(n28764), .B2(n28763), .A(n28762), .ZN(n28797) );
  OAI22_X1 U6237 ( .A1(n30157), .A2(n33828), .B1(n32754), .B2(n33827), .ZN(
        n30346) );
  OAI22_X1 U6238 ( .A1(n30157), .A2(n33827), .B1(n33322), .B2(n33828), .ZN(
        n23596) );
  XNOR2_X1 U6239 ( .A(n34610), .B(\fmem_data[12][7] ), .ZN(n33924) );
  OAI22_X1 U6240 ( .A1(n30158), .A2(n35019), .B1(n34035), .B2(n35018), .ZN(
        n30345) );
  NAND2_X1 U6241 ( .A1(n33202), .A2(n33201), .ZN(n33165) );
  OAI21_X1 U6242 ( .B1(n33202), .B2(n33201), .A(n33203), .ZN(n33166) );
  OAI22_X1 U6243 ( .A1(n30413), .A2(n34201), .B1(n33158), .B2(n34199), .ZN(
        n30467) );
  XNOR2_X1 U6244 ( .A(n31146), .B(n31145), .ZN(n3393) );
  XNOR2_X1 U6245 ( .A(n23575), .B(n23574), .ZN(n23576) );
  NAND2_X1 U6246 ( .A1(n8949), .A2(n3154), .ZN(n8950) );
  OR2_X1 U6247 ( .A1(n4048), .A2(n10972), .ZN(n4037) );
  OAI22_X1 U6248 ( .A1(n32008), .A2(n35705), .B1(n32007), .B2(n35704), .ZN(
        n32519) );
  OAI22_X1 U6249 ( .A1(n33790), .A2(n34437), .B1(n32613), .B2(n34435), .ZN(
        n32671) );
  NOR2_X1 U6250 ( .A1(n7599), .A2(n6169), .ZN(n3394) );
  OAI22_X1 U6251 ( .A1(n34100), .A2(n35011), .B1(n34099), .B2(n35010), .ZN(
        n34134) );
  XNOR2_X1 U6252 ( .A(n32131), .B(\fmem_data[4][5] ), .ZN(n34099) );
  NAND2_X1 U6253 ( .A1(n36260), .A2(n36259), .ZN(n32931) );
  OR2_X1 U6254 ( .A1(n37092), .A2(n37091), .ZN(n37295) );
  OAI22_X1 U6255 ( .A1(n31244), .A2(n34941), .B1(n31243), .B2(n34942), .ZN(
        n31565) );
  XNOR2_X1 U6256 ( .A(n36338), .B(\fmem_data[1][5] ), .ZN(n31244) );
  OAI22_X1 U6257 ( .A1(n30416), .A2(n33098), .B1(n33099), .B2(n33100), .ZN(
        n23595) );
  OAI22_X1 U6258 ( .A1(n33101), .A2(n33100), .B1(n33099), .B2(n33098), .ZN(
        n34994) );
  BUF_X1 U6259 ( .A(n6190), .Z(n3395) );
  XNOR2_X1 U6260 ( .A(n32328), .B(n32327), .ZN(n32330) );
  XNOR2_X1 U6261 ( .A(n32330), .B(n32329), .ZN(n32406) );
  OAI22_X1 U6262 ( .A1(n22775), .A2(n35497), .B1(n30358), .B2(n35498), .ZN(
        n34236) );
  XNOR2_X1 U6263 ( .A(n33553), .B(\fmem_data[5][7] ), .ZN(n22775) );
  XNOR2_X1 U6264 ( .A(n32360), .B(n32359), .ZN(n32378) );
  OAI22_X1 U6265 ( .A1(n31979), .A2(n34932), .B1(n32024), .B2(n34933), .ZN(
        n34258) );
  OAI22_X1 U6266 ( .A1(n30448), .A2(n35494), .B1(n30447), .B2(n35493), .ZN(
        n31734) );
  INV_X1 U6267 ( .A(n31801), .ZN(n35330) );
  AOI21_X1 U6268 ( .B1(n33956), .B2(n33954), .A(n33368), .ZN(n31801) );
  OAI22_X1 U6269 ( .A1(n24431), .A2(n35581), .B1(n31989), .B2(n35580), .ZN(
        n29536) );
  XNOR2_X1 U6270 ( .A(n31512), .B(\fmem_data[17][1] ), .ZN(n34528) );
  AND2_X1 U6271 ( .A1(n34343), .A2(n3578), .ZN(n3396) );
  NAND2_X1 U6272 ( .A1(\fmem_data[2][1] ), .A2(n3578), .ZN(n34343) );
  NAND4_X1 U6273 ( .A1(n3397), .A2(n3398), .A3(n3399), .A4(n3400), .ZN(n12785)
         );
  AND4_X1 U6274 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n3397) );
  AND4_X1 U6275 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n3398) );
  AND4_X1 U6276 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12760), .ZN(
        n3399) );
  AND4_X1 U6277 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n12764), .ZN(
        n3400) );
  NAND2_X1 U6278 ( .A1(n14001), .A2(n14000), .ZN(n35280) );
  OAI22_X1 U6279 ( .A1(n32752), .A2(n3678), .B1(n32164), .B2(n33725), .ZN(
        n30429) );
  XNOR2_X1 U6280 ( .A(n32319), .B(\fmem_data[29][5] ), .ZN(n24112) );
  XNOR2_X1 U6281 ( .A(n32319), .B(\fmem_data[29][1] ), .ZN(n32243) );
  XNOR2_X1 U6282 ( .A(n32319), .B(\fmem_data[29][7] ), .ZN(n33129) );
  AND2_X1 U6283 ( .A1(\xmem_data[28][3] ), .A2(n30674), .ZN(n3401) );
  NOR2_X1 U6284 ( .A1(n3401), .A2(n13441), .ZN(n13450) );
  AOI21_X1 U6285 ( .B1(n36114), .B2(n3561), .A(n32730), .ZN(n22360) );
  OAI22_X1 U6286 ( .A1(n32730), .A2(n3561), .B1(n32729), .B2(n36114), .ZN(
        n33207) );
  XNOR2_X1 U6287 ( .A(n32005), .B(\fmem_data[16][5] ), .ZN(n32564) );
  NAND3_X1 U6288 ( .A1(n12998), .A2(n12997), .A3(n12996), .ZN(n12999) );
  XNOR2_X1 U6289 ( .A(n31895), .B(\fmem_data[4][5] ), .ZN(n30418) );
  OAI22_X1 U6290 ( .A1(n30418), .A2(n35010), .B1(n31822), .B2(n35011), .ZN(
        n23923) );
  AOI21_X1 U6291 ( .B1(n35034), .B2(n35033), .A(n35032), .ZN(n35035) );
  BUF_X2 U6292 ( .A(n13476), .Z(n28334) );
  OR2_X1 U6293 ( .A1(n3354), .A2(n3691), .ZN(n33482) );
  OR2_X1 U6294 ( .A1(n3354), .A2(n3652), .ZN(n32605) );
  OR2_X1 U6295 ( .A1(n3353), .A2(n3620), .ZN(n33843) );
  AND2_X1 U6296 ( .A1(n3353), .A2(n32588), .ZN(n32786) );
  OR2_X1 U6297 ( .A1(n34611), .A2(n3624), .ZN(n29518) );
  AND2_X1 U6298 ( .A1(n3353), .A2(n31534), .ZN(n33464) );
  AND2_X1 U6299 ( .A1(n34611), .A2(n17079), .ZN(n26274) );
  OAI22_X1 U6300 ( .A1(n32527), .A2(n3578), .B1(n32526), .B2(n34343), .ZN(
        n32776) );
  XNOR2_X1 U6301 ( .A(n31885), .B(\fmem_data[5][3] ), .ZN(n33181) );
  XNOR2_X1 U6302 ( .A(n31885), .B(\fmem_data[5][7] ), .ZN(n35024) );
  NAND3_X1 U6303 ( .A1(n5568), .A2(n5566), .A3(n5567), .ZN(n31885) );
  XOR2_X1 U6304 ( .A(n27331), .B(n27332), .Z(n3403) );
  XOR2_X1 U6305 ( .A(n3403), .B(n27330), .Z(n30147) );
  NAND2_X1 U6306 ( .A1(n27330), .A2(n27331), .ZN(n3404) );
  NAND2_X1 U6307 ( .A1(n27330), .A2(n27332), .ZN(n3405) );
  NAND2_X1 U6308 ( .A1(n27331), .A2(n27332), .ZN(n3406) );
  NAND3_X1 U6309 ( .A1(n3404), .A2(n3405), .A3(n3406), .ZN(n26039) );
  OAI22_X1 U6310 ( .A1(n24726), .A2(n35182), .B1(n33163), .B2(n35181), .ZN(
        n27332) );
  OAI22_X1 U6311 ( .A1(n24727), .A2(n35749), .B1(n30408), .B2(n35748), .ZN(
        n27331) );
  XNOR2_X1 U6312 ( .A(n32596), .B(\fmem_data[18][7] ), .ZN(n33037) );
  OAI22_X1 U6313 ( .A1(n36121), .A2(n3575), .B1(n36245), .B2(n36120), .ZN(
        n36585) );
  OR2_X1 U6314 ( .A1(n36245), .A2(n3660), .ZN(n34595) );
  OR2_X1 U6315 ( .A1(n36245), .A2(n3588), .ZN(n32237) );
  XNOR2_X1 U6316 ( .A(n36245), .B(\fmem_data[29][7] ), .ZN(n32650) );
  AND2_X1 U6317 ( .A1(n36245), .A2(\fmem_data[29][0] ), .ZN(n36718) );
  AND2_X1 U6318 ( .A1(n36245), .A2(n32220), .ZN(n32264) );
  AND2_X1 U6319 ( .A1(n36245), .A2(n28532), .ZN(n31510) );
  XNOR2_X1 U6320 ( .A(n36245), .B(\fmem_data[29][5] ), .ZN(n31172) );
  AND2_X1 U6321 ( .A1(n36245), .A2(n33727), .ZN(n34604) );
  XNOR2_X1 U6322 ( .A(n36245), .B(\fmem_data[29][3] ), .ZN(n33595) );
  OR2_X1 U6323 ( .A1(n36245), .A2(n3587), .ZN(n31505) );
  OR2_X1 U6324 ( .A1(n36245), .A2(n3602), .ZN(n33951) );
  OR2_X1 U6325 ( .A1(n29470), .A2(n29469), .ZN(n29472) );
  NAND3_X1 U6326 ( .A1(n5189), .A2(n5188), .A3(n5187), .ZN(n5190) );
  NAND3_X1 U6327 ( .A1(n16075), .A2(n16074), .A3(n16073), .ZN(n16076) );
  NOR4_X1 U6328 ( .A1(n24478), .A2(n24477), .A3(n24476), .A4(n24475), .ZN(
        n24480) );
  NAND2_X1 U6329 ( .A1(n6993), .A2(load_xaddr_val[5]), .ZN(n6991) );
  NAND4_X2 U6330 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n35145)
         );
  NAND2_X1 U6331 ( .A1(n34966), .A2(n34965), .ZN(n34967) );
  OAI22_X1 U6332 ( .A1(n33184), .A2(n33642), .B1(n33183), .B2(n33643), .ZN(
        n33192) );
  OAI22_X1 U6333 ( .A1(n33184), .A2(n33643), .B1(n32562), .B2(n33642), .ZN(
        n26269) );
  BUF_X4 U6334 ( .A(n11489), .Z(n27710) );
  XNOR2_X1 U6335 ( .A(n31659), .B(\fmem_data[30][3] ), .ZN(n31997) );
  OR2_X1 U6336 ( .A1(n33036), .A2(n3870), .ZN(n31645) );
  XNOR2_X1 U6337 ( .A(n31511), .B(\fmem_data[16][7] ), .ZN(n33226) );
  OAI22_X1 U6338 ( .A1(n33226), .A2(n35753), .B1(n17851), .B2(n35752), .ZN(
        n19511) );
  XNOR2_X1 U6339 ( .A(n32898), .B(\fmem_data[8][7] ), .ZN(n31994) );
  OAI22_X1 U6340 ( .A1(n33964), .A2(n33961), .B1(n31993), .B2(n33963), .ZN(
        n32011) );
  OAI22_X1 U6341 ( .A1(n31994), .A2(n35729), .B1(n33256), .B2(n35730), .ZN(
        n32010) );
  XNOR2_X1 U6342 ( .A(n32899), .B(\fmem_data[8][7] ), .ZN(n33256) );
  OAI22_X1 U6343 ( .A1(n31951), .A2(n35760), .B1(n31950), .B2(n35761), .ZN(
        n32710) );
  OAI22_X1 U6344 ( .A1(n31443), .A2(n33059), .B1(n32079), .B2(n33057), .ZN(
        n31919) );
  OAI22_X1 U6345 ( .A1(n33164), .A2(n35182), .B1(n30815), .B2(n35181), .ZN(
        n22781) );
  OAI22_X1 U6346 ( .A1(n33946), .A2(n3577), .B1(n33778), .B2(n36196), .ZN(
        n31610) );
  BUF_X2 U6347 ( .A(n11561), .Z(n29667) );
  NAND2_X1 U6348 ( .A1(n35096), .A2(n35095), .ZN(n35097) );
  OAI22_X1 U6349 ( .A1(n30379), .A2(n33855), .B1(n32643), .B2(n33853), .ZN(
        n30454) );
  AOI21_X1 U6350 ( .B1(n33855), .B2(n33853), .A(n30379), .ZN(n5766) );
  OAI22_X1 U6351 ( .A1(n32725), .A2(n34941), .B1(n32724), .B2(n34942), .ZN(
        n32760) );
  XNOR2_X1 U6352 ( .A(n32938), .B(\fmem_data[1][5] ), .ZN(n32725) );
  XNOR2_X1 U6353 ( .A(n33150), .B(n34958), .ZN(n35059) );
  BUF_X4 U6354 ( .A(n11489), .Z(n29433) );
  OR2_X2 U6355 ( .A1(n7215), .A2(n10288), .ZN(n7421) );
  OAI21_X2 U6356 ( .B1(n7215), .B2(n6990), .A(n10589), .ZN(n8020) );
  NAND2_X1 U6357 ( .A1(n31838), .A2(n31837), .ZN(n31839) );
  OAI22_X1 U6358 ( .A1(n32021), .A2(n32780), .B1(n32020), .B2(n32779), .ZN(
        n33048) );
  XNOR2_X1 U6359 ( .A(n34982), .B(\fmem_data[25][7] ), .ZN(n35327) );
  NAND4_X1 U6360 ( .A1(n3407), .A2(n3408), .A3(n3409), .A4(n3410), .ZN(n29599)
         );
  AND4_X1 U6361 ( .A1(n29572), .A2(n29571), .A3(n29570), .A4(n29569), .ZN(
        n3407) );
  AND4_X1 U6362 ( .A1(n29578), .A2(n29577), .A3(n29576), .A4(n29575), .ZN(
        n3408) );
  AND4_X1 U6363 ( .A1(n29588), .A2(n29587), .A3(n29586), .A4(n29585), .ZN(
        n3409) );
  AND4_X1 U6364 ( .A1(n29597), .A2(n29596), .A3(n29595), .A4(n29594), .ZN(
        n3410) );
  XNOR2_X1 U6365 ( .A(n34630), .B(\fmem_data[14][5] ), .ZN(n32202) );
  XNOR2_X1 U6366 ( .A(n34630), .B(\fmem_data[14][3] ), .ZN(n33604) );
  XNOR2_X1 U6367 ( .A(n32317), .B(\fmem_data[4][5] ), .ZN(n34100) );
  OAI22_X1 U6368 ( .A1(n34100), .A2(n35010), .B1(n32318), .B2(n35011), .ZN(
        n33068) );
  OAI22_X1 U6369 ( .A1(n33950), .A2(n3566), .B1(n33949), .B2(n34529), .ZN(
        n34081) );
  XNOR2_X1 U6370 ( .A(n33555), .B(\fmem_data[21][5] ), .ZN(n34196) );
  INV_X1 U6371 ( .A(n3411), .ZN(n3412) );
  OR2_X1 U6372 ( .A1(n33844), .A2(n3689), .ZN(n32954) );
  AND2_X1 U6373 ( .A1(n3365), .A2(\fmem_data[9][0] ), .ZN(n36526) );
  OR2_X1 U6374 ( .A1(n33844), .A2(n3607), .ZN(n32431) );
  AND2_X1 U6375 ( .A1(n3365), .A2(n32577), .ZN(n32693) );
  AND2_X1 U6376 ( .A1(n33844), .A2(n31527), .ZN(n32962) );
  OR2_X1 U6377 ( .A1(n33844), .A2(n3608), .ZN(n33784) );
  OR2_X1 U6378 ( .A1(n3365), .A2(n3625), .ZN(n30493) );
  AND2_X1 U6379 ( .A1(n33844), .A2(n21394), .ZN(n33941) );
  OAI22_X1 U6380 ( .A1(n33966), .A2(n34422), .B1(n33965), .B2(n34424), .ZN(
        n34061) );
  NAND4_X1 U6381 ( .A1(n3415), .A2(n3416), .A3(n3417), .A4(n3418), .ZN(n12784)
         );
  AND4_X1 U6382 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n3415) );
  AND4_X1 U6383 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n3416) );
  AND4_X1 U6384 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n3417) );
  AND4_X1 U6385 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n3418) );
  OAI22_X1 U6386 ( .A1(n31671), .A2(n35712), .B1(n35711), .B2(n25146), .ZN(
        n31829) );
  NAND3_X1 U6387 ( .A1(n9173), .A2(n9172), .A3(n9171), .ZN(n9174) );
  XNOR2_X1 U6388 ( .A(n34670), .B(n34854), .ZN(n3419) );
  OR2_X2 U6389 ( .A1(n7215), .A2(n6992), .ZN(n6183) );
  BUF_X1 U6390 ( .A(n30259), .Z(n3421) );
  NOR2_X1 U6391 ( .A1(n6202), .A2(n3246), .ZN(n30259) );
  NAND2_X1 U6392 ( .A1(n16064), .A2(n16063), .ZN(n34982) );
  NAND2_X1 U6393 ( .A1(n35480), .A2(n35479), .ZN(n3422) );
  NAND2_X1 U6394 ( .A1(n37150), .A2(n37149), .ZN(n37218) );
  AOI22_X1 U6395 ( .A1(n28700), .A2(\xmem_data[50][5] ), .B1(n28137), .B2(
        \xmem_data[51][5] ), .ZN(n11959) );
  XNOR2_X1 U6396 ( .A(n32582), .B(\fmem_data[10][5] ), .ZN(n31999) );
  XNOR2_X1 U6397 ( .A(n33483), .B(\fmem_data[31][5] ), .ZN(n33880) );
  XNOR2_X1 U6398 ( .A(n33483), .B(\fmem_data[31][3] ), .ZN(n34471) );
  OAI22_X1 U6399 ( .A1(n30437), .A2(n35591), .B1(n33132), .B2(n35592), .ZN(
        n26029) );
  OAI22_X1 U6400 ( .A1(n33133), .A2(n35592), .B1(n33132), .B2(n35591), .ZN(
        n35045) );
  OAI22_X1 U6401 ( .A1(n34190), .A2(n36240), .B1(n34189), .B2(n3482), .ZN(
        n34310) );
  NAND4_X1 U6402 ( .A1(n18343), .A2(n18344), .A3(n18345), .A4(n18342), .ZN(
        n3425) );
  NAND4_X1 U6403 ( .A1(n18343), .A2(n18344), .A3(n18345), .A4(n18342), .ZN(
        n31513) );
  XOR2_X1 U6404 ( .A(n32767), .B(n32766), .Z(n3426) );
  XOR2_X1 U6405 ( .A(n32765), .B(n3426), .Z(n32824) );
  NAND2_X1 U6406 ( .A1(n32765), .A2(n32767), .ZN(n3427) );
  NAND2_X1 U6407 ( .A1(n32765), .A2(n32766), .ZN(n3428) );
  NAND2_X1 U6408 ( .A1(n32767), .A2(n32766), .ZN(n3429) );
  NAND3_X1 U6409 ( .A1(n3427), .A2(n3428), .A3(n3429), .ZN(n33290) );
  NAND3_X1 U6410 ( .A1(n17711), .A2(n17710), .A3(n17709), .ZN(n17712) );
  OAI22_X1 U6411 ( .A1(n32572), .A2(n34736), .B1(n32571), .B2(n33690), .ZN(
        n32800) );
  NAND2_X1 U6412 ( .A1(n32737), .A2(n32736), .ZN(n32738) );
  NOR2_X1 U6413 ( .A1(n37140), .A2(n37141), .ZN(n3435) );
  NOR2_X1 U6414 ( .A1(n37140), .A2(n37141), .ZN(n37259) );
  XOR2_X1 U6415 ( .A(n35784), .B(n35783), .Z(n3436) );
  OAI22_X1 U6416 ( .A1(n36297), .A2(n3564), .B1(n36296), .B2(n36295), .ZN(
        n36717) );
  XNOR2_X1 U6417 ( .A(n36296), .B(\fmem_data[0][7] ), .ZN(n31013) );
  AND2_X1 U6418 ( .A1(n36296), .A2(n32589), .ZN(n32785) );
  AND2_X1 U6419 ( .A1(n36296), .A2(\fmem_data[0][0] ), .ZN(n36558) );
  AND2_X1 U6420 ( .A1(n36296), .A2(n31535), .ZN(n33463) );
  AND2_X1 U6421 ( .A1(n36296), .A2(n17180), .ZN(n26273) );
  NAND4_X2 U6422 ( .A1(n17179), .A2(n17178), .A3(n17177), .A4(n17176), .ZN(
        n36296) );
  XNOR2_X1 U6423 ( .A(n32937), .B(\fmem_data[19][5] ), .ZN(n31395) );
  XNOR2_X1 U6424 ( .A(n35114), .B(\fmem_data[23][7] ), .ZN(n35259) );
  NAND2_X1 U6425 ( .A1(n4021), .A2(n4391), .ZN(n4058) );
  NAND2_X1 U6426 ( .A1(n33824), .A2(n33823), .ZN(n34115) );
  NAND4_X2 U6427 ( .A1(n27697), .A2(n27696), .A3(n27695), .A4(n27694), .ZN(
        n36311) );
  XNOR2_X1 U6428 ( .A(n8417), .B(n3402), .ZN(n8423) );
  AND2_X1 U6429 ( .A1(n8410), .A2(N345), .ZN(n4024) );
  XNOR2_X1 U6430 ( .A(n35326), .B(\fmem_data[25][7] ), .ZN(n35743) );
  OAI22_X1 U6431 ( .A1(n32514), .A2(n34986), .B1(n34047), .B2(n34985), .ZN(
        n33173) );
  XNOR2_X1 U6432 ( .A(n32513), .B(\fmem_data[25][5] ), .ZN(n34047) );
  NAND4_X1 U6433 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        n32513) );
  OAI22_X1 U6434 ( .A1(n33873), .A2(n33876), .B1(n31394), .B2(n33875), .ZN(
        n31577) );
  AND2_X1 U6435 ( .A1(n8933), .A2(n8934), .ZN(n8935) );
  NAND2_X1 U6436 ( .A1(n33885), .A2(n33884), .ZN(n34156) );
  OAI22_X1 U6437 ( .A1(n31976), .A2(n35655), .B1(n33135), .B2(n35656), .ZN(
        n33109) );
  NAND2_X1 U6438 ( .A1(n15585), .A2(n15584), .ZN(n32425) );
  OAI22_X1 U6439 ( .A1(n34112), .A2(n3931), .B1(n32439), .B2(n36216), .ZN(
        n31553) );
  OAI22_X1 U6440 ( .A1(n33702), .A2(n36216), .B1(n32439), .B2(n3931), .ZN(
        n32878) );
  OAI21_X1 U6441 ( .B1(n36773), .B2(n36775), .A(n36774), .ZN(n36179) );
  NAND2_X1 U6442 ( .A1(n36773), .A2(n36775), .ZN(n36178) );
  XNOR2_X1 U6443 ( .A(n3303), .B(\fmem_data[31][1] ), .ZN(n33702) );
  NAND4_X1 U6444 ( .A1(n3437), .A2(n3438), .A3(n3439), .A4(n3440), .ZN(n18382)
         );
  AND4_X1 U6445 ( .A1(n18369), .A2(n18368), .A3(n18367), .A4(n18366), .ZN(
        n3437) );
  AND4_X1 U6446 ( .A1(n18373), .A2(n18372), .A3(n18371), .A4(n18370), .ZN(
        n3438) );
  AND4_X1 U6447 ( .A1(n18377), .A2(n18376), .A3(n18375), .A4(n18374), .ZN(
        n3439) );
  AND4_X1 U6448 ( .A1(n18381), .A2(n18380), .A3(n18379), .A4(n18378), .ZN(
        n3440) );
  AND3_X1 U6449 ( .A1(n3441), .A2(n25005), .A3(n25006), .ZN(n25015) );
  AND4_X1 U6450 ( .A1(n25004), .A2(n25003), .A3(n25002), .A4(n25001), .ZN(
        n3441) );
  OAI21_X1 U6451 ( .B1(n34332), .B2(n34330), .A(n34331), .ZN(n33885) );
  OAI22_X1 U6452 ( .A1(n24335), .A2(n35515), .B1(n33315), .B2(n35516), .ZN(
        n11340) );
  XNOR2_X1 U6453 ( .A(n32586), .B(\fmem_data[12][7] ), .ZN(n33315) );
  XNOR2_X1 U6454 ( .A(n32025), .B(\fmem_data[12][7] ), .ZN(n24335) );
  XNOR2_X1 U6455 ( .A(n35336), .B(\fmem_data[2][7] ), .ZN(n35720) );
  XNOR2_X1 U6456 ( .A(n35336), .B(\fmem_data[2][1] ), .ZN(n33271) );
  OAI21_X1 U6457 ( .B1(n34682), .B2(n34683), .A(n34681), .ZN(n34685) );
  OAI22_X1 U6458 ( .A1(n34036), .A2(n35018), .B1(n34035), .B2(n35019), .ZN(
        n34244) );
  XNOR2_X1 U6459 ( .A(n31221), .B(\fmem_data[2][5] ), .ZN(n34035) );
  XNOR2_X1 U6460 ( .A(n33554), .B(\fmem_data[2][7] ), .ZN(n22777) );
  OAI22_X1 U6461 ( .A1(n31249), .A2(n34904), .B1(n31248), .B2(n34903), .ZN(
        n31563) );
  BUF_X2 U6462 ( .A(n11850), .Z(n27742) );
  OAI22_X1 U6463 ( .A1(n30442), .A2(n34420), .B1(n28403), .B2(n34418), .ZN(
        n17751) );
  OAI22_X1 U6464 ( .A1(n32195), .A2(n34418), .B1(n28403), .B2(n34420), .ZN(
        n28929) );
  OAI21_X1 U6465 ( .B1(n17749), .B2(n17750), .A(n17751), .ZN(n10945) );
  NAND4_X1 U6466 ( .A1(n21952), .A2(n21951), .A3(n21950), .A4(n21949), .ZN(
        n3442) );
  NAND4_X1 U6467 ( .A1(n21952), .A2(n21951), .A3(n21950), .A4(n21949), .ZN(
        n31383) );
  NAND2_X1 U6468 ( .A1(n24010), .A2(n27778), .ZN(n24011) );
  XNOR2_X1 U6469 ( .A(n3359), .B(\fmem_data[2][5] ), .ZN(n30158) );
  XNOR2_X1 U6470 ( .A(n3359), .B(\fmem_data[2][7] ), .ZN(n33325) );
  BUF_X2 U6471 ( .A(n7993), .Z(n3445) );
  BUF_X2 U6472 ( .A(n7993), .Z(n3446) );
  BUF_X2 U6473 ( .A(n7993), .Z(n3447) );
  NAND2_X1 U6474 ( .A1(n6189), .A2(n6196), .ZN(n7993) );
  AOI22_X1 U6475 ( .A1(n7445), .A2(n27737), .B1(n7444), .B2(n27778), .ZN(n7496) );
  NOR3_X1 U6476 ( .A1(n18250), .A2(n18249), .A3(n18248), .ZN(n18256) );
  NAND2_X1 U6477 ( .A1(n37270), .A2(n37269), .ZN(n37271) );
  XNOR2_X1 U6478 ( .A(n33756), .B(\fmem_data[28][5] ), .ZN(n32581) );
  XNOR2_X1 U6479 ( .A(n33756), .B(\fmem_data[28][3] ), .ZN(n33574) );
  XNOR2_X1 U6480 ( .A(n33756), .B(\fmem_data[28][7] ), .ZN(n31951) );
  OAI22_X1 U6481 ( .A1(n34020), .A2(n34412), .B1(n34413), .B2(n34410), .ZN(
        n31573) );
  NAND2_X1 U6482 ( .A1(n26251), .A2(n26250), .ZN(n33019) );
  NAND2_X1 U6483 ( .A1(n32560), .A2(n32557), .ZN(n3450) );
  NAND2_X1 U6484 ( .A1(n3275), .A2(n32557), .ZN(n3451) );
  NAND2_X1 U6485 ( .A1(n34174), .A2(n34173), .ZN(n34176) );
  XNOR2_X1 U6486 ( .A(n33676), .B(n33675), .ZN(n33818) );
  OAI22_X1 U6487 ( .A1(n34441), .A2(n34440), .B1(n34439), .B2(n3483), .ZN(
        n34522) );
  OAI22_X1 U6488 ( .A1(n32148), .A2(n3483), .B1(n34439), .B2(n34440), .ZN(
        n33889) );
  OAI22_X1 U6489 ( .A1(n33038), .A2(n35704), .B1(n31820), .B2(n35705), .ZN(
        n26026) );
  OAI22_X1 U6490 ( .A1(n33038), .A2(n35705), .B1(n33037), .B2(n35704), .ZN(
        n33063) );
  NAND2_X1 U6491 ( .A1(n33290), .A2(n33289), .ZN(n33291) );
  INV_X1 U6492 ( .A(n37216), .ZN(n37219) );
  NAND2_X1 U6493 ( .A1(n8100), .A2(n8099), .ZN(n3452) );
  OR2_X1 U6494 ( .A1(n26038), .A2(n26037), .ZN(n3453) );
  NAND2_X1 U6495 ( .A1(n3453), .A2(n26039), .ZN(n24837) );
  OAI22_X1 U6496 ( .A1(n31954), .A2(n35489), .B1(n31639), .B2(n35490), .ZN(
        n26037) );
  NAND2_X1 U6497 ( .A1(n35961), .A2(n35960), .ZN(n35951) );
  NOR2_X1 U6498 ( .A1(n35961), .A2(n35960), .ZN(n35953) );
  OAI22_X1 U6499 ( .A1(n33247), .A2(n35744), .B1(n35745), .B2(n34860), .ZN(
        n33379) );
  BUF_X1 U6500 ( .A(n6999), .Z(n8293) );
  NAND2_X1 U6501 ( .A1(n27305), .A2(n27304), .ZN(n27311) );
  OAI22_X1 U6502 ( .A1(n31197), .A2(n34908), .B1(n31196), .B2(n34909), .ZN(
        n31518) );
  XNOR2_X1 U6503 ( .A(n34361), .B(n3668), .ZN(n32141) );
  XNOR2_X1 U6504 ( .A(n34361), .B(n3674), .ZN(n34411) );
  NAND4_X1 U6505 ( .A1(n18531), .A2(n18530), .A3(n18529), .A4(n18528), .ZN(
        n3454) );
  NAND4_X1 U6506 ( .A1(n18531), .A2(n18530), .A3(n18529), .A4(n18528), .ZN(
        n31818) );
  OAI22_X1 U6507 ( .A1(n32154), .A2(n34919), .B1(n32153), .B2(n34918), .ZN(
        n32250) );
  NAND2_X1 U6508 ( .A1(n4031), .A2(n37199), .ZN(n4061) );
  XNOR2_X1 U6509 ( .A(n6173), .B(n37199), .ZN(n8422) );
  XNOR2_X1 U6510 ( .A(n3321), .B(\fmem_data[27][5] ), .ZN(n33168) );
  AOI22_X1 U6511 ( .A1(n30782), .A2(n7040), .B1(n30741), .B2(n7039), .ZN(n3455) );
  XNOR2_X1 U6512 ( .A(n34212), .B(n3323), .ZN(n34400) );
  OAI22_X1 U6513 ( .A1(n33968), .A2(n34208), .B1(n33061), .B2(n34206), .ZN(
        n32009) );
  NAND3_X1 U6514 ( .A1(n11120), .A2(n11119), .A3(n11118), .ZN(n11121) );
  OAI22_X1 U6515 ( .A1(n32016), .A2(n33328), .B1(n32006), .B2(n33326), .ZN(
        n30841) );
  OAI22_X1 U6516 ( .A1(n32006), .A2(n33328), .B1(n32564), .B2(n33326), .ZN(
        n32520) );
  NAND2_X1 U6517 ( .A1(n8732), .A2(n8731), .ZN(n32438) );
  XNOR2_X1 U6518 ( .A(n33009), .B(n33008), .ZN(n36149) );
  NAND2_X1 U6519 ( .A1(n31626), .A2(n31624), .ZN(n28925) );
  XNOR2_X1 U6520 ( .A(n31413), .B(n31412), .ZN(n31415) );
  OAI22_X1 U6521 ( .A1(n30347), .A2(n34505), .B1(n29542), .B2(n34503), .ZN(
        n34256) );
  NAND2_X1 U6522 ( .A1(n34715), .A2(n34714), .ZN(n34281) );
  BUF_X2 U6523 ( .A(n10861), .Z(n29753) );
  AOI21_X1 U6524 ( .B1(n30317), .B2(\xmem_data[61][4] ), .A(n6338), .ZN(n6340)
         );
  XNOR2_X1 U6525 ( .A(n33479), .B(\fmem_data[15][3] ), .ZN(n33731) );
  XNOR2_X1 U6526 ( .A(n32787), .B(\fmem_data[2][3] ), .ZN(n3456) );
  NAND2_X1 U6527 ( .A1(n31807), .A2(n31806), .ZN(n31808) );
  OAI22_X1 U6528 ( .A1(n33235), .A2(n35697), .B1(n33234), .B2(n35696), .ZN(
        n33332) );
  NAND3_X1 U6529 ( .A1(n6183), .A2(n3248), .A3(n6178), .ZN(n11362) );
  NAND2_X1 U6530 ( .A1(n8100), .A2(n8099), .ZN(n31246) );
  OAI22_X1 U6531 ( .A1(n30384), .A2(n34989), .B1(n23918), .B2(n34990), .ZN(
        n24840) );
  NAND2_X1 U6532 ( .A1(n36656), .A2(n36655), .ZN(n36444) );
  NAND2_X1 U6533 ( .A1(n33278), .A2(n33277), .ZN(n33279) );
  NOR2_X1 U6534 ( .A1(n4038), .A2(n9417), .ZN(n4039) );
  NAND2_X1 U6535 ( .A1(n8409), .A2(n4038), .ZN(n8417) );
  NAND2_X1 U6536 ( .A1(n4041), .A2(n4038), .ZN(n4080) );
  AND2_X1 U6537 ( .A1(n4038), .A2(N345), .ZN(n4031) );
  NAND2_X1 U6538 ( .A1(n34690), .A2(n34689), .ZN(n34889) );
  OAI21_X1 U6539 ( .B1(n34688), .B2(n34687), .A(n34686), .ZN(n34690) );
  NAND2_X1 U6540 ( .A1(n32919), .A2(n32918), .ZN(n32095) );
  NAND2_X1 U6541 ( .A1(n31769), .A2(n31768), .ZN(n31770) );
  NAND4_X1 U6542 ( .A1(n3458), .A2(n3459), .A3(n3460), .A4(n3461), .ZN(n10921)
         );
  AND4_X1 U6543 ( .A1(n10908), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n3458) );
  AND4_X1 U6544 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n3459) );
  AND4_X1 U6545 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n3460) );
  AND4_X1 U6546 ( .A1(n10920), .A2(n10919), .A3(n10918), .A4(n10917), .ZN(
        n3461) );
  NAND2_X1 U6547 ( .A1(n37148), .A2(n37147), .ZN(n37238) );
  AOI21_X1 U6548 ( .B1(n35619), .B2(n35618), .A(n35617), .ZN(n35620) );
  OAI22_X1 U6549 ( .A1(n35617), .A2(n35619), .B1(n35360), .B2(n35618), .ZN(
        n35735) );
  XNOR2_X1 U6550 ( .A(n35242), .B(\fmem_data[27][7] ), .ZN(n35640) );
  NAND2_X1 U6551 ( .A1(n3455), .A2(n7094), .ZN(n3462) );
  XNOR2_X1 U6552 ( .A(n33019), .B(\fmem_data[23][7] ), .ZN(n34240) );
  OAI22_X1 U6553 ( .A1(n34360), .A2(n36241), .B1(n3430), .B2(n3662), .ZN(
        n32874) );
  XNOR2_X1 U6554 ( .A(n36043), .B(n36042), .ZN(n36755) );
  OAI22_X1 U6555 ( .A1(n34240), .A2(n35651), .B1(n33020), .B2(n35652), .ZN(
        n33143) );
  NAND2_X1 U6556 ( .A1(n34123), .A2(n34122), .ZN(n33952) );
  AND2_X1 U6557 ( .A1(n7215), .A2(n4027), .ZN(n6169) );
  CLKBUF_X1 U6558 ( .A(n7215), .Z(n7423) );
  AOI21_X1 U6559 ( .B1(n30070), .B2(\xmem_data[102][1] ), .A(n23031), .ZN(
        n23032) );
  NAND2_X1 U6560 ( .A1(n31601), .A2(n31602), .ZN(n31237) );
  OAI22_X1 U6561 ( .A1(n35111), .A2(n35663), .B1(n31974), .B2(n35662), .ZN(
        n31679) );
  OAI22_X1 U6562 ( .A1(n35111), .A2(n35662), .B1(n35257), .B2(n35663), .ZN(
        n35139) );
  XNOR2_X1 U6563 ( .A(n32425), .B(\fmem_data[19][3] ), .ZN(n34192) );
  NAND2_X1 U6564 ( .A1(n36033), .A2(n36032), .ZN(n33016) );
  OAI22_X1 U6565 ( .A1(n35141), .A2(n35618), .B1(n35360), .B2(n35619), .ZN(
        n35169) );
  XNOR2_X1 U6566 ( .A(n33027), .B(\fmem_data[7][5] ), .ZN(n34233) );
  BUF_X1 U6567 ( .A(n34556), .Z(n3463) );
  BUF_X1 U6568 ( .A(n3464), .Z(n3465) );
  BUF_X1 U6569 ( .A(n29187), .Z(n3466) );
  NAND2_X1 U6570 ( .A1(n37101), .A2(n37100), .ZN(n37281) );
  NAND2_X1 U6571 ( .A1(n36728), .A2(n36727), .ZN(n36317) );
  XNOR2_X1 U6572 ( .A(n36728), .B(n36727), .ZN(n36730) );
  XNOR2_X1 U6573 ( .A(n36311), .B(\fmem_data[7][3] ), .ZN(n34504) );
  OR2_X1 U6574 ( .A1(n36311), .A2(n3648), .ZN(n31398) );
  OR2_X1 U6575 ( .A1(n36311), .A2(n3685), .ZN(n33722) );
  AND2_X1 U6576 ( .A1(n36311), .A2(n32881), .ZN(n36204) );
  AND2_X1 U6577 ( .A1(n36311), .A2(n27698), .ZN(n31216) );
  AND2_X1 U6578 ( .A1(n36311), .A2(\fmem_data[7][0] ), .ZN(n36726) );
  XNOR2_X1 U6579 ( .A(n34398), .B(n34397), .ZN(n34799) );
  OAI22_X1 U6580 ( .A1(n32732), .A2(n3575), .B1(n32731), .B2(n36120), .ZN(
        n33206) );
  XNOR2_X1 U6581 ( .A(n35357), .B(\fmem_data[29][1] ), .ZN(n32732) );
  NAND2_X1 U6582 ( .A1(n34180), .A2(n34179), .ZN(n27304) );
  OAI21_X1 U6583 ( .B1(n34180), .B2(n34179), .A(n34181), .ZN(n27305) );
  XNOR2_X1 U6584 ( .A(n36632), .B(n36631), .ZN(n36634) );
  OAI22_X1 U6585 ( .A1(n34484), .A2(n3576), .B1(n34623), .B2(n34483), .ZN(
        n36330) );
  OR2_X1 U6586 ( .A1(n34623), .A2(n3694), .ZN(n32956) );
  XNOR2_X1 U6587 ( .A(n34623), .B(\fmem_data[5][3] ), .ZN(n32423) );
  OR2_X1 U6588 ( .A1(n34623), .A2(n3623), .ZN(n27973) );
  XNOR2_X1 U6589 ( .A(n34623), .B(\fmem_data[5][5] ), .ZN(n33858) );
  AND2_X1 U6590 ( .A1(n34623), .A2(n33960), .ZN(n34068) );
  AND2_X1 U6591 ( .A1(n34623), .A2(n32121), .ZN(n32685) );
  AND2_X1 U6592 ( .A1(n34623), .A2(n31582), .ZN(n32957) );
  AND2_X1 U6593 ( .A1(n34623), .A2(\fmem_data[5][0] ), .ZN(n36521) );
  NAND4_X1 U6594 ( .A1(n3467), .A2(n3468), .A3(n3469), .A4(n3470), .ZN(n10938)
         );
  AND4_X1 U6595 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n3467) );
  AND4_X1 U6596 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n3468) );
  AND4_X1 U6597 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n3469) );
  AND4_X1 U6598 ( .A1(n10937), .A2(n10936), .A3(n10935), .A4(n10934), .ZN(
        n3470) );
  XNOR2_X1 U6599 ( .A(n35030), .B(\fmem_data[15][5] ), .ZN(n23918) );
  OAI22_X1 U6600 ( .A1(n34988), .A2(n34990), .B1(n23918), .B2(n34989), .ZN(
        n31785) );
  XNOR2_X1 U6601 ( .A(n31940), .B(\fmem_data[23][7] ), .ZN(n35115) );
  XNOR2_X1 U6602 ( .A(n31940), .B(\fmem_data[23][1] ), .ZN(n33905) );
  XNOR2_X1 U6603 ( .A(n31940), .B(\fmem_data[23][5] ), .ZN(n34235) );
  NAND2_X1 U6604 ( .A1(n7496), .A2(n7495), .ZN(n35242) );
  XNOR2_X1 U6605 ( .A(n35242), .B(\fmem_data[27][1] ), .ZN(n32168) );
  OR2_X1 U6606 ( .A1(n32168), .A2(n17754), .ZN(n23582) );
  OAI22_X1 U6607 ( .A1(n32168), .A2(n3482), .B1(n34189), .B2(n36240), .ZN(
        n32196) );
  NAND2_X1 U6608 ( .A1(n37250), .A2(n37252), .ZN(n37188) );
  INV_X1 U6609 ( .A(n37250), .ZN(n37251) );
  OAI22_X1 U6610 ( .A1(n36337), .A2(n36226), .B1(n3633), .B2(n36225), .ZN(
        n36693) );
  OR2_X1 U6611 ( .A1(n36337), .A2(n3717), .ZN(n36214) );
  OR2_X1 U6612 ( .A1(n36337), .A2(n3686), .ZN(n34337) );
  AND2_X1 U6613 ( .A1(n36337), .A2(n32901), .ZN(n36236) );
  XNOR2_X1 U6614 ( .A(n36337), .B(\fmem_data[19][5] ), .ZN(n31396) );
  OR2_X1 U6615 ( .A1(n36337), .A2(n3606), .ZN(n31225) );
  OR2_X1 U6616 ( .A1(n36337), .A2(n3640), .ZN(n32106) );
  AND2_X1 U6617 ( .A1(n36337), .A2(n33830), .ZN(n34509) );
  AND2_X1 U6618 ( .A1(n36337), .A2(n29844), .ZN(n31135) );
  NAND2_X1 U6619 ( .A1(n35304), .A2(n35303), .ZN(n35306) );
  XNOR2_X1 U6620 ( .A(n35911), .B(n35539), .ZN(n35950) );
  XNOR2_X1 U6621 ( .A(n33246), .B(\fmem_data[25][1] ), .ZN(n34439) );
  NOR2_X2 U6622 ( .A1(n3457), .A2(n7408), .ZN(n8700) );
  OAI22_X1 U6623 ( .A1(n32514), .A2(n34985), .B1(n33041), .B2(n34986), .ZN(
        n31006) );
  BUF_X2 U6624 ( .A(n25604), .Z(n30885) );
  NOR2_X2 U6625 ( .A1(n4058), .A2(n10972), .ZN(n4478) );
  INV_X2 U6626 ( .A(n4399), .ZN(n14976) );
  BUF_X2 U6627 ( .A(n14976), .Z(n20782) );
  BUF_X2 U6628 ( .A(n14976), .Z(n20734) );
  BUF_X2 U6629 ( .A(n13415), .Z(n25398) );
  BUF_X2 U6630 ( .A(n13486), .Z(n25582) );
  BUF_X2 U6631 ( .A(n13486), .Z(n24685) );
  BUF_X2 U6632 ( .A(n14883), .Z(n28098) );
  BUF_X2 U6633 ( .A(n14981), .Z(n27526) );
  BUF_X2 U6634 ( .A(n4158), .Z(n28428) );
  BUF_X2 U6635 ( .A(n13436), .Z(n30514) );
  BUF_X2 U6636 ( .A(n13436), .Z(n31268) );
  BUF_X2 U6637 ( .A(n13476), .Z(n17041) );
  BUF_X2 U6638 ( .A(n13149), .Z(n23717) );
  BUF_X2 U6639 ( .A(n14937), .Z(n24509) );
  BUF_X2 U6640 ( .A(n14937), .Z(n20585) );
  BUF_X2 U6641 ( .A(n14925), .Z(n23739) );
  BUF_X1 U6642 ( .A(n4236), .Z(n10977) );
  BUF_X2 U6643 ( .A(n13469), .Z(n24695) );
  BUF_X2 U6644 ( .A(n13469), .Z(n20500) );
  BUF_X2 U6645 ( .A(n14989), .Z(n20723) );
  NOR2_X1 U6646 ( .A1(n8005), .A2(n11358), .ZN(n8073) );
  BUF_X2 U6647 ( .A(n13486), .Z(n29325) );
  BUF_X2 U6648 ( .A(n14926), .Z(n27938) );
  BUF_X1 U6649 ( .A(n14934), .Z(n28416) );
  BUF_X1 U6650 ( .A(n4177), .Z(n13435) );
  BUF_X1 U6651 ( .A(n14934), .Z(n28515) );
  BUF_X2 U6652 ( .A(n13420), .Z(n29298) );
  INV_X2 U6653 ( .A(n4444), .ZN(n13188) );
  BUF_X2 U6654 ( .A(n14913), .Z(n29238) );
  NOR2_X1 U6655 ( .A1(n8005), .A2(n11359), .ZN(n8074) );
  BUF_X2 U6656 ( .A(n14882), .Z(n23778) );
  BUF_X2 U6657 ( .A(n14999), .Z(n22703) );
  BUF_X2 U6658 ( .A(n14898), .Z(n24160) );
  BUF_X2 U6659 ( .A(n28947), .Z(n28037) );
  INV_X2 U6660 ( .A(n4368), .ZN(n28947) );
  AND4_X1 U6661 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n3471) );
  AND4_X1 U6662 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n3472) );
  BUF_X2 U6663 ( .A(n4478), .Z(n27551) );
  BUF_X2 U6664 ( .A(n14883), .Z(n24622) );
  INV_X2 U6665 ( .A(n4489), .ZN(n14975) );
  BUF_X2 U6666 ( .A(n14970), .Z(n29048) );
  BUF_X2 U6667 ( .A(n13468), .Z(n31347) );
  BUF_X1 U6668 ( .A(n3324), .Z(n24220) );
  BUF_X1 U6669 ( .A(n28947), .Z(n22752) );
  BUF_X2 U6670 ( .A(n28947), .Z(n29118) );
  AND4_X1 U6671 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n3473) );
  AND4_X1 U6672 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n3474) );
  AND4_X1 U6673 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n3475) );
  AND4_X1 U6674 ( .A1(n8085), .A2(n8084), .A3(n8083), .A4(n8082), .ZN(n3476)
         );
  AND4_X1 U6675 ( .A1(n26834), .A2(n26833), .A3(n26832), .A4(n26831), .ZN(
        n3477) );
  AND4_X1 U6676 ( .A1(n27077), .A2(n27082), .A3(n27081), .A4(n3548), .ZN(n3478) );
  AND4_X1 U6677 ( .A1(n15586), .A2(n15591), .A3(n15590), .A4(n3547), .ZN(n3479) );
  AND4_X1 U6678 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n3480)
         );
  AND3_X1 U6679 ( .A1(n24875), .A2(n24874), .A3(n24873), .ZN(n3481) );
  BUF_X2 U6680 ( .A(n13149), .Z(n21007) );
  INV_X2 U6681 ( .A(n4399), .ZN(n13486) );
  BUF_X2 U6682 ( .A(n26543), .Z(n30664) );
  BUF_X2 U6683 ( .A(n11484), .Z(n30280) );
  BUF_X2 U6684 ( .A(n14989), .Z(n25562) );
  BUF_X2 U6685 ( .A(n14875), .Z(n25360) );
  BUF_X2 U6686 ( .A(n14890), .Z(n30882) );
  BUF_X2 U6687 ( .A(n10456), .Z(n20769) );
  BUF_X2 U6688 ( .A(n14875), .Z(n27437) );
  INV_X2 U6689 ( .A(n4178), .ZN(n14937) );
  BUF_X2 U6690 ( .A(n4478), .Z(n23813) );
  BUF_X2 U6691 ( .A(n4478), .Z(n28374) );
  BUF_X2 U6692 ( .A(n14983), .Z(n30589) );
  BUF_X2 U6693 ( .A(n11780), .Z(n30293) );
  BUF_X2 U6694 ( .A(n4527), .Z(n14982) );
  BUF_X1 U6695 ( .A(n13420), .Z(n27568) );
  BUF_X2 U6696 ( .A(n14982), .Z(n30674) );
  BUF_X2 U6697 ( .A(n14982), .Z(n21060) );
  BUF_X1 U6698 ( .A(n14881), .Z(n29189) );
  BUF_X2 U6699 ( .A(n8088), .Z(n29786) );
  BUF_X1 U6700 ( .A(n3324), .Z(n24190) );
  BUF_X1 U6701 ( .A(n3324), .Z(n28460) );
  BUF_X2 U6702 ( .A(n14933), .Z(n28415) );
  BUF_X2 U6703 ( .A(n14933), .Z(n27943) );
  BUF_X2 U6704 ( .A(n14996), .Z(n29180) );
  BUF_X2 U6705 ( .A(n28974), .Z(n28317) );
  BUF_X1 U6706 ( .A(n28974), .Z(n24525) );
  INV_X2 U6707 ( .A(n8410), .ZN(n6173) );
  INV_X1 U6708 ( .A(n35739), .ZN(n27324) );
  OR2_X1 U6709 ( .A1(n33056), .A2(n3835), .ZN(n3491) );
  OR2_X1 U6710 ( .A1(n30353), .A2(n3872), .ZN(n3492) );
  OR2_X1 U6711 ( .A1(n32013), .A2(n3871), .ZN(n3493) );
  AND2_X1 U6712 ( .A1(n33576), .A2(n31491), .ZN(n3494) );
  OR2_X1 U6713 ( .A1(n32015), .A2(n3878), .ZN(n3495) );
  OR2_X1 U6714 ( .A1(n34837), .A2(n3876), .ZN(n3496) );
  AND4_X1 U6715 ( .A1(n11704), .A2(n11703), .A3(n11702), .A4(n11701), .ZN(
        n3497) );
  AND2_X1 U6716 ( .A1(n28510), .A2(\xmem_data[119][3] ), .ZN(n3498) );
  AND2_X1 U6717 ( .A1(n28510), .A2(\xmem_data[14][5] ), .ZN(n3499) );
  AND4_X1 U6718 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n3500)
         );
  AND4_X1 U6719 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n3501)
         );
  AND4_X1 U6720 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(n3502)
         );
  AND4_X1 U6721 ( .A1(n15874), .A2(n15873), .A3(n15872), .A4(n15871), .ZN(
        n3503) );
  AND2_X1 U6722 ( .A1(n25425), .A2(\xmem_data[12][5] ), .ZN(n3504) );
  AND4_X1 U6723 ( .A1(n16994), .A2(n16993), .A3(n16992), .A4(n16991), .ZN(
        n3505) );
  AND4_X1 U6724 ( .A1(n27373), .A2(n27372), .A3(n27371), .A4(n27370), .ZN(
        n3506) );
  AND4_X1 U6725 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n3507)
         );
  AND4_X1 U6726 ( .A1(n24777), .A2(n24776), .A3(n24775), .A4(n24774), .ZN(
        n3508) );
  AND4_X1 U6727 ( .A1(n6617), .A2(n6618), .A3(n6616), .A4(n6615), .ZN(n3509)
         );
  AND4_X1 U6728 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n3510)
         );
  AND4_X1 U6729 ( .A1(n17690), .A2(n17689), .A3(n17688), .A4(n17687), .ZN(
        n3511) );
  AND4_X1 U6730 ( .A1(n27734), .A2(n27733), .A3(n27732), .A4(n27731), .ZN(
        n3512) );
  AND4_X1 U6731 ( .A1(n29720), .A2(n29719), .A3(n29718), .A4(n29717), .ZN(
        n3513) );
  AND4_X1 U6732 ( .A1(n24505), .A2(n24504), .A3(n24503), .A4(n24502), .ZN(
        n3514) );
  AND4_X1 U6733 ( .A1(n28792), .A2(n28791), .A3(n28790), .A4(n28789), .ZN(
        n3515) );
  AND4_X1 U6734 ( .A1(n29140), .A2(n29139), .A3(n29138), .A4(n29137), .ZN(
        n3516) );
  AND4_X1 U6735 ( .A1(n14844), .A2(n14843), .A3(n14842), .A4(n14841), .ZN(
        n3517) );
  AND4_X1 U6736 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n3518)
         );
  AND4_X1 U6737 ( .A1(n7931), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n3519)
         );
  AND4_X1 U6738 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n3520)
         );
  AND4_X1 U6739 ( .A1(n24822), .A2(n24821), .A3(n24820), .A4(n24819), .ZN(
        n3521) );
  AND4_X1 U6740 ( .A1(n14484), .A2(n14483), .A3(n14482), .A4(n14481), .ZN(
        n3522) );
  AND4_X1 U6741 ( .A1(n27775), .A2(n27774), .A3(n27773), .A4(n27772), .ZN(
        n3523) );
  AND4_X1 U6742 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n3524)
         );
  AND4_X1 U6743 ( .A1(n28200), .A2(n28199), .A3(n28198), .A4(n28197), .ZN(
        n3525) );
  AND4_X1 U6744 ( .A1(n7560), .A2(n7559), .A3(n7558), .A4(n7557), .ZN(n3526)
         );
  AND4_X1 U6745 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n3527)
         );
  AND4_X1 U6746 ( .A1(n16081), .A2(n16080), .A3(n16079), .A4(n16078), .ZN(
        n3528) );
  AND4_X1 U6747 ( .A1(n26820), .A2(n26819), .A3(n26818), .A4(n26817), .ZN(
        n3529) );
  AND4_X1 U6748 ( .A1(n9179), .A2(n9178), .A3(n9177), .A4(n9176), .ZN(n3530)
         );
  AND4_X1 U6749 ( .A1(n21301), .A2(n21300), .A3(n21299), .A4(n21298), .ZN(
        n3531) );
  AND4_X1 U6750 ( .A1(n21994), .A2(n21993), .A3(n21992), .A4(n21991), .ZN(
        n3532) );
  AND4_X1 U6751 ( .A1(n23125), .A2(n23124), .A3(n23123), .A4(n23122), .ZN(
        n3533) );
  AND4_X1 U6752 ( .A1(n7579), .A2(n7578), .A3(n7577), .A4(n7576), .ZN(n3534)
         );
  AND4_X1 U6753 ( .A1(n13769), .A2(n13768), .A3(n13767), .A4(n13766), .ZN(
        n3535) );
  AND4_X1 U6754 ( .A1(n29653), .A2(n29652), .A3(n29651), .A4(n29650), .ZN(
        n3536) );
  AND4_X1 U6755 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n3537) );
  AND4_X1 U6756 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n3538) );
  AND4_X1 U6757 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n3539) );
  AND4_X1 U6758 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n3540) );
  AND4_X1 U6759 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n3541)
         );
  AND4_X1 U6760 ( .A1(n16487), .A2(n16486), .A3(n16485), .A4(n16484), .ZN(
        n3542) );
  AND4_X1 U6761 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n3543) );
  AND4_X1 U6762 ( .A1(n18198), .A2(n18197), .A3(n18196), .A4(n18195), .ZN(
        n3544) );
  AND4_X1 U6763 ( .A1(n22255), .A2(n22254), .A3(n22253), .A4(n22252), .ZN(
        n3545) );
  AND4_X1 U6764 ( .A1(n15837), .A2(n15836), .A3(n15835), .A4(n15834), .ZN(
        n3546) );
  AND3_X1 U6765 ( .A1(n15589), .A2(n15588), .A3(n15587), .ZN(n3547) );
  AND3_X1 U6766 ( .A1(n27080), .A2(n27079), .A3(n27078), .ZN(n3548) );
  NOR3_X1 U6767 ( .A1(n20658), .A2(n20657), .A3(n3911), .ZN(n3549) );
  AND3_X1 U6768 ( .A1(n18227), .A2(n18226), .A3(n18225), .ZN(n3550) );
  AND3_X1 U6769 ( .A1(n3525), .A2(n28204), .A3(n28203), .ZN(n3551) );
  AND2_X1 U6770 ( .A1(n15595), .A2(n15594), .ZN(n3552) );
  AND2_X1 U6771 ( .A1(n4682), .A2(n4681), .ZN(n3553) );
  AND3_X1 U6772 ( .A1(n24880), .A2(n24879), .A3(n24878), .ZN(n3554) );
  NAND2_X1 U6773 ( .A1(\fmem_data[21][1] ), .A2(n3570), .ZN(n34613) );
  NAND2_X1 U6774 ( .A1(n28373), .A2(\xmem_data[15][0] ), .ZN(n3555) );
  NAND2_X1 U6775 ( .A1(n29350), .A2(\xmem_data[8][3] ), .ZN(n3556) );
  AND3_X1 U6776 ( .A1(n20309), .A2(n20308), .A3(n20307), .ZN(n3557) );
  BUF_X2 U6777 ( .A(n14990), .Z(n20725) );
  BUF_X2 U6778 ( .A(n4078), .Z(n14990) );
  BUF_X2 U6779 ( .A(n6309), .Z(n30258) );
  BUF_X2 U6780 ( .A(n6281), .Z(n30304) );
  INV_X2 U6781 ( .A(n4178), .ZN(n13149) );
  BUF_X2 U6782 ( .A(n15011), .Z(n29103) );
  INV_X1 U6783 ( .A(n4242), .ZN(n14913) );
  BUF_X2 U6784 ( .A(n14981), .Z(n28468) );
  BUF_X2 U6785 ( .A(n14919), .Z(n28500) );
  BUF_X1 U6786 ( .A(n14981), .Z(n25527) );
  BUF_X1 U6787 ( .A(n4527), .Z(n13127) );
  BUF_X1 U6788 ( .A(n28947), .Z(n25357) );
  BUF_X1 U6789 ( .A(n11437), .Z(n30730) );
  BUF_X1 U6790 ( .A(n11437), .Z(n28145) );
  OR2_X1 U6791 ( .A1(n32178), .A2(n16358), .ZN(n3586) );
  BUF_X1 U6792 ( .A(n11780), .Z(n29798) );
  OR2_X1 U6793 ( .A1(n33170), .A2(n24114), .ZN(n3618) );
  BUF_X1 U6794 ( .A(n3324), .Z(n20593) );
  BUF_X1 U6795 ( .A(n10999), .Z(n30854) );
  INV_X2 U6796 ( .A(n4536), .ZN(n13475) );
  BUF_X1 U6797 ( .A(n10977), .Z(n29023) );
  BUF_X1 U6798 ( .A(n15000), .Z(n20586) );
  BUF_X1 U6799 ( .A(n14936), .Z(n20543) );
  BUF_X1 U6800 ( .A(n15000), .Z(n25383) );
  BUF_X1 U6801 ( .A(n15000), .Z(n30615) );
  OR2_X1 U6802 ( .A1(n4050), .A2(n4058), .ZN(n3676) );
  BUF_X1 U6803 ( .A(n8293), .Z(n30775) );
  AND4_X1 U6804 ( .A1(n17668), .A2(n17667), .A3(n17666), .A4(n17665), .ZN(
        n3702) );
  AND4_X1 U6805 ( .A1(n16312), .A2(n16311), .A3(n16310), .A4(n16309), .ZN(
        n3703) );
  OR2_X1 U6806 ( .A1(n30446), .A2(n4157), .ZN(n3704) );
  OR2_X1 U6807 ( .A1(n33196), .A2(n33195), .ZN(n3705) );
  AND4_X1 U6808 ( .A1(n24269), .A2(n24268), .A3(n24267), .A4(n24266), .ZN(
        n3706) );
  OR2_X1 U6809 ( .A1(n31943), .A2(n31942), .ZN(n3707) );
  OR2_X1 U6810 ( .A1(n37099), .A2(n37098), .ZN(n3708) );
  AND4_X1 U6811 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n3709) );
  AND2_X1 U6812 ( .A1(n10455), .A2(n10454), .ZN(n3710) );
  AND4_X1 U6813 ( .A1(n29194), .A2(n29193), .A3(n29192), .A4(n29191), .ZN(
        n3711) );
  AND4_X1 U6814 ( .A1(n5624), .A2(n5623), .A3(n5622), .A4(n5621), .ZN(n3712)
         );
  AND4_X1 U6815 ( .A1(n21984), .A2(n21983), .A3(n21982), .A4(n21981), .ZN(
        n3713) );
  OR2_X1 U6816 ( .A1(n34947), .A2(n34946), .ZN(n3714) );
  NOR4_X1 U6817 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n3715) );
  OR2_X1 U6818 ( .A1(n11213), .A2(n27573), .ZN(n3716) );
  OR2_X1 U6819 ( .A1(n29305), .A2(n29341), .ZN(n3718) );
  OR2_X1 U6820 ( .A1(n28826), .A2(n30879), .ZN(n3719) );
  OR2_X1 U6821 ( .A1(n12152), .A2(n12151), .ZN(n3720) );
  NAND2_X1 U6822 ( .A1(n6011), .A2(n24236), .ZN(n3721) );
  OR3_X1 U6823 ( .A1(n17138), .A2(n17137), .A3(n17136), .ZN(n3722) );
  OR2_X1 U6824 ( .A1(n14911), .A2(n15043), .ZN(n3723) );
  OR2_X1 U6825 ( .A1(n17089), .A2(n17088), .ZN(n3724) );
  AND2_X1 U6826 ( .A1(n24657), .A2(\xmem_data[30][6] ), .ZN(n3725) );
  NAND2_X1 U6827 ( .A1(n3222), .A2(\xmem_data[3][3] ), .ZN(n3726) );
  AND4_X1 U6828 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n3727) );
  OR2_X1 U6829 ( .A1(n30364), .A2(n30363), .ZN(n3728) );
  OR2_X1 U6830 ( .A1(n32181), .A2(n22456), .ZN(n3729) );
  OR2_X1 U6831 ( .A1(n33062), .A2(n25839), .ZN(n3730) );
  NAND2_X1 U6832 ( .A1(n13434), .A2(n24508), .ZN(n3731) );
  AND2_X1 U6833 ( .A1(n24443), .A2(\xmem_data[2][4] ), .ZN(n3733) );
  AND2_X1 U6834 ( .A1(n29103), .A2(\xmem_data[1][6] ), .ZN(n3734) );
  AND2_X1 U6835 ( .A1(n3231), .A2(\xmem_data[3][0] ), .ZN(n3736) );
  AND2_X1 U6836 ( .A1(n3433), .A2(\xmem_data[9][4] ), .ZN(n3737) );
  AND4_X1 U6837 ( .A1(n25479), .A2(n25478), .A3(n25477), .A4(n25476), .ZN(
        n3738) );
  AND2_X1 U6838 ( .A1(n29173), .A2(\xmem_data[10][0] ), .ZN(n3739) );
  AND2_X1 U6839 ( .A1(n30309), .A2(\xmem_data[51][3] ), .ZN(n3741) );
  AND2_X1 U6840 ( .A1(n27547), .A2(\xmem_data[21][0] ), .ZN(n3742) );
  AND4_X1 U6841 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n3743)
         );
  AND4_X1 U6842 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        n3744) );
  AND4_X1 U6843 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n13264), .ZN(
        n3745) );
  AND4_X1 U6844 ( .A1(n15024), .A2(n15023), .A3(n15022), .A4(n15021), .ZN(
        n3746) );
  AND4_X1 U6845 ( .A1(n28553), .A2(n28552), .A3(n28551), .A4(n28550), .ZN(
        n3747) );
  AND4_X1 U6846 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n3748) );
  AND4_X1 U6847 ( .A1(n28413), .A2(n28412), .A3(n28411), .A4(n28410), .ZN(
        n3749) );
  AND4_X1 U6848 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n3750) );
  AND4_X1 U6849 ( .A1(n5518), .A2(n5517), .A3(n5516), .A4(n5515), .ZN(n3751)
         );
  AND4_X1 U6850 ( .A1(n11135), .A2(n11134), .A3(n11133), .A4(n11132), .ZN(
        n3752) );
  AND4_X1 U6851 ( .A1(n8753), .A2(n8752), .A3(n8751), .A4(n8750), .ZN(n3753)
         );
  AND4_X1 U6852 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n3754) );
  AND4_X1 U6853 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n3755)
         );
  AND4_X1 U6854 ( .A1(n18269), .A2(n18268), .A3(n18267), .A4(n18266), .ZN(
        n3756) );
  AND4_X1 U6855 ( .A1(n29444), .A2(n29443), .A3(n29442), .A4(n29441), .ZN(
        n3757) );
  AND4_X1 U6856 ( .A1(n19835), .A2(n19834), .A3(n19833), .A4(n19832), .ZN(
        n3758) );
  AND4_X1 U6857 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n3759)
         );
  AND4_X1 U6858 ( .A1(n16292), .A2(n16291), .A3(n16290), .A4(n16289), .ZN(
        n3760) );
  AND4_X1 U6859 ( .A1(n14819), .A2(n14818), .A3(n14817), .A4(n14816), .ZN(
        n3761) );
  AND4_X1 U6860 ( .A1(n24804), .A2(n24803), .A3(n24802), .A4(n24801), .ZN(
        n3762) );
  AND4_X1 U6861 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n3763) );
  AND4_X1 U6862 ( .A1(n24751), .A2(n24750), .A3(n24749), .A4(n24748), .ZN(
        n3764) );
  AND4_X1 U6863 ( .A1(n26450), .A2(n26449), .A3(n26448), .A4(n26447), .ZN(
        n3765) );
  AND4_X1 U6864 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n3766)
         );
  AND4_X1 U6865 ( .A1(n20479), .A2(n20478), .A3(n20477), .A4(n20476), .ZN(
        n3767) );
  AND4_X1 U6866 ( .A1(n7312), .A2(n7311), .A3(n7310), .A4(n7309), .ZN(n3768)
         );
  AND4_X1 U6867 ( .A1(n29730), .A2(n29729), .A3(n29728), .A4(n29727), .ZN(
        n3769) );
  AND4_X1 U6868 ( .A1(n26571), .A2(n26570), .A3(n26569), .A4(n26568), .ZN(
        n3770) );
  AND4_X1 U6869 ( .A1(n7532), .A2(n7531), .A3(n7530), .A4(n7529), .ZN(n3771)
         );
  AND4_X1 U6870 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n3772)
         );
  AND4_X1 U6871 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n3773)
         );
  AND4_X1 U6872 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n3774)
         );
  AND4_X1 U6873 ( .A1(n10876), .A2(n10875), .A3(n10874), .A4(n10873), .ZN(
        n3775) );
  AND4_X1 U6874 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n3776) );
  AND4_X1 U6875 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n3777) );
  AND4_X1 U6876 ( .A1(n15810), .A2(n15809), .A3(n15808), .A4(n15807), .ZN(
        n3778) );
  AND4_X1 U6877 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n3779)
         );
  AND4_X1 U6878 ( .A1(n29493), .A2(n29492), .A3(n29491), .A4(n29490), .ZN(
        n3780) );
  AND4_X1 U6879 ( .A1(n8363), .A2(n8362), .A3(n8361), .A4(n8360), .ZN(n3781)
         );
  AND4_X1 U6880 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n3782)
         );
  AND4_X1 U6881 ( .A1(n26866), .A2(n26865), .A3(n26864), .A4(n26863), .ZN(
        n3783) );
  AND4_X1 U6882 ( .A1(n9510), .A2(n9509), .A3(n9508), .A4(n9507), .ZN(n3784)
         );
  AND4_X1 U6883 ( .A1(n26345), .A2(n26344), .A3(n26343), .A4(n26342), .ZN(
        n3785) );
  AND4_X1 U6884 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n3786) );
  AND4_X1 U6885 ( .A1(n17171), .A2(n17170), .A3(n17169), .A4(n17168), .ZN(
        n3787) );
  AND4_X1 U6886 ( .A1(n21321), .A2(n21320), .A3(n21319), .A4(n21318), .ZN(
        n3788) );
  AND4_X1 U6887 ( .A1(n24773), .A2(n24772), .A3(n24771), .A4(n24770), .ZN(
        n3789) );
  AND4_X1 U6888 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n3790)
         );
  AND4_X1 U6889 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n8813), .ZN(n3791)
         );
  AND4_X1 U6890 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n3792) );
  AND4_X1 U6891 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n3793)
         );
  AND4_X1 U6892 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n3794)
         );
  AND4_X1 U6893 ( .A1(n14840), .A2(n14839), .A3(n14838), .A4(n14837), .ZN(
        n3795) );
  AND4_X1 U6894 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n3796)
         );
  AND4_X1 U6895 ( .A1(n27792), .A2(n27791), .A3(n27790), .A4(n27789), .ZN(
        n3797) );
  AND4_X1 U6896 ( .A1(n7731), .A2(n7730), .A3(n7729), .A4(n7728), .ZN(n3798)
         );
  AND4_X1 U6897 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n3799) );
  AND4_X1 U6898 ( .A1(n26816), .A2(n26815), .A3(n26814), .A4(n26813), .ZN(
        n3800) );
  AND4_X1 U6899 ( .A1(n16343), .A2(n16342), .A3(n16341), .A4(n16340), .ZN(
        n3801) );
  AND4_X1 U6900 ( .A1(n25874), .A2(n25873), .A3(n25872), .A4(n25871), .ZN(
        n3802) );
  AND4_X1 U6901 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n3803) );
  AND4_X1 U6902 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n3804) );
  AND2_X1 U6903 ( .A1(n25492), .A2(\xmem_data[10][2] ), .ZN(n3805) );
  AND4_X1 U6904 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n3806)
         );
  AND4_X1 U6905 ( .A1(n17704), .A2(n17703), .A3(n17702), .A4(n17701), .ZN(
        n3807) );
  AND4_X1 U6906 ( .A1(n29099), .A2(n29098), .A3(n29097), .A4(n29096), .ZN(
        n3808) );
  AND4_X1 U6907 ( .A1(n27722), .A2(n27721), .A3(n27720), .A4(n27719), .ZN(
        n3809) );
  AND4_X1 U6908 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(
        n3810) );
  AND4_X1 U6909 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n3811) );
  AND4_X1 U6910 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n3812)
         );
  AND4_X1 U6911 ( .A1(n7927), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n3813)
         );
  AND4_X1 U6912 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n3814) );
  AND4_X1 U6913 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n3815) );
  AND4_X1 U6914 ( .A1(n15655), .A2(n15654), .A3(n15653), .A4(n15652), .ZN(
        n3816) );
  AND4_X1 U6915 ( .A1(n27993), .A2(n27992), .A3(n27991), .A4(n27990), .ZN(
        n3817) );
  AND4_X1 U6916 ( .A1(n24501), .A2(n24500), .A3(n24499), .A4(n24498), .ZN(
        n3818) );
  AND4_X1 U6917 ( .A1(n17627), .A2(n17626), .A3(n17625), .A4(n17624), .ZN(
        n3819) );
  AND4_X1 U6918 ( .A1(n23055), .A2(n23054), .A3(n23053), .A4(n23052), .ZN(
        n3820) );
  AND4_X1 U6919 ( .A1(n24818), .A2(n24817), .A3(n24816), .A4(n24815), .ZN(
        n3821) );
  AND4_X1 U6920 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n3822) );
  AND4_X1 U6921 ( .A1(n26420), .A2(n26419), .A3(n26418), .A4(n26417), .ZN(
        n3823) );
  AND4_X1 U6922 ( .A1(n28184), .A2(n28183), .A3(n28182), .A4(n28181), .ZN(
        n3824) );
  AND4_X1 U6923 ( .A1(n19679), .A2(n19678), .A3(n19677), .A4(n19676), .ZN(
        n3825) );
  AND4_X1 U6924 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n3826)
         );
  AND4_X1 U6925 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n3827)
         );
  AND4_X1 U6926 ( .A1(n8334), .A2(n8333), .A3(n8332), .A4(n8331), .ZN(n3828)
         );
  AND4_X1 U6927 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        n3829) );
  AND4_X1 U6928 ( .A1(n18174), .A2(n18173), .A3(n18172), .A4(n18171), .ZN(
        n3830) );
  AND4_X1 U6929 ( .A1(n23121), .A2(n23120), .A3(n23119), .A4(n23118), .ZN(
        n3831) );
  AND4_X1 U6930 ( .A1(n13722), .A2(n13721), .A3(n13720), .A4(n13719), .ZN(
        n3832) );
  AND4_X1 U6931 ( .A1(n7224), .A2(n7223), .A3(n7222), .A4(n7221), .ZN(n3833)
         );
  AND2_X1 U6932 ( .A1(n6280), .A2(n30329), .ZN(n3834) );
  AND2_X1 U6933 ( .A1(n33176), .A2(n33174), .ZN(n3835) );
  BUF_X1 U6934 ( .A(n4026), .Z(n8409) );
  AND4_X1 U6935 ( .A1(n16971), .A2(n16970), .A3(n16969), .A4(n16968), .ZN(
        n3836) );
  AND4_X1 U6936 ( .A1(n27363), .A2(n27362), .A3(n27361), .A4(n27360), .ZN(
        n3837) );
  AND4_X1 U6937 ( .A1(n18483), .A2(n18482), .A3(n18481), .A4(n18480), .ZN(
        n3838) );
  AND4_X1 U6938 ( .A1(n27810), .A2(n27809), .A3(n27808), .A4(n27807), .ZN(
        n3839) );
  AND4_X1 U6939 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n3840)
         );
  AND4_X1 U6940 ( .A1(n18059), .A2(n18058), .A3(n18057), .A4(n18056), .ZN(
        n3841) );
  AND4_X1 U6941 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), .ZN(n3842)
         );
  AND4_X1 U6942 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n3843) );
  AND4_X1 U6943 ( .A1(n27337), .A2(n27336), .A3(n27335), .A4(n27334), .ZN(
        n3844) );
  AND4_X1 U6944 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n3845)
         );
  AND4_X1 U6945 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n3846)
         );
  AND4_X1 U6946 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n3847)
         );
  AND4_X1 U6947 ( .A1(n7325), .A2(n7324), .A3(n7323), .A4(n7322), .ZN(n3848)
         );
  AND4_X1 U6948 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n3849) );
  AND4_X1 U6949 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n3850) );
  AND4_X1 U6950 ( .A1(n16646), .A2(n16645), .A3(n16644), .A4(n16643), .ZN(
        n3851) );
  AND4_X1 U6951 ( .A1(n16873), .A2(n16872), .A3(n16871), .A4(n16870), .ZN(
        n3852) );
  AND4_X1 U6952 ( .A1(n19785), .A2(n19784), .A3(n19783), .A4(n19782), .ZN(
        n3853) );
  AND4_X1 U6953 ( .A1(n22028), .A2(n22027), .A3(n22026), .A4(n22025), .ZN(
        n3854) );
  AND4_X1 U6954 ( .A1(n24951), .A2(n24950), .A3(n24949), .A4(n24948), .ZN(
        n3855) );
  AND4_X1 U6955 ( .A1(n26755), .A2(n26754), .A3(n26753), .A4(n26752), .ZN(
        n3856) );
  AND4_X1 U6956 ( .A1(n28770), .A2(n28769), .A3(n28768), .A4(n28767), .ZN(
        n3857) );
  AND4_X1 U6957 ( .A1(n29645), .A2(n29644), .A3(n29643), .A4(n29642), .ZN(
        n3858) );
  AND4_X1 U6958 ( .A1(n18455), .A2(n18454), .A3(n18453), .A4(n18452), .ZN(
        n3859) );
  AND4_X1 U6959 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n3860)
         );
  AND2_X1 U6960 ( .A1(n30730), .A2(\xmem_data[53][2] ), .ZN(n3861) );
  AND4_X1 U6961 ( .A1(n21990), .A2(n21989), .A3(n21988), .A4(n21987), .ZN(
        n3862) );
  AND4_X1 U6962 ( .A1(n26098), .A2(n26097), .A3(n26096), .A4(n26095), .ZN(
        n3863) );
  AND4_X1 U6963 ( .A1(n9166), .A2(n9165), .A3(n9164), .A4(n9163), .ZN(n3864)
         );
  AND4_X1 U6964 ( .A1(n16068), .A2(n16067), .A3(n16066), .A4(n16065), .ZN(
        n3865) );
  AND4_X1 U6965 ( .A1(n16111), .A2(n16110), .A3(n16109), .A4(n16108), .ZN(
        n3866) );
  AND4_X1 U6966 ( .A1(n26877), .A2(n26876), .A3(n26875), .A4(n26874), .ZN(
        n3867) );
  AND4_X1 U6967 ( .A1(n29122), .A2(n29121), .A3(n29120), .A4(n29119), .ZN(
        n3868) );
  AND4_X1 U6968 ( .A1(n26498), .A2(n26497), .A3(n26496), .A4(n26495), .ZN(
        n3869) );
  AND2_X1 U6969 ( .A1(n33679), .A2(n33681), .ZN(n3870) );
  AND2_X1 U6970 ( .A1(n34495), .A2(n34497), .ZN(n3871) );
  AND2_X1 U6971 ( .A1(n34429), .A2(n34533), .ZN(n3872) );
  AND2_X1 U6972 ( .A1(n30877), .A2(\xmem_data[17][7] ), .ZN(n3873) );
  AND2_X1 U6973 ( .A1(n27547), .A2(\xmem_data[21][7] ), .ZN(n3874) );
  AND4_X1 U6974 ( .A1(n27752), .A2(n27751), .A3(n27750), .A4(n27749), .ZN(
        n3875) );
  AND2_X1 U6975 ( .A1(n34836), .A2(n34835), .ZN(n3876) );
  AND2_X1 U6976 ( .A1(n29103), .A2(\xmem_data[25][4] ), .ZN(n3877) );
  AND2_X1 U6977 ( .A1(n33796), .A2(n33797), .ZN(n3878) );
  OR2_X1 U6978 ( .A1(n35086), .A2(n35085), .ZN(n3879) );
  AND2_X1 U6979 ( .A1(n24131), .A2(\xmem_data[18][5] ), .ZN(n3880) );
  AND2_X1 U6980 ( .A1(n30877), .A2(n22179), .ZN(n3881) );
  AND2_X1 U6981 ( .A1(n27547), .A2(n5564), .ZN(n3882) );
  AND2_X1 U6982 ( .A1(n29306), .A2(n12688), .ZN(n3883) );
  AND2_X1 U6983 ( .A1(n25450), .A2(n22023), .ZN(n3884) );
  AND2_X1 U6984 ( .A1(n28510), .A2(\xmem_data[31][2] ), .ZN(n3885) );
  AND2_X1 U6985 ( .A1(n28007), .A2(\xmem_data[31][1] ), .ZN(n3886) );
  AND3_X1 U6986 ( .A1(n13702), .A2(n13701), .A3(n13700), .ZN(n3887) );
  AND2_X1 U6987 ( .A1(n27547), .A2(n17966), .ZN(n3888) );
  AND2_X1 U6988 ( .A1(n28343), .A2(n18090), .ZN(n3889) );
  AND2_X1 U6989 ( .A1(n30877), .A2(n15012), .ZN(n3890) );
  AND2_X1 U6990 ( .A1(n28343), .A2(n19754), .ZN(n3891) );
  AND2_X1 U6991 ( .A1(n24657), .A2(n20461), .ZN(n3892) );
  AND2_X1 U6992 ( .A1(n25492), .A2(n22299), .ZN(n3893) );
  AND2_X1 U6993 ( .A1(n29306), .A2(n28889), .ZN(n3894) );
  AND2_X1 U6994 ( .A1(n24657), .A2(n9681), .ZN(n3895) );
  AND2_X1 U6995 ( .A1(n29103), .A2(n20189), .ZN(n3896) );
  AND2_X1 U6996 ( .A1(n23771), .A2(n11234), .ZN(n3897) );
  NOR3_X1 U6997 ( .A1(n22273), .A2(n22272), .A3(n22271), .ZN(n3898) );
  AND2_X1 U6998 ( .A1(n3231), .A2(n14309), .ZN(n3899) );
  AND3_X1 U6999 ( .A1(n18287), .A2(n18286), .A3(n18285), .ZN(n3900) );
  NAND2_X1 U7000 ( .A1(n39054), .A2(n39035), .ZN(n4050) );
  INV_X1 U7001 ( .A(n4050), .ZN(n4049) );
  AND2_X1 U7002 ( .A1(n25492), .A2(n19184), .ZN(n3901) );
  AND2_X1 U7003 ( .A1(n31252), .A2(n29342), .ZN(n3902) );
  AND3_X1 U7004 ( .A1(n21289), .A2(n21288), .A3(n21287), .ZN(n3903) );
  AND4_X1 U7005 ( .A1(n21305), .A2(n21304), .A3(n21303), .A4(n21302), .ZN(
        n3904) );
  AND4_X1 U7006 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n3905) );
  OR2_X1 U7007 ( .A1(n30471), .A2(n10364), .ZN(n3906) );
  AND3_X1 U7008 ( .A1(n13439), .A2(n13438), .A3(n13437), .ZN(n3907) );
  AND2_X1 U7009 ( .A1(n30882), .A2(\xmem_data[16][0] ), .ZN(n3908) );
  AND4_X1 U7010 ( .A1(n21386), .A2(n21385), .A3(n21384), .A4(n21383), .ZN(
        n3909) );
  AND3_X1 U7011 ( .A1(n25363), .A2(n25362), .A3(n25361), .ZN(n3910) );
  AND2_X1 U7012 ( .A1(n28510), .A2(\xmem_data[31][6] ), .ZN(n3911) );
  AND4_X1 U7013 ( .A1(n17686), .A2(n17685), .A3(n17684), .A4(n17683), .ZN(
        n3912) );
  AND2_X1 U7014 ( .A1(n30106), .A2(\xmem_data[45][0] ), .ZN(n3913) );
  AND2_X1 U7015 ( .A1(n3231), .A2(\xmem_data[14][2] ), .ZN(n3914) );
  AND4_X1 U7016 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n3915)
         );
  AND2_X1 U7017 ( .A1(n28108), .A2(n28107), .ZN(n3916) );
  AND3_X1 U7018 ( .A1(n14499), .A2(n14498), .A3(n14497), .ZN(n3917) );
  OR3_X1 U7019 ( .A1(n14099), .A2(n14098), .A3(n14097), .ZN(n3918) );
  OR3_X1 U7020 ( .A1(n15651), .A2(n15650), .A3(n15649), .ZN(n3919) );
  INV_X1 U7021 ( .A(n3402), .ZN(n8416) );
  AND2_X1 U7022 ( .A1(n29045), .A2(\xmem_data[82][1] ), .ZN(n3920) );
  AND2_X1 U7023 ( .A1(n15813), .A2(n15812), .ZN(n3921) );
  AND2_X1 U7024 ( .A1(n15855), .A2(n15854), .ZN(n3922) );
  NOR2_X1 U7025 ( .A1(n33928), .A2(n30425), .ZN(n30426) );
  AND2_X1 U7026 ( .A1(n16491), .A2(n16490), .ZN(n3923) );
  AND2_X1 U7027 ( .A1(n24657), .A2(\xmem_data[57][1] ), .ZN(n3924) );
  AND2_X1 U7028 ( .A1(n10473), .A2(n10472), .ZN(n3925) );
  AND2_X1 U7029 ( .A1(n26698), .A2(n26697), .ZN(n3926) );
  AND2_X1 U7030 ( .A1(n13636), .A2(n29143), .ZN(n3927) );
  AND2_X1 U7031 ( .A1(n3231), .A2(\xmem_data[25][2] ), .ZN(n3928) );
  AND2_X1 U7032 ( .A1(n7581), .A2(n7580), .ZN(n3929) );
  AND2_X1 U7033 ( .A1(n15618), .A2(n15617), .ZN(n3930) );
  AND2_X1 U7034 ( .A1(n29045), .A2(\xmem_data[45][5] ), .ZN(n3932) );
  AND2_X1 U7035 ( .A1(n15870), .A2(n15869), .ZN(n3933) );
  AND2_X1 U7036 ( .A1(n7844), .A2(n7843), .ZN(n3934) );
  AND3_X1 U7037 ( .A1(n15641), .A2(n15640), .A3(n15639), .ZN(n3935) );
  AND2_X1 U7038 ( .A1(n15670), .A2(n15669), .ZN(n3936) );
  AND2_X1 U7039 ( .A1(n35004), .A2(n35003), .ZN(n3937) );
  AND2_X1 U7040 ( .A1(n4673), .A2(n4672), .ZN(n3938) );
  NOR2_X1 U7041 ( .A1(n11112), .A2(n11111), .ZN(n3939) );
  NOR2_X1 U7042 ( .A1(n25622), .A2(n25621), .ZN(n3940) );
  AND2_X1 U7043 ( .A1(n11382), .A2(n39041), .ZN(n3941) );
  AND2_X1 U7044 ( .A1(n28149), .A2(n28148), .ZN(n3942) );
  AND2_X1 U7045 ( .A1(n34043), .A2(n34045), .ZN(n3943) );
  OR2_X1 U7046 ( .A1(n6171), .A2(n6170), .ZN(n3944) );
  INV_X1 U7047 ( .A(n31823), .ZN(n35134) );
  AOI21_X1 U7048 ( .B1(n33105), .B2(n33103), .A(n33106), .ZN(n31823) );
  AND2_X1 U7049 ( .A1(n35037), .A2(n35036), .ZN(n3946) );
  AND2_X1 U7050 ( .A1(n25514), .A2(\xmem_data[7][5] ), .ZN(n3947) );
  AND2_X1 U7051 ( .A1(n35007), .A2(n35006), .ZN(n3948) );
  AND3_X1 U7052 ( .A1(n6448), .A2(n6447), .A3(n6446), .ZN(n3949) );
  NAND2_X1 U7053 ( .A1(n30295), .A2(\xmem_data[2][5] ), .ZN(n3950) );
  OR2_X1 U7054 ( .A1(n28992), .A2(n28991), .ZN(n3951) );
  AND3_X1 U7055 ( .A1(n19321), .A2(n19320), .A3(n19319), .ZN(n3952) );
  NAND2_X1 U7056 ( .A1(n22879), .A2(n23822), .ZN(n3953) );
  AND2_X1 U7057 ( .A1(n24877), .A2(n24876), .ZN(n3954) );
  NAND2_X1 U7058 ( .A1(n16465), .A2(n25396), .ZN(n3955) );
  AND2_X1 U7059 ( .A1(n32779), .A2(n32780), .ZN(n3956) );
  INV_X1 U7060 ( .A(n30443), .ZN(n31689) );
  AND2_X1 U7061 ( .A1(n28307), .A2(\xmem_data[7][0] ), .ZN(n3957) );
  AND2_X1 U7062 ( .A1(n13474), .A2(\xmem_data[9][0] ), .ZN(n3958) );
  OR2_X1 U7063 ( .A1(n25381), .A2(n25380), .ZN(n3959) );
  AND2_X1 U7064 ( .A1(n29103), .A2(\xmem_data[15][0] ), .ZN(n3960) );
  OR2_X1 U7065 ( .A1(n21332), .A2(n21331), .ZN(n3961) );
  AND2_X1 U7066 ( .A1(n31252), .A2(n17319), .ZN(n3962) );
  OR2_X1 U7067 ( .A1(n16383), .A2(n16382), .ZN(n3963) );
  OR2_X1 U7068 ( .A1(n20203), .A2(n20202), .ZN(n3964) );
  OR2_X1 U7069 ( .A1(n24485), .A2(n24484), .ZN(n3965) );
  AND2_X1 U7070 ( .A1(n31252), .A2(\xmem_data[15][4] ), .ZN(n3966) );
  OR2_X1 U7071 ( .A1(n5089), .A2(n5088), .ZN(n3967) );
  OR2_X1 U7072 ( .A1(n13645), .A2(n13644), .ZN(n3968) );
  AND2_X1 U7073 ( .A1(n31252), .A2(\xmem_data[25][7] ), .ZN(n3969) );
  NAND4_X1 U7074 ( .A1(n25851), .A2(n25850), .A3(n25849), .A4(n25848), .ZN(
        n3970) );
  OR3_X1 U7075 ( .A1(n14510), .A2(n14509), .A3(n14508), .ZN(n3971) );
  AND2_X1 U7076 ( .A1(n28045), .A2(\xmem_data[23][0] ), .ZN(n3972) );
  OR2_X1 U7077 ( .A1(n27648), .A2(n27647), .ZN(n3973) );
  AND2_X1 U7078 ( .A1(n28343), .A2(\xmem_data[14][6] ), .ZN(n3974) );
  NAND2_X1 U7079 ( .A1(n29086), .A2(\xmem_data[36][0] ), .ZN(n3975) );
  AND2_X1 U7080 ( .A1(n28045), .A2(\xmem_data[13][4] ), .ZN(n3976) );
  AND2_X1 U7081 ( .A1(n28007), .A2(\xmem_data[13][6] ), .ZN(n3977) );
  NAND4_X1 U7082 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n3978)
         );
  OR2_X1 U7083 ( .A1(n19145), .A2(n19144), .ZN(n3979) );
  NAND2_X1 U7084 ( .A1(n29439), .A2(\xmem_data[127][2] ), .ZN(n3980) );
  OR2_X1 U7085 ( .A1(n22263), .A2(n22262), .ZN(n3981) );
  OR2_X1 U7086 ( .A1(n13288), .A2(n3725), .ZN(n3982) );
  OR2_X1 U7087 ( .A1(n5576), .A2(n5575), .ZN(n3983) );
  OR2_X1 U7088 ( .A1(n5602), .A2(n5601), .ZN(n3984) );
  OR2_X1 U7089 ( .A1(n21292), .A2(n21291), .ZN(n3985) );
  OR2_X1 U7090 ( .A1(n10200), .A2(n10199), .ZN(n3986) );
  NAND3_X1 U7091 ( .A1(n19149), .A2(n19148), .A3(n19147), .ZN(n3988) );
  NAND4_X1 U7092 ( .A1(n19923), .A2(n19922), .A3(n19921), .A4(n19920), .ZN(
        n3989) );
  OR2_X1 U7093 ( .A1(n10451), .A2(n10450), .ZN(n3990) );
  OR2_X1 U7094 ( .A1(n17655), .A2(n17654), .ZN(n3991) );
  INV_X1 U7095 ( .A(n31491), .ZN(n33575) );
  AND2_X1 U7096 ( .A1(n36244), .A2(n31490), .ZN(n31491) );
  OR2_X1 U7097 ( .A1(n8736), .A2(n8735), .ZN(n3992) );
  OR2_X1 U7098 ( .A1(n18029), .A2(n18028), .ZN(n3993) );
  OR2_X1 U7099 ( .A1(n21543), .A2(n21542), .ZN(n3994) );
  OR2_X1 U7100 ( .A1(n18302), .A2(n3741), .ZN(n3995) );
  OR2_X1 U7101 ( .A1(n16373), .A2(n16372), .ZN(n3996) );
  NAND2_X1 U7102 ( .A1(n27551), .A2(\xmem_data[14][0] ), .ZN(n3997) );
  NAND3_X1 U7103 ( .A1(n26895), .A2(n26894), .A3(n26893), .ZN(n3998) );
  AND2_X1 U7104 ( .A1(n37239), .A2(n37238), .ZN(n4000) );
  NAND2_X1 U7105 ( .A1(n25358), .A2(\xmem_data[30][3] ), .ZN(n4001) );
  AND2_X1 U7106 ( .A1(n24553), .A2(\xmem_data[29][0] ), .ZN(n4002) );
  OR2_X1 U7107 ( .A1(n17919), .A2(n17918), .ZN(n4003) );
  OR2_X1 U7108 ( .A1(n24276), .A2(n24275), .ZN(n4004) );
  NAND2_X1 U7109 ( .A1(n27547), .A2(\xmem_data[31][3] ), .ZN(n4005) );
  NAND2_X1 U7110 ( .A1(n29674), .A2(\xmem_data[40][1] ), .ZN(n4006) );
  AND2_X1 U7111 ( .A1(n37205), .A2(n37234), .ZN(n4007) );
  AND2_X1 U7112 ( .A1(n18200), .A2(n18199), .ZN(n4008) );
  AND2_X1 U7113 ( .A1(n29406), .A2(n29405), .ZN(n4009) );
  AND2_X1 U7114 ( .A1(n20306), .A2(n20305), .ZN(n4010) );
  AND2_X1 U7115 ( .A1(n37256), .A2(n37255), .ZN(n4011) );
  OR2_X1 U7116 ( .A1(n33190), .A2(n25149), .ZN(n4012) );
  AND2_X1 U7117 ( .A1(n36012), .A2(n37229), .ZN(n4013) );
  BUF_X1 U7118 ( .A(n4063), .Z(n10288) );
  AND2_X1 U7119 ( .A1(n37248), .A2(n37247), .ZN(n4014) );
  AND2_X1 U7120 ( .A1(n25614), .A2(n25613), .ZN(n4015) );
  AND2_X1 U7121 ( .A1(n25383), .A2(\xmem_data[31][5] ), .ZN(n4016) );
  NAND4_X1 U7122 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4017)
         );
  NAND2_X1 U7123 ( .A1(\fmem_data[25][1] ), .A2(n3483), .ZN(n34440) );
  AND2_X1 U7124 ( .A1(n25492), .A2(\xmem_data[10][3] ), .ZN(n4019) );
  NAND2_X1 U7125 ( .A1(n37181), .A2(n37180), .ZN(n37241) );
  AND2_X1 U7126 ( .A1(n39052), .A2(n39053), .ZN(n4021) );
  BUF_X2 U7127 ( .A(N284), .Z(n4391) );
  INV_X4 U7128 ( .A(n3676), .ZN(n29064) );
  INV_X1 U7129 ( .A(n39052), .ZN(n4038) );
  NAND3_X1 U7130 ( .A1(n4391), .A2(n4038), .A3(n3346), .ZN(n4059) );
  NOR2_X1 U7131 ( .A1(n4059), .A2(n4050), .ZN(n4248) );
  AND2_X1 U7132 ( .A1(n3219), .A2(\xmem_data[25][7] ), .ZN(n4022) );
  AOI21_X1 U7133 ( .B1(n25354), .B2(\xmem_data[24][7] ), .A(n4022), .ZN(n4023)
         );
  INV_X1 U7134 ( .A(n4023), .ZN(n4036) );
  BUF_X1 U7135 ( .A(N284), .Z(n4026) );
  BUF_X1 U7136 ( .A(n14926), .Z(n25617) );
  AND2_X1 U7137 ( .A1(n4391), .A2(N345), .ZN(n4025) );
  NOR2_X1 U7138 ( .A1(n13132), .A2(n4050), .ZN(n4204) );
  BUF_X2 U7139 ( .A(n4204), .Z(n14927) );
  BUF_X1 U7140 ( .A(n14927), .Z(n25616) );
  AOI22_X1 U7141 ( .A1(n25617), .A2(\xmem_data[28][7] ), .B1(n25616), .B2(
        \xmem_data[29][7] ), .ZN(n4029) );
  NAND2_X2 U7142 ( .A1(n39054), .A2(N466), .ZN(n10972) );
  INV_X1 U7143 ( .A(n10972), .ZN(n4027) );
  NOR2_X2 U7144 ( .A1(n4026), .A2(\add_x_2/A[0] ), .ZN(n6171) );
  AND2_X2 U7145 ( .A1(n6171), .A2(n6586), .ZN(n6992) );
  AND2_X4 U7146 ( .A1(n6992), .A2(n4027), .ZN(n14991) );
  NAND2_X1 U7147 ( .A1(n3281), .A2(\xmem_data[30][7] ), .ZN(n4028) );
  NAND2_X1 U7148 ( .A1(n4029), .A2(n4028), .ZN(n4034) );
  AND2_X1 U7149 ( .A1(n39052), .A2(N345), .ZN(n4060) );
  NAND2_X1 U7150 ( .A1(n39010), .A2(n4060), .ZN(n4048) );
  INV_X1 U7151 ( .A(n4048), .ZN(n4030) );
  AND2_X4 U7152 ( .A1(n4030), .A2(n4049), .ZN(n14988) );
  BUF_X1 U7153 ( .A(n14988), .Z(n25612) );
  NOR2_X1 U7154 ( .A1(n4061), .A2(n4050), .ZN(n4253) );
  AOI22_X1 U7155 ( .A1(n25612), .A2(\xmem_data[26][7] ), .B1(n20500), .B2(
        \xmem_data[27][7] ), .ZN(n4032) );
  INV_X1 U7156 ( .A(n4032), .ZN(n4033) );
  OR2_X1 U7157 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  NOR2_X1 U7158 ( .A1(n4036), .A2(n4035), .ZN(n4047) );
  AOI22_X1 U7159 ( .A1(n25604), .A2(\xmem_data[0][7] ), .B1(n27943), .B2(
        \xmem_data[1][7] ), .ZN(n4045) );
  NOR2_X1 U7160 ( .A1(n4061), .A2(n10972), .ZN(n4177) );
  BUF_X1 U7161 ( .A(n13435), .Z(n25605) );
  AOI22_X1 U7162 ( .A1(n28743), .A2(\xmem_data[2][7] ), .B1(n25605), .B2(
        \xmem_data[3][7] ), .ZN(n4044) );
  NOR2_X1 U7163 ( .A1(n13132), .A2(n10972), .ZN(n4404) );
  BUF_X2 U7164 ( .A(n4404), .Z(n14898) );
  BUF_X1 U7165 ( .A(n14898), .Z(n25606) );
  AOI22_X1 U7166 ( .A1(n31268), .A2(\xmem_data[4][7] ), .B1(n25606), .B2(
        \xmem_data[5][7] ), .ZN(n4043) );
  NAND2_X1 U7167 ( .A1(n39035), .A2(n38997), .ZN(n4063) );
  INV_X1 U7168 ( .A(n4063), .ZN(n4040) );
  NAND2_X1 U7169 ( .A1(n39053), .A2(n39010), .ZN(n9417) );
  BUF_X1 U7170 ( .A(n3464), .Z(n25607) );
  AND2_X1 U7171 ( .A1(n39053), .A2(n39010), .ZN(n4041) );
  AOI22_X1 U7172 ( .A1(n20776), .A2(\xmem_data[6][7] ), .B1(n3208), .B2(
        \xmem_data[7][7] ), .ZN(n4042) );
  AND4_X1 U7173 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  NAND2_X1 U7174 ( .A1(n4047), .A2(n4046), .ZN(n4073) );
  NAND2_X1 U7175 ( .A1(n38997), .A2(N466), .ZN(n4065) );
  INV_X1 U7176 ( .A(n4065), .ZN(n4064) );
  BUF_X1 U7177 ( .A(n31263), .Z(n25630) );
  OR2_X1 U7178 ( .A1(n13132), .A2(n4065), .ZN(n4368) );
  INV_X1 U7179 ( .A(n4368), .ZN(n28974) );
  BUF_X1 U7180 ( .A(n28974), .Z(n25629) );
  AOI22_X1 U7181 ( .A1(n25630), .A2(\xmem_data[20][7] ), .B1(n25629), .B2(
        \xmem_data[21][7] ), .ZN(n4057) );
  NOR2_X1 U7182 ( .A1(n4048), .A2(n4065), .ZN(n4527) );
  BUF_X1 U7183 ( .A(n13127), .Z(n25628) );
  AND2_X4 U7184 ( .A1(n6992), .A2(n4049), .ZN(n28973) );
  BUF_X1 U7185 ( .A(n28973), .Z(n25624) );
  NOR2_X1 U7186 ( .A1(n4080), .A2(n4050), .ZN(n4247) );
  BUF_X1 U7187 ( .A(n4247), .Z(n14983) );
  AOI22_X1 U7188 ( .A1(n25624), .A2(\xmem_data[22][7] ), .B1(n3247), .B2(
        \xmem_data[23][7] ), .ZN(n4052) );
  OR2_X1 U7189 ( .A1(n4061), .A2(n4065), .ZN(n4456) );
  INV_X1 U7190 ( .A(n4456), .ZN(n10456) );
  NAND2_X1 U7191 ( .A1(n10456), .A2(\xmem_data[19][7] ), .ZN(n4051) );
  NAND2_X1 U7192 ( .A1(n4052), .A2(n4051), .ZN(n4055) );
  NOR2_X1 U7193 ( .A1(n4059), .A2(n4065), .ZN(n4526) );
  AOI22_X1 U7194 ( .A1(n14976), .A2(\xmem_data[16][7] ), .B1(n23725), .B2(
        \xmem_data[17][7] ), .ZN(n4053) );
  INV_X1 U7195 ( .A(n4053), .ZN(n4054) );
  AOI211_X1 U7196 ( .C1(n25628), .C2(\xmem_data[18][7] ), .A(n4055), .B(n4054), 
        .ZN(n4056) );
  NAND2_X1 U7197 ( .A1(n4057), .A2(n4056), .ZN(n4071) );
  OR2_X1 U7198 ( .A1(n4058), .A2(n4063), .ZN(n4178) );
  BUF_X1 U7199 ( .A(n14937), .Z(n25635) );
  OR2_X1 U7200 ( .A1(n4059), .A2(n4063), .ZN(n4237) );
  INV_X1 U7201 ( .A(n4237), .ZN(n13415) );
  AOI22_X1 U7202 ( .A1(n25635), .A2(\xmem_data[8][7] ), .B1(n25715), .B2(
        \xmem_data[9][7] ), .ZN(n4069) );
  AND3_X4 U7203 ( .A1(n39010), .A2(n4060), .A3(n4040), .ZN(n14971) );
  AOI22_X1 U7204 ( .A1(n27855), .A2(\xmem_data[10][7] ), .B1(n31360), .B2(
        \xmem_data[11][7] ), .ZN(n4068) );
  BUF_X1 U7205 ( .A(n14972), .Z(n25632) );
  OR2_X1 U7206 ( .A1(n13132), .A2(n4063), .ZN(n4516) );
  AOI22_X1 U7207 ( .A1(n25632), .A2(\xmem_data[12][7] ), .B1(n27856), .B2(
        \xmem_data[13][7] ), .ZN(n4067) );
  AND2_X4 U7208 ( .A1(n6992), .A2(n4064), .ZN(n14974) );
  BUF_X1 U7209 ( .A(n14974), .Z(n25636) );
  OR2_X1 U7210 ( .A1(n4080), .A2(n4065), .ZN(n4489) );
  AOI22_X1 U7211 ( .A1(n25636), .A2(\xmem_data[14][7] ), .B1(n25583), .B2(
        \xmem_data[15][7] ), .ZN(n4066) );
  NAND4_X1 U7212 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OR2_X1 U7213 ( .A1(n4071), .A2(n4070), .ZN(n4072) );
  NOR2_X1 U7214 ( .A1(n4073), .A2(n4072), .ZN(n4076) );
  INV_X1 U7215 ( .A(n10972), .ZN(n7216) );
  NAND2_X1 U7216 ( .A1(n7216), .A2(n9417), .ZN(n4074) );
  NOR2_X1 U7217 ( .A1(n39041), .A2(n4074), .ZN(n4075) );
  AOI21_X1 U7218 ( .B1(n39041), .B2(n4074), .A(n4075), .ZN(n4130) );
  BUF_X2 U7219 ( .A(N466), .Z(n6990) );
  NAND2_X1 U7220 ( .A1(n9417), .A2(n6990), .ZN(n4497) );
  NOR2_X1 U7221 ( .A1(n39041), .A2(load_xaddr_val[6]), .ZN(n20311) );
  BUF_X4 U7222 ( .A(n39054), .Z(n10589) );
  NAND2_X1 U7223 ( .A1(n20311), .A2(n10589), .ZN(n13431) );
  OAI22_X1 U7224 ( .A1(n4075), .A2(n39040), .B1(n4497), .B2(n13431), .ZN(n4108) );
  NOR2_X1 U7225 ( .A1(n4130), .A2(n4108), .ZN(n19018) );
  INV_X1 U7226 ( .A(n19018), .ZN(n25647) );
  NOR2_X1 U7227 ( .A1(n4076), .A2(n25647), .ZN(n4106) );
  BUF_X1 U7228 ( .A(n29064), .Z(n25730) );
  AND2_X1 U7229 ( .A1(n3220), .A2(\xmem_data[57][7] ), .ZN(n4077) );
  AOI21_X1 U7230 ( .B1(n25730), .B2(\xmem_data[56][7] ), .A(n4077), .ZN(n4086)
         );
  AOI22_X1 U7231 ( .A1(n27938), .A2(\xmem_data[60][7] ), .B1(n20993), .B2(
        \xmem_data[61][7] ), .ZN(n4079) );
  INV_X1 U7232 ( .A(n4079), .ZN(n4084) );
  BUF_X1 U7233 ( .A(n14988), .Z(n25731) );
  AOI22_X1 U7234 ( .A1(n25731), .A2(\xmem_data[58][7] ), .B1(n27869), .B2(
        \xmem_data[59][7] ), .ZN(n4082) );
  BUF_X1 U7235 ( .A(n14991), .Z(n25732) );
  OR2_X2 U7236 ( .A1(n10972), .A2(n4080), .ZN(n4254) );
  AOI22_X1 U7237 ( .A1(n25732), .A2(\xmem_data[62][7] ), .B1(n15011), .B2(
        \xmem_data[63][7] ), .ZN(n4081) );
  NAND2_X1 U7238 ( .A1(n4082), .A2(n4081), .ZN(n4083) );
  NOR2_X1 U7239 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  NAND2_X1 U7240 ( .A1(n4086), .A2(n4085), .ZN(n4103) );
  BUF_X1 U7241 ( .A(n4526), .Z(n14919) );
  BUF_X1 U7242 ( .A(n14919), .Z(n25723) );
  AOI22_X1 U7243 ( .A1(n3209), .A2(\xmem_data[48][7] ), .B1(n25723), .B2(
        \xmem_data[49][7] ), .ZN(n4091) );
  AND2_X1 U7244 ( .A1(n10456), .A2(\xmem_data[51][7] ), .ZN(n4087) );
  AOI21_X1 U7245 ( .B1(n17051), .B2(\xmem_data[50][7] ), .A(n4087), .ZN(n4090)
         );
  BUF_X1 U7246 ( .A(n31263), .Z(n25724) );
  AOI22_X1 U7247 ( .A1(n25724), .A2(\xmem_data[52][7] ), .B1(n20709), .B2(
        \xmem_data[53][7] ), .ZN(n4089) );
  BUF_X1 U7248 ( .A(n28973), .Z(n25725) );
  AOI22_X1 U7249 ( .A1(n25725), .A2(\xmem_data[54][7] ), .B1(n24439), .B2(
        \xmem_data[55][7] ), .ZN(n4088) );
  NAND4_X1 U7250 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4102)
         );
  AOI22_X1 U7251 ( .A1(n25707), .A2(\xmem_data[32][7] ), .B1(n24590), .B2(
        \xmem_data[33][7] ), .ZN(n4095) );
  BUF_X1 U7252 ( .A(n14997), .Z(n25708) );
  BUF_X2 U7253 ( .A(n4177), .Z(n13168) );
  AOI22_X1 U7254 ( .A1(n25708), .A2(\xmem_data[34][7] ), .B1(n13168), .B2(
        \xmem_data[35][7] ), .ZN(n4094) );
  BUF_X1 U7255 ( .A(n10977), .Z(n25710) );
  BUF_X2 U7256 ( .A(n4404), .Z(n14935) );
  BUF_X1 U7257 ( .A(n14935), .Z(n25709) );
  AOI22_X1 U7258 ( .A1(n28980), .A2(\xmem_data[36][7] ), .B1(n25709), .B2(
        \xmem_data[37][7] ), .ZN(n4093) );
  AOI22_X1 U7259 ( .A1(n25519), .A2(\xmem_data[38][7] ), .B1(n30615), .B2(
        \xmem_data[39][7] ), .ZN(n4092) );
  NAND4_X1 U7260 ( .A1(n4095), .A2(n4094), .A3(n4093), .A4(n4092), .ZN(n4101)
         );
  BUF_X1 U7261 ( .A(n13415), .Z(n25715) );
  AOI22_X1 U7262 ( .A1(n25573), .A2(\xmem_data[40][7] ), .B1(n25715), .B2(
        \xmem_data[41][7] ), .ZN(n4099) );
  AOI22_X1 U7263 ( .A1(n23802), .A2(\xmem_data[42][7] ), .B1(n31254), .B2(
        \xmem_data[43][7] ), .ZN(n4098) );
  BUF_X1 U7264 ( .A(n3324), .Z(n25717) );
  BUF_X1 U7265 ( .A(n14882), .Z(n25716) );
  AOI22_X1 U7266 ( .A1(n24548), .A2(\xmem_data[44][7] ), .B1(n25581), .B2(
        \xmem_data[45][7] ), .ZN(n4097) );
  BUF_X1 U7267 ( .A(n14974), .Z(n25718) );
  INV_X1 U7268 ( .A(n4489), .ZN(n14914) );
  AOI22_X1 U7269 ( .A1(n25718), .A2(\xmem_data[46][7] ), .B1(n31314), .B2(
        \xmem_data[47][7] ), .ZN(n4096) );
  NAND4_X1 U7270 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4100)
         );
  OR4_X1 U7271 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104) );
  INV_X1 U7272 ( .A(n4108), .ZN(n4129) );
  AND2_X1 U7273 ( .A1(n4104), .A2(n25741), .ZN(n4105) );
  NOR2_X1 U7274 ( .A1(n4106), .A2(n4105), .ZN(n4155) );
  INV_X1 U7275 ( .A(n4254), .ZN(n15011) );
  NOR2_X1 U7276 ( .A1(n25647), .A2(n39024), .ZN(n4107) );
  NAND2_X1 U7277 ( .A1(n25514), .A2(n4107), .ZN(n4154) );
  AND2_X1 U7278 ( .A1(n4130), .A2(n4108), .ZN(n25706) );
  BUF_X1 U7279 ( .A(n31276), .Z(n25670) );
  AOI22_X1 U7280 ( .A1(n25670), .A2(\xmem_data[96][7] ), .B1(n24158), .B2(
        \xmem_data[97][7] ), .ZN(n4112) );
  AOI22_X1 U7281 ( .A1(n24640), .A2(\xmem_data[98][7] ), .B1(n30552), .B2(
        \xmem_data[99][7] ), .ZN(n4111) );
  BUF_X1 U7282 ( .A(n14935), .Z(n25671) );
  AOI22_X1 U7283 ( .A1(n17041), .A2(\xmem_data[100][7] ), .B1(n25671), .B2(
        \xmem_data[101][7] ), .ZN(n4110) );
  BUF_X1 U7284 ( .A(n3464), .Z(n25672) );
  AOI22_X1 U7285 ( .A1(n25672), .A2(\xmem_data[102][7] ), .B1(n25574), .B2(
        \xmem_data[103][7] ), .ZN(n4109) );
  NAND4_X1 U7286 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(n4128)
         );
  BUF_X1 U7287 ( .A(n14912), .Z(n25677) );
  AOI22_X1 U7288 ( .A1(n14937), .A2(\xmem_data[104][7] ), .B1(n25677), .B2(
        \xmem_data[105][7] ), .ZN(n4116) );
  BUF_X1 U7289 ( .A(n14971), .Z(n25678) );
  AOI22_X1 U7290 ( .A1(n25678), .A2(\xmem_data[106][7] ), .B1(n24221), .B2(
        \xmem_data[107][7] ), .ZN(n4115) );
  BUF_X1 U7291 ( .A(n14882), .Z(n25679) );
  AOI22_X1 U7292 ( .A1(n17002), .A2(\xmem_data[108][7] ), .B1(n30598), .B2(
        \xmem_data[109][7] ), .ZN(n4114) );
  AOI22_X1 U7293 ( .A1(n3151), .A2(\xmem_data[110][7] ), .B1(n24622), .B2(
        \xmem_data[111][7] ), .ZN(n4113) );
  NAND4_X1 U7294 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4127)
         );
  AOI22_X1 U7295 ( .A1(n20782), .A2(\xmem_data[112][7] ), .B1(n20733), .B2(
        \xmem_data[113][7] ), .ZN(n4120) );
  BUF_X1 U7296 ( .A(n13127), .Z(n25684) );
  AOI22_X1 U7297 ( .A1(n25684), .A2(\xmem_data[114][7] ), .B1(n17050), .B2(
        \xmem_data[115][7] ), .ZN(n4119) );
  BUF_X1 U7298 ( .A(n31263), .Z(n25686) );
  BUF_X1 U7299 ( .A(n28974), .Z(n25685) );
  AOI22_X1 U7300 ( .A1(n25686), .A2(\xmem_data[116][7] ), .B1(n25685), .B2(
        \xmem_data[117][7] ), .ZN(n4118) );
  BUF_X1 U7301 ( .A(n4247), .Z(n13468) );
  BUF_X1 U7302 ( .A(n13468), .Z(n25687) );
  AOI22_X1 U7303 ( .A1(n3317), .A2(\xmem_data[118][7] ), .B1(n25687), .B2(
        \xmem_data[119][7] ), .ZN(n4117) );
  NAND4_X1 U7304 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4126)
         );
  BUF_X1 U7305 ( .A(n29064), .Z(n25692) );
  AOI22_X1 U7306 ( .A1(n25692), .A2(\xmem_data[120][7] ), .B1(n3217), .B2(
        \xmem_data[121][7] ), .ZN(n4124) );
  BUF_X1 U7307 ( .A(n14988), .Z(n25693) );
  AOI22_X1 U7308 ( .A1(n25693), .A2(\xmem_data[122][7] ), .B1(n23769), .B2(
        \xmem_data[123][7] ), .ZN(n4123) );
  BUF_X1 U7309 ( .A(n14926), .Z(n25694) );
  AOI22_X1 U7310 ( .A1(n25694), .A2(\xmem_data[124][7] ), .B1(n13444), .B2(
        \xmem_data[125][7] ), .ZN(n4122) );
  AOI22_X1 U7311 ( .A1(n28084), .A2(\xmem_data[126][7] ), .B1(n13474), .B2(
        \xmem_data[127][7] ), .ZN(n4121) );
  NAND4_X1 U7312 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4125)
         );
  OR4_X1 U7313 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), .ZN(n4152) );
  NOR2_X1 U7314 ( .A1(n4130), .A2(n4129), .ZN(n25704) );
  AOI22_X1 U7315 ( .A1(n25707), .A2(\xmem_data[64][7] ), .B1(n28415), .B2(
        \xmem_data[65][7] ), .ZN(n4134) );
  AOI22_X1 U7316 ( .A1(n25708), .A2(\xmem_data[66][7] ), .B1(n28515), .B2(
        \xmem_data[67][7] ), .ZN(n4133) );
  AOI22_X1 U7317 ( .A1(n28980), .A2(\xmem_data[68][7] ), .B1(n25709), .B2(
        \xmem_data[69][7] ), .ZN(n4132) );
  AOI22_X1 U7318 ( .A1(n29807), .A2(\xmem_data[70][7] ), .B1(n3208), .B2(
        \xmem_data[71][7] ), .ZN(n4131) );
  NAND4_X1 U7319 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4150)
         );
  AOI22_X1 U7320 ( .A1(n25573), .A2(\xmem_data[72][7] ), .B1(n25715), .B2(
        \xmem_data[73][7] ), .ZN(n4138) );
  AOI22_X1 U7321 ( .A1(n16990), .A2(\xmem_data[74][7] ), .B1(n25367), .B2(
        \xmem_data[75][7] ), .ZN(n4137) );
  AOI22_X1 U7322 ( .A1(n30899), .A2(\xmem_data[76][7] ), .B1(n29055), .B2(
        \xmem_data[77][7] ), .ZN(n4136) );
  AOI22_X1 U7323 ( .A1(n25718), .A2(\xmem_data[78][7] ), .B1(n27525), .B2(
        \xmem_data[79][7] ), .ZN(n4135) );
  NAND4_X1 U7324 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4149)
         );
  AOI22_X1 U7325 ( .A1(n3179), .A2(\xmem_data[80][7] ), .B1(n25723), .B2(
        \xmem_data[81][7] ), .ZN(n4142) );
  AOI22_X1 U7326 ( .A1(n25584), .A2(\xmem_data[82][7] ), .B1(n21059), .B2(
        \xmem_data[83][7] ), .ZN(n4141) );
  AOI22_X1 U7327 ( .A1(n25724), .A2(\xmem_data[84][7] ), .B1(n28366), .B2(
        \xmem_data[85][7] ), .ZN(n4140) );
  AOI22_X1 U7328 ( .A1(n25725), .A2(\xmem_data[86][7] ), .B1(n25360), .B2(
        \xmem_data[87][7] ), .ZN(n4139) );
  NAND4_X1 U7329 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4148)
         );
  AOI22_X1 U7330 ( .A1(n25730), .A2(\xmem_data[88][7] ), .B1(n3219), .B2(
        \xmem_data[89][7] ), .ZN(n4146) );
  AOI22_X1 U7331 ( .A1(n25731), .A2(\xmem_data[90][7] ), .B1(n24207), .B2(
        \xmem_data[91][7] ), .ZN(n4145) );
  AOI22_X1 U7332 ( .A1(n27938), .A2(\xmem_data[92][7] ), .B1(n29181), .B2(
        \xmem_data[93][7] ), .ZN(n4144) );
  AOI22_X1 U7333 ( .A1(n25732), .A2(\xmem_data[94][7] ), .B1(n3231), .B2(
        \xmem_data[95][7] ), .ZN(n4143) );
  NAND4_X1 U7334 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4147)
         );
  OR4_X1 U7335 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151) );
  AOI22_X1 U7336 ( .A1(n25706), .A2(n4152), .B1(n25704), .B2(n4151), .ZN(n4153) );
  XNOR2_X1 U7337 ( .A(n35120), .B(\fmem_data[6][3] ), .ZN(n30446) );
  XOR2_X1 U7338 ( .A(\fmem_data[6][3] ), .B(\fmem_data[6][2] ), .Z(n4156) );
  AND2_X1 U7339 ( .A1(n33598), .A2(n33596), .ZN(n4157) );
  NAND2_X1 U7340 ( .A1(n13474), .A2(\xmem_data[29][3] ), .ZN(n4190) );
  BUF_X1 U7341 ( .A(n14971), .Z(n23802) );
  BUF_X1 U7342 ( .A(n13452), .Z(n23801) );
  AOI22_X1 U7343 ( .A1(n23802), .A2(\xmem_data[8][3] ), .B1(n23801), .B2(
        \xmem_data[9][3] ), .ZN(n4162) );
  AOI22_X1 U7344 ( .A1(n29240), .A2(\xmem_data[10][3] ), .B1(n25581), .B2(
        \xmem_data[11][3] ), .ZN(n4161) );
  AOI22_X1 U7345 ( .A1(n29324), .A2(\xmem_data[12][3] ), .B1(n29126), .B2(
        \xmem_data[13][3] ), .ZN(n4160) );
  AOI22_X1 U7346 ( .A1(n24166), .A2(\xmem_data[14][3] ), .B1(n14981), .B2(
        \xmem_data[15][3] ), .ZN(n4159) );
  NAND4_X1 U7347 ( .A1(n4162), .A2(n4161), .A3(n4160), .A4(n4159), .ZN(n4165)
         );
  AOI22_X1 U7348 ( .A1(n16980), .A2(\xmem_data[20][3] ), .B1(n14875), .B2(
        \xmem_data[21][3] ), .ZN(n4163) );
  INV_X1 U7349 ( .A(n4163), .ZN(n4164) );
  NOR2_X1 U7350 ( .A1(n4165), .A2(n4164), .ZN(n4169) );
  AOI22_X1 U7351 ( .A1(n24694), .A2(\xmem_data[22][3] ), .B1(n3220), .B2(
        \xmem_data[23][3] ), .ZN(n4168) );
  AOI22_X1 U7352 ( .A1(n3380), .A2(\xmem_data[18][3] ), .B1(n30571), .B2(
        \xmem_data[19][3] ), .ZN(n4167) );
  AOI22_X1 U7353 ( .A1(n4527), .A2(\xmem_data[16][3] ), .B1(n17050), .B2(
        \xmem_data[17][3] ), .ZN(n4166) );
  NAND4_X1 U7354 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4186)
         );
  AOI22_X1 U7355 ( .A1(n17033), .A2(\xmem_data[24][3] ), .B1(n28476), .B2(
        \xmem_data[25][3] ), .ZN(n4176) );
  BUF_X1 U7356 ( .A(n14926), .Z(n23812) );
  BUF_X2 U7357 ( .A(n4204), .Z(n14890) );
  BUF_X1 U7358 ( .A(n14890), .Z(n23811) );
  AOI22_X1 U7359 ( .A1(n23812), .A2(\xmem_data[26][3] ), .B1(n23811), .B2(
        \xmem_data[27][3] ), .ZN(n4170) );
  INV_X1 U7360 ( .A(n4170), .ZN(n4174) );
  AOI22_X1 U7361 ( .A1(n23813), .A2(\xmem_data[30][3] ), .B1(n13475), .B2(
        \xmem_data[31][3] ), .ZN(n4172) );
  NAND2_X1 U7362 ( .A1(n20962), .A2(\xmem_data[28][3] ), .ZN(n4171) );
  NAND2_X1 U7363 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  NOR2_X1 U7364 ( .A1(n4174), .A2(n4173), .ZN(n4175) );
  NAND2_X1 U7365 ( .A1(n4176), .A2(n4175), .ZN(n4184) );
  BUF_X1 U7366 ( .A(n14997), .Z(n23792) );
  AOI22_X1 U7367 ( .A1(n23792), .A2(\xmem_data[0][3] ), .B1(n17012), .B2(
        \xmem_data[1][3] ), .ZN(n4182) );
  BUF_X1 U7368 ( .A(n14935), .Z(n23793) );
  AOI22_X1 U7369 ( .A1(n29272), .A2(\xmem_data[2][3] ), .B1(n23793), .B2(
        \xmem_data[3][3] ), .ZN(n4181) );
  BUF_X1 U7370 ( .A(n29187), .Z(n23795) );
  INV_X1 U7371 ( .A(n4444), .ZN(n14936) );
  BUF_X1 U7372 ( .A(n14936), .Z(n23794) );
  AOI22_X1 U7373 ( .A1(n28053), .A2(\xmem_data[4][3] ), .B1(n3208), .B2(
        \xmem_data[5][3] ), .ZN(n4180) );
  BUF_X1 U7374 ( .A(n13415), .Z(n23796) );
  AOI22_X1 U7375 ( .A1(n31330), .A2(\xmem_data[6][3] ), .B1(n23796), .B2(
        \xmem_data[7][3] ), .ZN(n4179) );
  NAND4_X1 U7376 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4183)
         );
  OR2_X1 U7377 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  NOR2_X1 U7378 ( .A1(n4186), .A2(n4185), .ZN(n4189) );
  NOR2_X1 U7379 ( .A1(n39053), .A2(n39035), .ZN(n10590) );
  NAND2_X1 U7380 ( .A1(n10590), .A2(n10589), .ZN(n4187) );
  NOR2_X1 U7381 ( .A1(n39041), .A2(n10972), .ZN(n10973) );
  INV_X1 U7382 ( .A(n10973), .ZN(n11381) );
  NOR2_X1 U7383 ( .A1(n8416), .A2(n11381), .ZN(n4188) );
  AOI21_X1 U7384 ( .B1(n39041), .B2(n4187), .A(n4188), .ZN(n4263) );
  XOR2_X1 U7385 ( .A(load_xaddr_val[6]), .B(n4188), .Z(n4213) );
  NOR2_X1 U7386 ( .A1(n4263), .A2(n4213), .ZN(n23822) );
  AOI21_X1 U7387 ( .B1(n4190), .B2(n4189), .A(n22877), .ZN(n4191) );
  INV_X1 U7388 ( .A(n4191), .ZN(n4268) );
  AND2_X1 U7389 ( .A1(n4263), .A2(n4213), .ZN(n23751) );
  AOI22_X1 U7390 ( .A1(n23792), .A2(\xmem_data[96][3] ), .B1(n24212), .B2(
        \xmem_data[97][3] ), .ZN(n4195) );
  BUF_X1 U7391 ( .A(n14898), .Z(n23715) );
  AOI22_X1 U7392 ( .A1(n28298), .A2(\xmem_data[98][3] ), .B1(n23715), .B2(
        \xmem_data[99][3] ), .ZN(n4194) );
  BUF_X2 U7393 ( .A(n14936), .Z(n23716) );
  AOI22_X1 U7394 ( .A1(n31354), .A2(\xmem_data[100][3] ), .B1(n23716), .B2(
        \xmem_data[101][3] ), .ZN(n4193) );
  AOI22_X1 U7395 ( .A1(n23717), .A2(\xmem_data[102][3] ), .B1(n31329), .B2(
        \xmem_data[103][3] ), .ZN(n4192) );
  NAND4_X1 U7396 ( .A1(n4195), .A2(n4194), .A3(n4193), .A4(n4192), .ZN(n4212)
         );
  BUF_X1 U7397 ( .A(n14971), .Z(n23722) );
  AOI22_X1 U7398 ( .A1(n23722), .A2(\xmem_data[104][3] ), .B1(n25435), .B2(
        \xmem_data[105][3] ), .ZN(n4199) );
  AOI22_X1 U7399 ( .A1(n24190), .A2(\xmem_data[106][3] ), .B1(n31361), .B2(
        \xmem_data[107][3] ), .ZN(n4198) );
  BUF_X1 U7400 ( .A(n14974), .Z(n23724) );
  BUF_X1 U7401 ( .A(n14914), .Z(n23723) );
  AOI22_X1 U7402 ( .A1(n23724), .A2(\xmem_data[108][3] ), .B1(n23723), .B2(
        \xmem_data[109][3] ), .ZN(n4197) );
  BUF_X1 U7403 ( .A(n14981), .Z(n23725) );
  AOI22_X1 U7404 ( .A1(n20734), .A2(\xmem_data[110][3] ), .B1(n23725), .B2(
        \xmem_data[111][3] ), .ZN(n4196) );
  NAND4_X1 U7405 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4211)
         );
  BUF_X1 U7406 ( .A(n13127), .Z(n23730) );
  AOI22_X1 U7407 ( .A1(n23730), .A2(\xmem_data[112][3] ), .B1(n20579), .B2(
        \xmem_data[113][3] ), .ZN(n4203) );
  AOI22_X1 U7408 ( .A1(n29124), .A2(\xmem_data[114][3] ), .B1(n30571), .B2(
        \xmem_data[115][3] ), .ZN(n4202) );
  BUF_X1 U7409 ( .A(n28973), .Z(n23732) );
  BUF_X1 U7410 ( .A(n13468), .Z(n23731) );
  AOI22_X1 U7411 ( .A1(n23732), .A2(\xmem_data[116][3] ), .B1(n23731), .B2(
        \xmem_data[117][3] ), .ZN(n4201) );
  BUF_X1 U7412 ( .A(n29064), .Z(n23734) );
  AOI22_X1 U7413 ( .A1(n23734), .A2(\xmem_data[118][3] ), .B1(n3217), .B2(
        \xmem_data[119][3] ), .ZN(n4200) );
  NAND4_X1 U7414 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4210)
         );
  BUF_X1 U7415 ( .A(n14988), .Z(n23740) );
  AOI22_X1 U7416 ( .A1(n23740), .A2(\xmem_data[120][3] ), .B1(n23739), .B2(
        \xmem_data[121][3] ), .ZN(n4208) );
  BUF_X1 U7417 ( .A(n14990), .Z(n23741) );
  BUF_X2 U7418 ( .A(n4204), .Z(n13444) );
  AOI22_X1 U7419 ( .A1(n23741), .A2(\xmem_data[122][3] ), .B1(n3256), .B2(
        \xmem_data[123][3] ), .ZN(n4207) );
  BUF_X1 U7420 ( .A(n14991), .Z(n23742) );
  AOI22_X1 U7421 ( .A1(n23742), .A2(\xmem_data[124][3] ), .B1(n27547), .B2(
        \xmem_data[125][3] ), .ZN(n4206) );
  AOI22_X1 U7422 ( .A1(n27447), .A2(\xmem_data[126][3] ), .B1(n13475), .B2(
        \xmem_data[127][3] ), .ZN(n4205) );
  NAND4_X1 U7423 ( .A1(n4208), .A2(n4207), .A3(n4206), .A4(n4205), .ZN(n4209)
         );
  OR4_X1 U7424 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4235) );
  INV_X1 U7425 ( .A(n4213), .ZN(n4264) );
  NOR2_X1 U7426 ( .A1(n4263), .A2(n4264), .ZN(n23713) );
  AOI22_X1 U7427 ( .A1(n24556), .A2(\xmem_data[64][3] ), .B1(n24132), .B2(
        \xmem_data[65][3] ), .ZN(n4217) );
  AOI22_X1 U7428 ( .A1(n3176), .A2(\xmem_data[66][3] ), .B1(n23715), .B2(
        \xmem_data[67][3] ), .ZN(n4216) );
  AOI22_X1 U7429 ( .A1(n25672), .A2(\xmem_data[68][3] ), .B1(n23716), .B2(
        \xmem_data[69][3] ), .ZN(n4215) );
  AOI22_X1 U7430 ( .A1(n23717), .A2(\xmem_data[70][3] ), .B1(n21006), .B2(
        \xmem_data[71][3] ), .ZN(n4214) );
  NAND4_X1 U7431 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4233)
         );
  AOI22_X1 U7432 ( .A1(n23722), .A2(\xmem_data[72][3] ), .B1(n24510), .B2(
        \xmem_data[73][3] ), .ZN(n4221) );
  AOI22_X1 U7433 ( .A1(n20593), .A2(\xmem_data[74][3] ), .B1(n23778), .B2(
        \xmem_data[75][3] ), .ZN(n4220) );
  AOI22_X1 U7434 ( .A1(n23724), .A2(\xmem_data[76][3] ), .B1(n23723), .B2(
        \xmem_data[77][3] ), .ZN(n4219) );
  AOI22_X1 U7435 ( .A1(n20818), .A2(\xmem_data[78][3] ), .B1(n23725), .B2(
        \xmem_data[79][3] ), .ZN(n4218) );
  NAND4_X1 U7436 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4232)
         );
  AOI22_X1 U7437 ( .A1(n23730), .A2(\xmem_data[80][3] ), .B1(n29125), .B2(
        \xmem_data[81][3] ), .ZN(n4225) );
  AOI22_X1 U7438 ( .A1(n20953), .A2(\xmem_data[82][3] ), .B1(n12471), .B2(
        \xmem_data[83][3] ), .ZN(n4224) );
  AOI22_X1 U7439 ( .A1(n23732), .A2(\xmem_data[84][3] ), .B1(n23731), .B2(
        \xmem_data[85][3] ), .ZN(n4223) );
  AOI22_X1 U7440 ( .A1(n23734), .A2(\xmem_data[86][3] ), .B1(n3220), .B2(
        \xmem_data[87][3] ), .ZN(n4222) );
  NAND4_X1 U7441 ( .A1(n4225), .A2(n4224), .A3(n4223), .A4(n4222), .ZN(n4231)
         );
  AOI22_X1 U7442 ( .A1(n23740), .A2(\xmem_data[88][3] ), .B1(n23739), .B2(
        \xmem_data[89][3] ), .ZN(n4229) );
  AOI22_X1 U7443 ( .A1(n23741), .A2(\xmem_data[90][3] ), .B1(n27994), .B2(
        \xmem_data[91][3] ), .ZN(n4228) );
  AOI22_X1 U7444 ( .A1(n23742), .A2(\xmem_data[92][3] ), .B1(n29045), .B2(
        \xmem_data[93][3] ), .ZN(n4227) );
  AOI22_X1 U7445 ( .A1(n27447), .A2(\xmem_data[94][3] ), .B1(n13475), .B2(
        \xmem_data[95][3] ), .ZN(n4226) );
  NAND4_X1 U7446 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230)
         );
  OR4_X1 U7447 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4234) );
  AOI22_X1 U7448 ( .A1(n23751), .A2(n4235), .B1(n23713), .B2(n4234), .ZN(n4267) );
  BUF_X1 U7449 ( .A(n14997), .Z(n23762) );
  BUF_X1 U7450 ( .A(n14934), .Z(n23761) );
  AOI22_X1 U7451 ( .A1(n23762), .A2(\xmem_data[32][3] ), .B1(n23761), .B2(
        \xmem_data[33][3] ), .ZN(n4241) );
  BUF_X2 U7452 ( .A(n4236), .Z(n13436) );
  BUF_X1 U7453 ( .A(n13436), .Z(n23763) );
  AOI22_X1 U7454 ( .A1(n23763), .A2(\xmem_data[34][3] ), .B1(n29309), .B2(
        \xmem_data[35][3] ), .ZN(n4240) );
  AOI22_X1 U7455 ( .A1(n28091), .A2(\xmem_data[36][3] ), .B1(n20586), .B2(
        \xmem_data[37][3] ), .ZN(n4239) );
  BUF_X1 U7456 ( .A(n13149), .Z(n23764) );
  AOI22_X1 U7457 ( .A1(n23764), .A2(\xmem_data[38][3] ), .B1(n25677), .B2(
        \xmem_data[39][3] ), .ZN(n4238) );
  NAND4_X1 U7458 ( .A1(n4241), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(n4262)
         );
  BUF_X1 U7459 ( .A(n14971), .Z(n23777) );
  BUF_X1 U7460 ( .A(n14913), .Z(n23776) );
  AOI22_X1 U7461 ( .A1(n23777), .A2(\xmem_data[40][3] ), .B1(n23776), .B2(
        \xmem_data[41][3] ), .ZN(n4246) );
  AOI22_X1 U7462 ( .A1(n28385), .A2(\xmem_data[42][3] ), .B1(n23778), .B2(
        \xmem_data[43][3] ), .ZN(n4245) );
  BUF_X1 U7463 ( .A(n14974), .Z(n23780) );
  BUF_X1 U7464 ( .A(n14914), .Z(n23779) );
  AOI22_X1 U7465 ( .A1(n23780), .A2(\xmem_data[44][3] ), .B1(n23779), .B2(
        \xmem_data[45][3] ), .ZN(n4244) );
  BUF_X1 U7466 ( .A(n14981), .Z(n23781) );
  AOI22_X1 U7467 ( .A1(n24606), .A2(\xmem_data[46][3] ), .B1(n23781), .B2(
        \xmem_data[47][3] ), .ZN(n4243) );
  NAND4_X1 U7468 ( .A1(n4246), .A2(n4245), .A3(n4244), .A4(n4243), .ZN(n4261)
         );
  BUF_X1 U7469 ( .A(n13127), .Z(n23753) );
  AOI22_X1 U7470 ( .A1(n23753), .A2(\xmem_data[48][3] ), .B1(n29125), .B2(
        \xmem_data[49][3] ), .ZN(n4252) );
  AOI22_X1 U7471 ( .A1(n25724), .A2(\xmem_data[50][3] ), .B1(n25357), .B2(
        \xmem_data[51][3] ), .ZN(n4251) );
  BUF_X1 U7472 ( .A(n28973), .Z(n23754) );
  AOI22_X1 U7473 ( .A1(n23754), .A2(\xmem_data[52][3] ), .B1(n28501), .B2(
        \xmem_data[53][3] ), .ZN(n4250) );
  BUF_X1 U7474 ( .A(n29064), .Z(n23756) );
  AOI22_X1 U7475 ( .A1(n23756), .A2(\xmem_data[54][3] ), .B1(n3221), .B2(
        \xmem_data[55][3] ), .ZN(n4249) );
  NAND4_X1 U7476 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4260)
         );
  BUF_X1 U7477 ( .A(n14988), .Z(n23770) );
  BUF_X1 U7478 ( .A(n14989), .Z(n23769) );
  AOI22_X1 U7479 ( .A1(n23770), .A2(\xmem_data[56][3] ), .B1(n23769), .B2(
        \xmem_data[57][3] ), .ZN(n4258) );
  AOI22_X1 U7480 ( .A1(n20725), .A2(\xmem_data[58][3] ), .B1(n27903), .B2(
        \xmem_data[59][3] ), .ZN(n4257) );
  BUF_X1 U7481 ( .A(n14928), .Z(n23771) );
  AOI22_X1 U7482 ( .A1(n3135), .A2(\xmem_data[60][3] ), .B1(n31252), .B2(
        \xmem_data[61][3] ), .ZN(n4256) );
  AOI22_X1 U7483 ( .A1(n27447), .A2(\xmem_data[62][3] ), .B1(n24158), .B2(
        \xmem_data[63][3] ), .ZN(n4255) );
  NAND4_X1 U7484 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4259)
         );
  OR4_X1 U7485 ( .A1(n4262), .A2(n4261), .A3(n4260), .A4(n4259), .ZN(n4265) );
  AND2_X1 U7486 ( .A1(n4264), .A2(n4263), .ZN(n23790) );
  NAND2_X1 U7487 ( .A1(n4265), .A2(n23790), .ZN(n4266) );
  XNOR2_X1 U7488 ( .A(n32317), .B(\fmem_data[4][7] ), .ZN(n24727) );
  XOR2_X1 U7489 ( .A(\fmem_data[4][6] ), .B(\fmem_data[4][7] ), .Z(n4269) );
  AOI22_X1 U7490 ( .A1(n23753), .A2(\xmem_data[48][4] ), .B1(n20769), .B2(
        \xmem_data[49][4] ), .ZN(n4273) );
  AOI22_X1 U7491 ( .A1(n30909), .A2(\xmem_data[50][4] ), .B1(n28037), .B2(
        \xmem_data[51][4] ), .ZN(n4272) );
  AOI22_X1 U7492 ( .A1(n23754), .A2(\xmem_data[52][4] ), .B1(n30589), .B2(
        \xmem_data[53][4] ), .ZN(n4271) );
  AOI22_X1 U7493 ( .A1(n23756), .A2(\xmem_data[54][4] ), .B1(n3222), .B2(
        \xmem_data[55][4] ), .ZN(n4270) );
  NAND4_X1 U7494 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4290)
         );
  AOI22_X1 U7495 ( .A1(n23777), .A2(\xmem_data[40][4] ), .B1(n23776), .B2(
        \xmem_data[41][4] ), .ZN(n4277) );
  AOI22_X1 U7496 ( .A1(n25575), .A2(\xmem_data[42][4] ), .B1(n23778), .B2(
        \xmem_data[43][4] ), .ZN(n4276) );
  AOI22_X1 U7497 ( .A1(n23780), .A2(\xmem_data[44][4] ), .B1(n23779), .B2(
        \xmem_data[45][4] ), .ZN(n4275) );
  AOI22_X1 U7498 ( .A1(n3209), .A2(\xmem_data[46][4] ), .B1(n23781), .B2(
        \xmem_data[47][4] ), .ZN(n4274) );
  NAND4_X1 U7499 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4288)
         );
  AOI22_X1 U7500 ( .A1(n23770), .A2(\xmem_data[56][4] ), .B1(n23769), .B2(
        \xmem_data[57][4] ), .ZN(n4281) );
  AOI22_X1 U7501 ( .A1(n29174), .A2(\xmem_data[58][4] ), .B1(n22711), .B2(
        \xmem_data[59][4] ), .ZN(n4280) );
  AOI22_X1 U7502 ( .A1(n3137), .A2(\xmem_data[60][4] ), .B1(n25514), .B2(
        \xmem_data[61][4] ), .ZN(n4279) );
  AOI22_X1 U7503 ( .A1(n27447), .A2(\xmem_data[62][4] ), .B1(n25456), .B2(
        \xmem_data[63][4] ), .ZN(n4278) );
  NAND4_X1 U7504 ( .A1(n4281), .A2(n4280), .A3(n4279), .A4(n4278), .ZN(n4287)
         );
  AOI22_X1 U7505 ( .A1(n23762), .A2(\xmem_data[32][4] ), .B1(n23761), .B2(
        \xmem_data[33][4] ), .ZN(n4285) );
  AOI22_X1 U7506 ( .A1(n23763), .A2(\xmem_data[34][4] ), .B1(n28090), .B2(
        \xmem_data[35][4] ), .ZN(n4284) );
  AOI22_X1 U7507 ( .A1(n27818), .A2(\xmem_data[36][4] ), .B1(n15000), .B2(
        \xmem_data[37][4] ), .ZN(n4283) );
  AOI22_X1 U7508 ( .A1(n23764), .A2(\xmem_data[38][4] ), .B1(n14970), .B2(
        \xmem_data[39][4] ), .ZN(n4282) );
  NAND4_X1 U7509 ( .A1(n4285), .A2(n4284), .A3(n4283), .A4(n4282), .ZN(n4286)
         );
  OR3_X1 U7510 ( .A1(n4288), .A2(n4287), .A3(n4286), .ZN(n4289) );
  OAI21_X1 U7511 ( .B1(n4290), .B2(n4289), .A(n23790), .ZN(n4291) );
  INV_X1 U7512 ( .A(n4291), .ZN(n4340) );
  AOI22_X1 U7513 ( .A1(n23730), .A2(\xmem_data[112][4] ), .B1(n29248), .B2(
        \xmem_data[113][4] ), .ZN(n4296) );
  AOI22_X1 U7514 ( .A1(n3380), .A2(\xmem_data[114][4] ), .B1(n28366), .B2(
        \xmem_data[115][4] ), .ZN(n4295) );
  AOI22_X1 U7515 ( .A1(n23732), .A2(\xmem_data[116][4] ), .B1(n23731), .B2(
        \xmem_data[117][4] ), .ZN(n4294) );
  AND2_X1 U7516 ( .A1(n3218), .A2(\xmem_data[119][4] ), .ZN(n4292) );
  AOI21_X1 U7517 ( .B1(n23734), .B2(\xmem_data[118][4] ), .A(n4292), .ZN(n4293) );
  NAND4_X1 U7518 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), .ZN(n4313)
         );
  AOI22_X1 U7519 ( .A1(n23722), .A2(\xmem_data[104][4] ), .B1(n25435), .B2(
        \xmem_data[105][4] ), .ZN(n4300) );
  AOI22_X1 U7520 ( .A1(n30557), .A2(\xmem_data[106][4] ), .B1(n21009), .B2(
        \xmem_data[107][4] ), .ZN(n4299) );
  AOI22_X1 U7521 ( .A1(n23724), .A2(\xmem_data[108][4] ), .B1(n23723), .B2(
        \xmem_data[109][4] ), .ZN(n4298) );
  AOI22_X1 U7522 ( .A1(n31316), .A2(\xmem_data[110][4] ), .B1(n23725), .B2(
        \xmem_data[111][4] ), .ZN(n4297) );
  NAND4_X1 U7523 ( .A1(n4300), .A2(n4299), .A3(n4298), .A4(n4297), .ZN(n4311)
         );
  AOI22_X1 U7524 ( .A1(n23740), .A2(\xmem_data[120][4] ), .B1(n23739), .B2(
        \xmem_data[121][4] ), .ZN(n4304) );
  AOI22_X1 U7525 ( .A1(n23741), .A2(\xmem_data[122][4] ), .B1(n21068), .B2(
        \xmem_data[123][4] ), .ZN(n4303) );
  AOI22_X1 U7526 ( .A1(n23742), .A2(\xmem_data[124][4] ), .B1(n23771), .B2(
        \xmem_data[125][4] ), .ZN(n4302) );
  AOI22_X1 U7527 ( .A1(n27447), .A2(\xmem_data[126][4] ), .B1(n13475), .B2(
        \xmem_data[127][4] ), .ZN(n4301) );
  NAND4_X1 U7528 ( .A1(n4304), .A2(n4303), .A3(n4302), .A4(n4301), .ZN(n4310)
         );
  AOI22_X1 U7529 ( .A1(n28309), .A2(\xmem_data[96][4] ), .B1(n28375), .B2(
        \xmem_data[97][4] ), .ZN(n4308) );
  AOI22_X1 U7530 ( .A1(n28298), .A2(\xmem_data[98][4] ), .B1(n23715), .B2(
        \xmem_data[99][4] ), .ZN(n4307) );
  AOI22_X1 U7531 ( .A1(n21048), .A2(\xmem_data[100][4] ), .B1(n23716), .B2(
        \xmem_data[101][4] ), .ZN(n4306) );
  AOI22_X1 U7532 ( .A1(n23717), .A2(\xmem_data[102][4] ), .B1(n29048), .B2(
        \xmem_data[103][4] ), .ZN(n4305) );
  NAND4_X1 U7533 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), .ZN(n4309)
         );
  OR3_X1 U7534 ( .A1(n4311), .A2(n4310), .A3(n4309), .ZN(n4312) );
  OAI21_X1 U7535 ( .B1(n4313), .B2(n4312), .A(n23751), .ZN(n4314) );
  INV_X1 U7536 ( .A(n4314), .ZN(n4339) );
  AOI22_X1 U7537 ( .A1(n23753), .A2(\xmem_data[80][4] ), .B1(n20707), .B2(
        \xmem_data[81][4] ), .ZN(n4319) );
  AOI22_X1 U7538 ( .A1(n25630), .A2(\xmem_data[82][4] ), .B1(n22729), .B2(
        \xmem_data[83][4] ), .ZN(n4318) );
  AOI22_X1 U7539 ( .A1(n23754), .A2(\xmem_data[84][4] ), .B1(n25687), .B2(
        \xmem_data[85][4] ), .ZN(n4317) );
  AND2_X1 U7540 ( .A1(n3221), .A2(\xmem_data[87][4] ), .ZN(n4315) );
  AOI21_X1 U7541 ( .B1(n23756), .B2(\xmem_data[86][4] ), .A(n4315), .ZN(n4316)
         );
  NAND4_X1 U7542 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4336)
         );
  AOI22_X1 U7543 ( .A1(n23762), .A2(\xmem_data[64][4] ), .B1(n23761), .B2(
        \xmem_data[65][4] ), .ZN(n4323) );
  AOI22_X1 U7544 ( .A1(n23763), .A2(\xmem_data[66][4] ), .B1(n28052), .B2(
        \xmem_data[67][4] ), .ZN(n4322) );
  AOI22_X1 U7545 ( .A1(n27455), .A2(\xmem_data[68][4] ), .B1(n29162), .B2(
        \xmem_data[69][4] ), .ZN(n4321) );
  AOI22_X1 U7546 ( .A1(n23764), .A2(\xmem_data[70][4] ), .B1(n21006), .B2(
        \xmem_data[71][4] ), .ZN(n4320) );
  NAND4_X1 U7547 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4334)
         );
  AOI22_X1 U7548 ( .A1(n23770), .A2(\xmem_data[88][4] ), .B1(n23769), .B2(
        \xmem_data[89][4] ), .ZN(n4327) );
  AOI22_X1 U7549 ( .A1(n24141), .A2(\xmem_data[90][4] ), .B1(n25486), .B2(
        \xmem_data[91][4] ), .ZN(n4326) );
  AOI22_X1 U7550 ( .A1(n30698), .A2(\xmem_data[92][4] ), .B1(n28510), .B2(
        \xmem_data[93][4] ), .ZN(n4325) );
  AOI22_X1 U7551 ( .A1(n27447), .A2(\xmem_data[94][4] ), .B1(n3358), .B2(
        \xmem_data[95][4] ), .ZN(n4324) );
  NAND4_X1 U7552 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(n4333)
         );
  AOI22_X1 U7553 ( .A1(n23777), .A2(\xmem_data[72][4] ), .B1(n23776), .B2(
        \xmem_data[73][4] ), .ZN(n4331) );
  AOI22_X1 U7554 ( .A1(n25575), .A2(\xmem_data[74][4] ), .B1(n23778), .B2(
        \xmem_data[75][4] ), .ZN(n4330) );
  AOI22_X1 U7555 ( .A1(n23780), .A2(\xmem_data[76][4] ), .B1(n23779), .B2(
        \xmem_data[77][4] ), .ZN(n4329) );
  AOI22_X1 U7556 ( .A1(n22719), .A2(\xmem_data[78][4] ), .B1(n23781), .B2(
        \xmem_data[79][4] ), .ZN(n4328) );
  NAND4_X1 U7557 ( .A1(n4331), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n4332)
         );
  OR3_X1 U7558 ( .A1(n4334), .A2(n4333), .A3(n4332), .ZN(n4335) );
  OAI21_X1 U7559 ( .B1(n4336), .B2(n4335), .A(n23713), .ZN(n4337) );
  INV_X1 U7560 ( .A(n4337), .ZN(n4338) );
  NOR3_X1 U7561 ( .A1(n4340), .A2(n4339), .A3(n4338), .ZN(n4365) );
  AOI22_X1 U7562 ( .A1(n30698), .A2(\xmem_data[28][4] ), .B1(n24657), .B2(
        \xmem_data[29][4] ), .ZN(n4341) );
  INV_X1 U7563 ( .A(n4341), .ZN(n4362) );
  AOI22_X1 U7564 ( .A1(n28772), .A2(\xmem_data[16][4] ), .B1(n30601), .B2(
        \xmem_data[17][4] ), .ZN(n4345) );
  AOI22_X1 U7565 ( .A1(n30862), .A2(\xmem_data[18][4] ), .B1(n28037), .B2(
        \xmem_data[19][4] ), .ZN(n4344) );
  AOI22_X1 U7566 ( .A1(n24693), .A2(\xmem_data[20][4] ), .B1(n31347), .B2(
        \xmem_data[21][4] ), .ZN(n4343) );
  AOI22_X1 U7567 ( .A1(n25508), .A2(\xmem_data[22][4] ), .B1(n3220), .B2(
        \xmem_data[23][4] ), .ZN(n4342) );
  NAND4_X1 U7568 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4360)
         );
  AOI22_X1 U7569 ( .A1(n23802), .A2(\xmem_data[8][4] ), .B1(n23801), .B2(
        \xmem_data[9][4] ), .ZN(n4349) );
  AOI22_X1 U7570 ( .A1(n28460), .A2(\xmem_data[10][4] ), .B1(n24117), .B2(
        \xmem_data[11][4] ), .ZN(n4348) );
  AOI22_X1 U7571 ( .A1(n30686), .A2(\xmem_data[12][4] ), .B1(n20781), .B2(
        \xmem_data[13][4] ), .ZN(n4347) );
  AOI22_X1 U7572 ( .A1(n24467), .A2(\xmem_data[14][4] ), .B1(n25359), .B2(
        \xmem_data[15][4] ), .ZN(n4346) );
  NAND4_X1 U7573 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(n4359)
         );
  AOI22_X1 U7574 ( .A1(n23792), .A2(\xmem_data[0][4] ), .B1(n24212), .B2(
        \xmem_data[1][4] ), .ZN(n4353) );
  AOI22_X1 U7575 ( .A1(n17041), .A2(\xmem_data[2][4] ), .B1(n23793), .B2(
        \xmem_data[3][4] ), .ZN(n4352) );
  AOI22_X1 U7576 ( .A1(n24213), .A2(\xmem_data[4][4] ), .B1(n3208), .B2(
        \xmem_data[5][4] ), .ZN(n4351) );
  AOI22_X1 U7577 ( .A1(n24214), .A2(\xmem_data[6][4] ), .B1(n23796), .B2(
        \xmem_data[7][4] ), .ZN(n4350) );
  NAND4_X1 U7578 ( .A1(n4353), .A2(n4352), .A3(n4351), .A4(n4350), .ZN(n4358)
         );
  AOI22_X1 U7579 ( .A1(n23812), .A2(\xmem_data[26][4] ), .B1(n23811), .B2(
        \xmem_data[27][4] ), .ZN(n4356) );
  AOI22_X1 U7580 ( .A1(n23813), .A2(\xmem_data[30][4] ), .B1(n13475), .B2(
        \xmem_data[31][4] ), .ZN(n4355) );
  AOI22_X1 U7581 ( .A1(n23770), .A2(\xmem_data[24][4] ), .B1(n27444), .B2(
        \xmem_data[25][4] ), .ZN(n4354) );
  NAND3_X1 U7582 ( .A1(n4356), .A2(n4355), .A3(n4354), .ZN(n4357) );
  OR4_X1 U7583 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4361) );
  NOR2_X1 U7584 ( .A1(n4362), .A2(n4361), .ZN(n4363) );
  NAND2_X1 U7585 ( .A1(n4365), .A2(n4364), .ZN(n32584) );
  XNOR2_X1 U7586 ( .A(n32584), .B(\fmem_data[4][7] ), .ZN(n33305) );
  OAI22_X1 U7587 ( .A1(n24727), .A2(n35748), .B1(n33305), .B2(n35749), .ZN(
        n34669) );
  BUF_X1 U7588 ( .A(n14919), .Z(n22751) );
  AND2_X1 U7589 ( .A1(n22751), .A2(\xmem_data[16][7] ), .ZN(n4367) );
  AOI21_X1 U7590 ( .B1(n28192), .B2(\xmem_data[17][7] ), .A(n4367), .ZN(n4372)
         );
  INV_X1 U7591 ( .A(n4456), .ZN(n13457) );
  AOI22_X1 U7592 ( .A1(n17050), .A2(\xmem_data[18][7] ), .B1(n24607), .B2(
        \xmem_data[19][7] ), .ZN(n4371) );
  AOI22_X1 U7593 ( .A1(n22752), .A2(\xmem_data[20][7] ), .B1(n3414), .B2(
        \xmem_data[21][7] ), .ZN(n4370) );
  BUF_X1 U7594 ( .A(n13468), .Z(n22753) );
  AOI22_X1 U7595 ( .A1(n22753), .A2(\xmem_data[22][7] ), .B1(n29064), .B2(
        \xmem_data[23][7] ), .ZN(n4369) );
  NAND4_X1 U7596 ( .A1(n4372), .A2(n4371), .A3(n4370), .A4(n4369), .ZN(n4387)
         );
  AOI22_X1 U7597 ( .A1(n27918), .A2(\xmem_data[8][7] ), .B1(n21008), .B2(
        \xmem_data[9][7] ), .ZN(n4376) );
  AOI22_X1 U7598 ( .A1(n29238), .A2(\xmem_data[10][7] ), .B1(n3177), .B2(
        \xmem_data[11][7] ), .ZN(n4375) );
  AOI22_X1 U7599 ( .A1(n25581), .A2(\xmem_data[12][7] ), .B1(n3337), .B2(
        \xmem_data[13][7] ), .ZN(n4374) );
  AOI22_X1 U7600 ( .A1(n28983), .A2(\xmem_data[14][7] ), .B1(n3171), .B2(
        \xmem_data[15][7] ), .ZN(n4373) );
  NAND4_X1 U7601 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4386)
         );
  BUF_X1 U7602 ( .A(n14935), .Z(n22741) );
  AOI22_X1 U7603 ( .A1(n22741), .A2(\xmem_data[4][7] ), .B1(n28154), .B2(
        \xmem_data[5][7] ), .ZN(n4380) );
  BUF_X1 U7604 ( .A(n14934), .Z(n22740) );
  AOI22_X1 U7605 ( .A1(n22740), .A2(\xmem_data[2][7] ), .B1(n29023), .B2(
        \xmem_data[3][7] ), .ZN(n4379) );
  INV_X1 U7606 ( .A(n4536), .ZN(n10999) );
  BUF_X1 U7607 ( .A(n10999), .Z(n22739) );
  BUF_X1 U7608 ( .A(n14997), .Z(n22738) );
  AOI22_X1 U7609 ( .A1(n22739), .A2(\xmem_data[0][7] ), .B1(n22738), .B2(
        \xmem_data[1][7] ), .ZN(n4378) );
  BUF_X1 U7610 ( .A(n14936), .Z(n22742) );
  AOI22_X1 U7611 ( .A1(n22742), .A2(\xmem_data[6][7] ), .B1(n25635), .B2(
        \xmem_data[7][7] ), .ZN(n4377) );
  NAND4_X1 U7612 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(n4385)
         );
  BUF_X1 U7613 ( .A(n14890), .Z(n22759) );
  AOI22_X1 U7614 ( .A1(n22759), .A2(\xmem_data[28][7] ), .B1(n20962), .B2(
        \xmem_data[29][7] ), .ZN(n4383) );
  BUF_X1 U7615 ( .A(n14926), .Z(n22758) );
  AOI22_X1 U7616 ( .A1(n27507), .A2(\xmem_data[26][7] ), .B1(n22758), .B2(
        \xmem_data[27][7] ), .ZN(n4382) );
  AOI22_X1 U7617 ( .A1(n3218), .A2(\xmem_data[24][7] ), .B1(n28367), .B2(
        \xmem_data[25][7] ), .ZN(n4381) );
  NAND3_X1 U7618 ( .A1(n4383), .A2(n4382), .A3(n4381), .ZN(n4384) );
  NOR4_X1 U7619 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(n4390)
         );
  NAND2_X1 U7620 ( .A1(n25670), .A2(\xmem_data[31][7] ), .ZN(n4388) );
  NAND3_X1 U7621 ( .A1(n4390), .A2(n4389), .A3(n4388), .ZN(n4394) );
  NOR2_X1 U7622 ( .A1(n3402), .A2(n6172), .ZN(n14907) );
  INV_X1 U7623 ( .A(n14907), .ZN(n5090) );
  NAND2_X1 U7624 ( .A1(n7216), .A2(n5090), .ZN(n4392) );
  NOR2_X1 U7625 ( .A1(n39041), .A2(n4392), .ZN(n4393) );
  AOI21_X1 U7626 ( .B1(n4499), .B2(n4392), .A(n4393), .ZN(n4463) );
  INV_X1 U7627 ( .A(n20311), .ZN(n20978) );
  OAI22_X1 U7628 ( .A1(n4393), .A2(n39040), .B1(n20978), .B2(n4392), .ZN(n4462) );
  NOR2_X1 U7629 ( .A1(n4463), .A2(n4462), .ZN(n22768) );
  AOI22_X1 U7630 ( .A1(n25723), .A2(\xmem_data[80][7] ), .B1(n21060), .B2(
        \xmem_data[81][7] ), .ZN(n4398) );
  BUF_X1 U7631 ( .A(n13457), .Z(n22727) );
  AOI22_X1 U7632 ( .A1(n22727), .A2(\xmem_data[82][7] ), .B1(n20710), .B2(
        \xmem_data[83][7] ), .ZN(n4397) );
  BUF_X1 U7633 ( .A(n28974), .Z(n22729) );
  BUF_X1 U7634 ( .A(n28973), .Z(n22728) );
  AOI22_X1 U7635 ( .A1(n22729), .A2(\xmem_data[84][7] ), .B1(n22728), .B2(
        \xmem_data[85][7] ), .ZN(n4396) );
  AOI22_X1 U7636 ( .A1(n24172), .A2(\xmem_data[86][7] ), .B1(n24631), .B2(
        \xmem_data[87][7] ), .ZN(n4395) );
  NAND4_X1 U7637 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(n4417)
         );
  BUF_X1 U7638 ( .A(n14912), .Z(n22718) );
  BUF_X1 U7639 ( .A(n14971), .Z(n22717) );
  AOI22_X1 U7640 ( .A1(n22718), .A2(\xmem_data[72][7] ), .B1(n22717), .B2(
        \xmem_data[73][7] ), .ZN(n4403) );
  AOI22_X1 U7641 ( .A1(n25367), .A2(\xmem_data[74][7] ), .B1(n27952), .B2(
        \xmem_data[75][7] ), .ZN(n4402) );
  AOI22_X1 U7642 ( .A1(n29089), .A2(\xmem_data[76][7] ), .B1(n3270), .B2(
        \xmem_data[77][7] ), .ZN(n4401) );
  BUF_X1 U7643 ( .A(n13486), .Z(n22719) );
  AOI22_X1 U7644 ( .A1(n24622), .A2(\xmem_data[78][7] ), .B1(n22719), .B2(
        \xmem_data[79][7] ), .ZN(n4400) );
  NAND4_X1 U7645 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(n4415)
         );
  BUF_X1 U7646 ( .A(n10999), .Z(n22701) );
  AOI22_X1 U7647 ( .A1(n22701), .A2(\xmem_data[64][7] ), .B1(n28051), .B2(
        \xmem_data[65][7] ), .ZN(n4408) );
  BUF_X1 U7648 ( .A(n14934), .Z(n22702) );
  AOI22_X1 U7649 ( .A1(n22702), .A2(\xmem_data[66][7] ), .B1(n30514), .B2(
        \xmem_data[67][7] ), .ZN(n4407) );
  AOI22_X1 U7650 ( .A1(n22703), .A2(\xmem_data[68][7] ), .B1(n17018), .B2(
        \xmem_data[69][7] ), .ZN(n4406) );
  AOI22_X1 U7651 ( .A1(n20543), .A2(\xmem_data[70][7] ), .B1(n21007), .B2(
        \xmem_data[71][7] ), .ZN(n4405) );
  NAND4_X1 U7652 ( .A1(n4408), .A2(n4407), .A3(n4406), .A4(n4405), .ZN(n4414)
         );
  BUF_X1 U7653 ( .A(n14988), .Z(n22708) );
  AOI22_X1 U7654 ( .A1(n3219), .A2(\xmem_data[88][7] ), .B1(n22708), .B2(
        \xmem_data[89][7] ), .ZN(n4412) );
  BUF_X1 U7655 ( .A(n14989), .Z(n22710) );
  BUF_X1 U7656 ( .A(n14990), .Z(n22709) );
  AOI22_X1 U7657 ( .A1(n22710), .A2(\xmem_data[90][7] ), .B1(n22709), .B2(
        \xmem_data[91][7] ), .ZN(n4411) );
  BUF_X1 U7658 ( .A(n14927), .Z(n22711) );
  AOI22_X1 U7659 ( .A1(n22711), .A2(\xmem_data[92][7] ), .B1(n29157), .B2(
        \xmem_data[93][7] ), .ZN(n4410) );
  BUF_X1 U7660 ( .A(n25604), .Z(n22712) );
  AOI22_X1 U7661 ( .A1(n27547), .A2(\xmem_data[94][7] ), .B1(n22712), .B2(
        \xmem_data[95][7] ), .ZN(n4409) );
  NAND4_X1 U7662 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4413)
         );
  INV_X1 U7663 ( .A(n4462), .ZN(n4437) );
  NOR2_X1 U7664 ( .A1(n4463), .A2(n4437), .ZN(n22663) );
  AOI22_X1 U7665 ( .A1(n25723), .A2(\xmem_data[48][7] ), .B1(n28192), .B2(
        \xmem_data[49][7] ), .ZN(n4421) );
  AOI22_X1 U7666 ( .A1(n22727), .A2(\xmem_data[50][7] ), .B1(n25408), .B2(
        \xmem_data[51][7] ), .ZN(n4420) );
  AOI22_X1 U7667 ( .A1(n22729), .A2(\xmem_data[52][7] ), .B1(n22728), .B2(
        \xmem_data[53][7] ), .ZN(n4419) );
  AOI22_X1 U7668 ( .A1(n30589), .A2(\xmem_data[54][7] ), .B1(n28044), .B2(
        \xmem_data[55][7] ), .ZN(n4418) );
  NAND4_X1 U7669 ( .A1(n4421), .A2(n4420), .A3(n4419), .A4(n4418), .ZN(n4439)
         );
  AOI22_X1 U7670 ( .A1(n22718), .A2(\xmem_data[40][7] ), .B1(n22717), .B2(
        \xmem_data[41][7] ), .ZN(n4425) );
  AOI22_X1 U7671 ( .A1(n24510), .A2(\xmem_data[42][7] ), .B1(n30849), .B2(
        \xmem_data[43][7] ), .ZN(n4424) );
  AOI22_X1 U7672 ( .A1(n31361), .A2(\xmem_data[44][7] ), .B1(n3329), .B2(
        \xmem_data[45][7] ), .ZN(n4423) );
  AOI22_X1 U7673 ( .A1(n31314), .A2(\xmem_data[46][7] ), .B1(n22719), .B2(
        \xmem_data[47][7] ), .ZN(n4422) );
  NAND4_X1 U7674 ( .A1(n4425), .A2(n4424), .A3(n4423), .A4(n4422), .ZN(n4436)
         );
  AOI22_X1 U7675 ( .A1(n22701), .A2(\xmem_data[32][7] ), .B1(n24640), .B2(
        \xmem_data[33][7] ), .ZN(n4429) );
  AOI22_X1 U7676 ( .A1(n22702), .A2(\xmem_data[34][7] ), .B1(n23763), .B2(
        \xmem_data[35][7] ), .ZN(n4428) );
  AOI22_X1 U7677 ( .A1(n22703), .A2(\xmem_data[36][7] ), .B1(n24458), .B2(
        \xmem_data[37][7] ), .ZN(n4427) );
  AOI22_X1 U7678 ( .A1(n24134), .A2(\xmem_data[38][7] ), .B1(n20542), .B2(
        \xmem_data[39][7] ), .ZN(n4426) );
  NAND4_X1 U7679 ( .A1(n4429), .A2(n4428), .A3(n4427), .A4(n4426), .ZN(n4435)
         );
  AOI22_X1 U7680 ( .A1(n3222), .A2(\xmem_data[56][7] ), .B1(n22708), .B2(
        \xmem_data[57][7] ), .ZN(n4433) );
  AOI22_X1 U7681 ( .A1(n22710), .A2(\xmem_data[58][7] ), .B1(n22709), .B2(
        \xmem_data[59][7] ), .ZN(n4432) );
  AOI22_X1 U7682 ( .A1(n22711), .A2(\xmem_data[60][7] ), .B1(n25377), .B2(
        \xmem_data[61][7] ), .ZN(n4431) );
  AOI22_X1 U7683 ( .A1(n28343), .A2(\xmem_data[62][7] ), .B1(n22712), .B2(
        \xmem_data[63][7] ), .ZN(n4430) );
  NAND4_X1 U7684 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4434)
         );
  BUF_X1 U7685 ( .A(n14971), .Z(n22682) );
  AOI22_X1 U7686 ( .A1(n29048), .A2(\xmem_data[104][7] ), .B1(n22682), .B2(
        \xmem_data[105][7] ), .ZN(n4443) );
  BUF_X1 U7687 ( .A(n14972), .Z(n22683) );
  AOI22_X1 U7688 ( .A1(n31360), .A2(\xmem_data[106][7] ), .B1(n22683), .B2(
        \xmem_data[107][7] ), .ZN(n4442) );
  AOI22_X1 U7689 ( .A1(n29089), .A2(\xmem_data[108][7] ), .B1(n24571), .B2(
        \xmem_data[109][7] ), .ZN(n4441) );
  BUF_X1 U7690 ( .A(n14914), .Z(n22685) );
  BUF_X1 U7691 ( .A(n13486), .Z(n22684) );
  AOI22_X1 U7692 ( .A1(n22685), .A2(\xmem_data[110][7] ), .B1(n22684), .B2(
        \xmem_data[111][7] ), .ZN(n4440) );
  NAND4_X1 U7693 ( .A1(n4443), .A2(n4442), .A3(n4441), .A4(n4440), .ZN(n4455)
         );
  AOI22_X1 U7694 ( .A1(n3357), .A2(\xmem_data[96][7] ), .B1(n25424), .B2(
        \xmem_data[97][7] ), .ZN(n4448) );
  BUF_X1 U7695 ( .A(n14934), .Z(n22675) );
  AOI22_X1 U7696 ( .A1(n22675), .A2(\xmem_data[98][7] ), .B1(n25567), .B2(
        \xmem_data[99][7] ), .ZN(n4447) );
  BUF_X1 U7697 ( .A(n14898), .Z(n22674) );
  AOI22_X1 U7698 ( .A1(n22674), .A2(\xmem_data[100][7] ), .B1(n24458), .B2(
        \xmem_data[101][7] ), .ZN(n4446) );
  BUF_X1 U7699 ( .A(n13188), .Z(n22677) );
  BUF_X1 U7700 ( .A(n13149), .Z(n22676) );
  AOI22_X1 U7701 ( .A1(n22677), .A2(\xmem_data[102][7] ), .B1(n22676), .B2(
        \xmem_data[103][7] ), .ZN(n4445) );
  NAND4_X1 U7702 ( .A1(n4448), .A2(n4447), .A3(n4446), .A4(n4445), .ZN(n4454)
         );
  AOI22_X1 U7703 ( .A1(n3222), .A2(\xmem_data[120][7] ), .B1(n23770), .B2(
        \xmem_data[121][7] ), .ZN(n4452) );
  BUF_X1 U7704 ( .A(n14989), .Z(n22667) );
  BUF_X1 U7705 ( .A(n14990), .Z(n22666) );
  AOI22_X1 U7706 ( .A1(n22667), .A2(\xmem_data[122][7] ), .B1(n22666), .B2(
        \xmem_data[123][7] ), .ZN(n4451) );
  BUF_X1 U7707 ( .A(n14927), .Z(n22669) );
  BUF_X1 U7708 ( .A(n14991), .Z(n22668) );
  AOI22_X1 U7709 ( .A1(n22669), .A2(\xmem_data[124][7] ), .B1(n22668), .B2(
        \xmem_data[125][7] ), .ZN(n4450) );
  AOI22_X1 U7710 ( .A1(n28343), .A2(\xmem_data[126][7] ), .B1(n28374), .B2(
        \xmem_data[127][7] ), .ZN(n4449) );
  NAND4_X1 U7711 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n4449), .ZN(n4453)
         );
  AOI22_X1 U7712 ( .A1(n28468), .A2(\xmem_data[112][7] ), .B1(n30257), .B2(
        \xmem_data[113][7] ), .ZN(n4461) );
  AOI22_X1 U7713 ( .A1(n30524), .A2(\xmem_data[114][7] ), .B1(n28038), .B2(
        \xmem_data[115][7] ), .ZN(n4460) );
  AOI22_X1 U7714 ( .A1(n24573), .A2(\xmem_data[116][7] ), .B1(n3414), .B2(
        \xmem_data[117][7] ), .ZN(n4459) );
  AND2_X1 U7715 ( .A1(n29173), .A2(\xmem_data[118][7] ), .ZN(n4457) );
  AOI21_X1 U7716 ( .B1(n29064), .B2(\xmem_data[119][7] ), .A(n4457), .ZN(n4458) );
  NAND4_X1 U7717 ( .A1(n4461), .A2(n4460), .A3(n4459), .A4(n4458), .ZN(n4464)
         );
  AND2_X1 U7718 ( .A1(n4463), .A2(n4462), .ZN(n22698) );
  XNOR2_X1 U7719 ( .A(n35405), .B(\fmem_data[5][3] ), .ZN(n30159) );
  INV_X1 U7720 ( .A(n4470), .ZN(n34668) );
  AOI22_X1 U7721 ( .A1(n29832), .A2(\xmem_data[10][4] ), .B1(n25562), .B2(
        \xmem_data[11][4] ), .ZN(n4477) );
  AOI22_X1 U7722 ( .A1(n25354), .A2(\xmem_data[8][4] ), .B1(n3222), .B2(
        \xmem_data[9][4] ), .ZN(n4471) );
  INV_X1 U7723 ( .A(n4471), .ZN(n4475) );
  BUF_X1 U7724 ( .A(n14927), .Z(n27994) );
  AOI22_X1 U7725 ( .A1(n27904), .A2(\xmem_data[12][4] ), .B1(n27994), .B2(
        \xmem_data[13][4] ), .ZN(n4473) );
  NAND2_X1 U7726 ( .A1(n3140), .A2(\xmem_data[14][4] ), .ZN(n4472) );
  NAND2_X1 U7727 ( .A1(n4473), .A2(n4472), .ZN(n4474) );
  NOR2_X1 U7728 ( .A1(n4475), .A2(n4474), .ZN(n4476) );
  NAND2_X1 U7729 ( .A1(n4477), .A2(n4476), .ZN(n4484) );
  BUF_X1 U7730 ( .A(n10999), .Z(n27988) );
  AOI22_X1 U7731 ( .A1(n25670), .A2(\xmem_data[16][4] ), .B1(n27988), .B2(
        \xmem_data[17][4] ), .ZN(n4482) );
  AOI22_X1 U7732 ( .A1(n30608), .A2(\xmem_data[18][4] ), .B1(n21075), .B2(
        \xmem_data[19][4] ), .ZN(n4481) );
  AOI22_X1 U7733 ( .A1(n25425), .A2(\xmem_data[20][4] ), .B1(n29271), .B2(
        \xmem_data[21][4] ), .ZN(n4480) );
  BUF_X1 U7734 ( .A(n14936), .Z(n27989) );
  AOI22_X1 U7735 ( .A1(n24545), .A2(\xmem_data[22][4] ), .B1(n27989), .B2(
        \xmem_data[23][4] ), .ZN(n4479) );
  NAND4_X1 U7736 ( .A1(n4482), .A2(n4481), .A3(n4480), .A4(n4479), .ZN(n4483)
         );
  OR2_X1 U7737 ( .A1(n4484), .A2(n4483), .ZN(n4503) );
  BUF_X1 U7738 ( .A(n14919), .Z(n27981) );
  AOI22_X1 U7739 ( .A1(n30497), .A2(\xmem_data[0][4] ), .B1(n27981), .B2(
        \xmem_data[1][4] ), .ZN(n4488) );
  AOI22_X1 U7740 ( .A1(n20985), .A2(\xmem_data[2][4] ), .B1(n20579), .B2(
        \xmem_data[3][4] ), .ZN(n4487) );
  AOI22_X1 U7741 ( .A1(n24607), .A2(\xmem_data[4][4] ), .B1(n20578), .B2(
        \xmem_data[5][4] ), .ZN(n4486) );
  AOI22_X1 U7742 ( .A1(n3449), .A2(\xmem_data[6][4] ), .B1(n25360), .B2(
        \xmem_data[7][4] ), .ZN(n4485) );
  NAND4_X1 U7743 ( .A1(n4488), .A2(n4487), .A3(n4486), .A4(n4485), .ZN(n4496)
         );
  AOI22_X1 U7744 ( .A1(n30949), .A2(\xmem_data[24][4] ), .B1(n25398), .B2(
        \xmem_data[25][4] ), .ZN(n4493) );
  AOI22_X1 U7745 ( .A1(n30309), .A2(\xmem_data[26][4] ), .B1(n13452), .B2(
        \xmem_data[27][4] ), .ZN(n4492) );
  BUF_X1 U7746 ( .A(n14881), .Z(n27974) );
  AOI22_X1 U7747 ( .A1(n27974), .A2(\xmem_data[28][4] ), .B1(n20816), .B2(
        \xmem_data[29][4] ), .ZN(n4491) );
  BUF_X1 U7748 ( .A(n14974), .Z(n27976) );
  BUF_X1 U7749 ( .A(n14883), .Z(n27975) );
  AOI22_X1 U7750 ( .A1(n3330), .A2(\xmem_data[30][4] ), .B1(n27975), .B2(
        \xmem_data[31][4] ), .ZN(n4490) );
  NAND4_X1 U7751 ( .A1(n4493), .A2(n4492), .A3(n4491), .A4(n4490), .ZN(n4494)
         );
  INV_X1 U7752 ( .A(n39041), .ZN(n37191) );
  NAND2_X1 U7753 ( .A1(n8414), .A2(n4497), .ZN(n4500) );
  INV_X1 U7754 ( .A(n4500), .ZN(n4498) );
  AOI22_X1 U7755 ( .A1(n37191), .A2(n4500), .B1(n4498), .B2(n4499), .ZN(n4571)
         );
  INV_X1 U7756 ( .A(load_xaddr_val[5]), .ZN(n4499) );
  NAND2_X1 U7757 ( .A1(load_xaddr_val[5]), .A2(n4500), .ZN(n4501) );
  XOR2_X1 U7758 ( .A(n39040), .B(n4501), .Z(n4525) );
  NOR2_X1 U7759 ( .A1(n4571), .A2(n4525), .ZN(n25287) );
  INV_X1 U7760 ( .A(n25287), .ZN(n24043) );
  AOI22_X1 U7761 ( .A1(n3171), .A2(\xmem_data[96][4] ), .B1(n25406), .B2(
        \xmem_data[97][4] ), .ZN(n4507) );
  BUF_X1 U7762 ( .A(n13127), .Z(n28036) );
  BUF_X1 U7763 ( .A(n13457), .Z(n28035) );
  AOI22_X1 U7764 ( .A1(n28036), .A2(\xmem_data[98][4] ), .B1(n28035), .B2(
        \xmem_data[99][4] ), .ZN(n4506) );
  BUF_X1 U7765 ( .A(n31263), .Z(n28038) );
  AOI22_X1 U7766 ( .A1(n28038), .A2(\xmem_data[100][4] ), .B1(n28037), .B2(
        \xmem_data[101][4] ), .ZN(n4505) );
  BUF_X1 U7767 ( .A(n28973), .Z(n28039) );
  AOI22_X1 U7768 ( .A1(n28039), .A2(\xmem_data[102][4] ), .B1(n28501), .B2(
        \xmem_data[103][4] ), .ZN(n4504) );
  NAND4_X1 U7769 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(n4524)
         );
  BUF_X1 U7770 ( .A(n29064), .Z(n28044) );
  AOI22_X1 U7771 ( .A1(n28044), .A2(\xmem_data[104][4] ), .B1(n3221), .B2(
        \xmem_data[105][4] ), .ZN(n4511) );
  AOI22_X1 U7772 ( .A1(n27831), .A2(\xmem_data[106][4] ), .B1(n25562), .B2(
        \xmem_data[107][4] ), .ZN(n4510) );
  AOI22_X1 U7773 ( .A1(n24697), .A2(\xmem_data[108][4] ), .B1(n27994), .B2(
        \xmem_data[109][4] ), .ZN(n4509) );
  AOI22_X1 U7774 ( .A1(n30710), .A2(\xmem_data[110][4] ), .B1(n30877), .B2(
        \xmem_data[111][4] ), .ZN(n4508) );
  NAND4_X1 U7775 ( .A1(n4511), .A2(n4510), .A3(n4509), .A4(n4508), .ZN(n4523)
         );
  BUF_X1 U7776 ( .A(n4478), .Z(n28050) );
  AOI22_X1 U7777 ( .A1(n28050), .A2(\xmem_data[112][4] ), .B1(n3358), .B2(
        \xmem_data[113][4] ), .ZN(n4515) );
  BUF_X1 U7778 ( .A(n14997), .Z(n28051) );
  AOI22_X1 U7779 ( .A1(n28051), .A2(\xmem_data[114][4] ), .B1(n28515), .B2(
        \xmem_data[115][4] ), .ZN(n4514) );
  BUF_X1 U7780 ( .A(n14935), .Z(n28052) );
  AOI22_X1 U7781 ( .A1(n16986), .A2(\xmem_data[116][4] ), .B1(n28052), .B2(
        \xmem_data[117][4] ), .ZN(n4513) );
  BUF_X1 U7782 ( .A(n29187), .Z(n28053) );
  AOI22_X1 U7783 ( .A1(n21048), .A2(\xmem_data[118][4] ), .B1(n27989), .B2(
        \xmem_data[119][4] ), .ZN(n4512) );
  NAND4_X1 U7784 ( .A1(n4515), .A2(n4514), .A3(n4513), .A4(n4512), .ZN(n4522)
         );
  BUF_X1 U7785 ( .A(n14937), .Z(n28059) );
  BUF_X1 U7786 ( .A(n13415), .Z(n28058) );
  AOI22_X1 U7787 ( .A1(n28059), .A2(\xmem_data[120][4] ), .B1(n28058), .B2(
        \xmem_data[121][4] ), .ZN(n4520) );
  AOI22_X1 U7788 ( .A1(n23777), .A2(\xmem_data[122][4] ), .B1(n29280), .B2(
        \xmem_data[123][4] ), .ZN(n4519) );
  BUF_X1 U7789 ( .A(n4158), .Z(n28061) );
  BUF_X1 U7790 ( .A(n14973), .Z(n28060) );
  AOI22_X1 U7791 ( .A1(n28061), .A2(\xmem_data[124][4] ), .B1(n28060), .B2(
        \xmem_data[125][4] ), .ZN(n4518) );
  BUF_X1 U7792 ( .A(n14883), .Z(n28062) );
  AOI22_X1 U7793 ( .A1(n3338), .A2(\xmem_data[126][4] ), .B1(n28062), .B2(
        \xmem_data[127][4] ), .ZN(n4517) );
  NAND4_X1 U7794 ( .A1(n4520), .A2(n4519), .A3(n4518), .A4(n4517), .ZN(n4521)
         );
  OR4_X1 U7795 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), .ZN(n4550) );
  INV_X1 U7796 ( .A(n4525), .ZN(n4572) );
  NOR2_X1 U7797 ( .A1(n4571), .A2(n4572), .ZN(n28033) );
  AOI22_X1 U7798 ( .A1(n27847), .A2(\xmem_data[64][4] ), .B1(n20488), .B2(
        \xmem_data[65][4] ), .ZN(n4531) );
  AOI22_X1 U7799 ( .A1(n30901), .A2(\xmem_data[66][4] ), .B1(n27567), .B2(
        \xmem_data[67][4] ), .ZN(n4530) );
  BUF_X1 U7800 ( .A(n31263), .Z(n28076) );
  BUF_X1 U7801 ( .A(n28974), .Z(n28075) );
  AOI22_X1 U7802 ( .A1(n28076), .A2(\xmem_data[68][4] ), .B1(n28075), .B2(
        \xmem_data[69][4] ), .ZN(n4529) );
  AOI22_X1 U7803 ( .A1(n3434), .A2(\xmem_data[70][4] ), .B1(n3247), .B2(
        \xmem_data[71][4] ), .ZN(n4528) );
  NAND4_X1 U7804 ( .A1(n4531), .A2(n4530), .A3(n4529), .A4(n4528), .ZN(n4548)
         );
  BUF_X1 U7805 ( .A(n29064), .Z(n28082) );
  AOI22_X1 U7806 ( .A1(n28082), .A2(\xmem_data[72][4] ), .B1(n3217), .B2(
        \xmem_data[73][4] ), .ZN(n4535) );
  AOI22_X1 U7807 ( .A1(n29431), .A2(\xmem_data[74][4] ), .B1(n23739), .B2(
        \xmem_data[75][4] ), .ZN(n4534) );
  BUF_X1 U7808 ( .A(n14926), .Z(n28083) );
  AOI22_X1 U7809 ( .A1(n28083), .A2(\xmem_data[76][4] ), .B1(n13444), .B2(
        \xmem_data[77][4] ), .ZN(n4533) );
  BUF_X1 U7810 ( .A(n14991), .Z(n28084) );
  AOI22_X1 U7811 ( .A1(n28084), .A2(\xmem_data[78][4] ), .B1(n28045), .B2(
        \xmem_data[79][4] ), .ZN(n4532) );
  NAND4_X1 U7812 ( .A1(n4535), .A2(n4534), .A3(n4533), .A4(n4532), .ZN(n4547)
         );
  AOI22_X1 U7813 ( .A1(n27551), .A2(\xmem_data[80][4] ), .B1(n13475), .B2(
        \xmem_data[81][4] ), .ZN(n4540) );
  BUF_X1 U7814 ( .A(n14997), .Z(n28089) );
  AOI22_X1 U7815 ( .A1(n28089), .A2(\xmem_data[82][4] ), .B1(n24159), .B2(
        \xmem_data[83][4] ), .ZN(n4539) );
  BUF_X1 U7816 ( .A(n14935), .Z(n28090) );
  AOI22_X1 U7817 ( .A1(n30614), .A2(\xmem_data[84][4] ), .B1(n28090), .B2(
        \xmem_data[85][4] ), .ZN(n4538) );
  BUF_X1 U7818 ( .A(n29187), .Z(n28091) );
  AOI22_X1 U7819 ( .A1(n3120), .A2(\xmem_data[86][4] ), .B1(n28299), .B2(
        \xmem_data[87][4] ), .ZN(n4537) );
  NAND4_X1 U7820 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4546)
         );
  BUF_X1 U7821 ( .A(n14937), .Z(n28096) );
  AOI22_X1 U7822 ( .A1(n28096), .A2(\xmem_data[88][4] ), .B1(n31270), .B2(
        \xmem_data[89][4] ), .ZN(n4544) );
  BUF_X1 U7823 ( .A(n13452), .Z(n28097) );
  AOI22_X1 U7824 ( .A1(n23802), .A2(\xmem_data[90][4] ), .B1(n28097), .B2(
        \xmem_data[91][4] ), .ZN(n4543) );
  AOI22_X1 U7825 ( .A1(n24647), .A2(\xmem_data[92][4] ), .B1(n27951), .B2(
        \xmem_data[93][4] ), .ZN(n4542) );
  AOI22_X1 U7826 ( .A1(n28461), .A2(\xmem_data[94][4] ), .B1(n28098), .B2(
        \xmem_data[95][4] ), .ZN(n4541) );
  NAND4_X1 U7827 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  OR4_X1 U7828 ( .A1(n4548), .A2(n4547), .A3(n4546), .A4(n4545), .ZN(n4549) );
  AOI22_X1 U7829 ( .A1(n28071), .A2(n4550), .B1(n28033), .B2(n4549), .ZN(n4575) );
  AOI22_X1 U7830 ( .A1(n3171), .A2(\xmem_data[32][4] ), .B1(n25527), .B2(
        \xmem_data[33][4] ), .ZN(n4554) );
  AOI22_X1 U7831 ( .A1(n20952), .A2(\xmem_data[34][4] ), .B1(n31344), .B2(
        \xmem_data[35][4] ), .ZN(n4553) );
  AOI22_X1 U7832 ( .A1(n28076), .A2(\xmem_data[36][4] ), .B1(n28075), .B2(
        \xmem_data[37][4] ), .ZN(n4552) );
  AOI22_X1 U7833 ( .A1(n3434), .A2(\xmem_data[38][4] ), .B1(n3247), .B2(
        \xmem_data[39][4] ), .ZN(n4551) );
  NAND4_X1 U7834 ( .A1(n4554), .A2(n4553), .A3(n4552), .A4(n4551), .ZN(n4570)
         );
  AOI22_X1 U7835 ( .A1(n28082), .A2(\xmem_data[40][4] ), .B1(n3221), .B2(
        \xmem_data[41][4] ), .ZN(n4558) );
  AOI22_X1 U7836 ( .A1(n25448), .A2(\xmem_data[42][4] ), .B1(n20787), .B2(
        \xmem_data[43][4] ), .ZN(n4557) );
  AOI22_X1 U7837 ( .A1(n28083), .A2(\xmem_data[44][4] ), .B1(n24633), .B2(
        \xmem_data[45][4] ), .ZN(n4556) );
  AOI22_X1 U7838 ( .A1(n28084), .A2(\xmem_data[46][4] ), .B1(n31252), .B2(
        \xmem_data[47][4] ), .ZN(n4555) );
  NAND4_X1 U7839 ( .A1(n4558), .A2(n4557), .A3(n4556), .A4(n4555), .ZN(n4569)
         );
  AOI22_X1 U7840 ( .A1(n27551), .A2(\xmem_data[48][4] ), .B1(n13475), .B2(
        \xmem_data[49][4] ), .ZN(n4562) );
  AOI22_X1 U7841 ( .A1(n28089), .A2(\xmem_data[50][4] ), .B1(n17012), .B2(
        \xmem_data[51][4] ), .ZN(n4561) );
  AOI22_X1 U7842 ( .A1(n3175), .A2(\xmem_data[52][4] ), .B1(n28090), .B2(
        \xmem_data[53][4] ), .ZN(n4560) );
  AOI22_X1 U7843 ( .A1(n24545), .A2(\xmem_data[54][4] ), .B1(n20543), .B2(
        \xmem_data[55][4] ), .ZN(n4559) );
  NAND4_X1 U7844 ( .A1(n4562), .A2(n4561), .A3(n4560), .A4(n4559), .ZN(n4568)
         );
  AOI22_X1 U7845 ( .A1(n28096), .A2(\xmem_data[56][4] ), .B1(n28058), .B2(
        \xmem_data[57][4] ), .ZN(n4566) );
  AOI22_X1 U7846 ( .A1(n22682), .A2(\xmem_data[58][4] ), .B1(n28097), .B2(
        \xmem_data[59][4] ), .ZN(n4565) );
  AOI22_X1 U7847 ( .A1(n24647), .A2(\xmem_data[60][4] ), .B1(n25716), .B2(
        \xmem_data[61][4] ), .ZN(n4564) );
  AOI22_X1 U7848 ( .A1(n20817), .A2(\xmem_data[62][4] ), .B1(n28098), .B2(
        \xmem_data[63][4] ), .ZN(n4563) );
  NAND4_X1 U7849 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4567)
         );
  OR4_X1 U7850 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4573) );
  AND2_X1 U7851 ( .A1(n4572), .A2(n4571), .ZN(n28107) );
  XNOR2_X1 U7852 ( .A(n31161), .B(\fmem_data[22][7] ), .ZN(n31665) );
  XOR2_X1 U7853 ( .A(\fmem_data[22][6] ), .B(\fmem_data[22][7] ), .Z(n4577) );
  AOI22_X1 U7854 ( .A1(n3209), .A2(\xmem_data[96][3] ), .B1(n21057), .B2(
        \xmem_data[97][3] ), .ZN(n4581) );
  AOI22_X1 U7855 ( .A1(n28036), .A2(\xmem_data[98][3] ), .B1(n28035), .B2(
        \xmem_data[99][3] ), .ZN(n4580) );
  AOI22_X1 U7856 ( .A1(n28038), .A2(\xmem_data[100][3] ), .B1(n28037), .B2(
        \xmem_data[101][3] ), .ZN(n4579) );
  AOI22_X1 U7857 ( .A1(n28039), .A2(\xmem_data[102][3] ), .B1(n20568), .B2(
        \xmem_data[103][3] ), .ZN(n4578) );
  NAND4_X1 U7858 ( .A1(n4581), .A2(n4580), .A3(n4579), .A4(n4578), .ZN(n4597)
         );
  AOI22_X1 U7859 ( .A1(n28044), .A2(\xmem_data[104][3] ), .B1(n3218), .B2(
        \xmem_data[105][3] ), .ZN(n4585) );
  AOI22_X1 U7860 ( .A1(n25448), .A2(\xmem_data[106][3] ), .B1(n22710), .B2(
        \xmem_data[107][3] ), .ZN(n4584) );
  AOI22_X1 U7861 ( .A1(n22666), .A2(\xmem_data[108][3] ), .B1(n22669), .B2(
        \xmem_data[109][3] ), .ZN(n4583) );
  AOI22_X1 U7862 ( .A1(n28084), .A2(\xmem_data[110][3] ), .B1(n28343), .B2(
        \xmem_data[111][3] ), .ZN(n4582) );
  NAND4_X1 U7863 ( .A1(n4585), .A2(n4584), .A3(n4583), .A4(n4582), .ZN(n4596)
         );
  AOI22_X1 U7864 ( .A1(n28050), .A2(\xmem_data[112][3] ), .B1(n25481), .B2(
        \xmem_data[113][3] ), .ZN(n4589) );
  AOI22_X1 U7865 ( .A1(n28051), .A2(\xmem_data[114][3] ), .B1(n24132), .B2(
        \xmem_data[115][3] ), .ZN(n4588) );
  AOI22_X1 U7866 ( .A1(n30614), .A2(\xmem_data[116][3] ), .B1(n28052), .B2(
        \xmem_data[117][3] ), .ZN(n4587) );
  AOI22_X1 U7867 ( .A1(n25607), .A2(\xmem_data[118][3] ), .B1(n3208), .B2(
        \xmem_data[119][3] ), .ZN(n4586) );
  NAND4_X1 U7868 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4595)
         );
  AOI22_X1 U7869 ( .A1(n28059), .A2(\xmem_data[120][3] ), .B1(n28058), .B2(
        \xmem_data[121][3] ), .ZN(n4593) );
  AOI22_X1 U7870 ( .A1(n28994), .A2(\xmem_data[122][3] ), .B1(n25435), .B2(
        \xmem_data[123][3] ), .ZN(n4592) );
  AOI22_X1 U7871 ( .A1(n28061), .A2(\xmem_data[124][3] ), .B1(n28060), .B2(
        \xmem_data[125][3] ), .ZN(n4591) );
  AOI22_X1 U7872 ( .A1(n25718), .A2(\xmem_data[126][3] ), .B1(n28062), .B2(
        \xmem_data[127][3] ), .ZN(n4590) );
  NAND4_X1 U7873 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4594)
         );
  OR4_X1 U7874 ( .A1(n4597), .A2(n4596), .A3(n4595), .A4(n4594), .ZN(n4619) );
  AOI22_X1 U7875 ( .A1(n20782), .A2(\xmem_data[64][3] ), .B1(n29017), .B2(
        \xmem_data[65][3] ), .ZN(n4601) );
  AOI22_X1 U7876 ( .A1(n28036), .A2(\xmem_data[66][3] ), .B1(n28035), .B2(
        \xmem_data[67][3] ), .ZN(n4600) );
  AOI22_X1 U7877 ( .A1(n28038), .A2(\xmem_data[68][3] ), .B1(n28037), .B2(
        \xmem_data[69][3] ), .ZN(n4599) );
  AOI22_X1 U7878 ( .A1(n28039), .A2(\xmem_data[70][3] ), .B1(n24439), .B2(
        \xmem_data[71][3] ), .ZN(n4598) );
  NAND4_X1 U7879 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4617)
         );
  AOI22_X1 U7880 ( .A1(n28044), .A2(\xmem_data[72][3] ), .B1(n3218), .B2(
        \xmem_data[73][3] ), .ZN(n4605) );
  AOI22_X1 U7881 ( .A1(n22708), .A2(\xmem_data[74][3] ), .B1(n23769), .B2(
        \xmem_data[75][3] ), .ZN(n4604) );
  AOI22_X1 U7882 ( .A1(n24697), .A2(\xmem_data[76][3] ), .B1(n22711), .B2(
        \xmem_data[77][3] ), .ZN(n4603) );
  AOI22_X1 U7883 ( .A1(n28308), .A2(\xmem_data[78][3] ), .B1(n23771), .B2(
        \xmem_data[79][3] ), .ZN(n4602) );
  NAND4_X1 U7884 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4616)
         );
  AOI22_X1 U7885 ( .A1(n28050), .A2(\xmem_data[80][3] ), .B1(n3358), .B2(
        \xmem_data[81][3] ), .ZN(n4609) );
  AOI22_X1 U7886 ( .A1(n28051), .A2(\xmem_data[82][3] ), .B1(n22702), .B2(
        \xmem_data[83][3] ), .ZN(n4608) );
  AOI22_X1 U7887 ( .A1(n24131), .A2(\xmem_data[84][3] ), .B1(n28052), .B2(
        \xmem_data[85][3] ), .ZN(n4607) );
  AOI22_X1 U7888 ( .A1(n16988), .A2(\xmem_data[86][3] ), .B1(n22742), .B2(
        \xmem_data[87][3] ), .ZN(n4606) );
  NAND4_X1 U7889 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4615)
         );
  AOI22_X1 U7890 ( .A1(n28059), .A2(\xmem_data[88][3] ), .B1(n28058), .B2(
        \xmem_data[89][3] ), .ZN(n4613) );
  AOI22_X1 U7891 ( .A1(n27825), .A2(\xmem_data[90][3] ), .B1(n31360), .B2(
        \xmem_data[91][3] ), .ZN(n4612) );
  AOI22_X1 U7892 ( .A1(n28061), .A2(\xmem_data[92][3] ), .B1(n28060), .B2(
        \xmem_data[93][3] ), .ZN(n4611) );
  AOI22_X1 U7893 ( .A1(n20732), .A2(\xmem_data[94][3] ), .B1(n28062), .B2(
        \xmem_data[95][3] ), .ZN(n4610) );
  NAND4_X1 U7894 ( .A1(n4613), .A2(n4612), .A3(n4611), .A4(n4610), .ZN(n4614)
         );
  OR4_X1 U7895 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4618) );
  AOI22_X1 U7896 ( .A1(n28071), .A2(n4619), .B1(n28033), .B2(n4618), .ZN(n4671) );
  AOI22_X1 U7897 ( .A1(n13486), .A2(\xmem_data[0][3] ), .B1(n27981), .B2(
        \xmem_data[1][3] ), .ZN(n4623) );
  AOI22_X1 U7898 ( .A1(n20577), .A2(\xmem_data[2][3] ), .B1(n24624), .B2(
        \xmem_data[3][3] ), .ZN(n4622) );
  AOI22_X1 U7899 ( .A1(n25724), .A2(\xmem_data[4][3] ), .B1(n29118), .B2(
        \xmem_data[5][3] ), .ZN(n4621) );
  AOI22_X1 U7900 ( .A1(n3449), .A2(\xmem_data[6][3] ), .B1(n24172), .B2(
        \xmem_data[7][3] ), .ZN(n4620) );
  NAND4_X1 U7901 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4629)
         );
  AOI22_X1 U7902 ( .A1(n31330), .A2(\xmem_data[24][3] ), .B1(n14970), .B2(
        \xmem_data[25][3] ), .ZN(n4627) );
  AOI22_X1 U7903 ( .A1(n29439), .A2(\xmem_data[26][3] ), .B1(n24116), .B2(
        \xmem_data[27][3] ), .ZN(n4626) );
  AOI22_X1 U7904 ( .A1(n27974), .A2(\xmem_data[28][3] ), .B1(n20816), .B2(
        \xmem_data[29][3] ), .ZN(n4625) );
  AOI22_X1 U7905 ( .A1(n3329), .A2(\xmem_data[30][3] ), .B1(n27975), .B2(
        \xmem_data[31][3] ), .ZN(n4624) );
  NAND4_X1 U7906 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4628)
         );
  AOI22_X1 U7907 ( .A1(n27508), .A2(\xmem_data[16][3] ), .B1(n27988), .B2(
        \xmem_data[17][3] ), .ZN(n4633) );
  AOI22_X1 U7908 ( .A1(n17013), .A2(\xmem_data[18][3] ), .B1(n28416), .B2(
        \xmem_data[19][3] ), .ZN(n4632) );
  AOI22_X1 U7909 ( .A1(n10977), .A2(\xmem_data[20][3] ), .B1(n20717), .B2(
        \xmem_data[21][3] ), .ZN(n4631) );
  AOI22_X1 U7910 ( .A1(n25461), .A2(\xmem_data[22][3] ), .B1(n27989), .B2(
        \xmem_data[23][3] ), .ZN(n4630) );
  NAND4_X1 U7911 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4636)
         );
  AOI22_X1 U7912 ( .A1(n29789), .A2(\xmem_data[10][3] ), .B1(n28476), .B2(
        \xmem_data[11][3] ), .ZN(n4634) );
  AOI22_X1 U7913 ( .A1(n24532), .A2(\xmem_data[8][3] ), .B1(n3217), .B2(
        \xmem_data[9][3] ), .ZN(n4637) );
  INV_X1 U7914 ( .A(n4637), .ZN(n4641) );
  AOI22_X1 U7915 ( .A1(n23812), .A2(\xmem_data[12][3] ), .B1(n27994), .B2(
        \xmem_data[13][3] ), .ZN(n4639) );
  NAND2_X1 U7916 ( .A1(n3146), .A2(\xmem_data[14][3] ), .ZN(n4638) );
  NAND2_X1 U7917 ( .A1(n4639), .A2(n4638), .ZN(n4640) );
  NOR2_X1 U7918 ( .A1(n4641), .A2(n4640), .ZN(n4642) );
  NAND3_X1 U7919 ( .A1(n4644), .A2(n4643), .A3(n4642), .ZN(n4647) );
  NOR2_X1 U7920 ( .A1(n24043), .A2(n39021), .ZN(n4645) );
  AND2_X1 U7921 ( .A1(n28510), .A2(n4645), .ZN(n4646) );
  AOI22_X1 U7922 ( .A1(n25526), .A2(\xmem_data[32][3] ), .B1(n27526), .B2(
        \xmem_data[33][3] ), .ZN(n4651) );
  AOI22_X1 U7923 ( .A1(n30901), .A2(\xmem_data[34][3] ), .B1(n17050), .B2(
        \xmem_data[35][3] ), .ZN(n4650) );
  AOI22_X1 U7924 ( .A1(n28076), .A2(\xmem_data[36][3] ), .B1(n28075), .B2(
        \xmem_data[37][3] ), .ZN(n4649) );
  AOI22_X1 U7925 ( .A1(n3434), .A2(\xmem_data[38][3] ), .B1(n3247), .B2(
        \xmem_data[39][3] ), .ZN(n4648) );
  NAND4_X1 U7926 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n4667)
         );
  AOI22_X1 U7927 ( .A1(n28082), .A2(\xmem_data[40][3] ), .B1(n3218), .B2(
        \xmem_data[41][3] ), .ZN(n4655) );
  AOI22_X1 U7928 ( .A1(n21067), .A2(\xmem_data[42][3] ), .B1(n28508), .B2(
        \xmem_data[43][3] ), .ZN(n4654) );
  AOI22_X1 U7929 ( .A1(n28083), .A2(\xmem_data[44][3] ), .B1(n25486), .B2(
        \xmem_data[45][3] ), .ZN(n4653) );
  AOI22_X1 U7930 ( .A1(n28084), .A2(\xmem_data[46][3] ), .B1(n3231), .B2(
        \xmem_data[47][3] ), .ZN(n4652) );
  NAND4_X1 U7931 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4666)
         );
  AOI22_X1 U7932 ( .A1(n27551), .A2(\xmem_data[48][3] ), .B1(n13475), .B2(
        \xmem_data[49][3] ), .ZN(n4659) );
  AOI22_X1 U7933 ( .A1(n28089), .A2(\xmem_data[50][3] ), .B1(n27452), .B2(
        \xmem_data[51][3] ), .ZN(n4658) );
  AOI22_X1 U7934 ( .A1(n30891), .A2(\xmem_data[52][3] ), .B1(n28090), .B2(
        \xmem_data[53][3] ), .ZN(n4657) );
  AOI22_X1 U7935 ( .A1(n27755), .A2(\xmem_data[54][3] ), .B1(n31269), .B2(
        \xmem_data[55][3] ), .ZN(n4656) );
  NAND4_X1 U7936 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4665)
         );
  AOI22_X1 U7937 ( .A1(n28096), .A2(\xmem_data[56][3] ), .B1(n24707), .B2(
        \xmem_data[57][3] ), .ZN(n4663) );
  AOI22_X1 U7938 ( .A1(n30617), .A2(\xmem_data[58][3] ), .B1(n28097), .B2(
        \xmem_data[59][3] ), .ZN(n4662) );
  AOI22_X1 U7939 ( .A1(n28493), .A2(\xmem_data[60][3] ), .B1(n25581), .B2(
        \xmem_data[61][3] ), .ZN(n4661) );
  AOI22_X1 U7940 ( .A1(n24522), .A2(\xmem_data[62][3] ), .B1(n28098), .B2(
        \xmem_data[63][3] ), .ZN(n4660) );
  NAND4_X1 U7941 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4664)
         );
  OR4_X1 U7942 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4668) );
  NAND2_X1 U7943 ( .A1(n4668), .A2(n28107), .ZN(n4669) );
  XNOR2_X1 U7944 ( .A(n31992), .B(\fmem_data[22][7] ), .ZN(n24111) );
  OAI22_X1 U7945 ( .A1(n31665), .A2(n35585), .B1(n35584), .B2(n24111), .ZN(
        n33343) );
  AOI22_X1 U7946 ( .A1(n30891), .A2(\xmem_data[4][3] ), .B1(n25606), .B2(
        \xmem_data[5][3] ), .ZN(n4673) );
  AOI22_X1 U7947 ( .A1(n25632), .A2(\xmem_data[12][3] ), .B1(n31361), .B2(
        \xmem_data[13][3] ), .ZN(n4672) );
  AOI22_X1 U7948 ( .A1(n25630), .A2(\xmem_data[20][3] ), .B1(n25629), .B2(
        \xmem_data[21][3] ), .ZN(n4680) );
  AOI22_X1 U7949 ( .A1(n25628), .A2(\xmem_data[18][3] ), .B1(n24122), .B2(
        \xmem_data[19][3] ), .ZN(n4679) );
  AOI22_X1 U7950 ( .A1(n24606), .A2(\xmem_data[16][3] ), .B1(n17049), .B2(
        \xmem_data[17][3] ), .ZN(n4674) );
  INV_X1 U7951 ( .A(n4674), .ZN(n4677) );
  AOI22_X1 U7952 ( .A1(n25624), .A2(\xmem_data[22][3] ), .B1(n22753), .B2(
        \xmem_data[23][3] ), .ZN(n4675) );
  INV_X1 U7953 ( .A(n4675), .ZN(n4676) );
  NOR2_X1 U7954 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  NAND4_X1 U7955 ( .A1(n3938), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4701)
         );
  AOI22_X1 U7956 ( .A1(n25636), .A2(\xmem_data[14][3] ), .B1(n20507), .B2(
        \xmem_data[15][3] ), .ZN(n4682) );
  AOI22_X1 U7957 ( .A1(n27818), .A2(\xmem_data[6][3] ), .B1(n22742), .B2(
        \xmem_data[7][3] ), .ZN(n4681) );
  AOI22_X1 U7958 ( .A1(n29410), .A2(\xmem_data[10][3] ), .B1(n25367), .B2(
        \xmem_data[11][3] ), .ZN(n4683) );
  NAND2_X1 U7959 ( .A1(n4005), .A2(n4683), .ZN(n4687) );
  NAND2_X1 U7960 ( .A1(n30884), .A2(\xmem_data[1][3] ), .ZN(n4685) );
  NAND2_X1 U7961 ( .A1(n25604), .A2(\xmem_data[0][3] ), .ZN(n4684) );
  NAND2_X1 U7962 ( .A1(n4685), .A2(n4684), .ZN(n4686) );
  NOR2_X1 U7963 ( .A1(n4687), .A2(n4686), .ZN(n4690) );
  AOI22_X1 U7964 ( .A1(n28233), .A2(\xmem_data[2][3] ), .B1(n25605), .B2(
        \xmem_data[3][3] ), .ZN(n4689) );
  AOI22_X1 U7965 ( .A1(n25635), .A2(\xmem_data[8][3] ), .B1(n28492), .B2(
        \xmem_data[9][3] ), .ZN(n4688) );
  NAND4_X1 U7966 ( .A1(n3553), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4699)
         );
  AOI22_X1 U7967 ( .A1(n30503), .A2(\xmem_data[24][3] ), .B1(n3218), .B2(
        \xmem_data[25][3] ), .ZN(n4697) );
  AOI22_X1 U7968 ( .A1(n25617), .A2(\xmem_data[28][3] ), .B1(n25616), .B2(
        \xmem_data[29][3] ), .ZN(n4691) );
  INV_X1 U7969 ( .A(n4691), .ZN(n4695) );
  AOI22_X1 U7970 ( .A1(n25612), .A2(\xmem_data[26][3] ), .B1(n28476), .B2(
        \xmem_data[27][3] ), .ZN(n4693) );
  NAND2_X1 U7971 ( .A1(n3281), .A2(\xmem_data[30][3] ), .ZN(n4692) );
  NAND2_X1 U7972 ( .A1(n4693), .A2(n4692), .ZN(n4694) );
  NOR2_X1 U7973 ( .A1(n4695), .A2(n4694), .ZN(n4696) );
  NAND2_X1 U7974 ( .A1(n4697), .A2(n4696), .ZN(n4698) );
  OR2_X1 U7975 ( .A1(n4699), .A2(n4698), .ZN(n4700) );
  OAI21_X1 U7976 ( .B1(n4701), .B2(n4700), .A(n19018), .ZN(n4702) );
  INV_X1 U7977 ( .A(n4702), .ZN(n4771) );
  AOI22_X1 U7978 ( .A1(n25707), .A2(\xmem_data[32][3] ), .B1(n25456), .B2(
        \xmem_data[33][3] ), .ZN(n4706) );
  AOI22_X1 U7979 ( .A1(n25708), .A2(\xmem_data[34][3] ), .B1(n23761), .B2(
        \xmem_data[35][3] ), .ZN(n4705) );
  AOI22_X1 U7980 ( .A1(n30891), .A2(\xmem_data[36][3] ), .B1(n25709), .B2(
        \xmem_data[37][3] ), .ZN(n4704) );
  AOI22_X1 U7981 ( .A1(n27517), .A2(\xmem_data[38][3] ), .B1(n3213), .B2(
        \xmem_data[39][3] ), .ZN(n4703) );
  NAND4_X1 U7982 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4722)
         );
  AOI22_X1 U7983 ( .A1(n25573), .A2(\xmem_data[40][3] ), .B1(n25715), .B2(
        \xmem_data[41][3] ), .ZN(n4710) );
  AOI22_X1 U7984 ( .A1(n30872), .A2(\xmem_data[42][3] ), .B1(n30871), .B2(
        \xmem_data[43][3] ), .ZN(n4709) );
  AOI22_X1 U7985 ( .A1(n24548), .A2(\xmem_data[44][3] ), .B1(n29281), .B2(
        \xmem_data[45][3] ), .ZN(n4708) );
  AOI22_X1 U7986 ( .A1(n25718), .A2(\xmem_data[46][3] ), .B1(n30599), .B2(
        \xmem_data[47][3] ), .ZN(n4707) );
  NAND4_X1 U7987 ( .A1(n4710), .A2(n4709), .A3(n4708), .A4(n4707), .ZN(n4721)
         );
  AOI22_X1 U7988 ( .A1(n3179), .A2(\xmem_data[48][3] ), .B1(n25723), .B2(
        \xmem_data[49][3] ), .ZN(n4714) );
  AOI22_X1 U7989 ( .A1(n24687), .A2(\xmem_data[50][3] ), .B1(n24468), .B2(
        \xmem_data[51][3] ), .ZN(n4713) );
  AOI22_X1 U7990 ( .A1(n25724), .A2(\xmem_data[52][3] ), .B1(n29118), .B2(
        \xmem_data[53][3] ), .ZN(n4712) );
  AOI22_X1 U7991 ( .A1(n25725), .A2(\xmem_data[54][3] ), .B1(n30863), .B2(
        \xmem_data[55][3] ), .ZN(n4711) );
  NAND4_X1 U7992 ( .A1(n4714), .A2(n4713), .A3(n4712), .A4(n4711), .ZN(n4720)
         );
  AOI22_X1 U7993 ( .A1(n25730), .A2(\xmem_data[56][3] ), .B1(n3218), .B2(
        \xmem_data[57][3] ), .ZN(n4718) );
  AOI22_X1 U7994 ( .A1(n25731), .A2(\xmem_data[58][3] ), .B1(n25509), .B2(
        \xmem_data[59][3] ), .ZN(n4717) );
  AOI22_X1 U7995 ( .A1(n29027), .A2(\xmem_data[60][3] ), .B1(n27903), .B2(
        \xmem_data[61][3] ), .ZN(n4716) );
  AOI22_X1 U7996 ( .A1(n25732), .A2(\xmem_data[62][3] ), .B1(n23771), .B2(
        \xmem_data[63][3] ), .ZN(n4715) );
  NAND4_X1 U7997 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4719)
         );
  OR4_X1 U7998 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4723) );
  AND2_X1 U7999 ( .A1(n4723), .A2(n25741), .ZN(n4770) );
  AOI22_X1 U8000 ( .A1(n25670), .A2(\xmem_data[64][3] ), .B1(n30884), .B2(
        \xmem_data[65][3] ), .ZN(n4727) );
  AOI22_X1 U8001 ( .A1(n30744), .A2(\xmem_data[66][3] ), .B1(n27513), .B2(
        \xmem_data[67][3] ), .ZN(n4726) );
  AOI22_X1 U8002 ( .A1(n17041), .A2(\xmem_data[68][3] ), .B1(n25671), .B2(
        \xmem_data[69][3] ), .ZN(n4725) );
  AOI22_X1 U8003 ( .A1(n25672), .A2(\xmem_data[70][3] ), .B1(n3213), .B2(
        \xmem_data[71][3] ), .ZN(n4724) );
  NAND4_X1 U8004 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4744)
         );
  AOI22_X1 U8005 ( .A1(n23717), .A2(\xmem_data[72][3] ), .B1(n25677), .B2(
        \xmem_data[73][3] ), .ZN(n4731) );
  AOI22_X1 U8006 ( .A1(n25678), .A2(\xmem_data[74][3] ), .B1(n24165), .B2(
        \xmem_data[75][3] ), .ZN(n4730) );
  AOI22_X1 U8007 ( .A1(n29100), .A2(\xmem_data[76][3] ), .B1(n28429), .B2(
        \xmem_data[77][3] ), .ZN(n4729) );
  AOI22_X1 U8008 ( .A1(n3307), .A2(\xmem_data[78][3] ), .B1(n24622), .B2(
        \xmem_data[79][3] ), .ZN(n4728) );
  NAND4_X1 U8009 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4743)
         );
  AOI22_X1 U8010 ( .A1(n3209), .A2(\xmem_data[80][3] ), .B1(n25723), .B2(
        \xmem_data[81][3] ), .ZN(n4735) );
  AOI22_X1 U8011 ( .A1(n25684), .A2(\xmem_data[82][3] ), .B1(n24122), .B2(
        \xmem_data[83][3] ), .ZN(n4734) );
  AOI22_X1 U8012 ( .A1(n25686), .A2(\xmem_data[84][3] ), .B1(n25685), .B2(
        \xmem_data[85][3] ), .ZN(n4733) );
  AOI22_X1 U8013 ( .A1(n21308), .A2(\xmem_data[86][3] ), .B1(n25687), .B2(
        \xmem_data[87][3] ), .ZN(n4732) );
  NAND4_X1 U8014 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4742)
         );
  AND2_X1 U8015 ( .A1(n3218), .A2(\xmem_data[89][3] ), .ZN(n4736) );
  AOI21_X1 U8016 ( .B1(n25692), .B2(\xmem_data[88][3] ), .A(n4736), .ZN(n4740)
         );
  AOI22_X1 U8017 ( .A1(n25693), .A2(\xmem_data[90][3] ), .B1(n20500), .B2(
        \xmem_data[91][3] ), .ZN(n4739) );
  AOI22_X1 U8018 ( .A1(n25694), .A2(\xmem_data[92][3] ), .B1(n13444), .B2(
        \xmem_data[93][3] ), .ZN(n4738) );
  AOI22_X1 U8019 ( .A1(n3374), .A2(\xmem_data[94][3] ), .B1(n28343), .B2(
        \xmem_data[95][3] ), .ZN(n4737) );
  NAND4_X1 U8020 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4741)
         );
  OR4_X1 U8021 ( .A1(n4744), .A2(n4743), .A3(n4742), .A4(n4741), .ZN(n4745) );
  NAND2_X1 U8022 ( .A1(n4745), .A2(n25704), .ZN(n4768) );
  AOI22_X1 U8023 ( .A1(n25670), .A2(\xmem_data[96][3] ), .B1(n27863), .B2(
        \xmem_data[97][3] ), .ZN(n4749) );
  AOI22_X1 U8024 ( .A1(n27911), .A2(\xmem_data[98][3] ), .B1(n17012), .B2(
        \xmem_data[99][3] ), .ZN(n4748) );
  AOI22_X1 U8025 ( .A1(n27537), .A2(\xmem_data[100][3] ), .B1(n25671), .B2(
        \xmem_data[101][3] ), .ZN(n4747) );
  AOI22_X1 U8026 ( .A1(n25672), .A2(\xmem_data[102][3] ), .B1(n3208), .B2(
        \xmem_data[103][3] ), .ZN(n4746) );
  NAND4_X1 U8027 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4765)
         );
  AOI22_X1 U8028 ( .A1(n20542), .A2(\xmem_data[104][3] ), .B1(n25677), .B2(
        \xmem_data[105][3] ), .ZN(n4753) );
  AOI22_X1 U8029 ( .A1(n25678), .A2(\xmem_data[106][3] ), .B1(n23801), .B2(
        \xmem_data[107][3] ), .ZN(n4752) );
  AOI22_X1 U8030 ( .A1(n28428), .A2(\xmem_data[108][3] ), .B1(n29281), .B2(
        \xmem_data[109][3] ), .ZN(n4751) );
  AOI22_X1 U8031 ( .A1(n3269), .A2(\xmem_data[110][3] ), .B1(n14975), .B2(
        \xmem_data[111][3] ), .ZN(n4750) );
  NAND4_X1 U8032 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4764)
         );
  AOI22_X1 U8033 ( .A1(n24166), .A2(\xmem_data[112][3] ), .B1(n23725), .B2(
        \xmem_data[113][3] ), .ZN(n4757) );
  AOI22_X1 U8034 ( .A1(n25684), .A2(\xmem_data[114][3] ), .B1(n25440), .B2(
        \xmem_data[115][3] ), .ZN(n4756) );
  AOI22_X1 U8035 ( .A1(n25686), .A2(\xmem_data[116][3] ), .B1(n25685), .B2(
        \xmem_data[117][3] ), .ZN(n4755) );
  AOI22_X1 U8036 ( .A1(n3387), .A2(\xmem_data[118][3] ), .B1(n25687), .B2(
        \xmem_data[119][3] ), .ZN(n4754) );
  NAND4_X1 U8037 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4763)
         );
  AOI22_X1 U8038 ( .A1(n25692), .A2(\xmem_data[120][3] ), .B1(n3222), .B2(
        \xmem_data[121][3] ), .ZN(n4761) );
  AOI22_X1 U8039 ( .A1(n25693), .A2(\xmem_data[122][3] ), .B1(n20992), .B2(
        \xmem_data[123][3] ), .ZN(n4760) );
  AOI22_X1 U8040 ( .A1(n25694), .A2(\xmem_data[124][3] ), .B1(n13444), .B2(
        \xmem_data[125][3] ), .ZN(n4759) );
  AOI22_X1 U8041 ( .A1(n24702), .A2(\xmem_data[126][3] ), .B1(n27547), .B2(
        \xmem_data[127][3] ), .ZN(n4758) );
  NAND4_X1 U8042 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), .ZN(n4762)
         );
  OR4_X1 U8043 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), .ZN(n4766) );
  NAND2_X1 U8044 ( .A1(n4766), .A2(n25706), .ZN(n4767) );
  NAND2_X1 U8045 ( .A1(n4768), .A2(n4767), .ZN(n4769) );
  XNOR2_X1 U8046 ( .A(n31957), .B(\fmem_data[6][7] ), .ZN(n25746) );
  XOR2_X1 U8047 ( .A(\fmem_data[6][6] ), .B(\fmem_data[6][7] ), .Z(n4772) );
  AOI22_X1 U8048 ( .A1(n25635), .A2(\xmem_data[8][4] ), .B1(n25398), .B2(
        \xmem_data[9][4] ), .ZN(n4776) );
  AOI22_X1 U8049 ( .A1(n30309), .A2(\xmem_data[10][4] ), .B1(n29318), .B2(
        \xmem_data[11][4] ), .ZN(n4775) );
  AOI22_X1 U8050 ( .A1(n25632), .A2(\xmem_data[12][4] ), .B1(n28291), .B2(
        \xmem_data[13][4] ), .ZN(n4774) );
  AOI22_X1 U8051 ( .A1(n25636), .A2(\xmem_data[14][4] ), .B1(n24223), .B2(
        \xmem_data[15][4] ), .ZN(n4773) );
  NAND4_X1 U8052 ( .A1(n4776), .A2(n4775), .A3(n4774), .A4(n4773), .ZN(n4787)
         );
  AND2_X1 U8053 ( .A1(n17050), .A2(\xmem_data[19][4] ), .ZN(n4780) );
  AOI22_X1 U8054 ( .A1(n20734), .A2(\xmem_data[16][4] ), .B1(n25527), .B2(
        \xmem_data[17][4] ), .ZN(n4778) );
  AOI22_X1 U8055 ( .A1(n25624), .A2(\xmem_data[22][4] ), .B1(n30589), .B2(
        \xmem_data[23][4] ), .ZN(n4777) );
  NAND2_X1 U8056 ( .A1(n4778), .A2(n4777), .ZN(n4779) );
  AOI211_X1 U8057 ( .C1(\xmem_data[18][4] ), .C2(n25628), .A(n4780), .B(n4779), 
        .ZN(n4781) );
  AOI22_X1 U8058 ( .A1(n25604), .A2(\xmem_data[0][4] ), .B1(n27988), .B2(
        \xmem_data[1][4] ), .ZN(n4785) );
  AOI22_X1 U8059 ( .A1(n30943), .A2(\xmem_data[2][4] ), .B1(n25605), .B2(
        \xmem_data[3][4] ), .ZN(n4784) );
  AOI22_X1 U8060 ( .A1(n27515), .A2(\xmem_data[4][4] ), .B1(n25606), .B2(
        \xmem_data[5][4] ), .ZN(n4783) );
  AOI22_X1 U8061 ( .A1(n3158), .A2(\xmem_data[6][4] ), .B1(n28299), .B2(
        \xmem_data[7][4] ), .ZN(n4782) );
  NOR3_X1 U8062 ( .A1(n4787), .A2(n4786), .A3(n4017), .ZN(n4799) );
  NAND2_X1 U8063 ( .A1(n3375), .A2(\xmem_data[30][4] ), .ZN(n4789) );
  NAND2_X1 U8064 ( .A1(n3218), .A2(\xmem_data[25][4] ), .ZN(n4788) );
  NAND2_X1 U8065 ( .A1(n4789), .A2(n4788), .ZN(n4790) );
  AOI21_X1 U8066 ( .B1(n20991), .B2(\xmem_data[24][4] ), .A(n4790), .ZN(n4792)
         );
  AOI22_X1 U8067 ( .A1(n25617), .A2(\xmem_data[28][4] ), .B1(n25616), .B2(
        \xmem_data[29][4] ), .ZN(n4791) );
  NAND2_X1 U8068 ( .A1(n4792), .A2(n4791), .ZN(n4797) );
  AOI22_X1 U8069 ( .A1(n25630), .A2(\xmem_data[20][4] ), .B1(n25629), .B2(
        \xmem_data[21][4] ), .ZN(n4795) );
  NAND2_X1 U8070 ( .A1(n29103), .A2(\xmem_data[31][4] ), .ZN(n4794) );
  AOI22_X1 U8071 ( .A1(n25612), .A2(\xmem_data[26][4] ), .B1(n30963), .B2(
        \xmem_data[27][4] ), .ZN(n4793) );
  NAND3_X1 U8072 ( .A1(n4795), .A2(n4794), .A3(n4793), .ZN(n4796) );
  AOI21_X1 U8073 ( .B1(n4799), .B2(n4798), .A(n25647), .ZN(n4800) );
  INV_X1 U8074 ( .A(n4800), .ZN(n4866) );
  AOI22_X1 U8075 ( .A1(n25670), .A2(\xmem_data[96][4] ), .B1(n20546), .B2(
        \xmem_data[97][4] ), .ZN(n4804) );
  AOI22_X1 U8076 ( .A1(n25708), .A2(\xmem_data[98][4] ), .B1(n22740), .B2(
        \xmem_data[99][4] ), .ZN(n4803) );
  AOI22_X1 U8077 ( .A1(n16986), .A2(\xmem_data[100][4] ), .B1(n25671), .B2(
        \xmem_data[101][4] ), .ZN(n4802) );
  AOI22_X1 U8078 ( .A1(n25672), .A2(\xmem_data[102][4] ), .B1(n20543), .B2(
        \xmem_data[103][4] ), .ZN(n4801) );
  NAND4_X1 U8079 ( .A1(n4804), .A2(n4803), .A3(n4802), .A4(n4801), .ZN(n4820)
         );
  AOI22_X1 U8080 ( .A1(n21007), .A2(\xmem_data[104][4] ), .B1(n25677), .B2(
        \xmem_data[105][4] ), .ZN(n4808) );
  AOI22_X1 U8081 ( .A1(n25678), .A2(\xmem_data[106][4] ), .B1(n24646), .B2(
        \xmem_data[107][4] ), .ZN(n4807) );
  AOI22_X1 U8082 ( .A1(n20731), .A2(\xmem_data[108][4] ), .B1(n20551), .B2(
        \xmem_data[109][4] ), .ZN(n4806) );
  AOI22_X1 U8083 ( .A1(n3269), .A2(\xmem_data[110][4] ), .B1(n20781), .B2(
        \xmem_data[111][4] ), .ZN(n4805) );
  NAND4_X1 U8084 ( .A1(n4808), .A2(n4807), .A3(n4806), .A4(n4805), .ZN(n4819)
         );
  AOI22_X1 U8085 ( .A1(n31316), .A2(\xmem_data[112][4] ), .B1(n28292), .B2(
        \xmem_data[113][4] ), .ZN(n4812) );
  AOI22_X1 U8086 ( .A1(n25684), .A2(\xmem_data[114][4] ), .B1(n27957), .B2(
        \xmem_data[115][4] ), .ZN(n4811) );
  AOI22_X1 U8087 ( .A1(n25686), .A2(\xmem_data[116][4] ), .B1(n25685), .B2(
        \xmem_data[117][4] ), .ZN(n4810) );
  AOI22_X1 U8088 ( .A1(n3149), .A2(\xmem_data[118][4] ), .B1(n25687), .B2(
        \xmem_data[119][4] ), .ZN(n4809) );
  NAND4_X1 U8089 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(n4818)
         );
  AOI22_X1 U8090 ( .A1(n25692), .A2(\xmem_data[120][4] ), .B1(n3221), .B2(
        \xmem_data[121][4] ), .ZN(n4816) );
  AOI22_X1 U8091 ( .A1(n25693), .A2(\xmem_data[122][4] ), .B1(n24695), .B2(
        \xmem_data[123][4] ), .ZN(n4815) );
  AOI22_X1 U8092 ( .A1(n25694), .A2(\xmem_data[124][4] ), .B1(n3255), .B2(
        \xmem_data[125][4] ), .ZN(n4814) );
  AOI22_X1 U8093 ( .A1(n29706), .A2(\xmem_data[126][4] ), .B1(n29103), .B2(
        \xmem_data[127][4] ), .ZN(n4813) );
  NAND4_X1 U8094 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4817)
         );
  OR4_X1 U8095 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4842) );
  AOI22_X1 U8096 ( .A1(n25707), .A2(\xmem_data[64][4] ), .B1(n28415), .B2(
        \xmem_data[65][4] ), .ZN(n4824) );
  AOI22_X1 U8097 ( .A1(n25708), .A2(\xmem_data[66][4] ), .B1(n28515), .B2(
        \xmem_data[67][4] ), .ZN(n4823) );
  AOI22_X1 U8098 ( .A1(n24131), .A2(\xmem_data[68][4] ), .B1(n25709), .B2(
        \xmem_data[69][4] ), .ZN(n4822) );
  AOI22_X1 U8099 ( .A1(n27818), .A2(\xmem_data[70][4] ), .B1(n24134), .B2(
        \xmem_data[71][4] ), .ZN(n4821) );
  NAND4_X1 U8100 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .ZN(n4840)
         );
  AOI22_X1 U8101 ( .A1(n22676), .A2(\xmem_data[72][4] ), .B1(n25715), .B2(
        \xmem_data[73][4] ), .ZN(n4828) );
  AOI22_X1 U8102 ( .A1(n31255), .A2(\xmem_data[74][4] ), .B1(n30871), .B2(
        \xmem_data[75][4] ), .ZN(n4827) );
  AOI22_X1 U8103 ( .A1(n17002), .A2(\xmem_data[76][4] ), .B1(n25679), .B2(
        \xmem_data[77][4] ), .ZN(n4826) );
  AOI22_X1 U8104 ( .A1(n25718), .A2(\xmem_data[78][4] ), .B1(n24570), .B2(
        \xmem_data[79][4] ), .ZN(n4825) );
  NAND4_X1 U8105 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .ZN(n4839)
         );
  AOI22_X1 U8106 ( .A1(n24166), .A2(\xmem_data[80][4] ), .B1(n25723), .B2(
        \xmem_data[81][4] ), .ZN(n4832) );
  AOI22_X1 U8107 ( .A1(n20770), .A2(\xmem_data[82][4] ), .B1(n22727), .B2(
        \xmem_data[83][4] ), .ZN(n4831) );
  AOI22_X1 U8108 ( .A1(n25724), .A2(\xmem_data[84][4] ), .B1(n31346), .B2(
        \xmem_data[85][4] ), .ZN(n4830) );
  AOI22_X1 U8109 ( .A1(n25725), .A2(\xmem_data[86][4] ), .B1(n25360), .B2(
        \xmem_data[87][4] ), .ZN(n4829) );
  NAND4_X1 U8110 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .ZN(n4838)
         );
  AOI22_X1 U8111 ( .A1(n25730), .A2(\xmem_data[88][4] ), .B1(n3221), .B2(
        \xmem_data[89][4] ), .ZN(n4836) );
  AOI22_X1 U8112 ( .A1(n25731), .A2(\xmem_data[90][4] ), .B1(n25491), .B2(
        \xmem_data[91][4] ), .ZN(n4835) );
  AOI22_X1 U8113 ( .A1(n25449), .A2(\xmem_data[92][4] ), .B1(n30550), .B2(
        \xmem_data[93][4] ), .ZN(n4834) );
  AOI22_X1 U8114 ( .A1(n25732), .A2(\xmem_data[94][4] ), .B1(n29306), .B2(
        \xmem_data[95][4] ), .ZN(n4833) );
  NAND4_X1 U8115 ( .A1(n4836), .A2(n4835), .A3(n4834), .A4(n4833), .ZN(n4837)
         );
  OR4_X1 U8116 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4841) );
  AOI22_X1 U8117 ( .A1(n25706), .A2(n4842), .B1(n25704), .B2(n4841), .ZN(n4865) );
  AOI22_X1 U8118 ( .A1(n25707), .A2(\xmem_data[32][4] ), .B1(n27943), .B2(
        \xmem_data[33][4] ), .ZN(n4846) );
  AOI22_X1 U8119 ( .A1(n25708), .A2(\xmem_data[34][4] ), .B1(n31326), .B2(
        \xmem_data[35][4] ), .ZN(n4845) );
  AOI22_X1 U8120 ( .A1(n30891), .A2(\xmem_data[36][4] ), .B1(n25709), .B2(
        \xmem_data[37][4] ), .ZN(n4844) );
  AOI22_X1 U8121 ( .A1(n30746), .A2(\xmem_data[38][4] ), .B1(n31269), .B2(
        \xmem_data[39][4] ), .ZN(n4843) );
  NAND4_X1 U8122 ( .A1(n4846), .A2(n4845), .A3(n4844), .A4(n4843), .ZN(n4862)
         );
  AOI22_X1 U8123 ( .A1(n25573), .A2(\xmem_data[40][4] ), .B1(n25715), .B2(
        \xmem_data[41][4] ), .ZN(n4850) );
  AOI22_X1 U8124 ( .A1(n23722), .A2(\xmem_data[42][4] ), .B1(n29280), .B2(
        \xmem_data[43][4] ), .ZN(n4849) );
  AOI22_X1 U8125 ( .A1(n3326), .A2(\xmem_data[44][4] ), .B1(n21009), .B2(
        \xmem_data[45][4] ), .ZN(n4848) );
  AOI22_X1 U8126 ( .A1(n25718), .A2(\xmem_data[46][4] ), .B1(n22685), .B2(
        \xmem_data[47][4] ), .ZN(n4847) );
  NAND4_X1 U8127 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4861)
         );
  AOI22_X1 U8128 ( .A1(n3209), .A2(\xmem_data[48][4] ), .B1(n25723), .B2(
        \xmem_data[49][4] ), .ZN(n4854) );
  AOI22_X1 U8129 ( .A1(n28467), .A2(\xmem_data[50][4] ), .B1(n20769), .B2(
        \xmem_data[51][4] ), .ZN(n4853) );
  AOI22_X1 U8130 ( .A1(n25724), .A2(\xmem_data[52][4] ), .B1(n21309), .B2(
        \xmem_data[53][4] ), .ZN(n4852) );
  AOI22_X1 U8131 ( .A1(n25725), .A2(\xmem_data[54][4] ), .B1(n27501), .B2(
        \xmem_data[55][4] ), .ZN(n4851) );
  NAND4_X1 U8132 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n4860)
         );
  AOI22_X1 U8133 ( .A1(n25730), .A2(\xmem_data[56][4] ), .B1(n3219), .B2(
        \xmem_data[57][4] ), .ZN(n4858) );
  AOI22_X1 U8134 ( .A1(n25731), .A2(\xmem_data[58][4] ), .B1(n28508), .B2(
        \xmem_data[59][4] ), .ZN(n4857) );
  AOI22_X1 U8135 ( .A1(n22666), .A2(\xmem_data[60][4] ), .B1(n20559), .B2(
        \xmem_data[61][4] ), .ZN(n4856) );
  AOI22_X1 U8136 ( .A1(n25732), .A2(\xmem_data[62][4] ), .B1(n3231), .B2(
        \xmem_data[63][4] ), .ZN(n4855) );
  NAND4_X1 U8137 ( .A1(n4858), .A2(n4857), .A3(n4856), .A4(n4855), .ZN(n4859)
         );
  OR4_X1 U8138 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4863) );
  NAND2_X1 U8139 ( .A1(n4863), .A2(n25741), .ZN(n4864) );
  XNOR2_X1 U8140 ( .A(n31958), .B(\fmem_data[6][7] ), .ZN(n13912) );
  OAI22_X1 U8141 ( .A1(n25746), .A2(n35511), .B1(n13912), .B2(n35512), .ZN(
        n33342) );
  AOI22_X1 U8142 ( .A1(n25629), .A2(\xmem_data[96][3] ), .B1(n24693), .B2(
        \xmem_data[97][3] ), .ZN(n4870) );
  BUF_X1 U8143 ( .A(n29064), .Z(n25508) );
  AOI22_X1 U8144 ( .A1(n25360), .A2(\xmem_data[98][3] ), .B1(n25508), .B2(
        \xmem_data[99][3] ), .ZN(n4869) );
  AOI22_X1 U8145 ( .A1(n3219), .A2(\xmem_data[100][3] ), .B1(n28137), .B2(
        \xmem_data[101][3] ), .ZN(n4868) );
  BUF_X1 U8146 ( .A(n14925), .Z(n25509) );
  AOI22_X1 U8147 ( .A1(n25509), .A2(\xmem_data[102][3] ), .B1(n20725), .B2(
        \xmem_data[103][3] ), .ZN(n4867) );
  NAND4_X1 U8148 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(n4886)
         );
  AOI22_X1 U8149 ( .A1(n25486), .A2(\xmem_data[104][3] ), .B1(n3131), .B2(
        \xmem_data[105][3] ), .ZN(n4874) );
  AOI22_X1 U8150 ( .A1(n25514), .A2(\xmem_data[106][3] ), .B1(n27910), .B2(
        \xmem_data[107][3] ), .ZN(n4873) );
  AOI22_X1 U8151 ( .A1(n28481), .A2(\xmem_data[108][3] ), .B1(n20799), .B2(
        \xmem_data[109][3] ), .ZN(n4872) );
  AOI22_X1 U8152 ( .A1(n20775), .A2(\xmem_data[110][3] ), .B1(n29310), .B2(
        \xmem_data[111][3] ), .ZN(n4871) );
  NAND4_X1 U8153 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n4885)
         );
  BUF_X1 U8154 ( .A(n3464), .Z(n25519) );
  AOI22_X1 U8155 ( .A1(n21076), .A2(\xmem_data[112][3] ), .B1(n25519), .B2(
        \xmem_data[113][3] ), .ZN(n4878) );
  AOI22_X1 U8156 ( .A1(n20938), .A2(\xmem_data[114][3] ), .B1(n23717), .B2(
        \xmem_data[115][3] ), .ZN(n4877) );
  BUF_X1 U8157 ( .A(n13415), .Z(n25520) );
  AOI22_X1 U8158 ( .A1(n25520), .A2(\xmem_data[116][3] ), .B1(n29319), .B2(
        \xmem_data[117][3] ), .ZN(n4876) );
  BUF_X1 U8159 ( .A(n14881), .Z(n25521) );
  AOI22_X1 U8160 ( .A1(n20941), .A2(\xmem_data[118][3] ), .B1(n25521), .B2(
        \xmem_data[119][3] ), .ZN(n4875) );
  NAND4_X1 U8161 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4884)
         );
  AOI22_X1 U8162 ( .A1(n17001), .A2(\xmem_data[120][3] ), .B1(n25718), .B2(
        \xmem_data[121][3] ), .ZN(n4882) );
  BUF_X1 U8163 ( .A(n14976), .Z(n25526) );
  AOI22_X1 U8164 ( .A1(n20553), .A2(\xmem_data[122][3] ), .B1(n25526), .B2(
        \xmem_data[123][3] ), .ZN(n4881) );
  AOI22_X1 U8165 ( .A1(n25527), .A2(\xmem_data[124][3] ), .B1(n28036), .B2(
        \xmem_data[125][3] ), .ZN(n4880) );
  BUF_X1 U8166 ( .A(n13457), .Z(n25528) );
  AOI22_X1 U8167 ( .A1(n25528), .A2(\xmem_data[126][3] ), .B1(n28076), .B2(
        \xmem_data[127][3] ), .ZN(n4879) );
  NAND4_X1 U8168 ( .A1(n4882), .A2(n4881), .A3(n4880), .A4(n4879), .ZN(n4883)
         );
  OR4_X1 U8169 ( .A1(n4886), .A2(n4885), .A3(n4884), .A4(n4883), .ZN(n4890) );
  AOI21_X1 U8170 ( .B1(n6172), .B2(n10590), .A(n10589), .ZN(n4887) );
  INV_X1 U8171 ( .A(n4887), .ZN(n4888) );
  AOI22_X1 U8172 ( .A1(n37191), .A2(n4888), .B1(n4887), .B2(n4499), .ZN(n4959)
         );
  NAND2_X1 U8173 ( .A1(load_xaddr_val[5]), .A2(n4888), .ZN(n4889) );
  XOR2_X1 U8174 ( .A(n39040), .B(n4889), .Z(n4958) );
  AND2_X1 U8175 ( .A1(n4959), .A2(n4958), .ZN(n25560) );
  AND2_X1 U8176 ( .A1(n4890), .A2(n25560), .ZN(n4965) );
  BUF_X1 U8177 ( .A(n28974), .Z(n25561) );
  AOI22_X1 U8178 ( .A1(n25561), .A2(\xmem_data[32][3] ), .B1(n28164), .B2(
        \xmem_data[33][3] ), .ZN(n4894) );
  AOI22_X1 U8179 ( .A1(n27437), .A2(\xmem_data[34][3] ), .B1(n25413), .B2(
        \xmem_data[35][3] ), .ZN(n4893) );
  AOI22_X1 U8180 ( .A1(n3220), .A2(\xmem_data[36][3] ), .B1(n29431), .B2(
        \xmem_data[37][3] ), .ZN(n4892) );
  AOI22_X1 U8181 ( .A1(n25562), .A2(\xmem_data[38][3] ), .B1(n3342), .B2(
        \xmem_data[39][3] ), .ZN(n4891) );
  NAND4_X1 U8182 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n4910)
         );
  AOI22_X1 U8183 ( .A1(n27550), .A2(\xmem_data[40][3] ), .B1(n3146), .B2(
        \xmem_data[41][3] ), .ZN(n4898) );
  AOI22_X1 U8184 ( .A1(n30877), .A2(\xmem_data[42][3] ), .B1(n30885), .B2(
        \xmem_data[43][3] ), .ZN(n4897) );
  AOI22_X1 U8185 ( .A1(n3358), .A2(\xmem_data[44][3] ), .B1(n28089), .B2(
        \xmem_data[45][3] ), .ZN(n4896) );
  BUF_X1 U8186 ( .A(n13476), .Z(n25567) );
  AOI22_X1 U8187 ( .A1(n25423), .A2(\xmem_data[46][3] ), .B1(n25567), .B2(
        \xmem_data[47][3] ), .ZN(n4895) );
  NAND4_X1 U8188 ( .A1(n4898), .A2(n4897), .A3(n4896), .A4(n4895), .ZN(n4909)
         );
  BUF_X1 U8189 ( .A(n14999), .Z(n25572) );
  AOI22_X1 U8190 ( .A1(n25572), .A2(\xmem_data[48][3] ), .B1(n30746), .B2(
        \xmem_data[49][3] ), .ZN(n4902) );
  AOI22_X1 U8191 ( .A1(n25574), .A2(\xmem_data[50][3] ), .B1(n25573), .B2(
        \xmem_data[51][3] ), .ZN(n4901) );
  AOI22_X1 U8192 ( .A1(n29316), .A2(\xmem_data[52][3] ), .B1(n27855), .B2(
        \xmem_data[53][3] ), .ZN(n4900) );
  BUF_X1 U8193 ( .A(n13452), .Z(n25576) );
  BUF_X1 U8194 ( .A(n4158), .Z(n25575) );
  AOI22_X1 U8195 ( .A1(n25576), .A2(\xmem_data[54][3] ), .B1(n25575), .B2(
        \xmem_data[55][3] ), .ZN(n4899) );
  NAND4_X1 U8196 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4908)
         );
  AOI22_X1 U8197 ( .A1(n30598), .A2(\xmem_data[56][3] ), .B1(n3300), .B2(
        \xmem_data[57][3] ), .ZN(n4906) );
  BUF_X1 U8198 ( .A(n14914), .Z(n25583) );
  AOI22_X1 U8199 ( .A1(n25583), .A2(\xmem_data[58][3] ), .B1(n25582), .B2(
        \xmem_data[59][3] ), .ZN(n4905) );
  BUF_X1 U8200 ( .A(n13127), .Z(n25584) );
  AOI22_X1 U8201 ( .A1(n25527), .A2(\xmem_data[60][3] ), .B1(n25584), .B2(
        \xmem_data[61][3] ), .ZN(n4904) );
  AOI22_X1 U8202 ( .A1(n30498), .A2(\xmem_data[62][3] ), .B1(n20827), .B2(
        \xmem_data[63][3] ), .ZN(n4903) );
  NAND4_X1 U8203 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907)
         );
  OR4_X1 U8204 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n4911) );
  INV_X1 U8205 ( .A(n4958), .ZN(n4932) );
  AND2_X1 U8206 ( .A1(n4932), .A2(n4959), .ZN(n25593) );
  AND2_X1 U8207 ( .A1(n4911), .A2(n25593), .ZN(n4964) );
  AOI22_X1 U8208 ( .A1(n30863), .A2(\xmem_data[66][3] ), .B1(n25508), .B2(
        \xmem_data[67][3] ), .ZN(n4915) );
  AOI22_X1 U8209 ( .A1(n20489), .A2(\xmem_data[64][3] ), .B1(n27813), .B2(
        \xmem_data[65][3] ), .ZN(n4914) );
  AOI22_X1 U8210 ( .A1(n3221), .A2(\xmem_data[68][3] ), .B1(n20724), .B2(
        \xmem_data[69][3] ), .ZN(n4913) );
  AOI22_X1 U8211 ( .A1(n25509), .A2(\xmem_data[70][3] ), .B1(n28475), .B2(
        \xmem_data[71][3] ), .ZN(n4912) );
  NAND4_X1 U8212 ( .A1(n4915), .A2(n4914), .A3(n4913), .A4(n4912), .ZN(n4931)
         );
  AOI22_X1 U8213 ( .A1(n21068), .A2(\xmem_data[72][3] ), .B1(n30295), .B2(
        \xmem_data[73][3] ), .ZN(n4919) );
  AOI22_X1 U8214 ( .A1(n25514), .A2(\xmem_data[74][3] ), .B1(n24638), .B2(
        \xmem_data[75][3] ), .ZN(n4918) );
  AOI22_X1 U8215 ( .A1(n20588), .A2(\xmem_data[76][3] ), .B1(n25708), .B2(
        \xmem_data[77][3] ), .ZN(n4917) );
  AOI22_X1 U8216 ( .A1(n20775), .A2(\xmem_data[78][3] ), .B1(n31268), .B2(
        \xmem_data[79][3] ), .ZN(n4916) );
  NAND4_X1 U8217 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n4930)
         );
  AOI22_X1 U8218 ( .A1(n25709), .A2(\xmem_data[80][3] ), .B1(n25519), .B2(
        \xmem_data[81][3] ), .ZN(n4923) );
  AOI22_X1 U8219 ( .A1(n25574), .A2(\xmem_data[82][3] ), .B1(n21007), .B2(
        \xmem_data[83][3] ), .ZN(n4922) );
  AOI22_X1 U8220 ( .A1(n25520), .A2(\xmem_data[84][3] ), .B1(n25678), .B2(
        \xmem_data[85][3] ), .ZN(n4921) );
  AOI22_X1 U8221 ( .A1(n24165), .A2(\xmem_data[86][3] ), .B1(n25521), .B2(
        \xmem_data[87][3] ), .ZN(n4920) );
  NAND4_X1 U8222 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(n4929)
         );
  AOI22_X1 U8223 ( .A1(n28494), .A2(\xmem_data[88][3] ), .B1(n3271), .B2(
        \xmem_data[89][3] ), .ZN(n4927) );
  AOI22_X1 U8224 ( .A1(n28983), .A2(\xmem_data[90][3] ), .B1(n25526), .B2(
        \xmem_data[91][3] ), .ZN(n4926) );
  AOI22_X1 U8225 ( .A1(n25527), .A2(\xmem_data[92][3] ), .B1(n29327), .B2(
        \xmem_data[93][3] ), .ZN(n4925) );
  AOI22_X1 U8226 ( .A1(n25528), .A2(\xmem_data[94][3] ), .B1(n24688), .B2(
        \xmem_data[95][3] ), .ZN(n4924) );
  NAND4_X1 U8227 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n4928)
         );
  OR4_X1 U8228 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(n4933) );
  NOR2_X1 U8229 ( .A1(n4959), .A2(n4932), .ZN(n25558) );
  NAND2_X1 U8230 ( .A1(n4933), .A2(n25558), .ZN(n4962) );
  AOI22_X1 U8231 ( .A1(n20775), .A2(\xmem_data[14][3] ), .B1(n27537), .B2(
        \xmem_data[15][3] ), .ZN(n4935) );
  AOI22_X1 U8232 ( .A1(n24556), .A2(\xmem_data[13][3] ), .B1(\xmem_data[9][3] ), .B2(n29567), .ZN(n4934) );
  NAND2_X1 U8233 ( .A1(n4935), .A2(n4934), .ZN(n4939) );
  BUF_X1 U8234 ( .A(n15011), .Z(n25492) );
  BUF_X1 U8235 ( .A(n10999), .Z(n25481) );
  BUF_X1 U8236 ( .A(n14927), .Z(n25486) );
  NAND2_X1 U8237 ( .A1(n4937), .A2(n4936), .ZN(n4938) );
  OR3_X1 U8238 ( .A1(n4939), .A2(n4019), .A3(n4938), .ZN(n4957) );
  AOI22_X1 U8239 ( .A1(n20816), .A2(\xmem_data[24][3] ), .B1(n21056), .B2(
        \xmem_data[25][3] ), .ZN(n4943) );
  AOI22_X1 U8240 ( .A1(n20781), .A2(\xmem_data[26][3] ), .B1(n20734), .B2(
        \xmem_data[27][3] ), .ZN(n4942) );
  AOI22_X1 U8241 ( .A1(n23781), .A2(\xmem_data[28][3] ), .B1(n13420), .B2(
        \xmem_data[29][3] ), .ZN(n4941) );
  AOI22_X1 U8242 ( .A1(n10456), .A2(\xmem_data[30][3] ), .B1(n20986), .B2(
        \xmem_data[31][3] ), .ZN(n4940) );
  NAND4_X1 U8243 ( .A1(n4943), .A2(n4942), .A3(n4941), .A4(n4940), .ZN(n4945)
         );
  AND2_X1 U8244 ( .A1(n25670), .A2(\xmem_data[11][3] ), .ZN(n4944) );
  OR2_X1 U8245 ( .A1(n4945), .A2(n4944), .ZN(n4956) );
  AOI22_X1 U8246 ( .A1(n24573), .A2(\xmem_data[0][3] ), .B1(n3305), .B2(
        \xmem_data[1][3] ), .ZN(n4949) );
  BUF_X1 U8247 ( .A(n13468), .Z(n25485) );
  AOI22_X1 U8248 ( .A1(n25485), .A2(\xmem_data[2][3] ), .B1(n28364), .B2(
        \xmem_data[3][3] ), .ZN(n4948) );
  AOI22_X1 U8249 ( .A1(n3219), .A2(\xmem_data[4][3] ), .B1(n29494), .B2(
        \xmem_data[5][3] ), .ZN(n4947) );
  BUF_X1 U8250 ( .A(n14990), .Z(n25490) );
  AOI22_X1 U8251 ( .A1(n25491), .A2(\xmem_data[6][3] ), .B1(n25490), .B2(
        \xmem_data[7][3] ), .ZN(n4946) );
  NAND4_X1 U8252 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4955)
         );
  AOI22_X1 U8253 ( .A1(n25572), .A2(\xmem_data[16][3] ), .B1(n21005), .B2(
        \xmem_data[17][3] ), .ZN(n4953) );
  AOI22_X1 U8254 ( .A1(n27454), .A2(\xmem_data[18][3] ), .B1(n31330), .B2(
        \xmem_data[19][3] ), .ZN(n4952) );
  AOI22_X1 U8255 ( .A1(n28492), .A2(\xmem_data[20][3] ), .B1(n17044), .B2(
        \xmem_data[21][3] ), .ZN(n4951) );
  AOI22_X1 U8256 ( .A1(n29318), .A2(\xmem_data[22][3] ), .B1(n3326), .B2(
        \xmem_data[23][3] ), .ZN(n4950) );
  NAND4_X1 U8257 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4954)
         );
  OR4_X1 U8258 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n4960) );
  NOR2_X1 U8259 ( .A1(n4959), .A2(n4958), .ZN(n19110) );
  INV_X1 U8260 ( .A(n19110), .ZN(n25505) );
  NAND2_X1 U8261 ( .A1(n4960), .A2(n19110), .ZN(n4961) );
  NAND2_X1 U8262 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  XOR2_X1 U8263 ( .A(\fmem_data[17][6] ), .B(\fmem_data[17][7] ), .Z(n4966) );
  AOI22_X1 U8264 ( .A1(n25481), .A2(\xmem_data[12][4] ), .B1(n28671), .B2(
        \xmem_data[13][4] ), .ZN(n4967) );
  INV_X1 U8265 ( .A(n4967), .ZN(n4978) );
  AOI22_X1 U8266 ( .A1(n30598), .A2(\xmem_data[24][4] ), .B1(n23780), .B2(
        \xmem_data[25][4] ), .ZN(n4972) );
  AOI22_X1 U8267 ( .A1(n27525), .A2(\xmem_data[26][4] ), .B1(n27542), .B2(
        \xmem_data[27][4] ), .ZN(n4971) );
  AND2_X1 U8268 ( .A1(n23725), .A2(\xmem_data[28][4] ), .ZN(n4968) );
  AOI21_X1 U8269 ( .B1(n28192), .B2(\xmem_data[29][4] ), .A(n4968), .ZN(n4970)
         );
  AOI22_X1 U8270 ( .A1(n24122), .A2(\xmem_data[30][4] ), .B1(n25358), .B2(
        \xmem_data[31][4] ), .ZN(n4969) );
  NAND4_X1 U8271 ( .A1(n4972), .A2(n4971), .A3(n4970), .A4(n4969), .ZN(n4977)
         );
  AOI22_X1 U8272 ( .A1(n25486), .A2(\xmem_data[8][4] ), .B1(n3375), .B2(
        \xmem_data[9][4] ), .ZN(n4975) );
  AOI22_X1 U8273 ( .A1(n27513), .A2(\xmem_data[14][4] ), .B1(n16986), .B2(
        \xmem_data[15][4] ), .ZN(n4974) );
  NAND2_X1 U8274 ( .A1(n25422), .A2(\xmem_data[11][4] ), .ZN(n4973) );
  NAND3_X1 U8275 ( .A1(n4975), .A2(n4974), .A3(n4973), .ZN(n4976) );
  NOR3_X1 U8276 ( .A1(n4978), .A2(n4977), .A3(n4976), .ZN(n4989) );
  AND2_X1 U8277 ( .A1(n25485), .A2(\xmem_data[2][4] ), .ZN(n4979) );
  AOI21_X1 U8278 ( .B1(n28044), .B2(\xmem_data[3][4] ), .A(n4979), .ZN(n4983)
         );
  AOI22_X1 U8279 ( .A1(n25561), .A2(\xmem_data[0][4] ), .B1(n29661), .B2(
        \xmem_data[1][4] ), .ZN(n4982) );
  AOI22_X1 U8280 ( .A1(n3222), .A2(\xmem_data[4][4] ), .B1(n29422), .B2(
        \xmem_data[5][4] ), .ZN(n4981) );
  AOI22_X1 U8281 ( .A1(n25491), .A2(\xmem_data[6][4] ), .B1(n25490), .B2(
        \xmem_data[7][4] ), .ZN(n4980) );
  AND4_X1 U8282 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n4988)
         );
  AOI22_X1 U8283 ( .A1(n25572), .A2(\xmem_data[16][4] ), .B1(n27755), .B2(
        \xmem_data[17][4] ), .ZN(n4987) );
  AOI22_X1 U8284 ( .A1(n29279), .A2(\xmem_data[18][4] ), .B1(n25434), .B2(
        \xmem_data[19][4] ), .ZN(n4986) );
  AOI22_X1 U8285 ( .A1(n29048), .A2(\xmem_data[20][4] ), .B1(n28781), .B2(
        \xmem_data[21][4] ), .ZN(n4985) );
  AOI22_X1 U8286 ( .A1(n25435), .A2(\xmem_data[22][4] ), .B1(n28428), .B2(
        \xmem_data[23][4] ), .ZN(n4984) );
  AND3_X1 U8287 ( .A1(n4989), .A2(n4988), .A3(n3915), .ZN(n4991) );
  NAND2_X1 U8288 ( .A1(n25492), .A2(\xmem_data[10][4] ), .ZN(n4990) );
  AOI21_X1 U8289 ( .B1(n4991), .B2(n4990), .A(n25505), .ZN(n4992) );
  INV_X1 U8290 ( .A(n4992), .ZN(n5060) );
  AOI22_X1 U8291 ( .A1(n25561), .A2(\xmem_data[64][4] ), .B1(n3434), .B2(
        \xmem_data[65][4] ), .ZN(n4997) );
  AND2_X1 U8292 ( .A1(n25360), .A2(\xmem_data[66][4] ), .ZN(n4993) );
  AOI21_X1 U8293 ( .B1(n20576), .B2(\xmem_data[67][4] ), .A(n4993), .ZN(n4996)
         );
  AOI22_X1 U8294 ( .A1(n3218), .A2(\xmem_data[68][4] ), .B1(n27708), .B2(
        \xmem_data[69][4] ), .ZN(n4995) );
  AOI22_X1 U8295 ( .A1(n25562), .A2(\xmem_data[70][4] ), .B1(n3342), .B2(
        \xmem_data[71][4] ), .ZN(n4994) );
  NAND4_X1 U8296 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n5014)
         );
  AOI22_X1 U8297 ( .A1(n20559), .A2(\xmem_data[72][4] ), .B1(n3140), .B2(
        \xmem_data[73][4] ), .ZN(n5001) );
  AOI22_X1 U8298 ( .A1(n29306), .A2(\xmem_data[74][4] ), .B1(n27551), .B2(
        \xmem_data[75][4] ), .ZN(n5000) );
  AOI22_X1 U8299 ( .A1(n25481), .A2(\xmem_data[76][4] ), .B1(n20587), .B2(
        \xmem_data[77][4] ), .ZN(n4999) );
  AOI22_X1 U8300 ( .A1(n22740), .A2(\xmem_data[78][4] ), .B1(n25567), .B2(
        \xmem_data[79][4] ), .ZN(n4998) );
  NAND4_X1 U8301 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n5013)
         );
  AOI22_X1 U8302 ( .A1(n20584), .A2(\xmem_data[80][4] ), .B1(n29396), .B2(
        \xmem_data[81][4] ), .ZN(n5005) );
  AOI22_X1 U8303 ( .A1(n25574), .A2(\xmem_data[82][4] ), .B1(n25573), .B2(
        \xmem_data[83][4] ), .ZN(n5004) );
  AOI22_X1 U8304 ( .A1(n17043), .A2(\xmem_data[84][4] ), .B1(n25678), .B2(
        \xmem_data[85][4] ), .ZN(n5003) );
  AOI22_X1 U8305 ( .A1(n25576), .A2(\xmem_data[86][4] ), .B1(n25575), .B2(
        \xmem_data[87][4] ), .ZN(n5002) );
  NAND4_X1 U8306 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n5012)
         );
  AOI22_X1 U8307 ( .A1(n25581), .A2(\xmem_data[88][4] ), .B1(n3330), .B2(
        \xmem_data[89][4] ), .ZN(n5010) );
  AOI22_X1 U8308 ( .A1(n25583), .A2(\xmem_data[90][4] ), .B1(n25582), .B2(
        \xmem_data[91][4] ), .ZN(n5009) );
  AND2_X1 U8309 ( .A1(n25527), .A2(\xmem_data[92][4] ), .ZN(n5006) );
  AOI21_X1 U8310 ( .B1(n25584), .B2(\xmem_data[93][4] ), .A(n5006), .ZN(n5008)
         );
  AOI22_X1 U8311 ( .A1(n28329), .A2(\xmem_data[94][4] ), .B1(n27925), .B2(
        \xmem_data[95][4] ), .ZN(n5007) );
  NAND4_X1 U8312 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n5011)
         );
  OR4_X1 U8313 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n5036) );
  AOI22_X1 U8314 ( .A1(n20489), .A2(\xmem_data[96][4] ), .B1(n23754), .B2(
        \xmem_data[97][4] ), .ZN(n5018) );
  AOI22_X1 U8315 ( .A1(n27501), .A2(\xmem_data[98][4] ), .B1(n25508), .B2(
        \xmem_data[99][4] ), .ZN(n5017) );
  AOI22_X1 U8316 ( .A1(n3219), .A2(\xmem_data[100][4] ), .B1(n29789), .B2(
        \xmem_data[101][4] ), .ZN(n5016) );
  AOI22_X1 U8317 ( .A1(n25509), .A2(\xmem_data[102][4] ), .B1(n25416), .B2(
        \xmem_data[103][4] ), .ZN(n5015) );
  NAND4_X1 U8318 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n5034)
         );
  AOI22_X1 U8319 ( .A1(n27903), .A2(\xmem_data[104][4] ), .B1(n29706), .B2(
        \xmem_data[105][4] ), .ZN(n5022) );
  AOI22_X1 U8320 ( .A1(n25514), .A2(\xmem_data[106][4] ), .B1(n23813), .B2(
        \xmem_data[107][4] ), .ZN(n5021) );
  AOI22_X1 U8321 ( .A1(n25456), .A2(\xmem_data[108][4] ), .B1(n30508), .B2(
        \xmem_data[109][4] ), .ZN(n5020) );
  AOI22_X1 U8322 ( .A1(n27452), .A2(\xmem_data[110][4] ), .B1(n28980), .B2(
        \xmem_data[111][4] ), .ZN(n5019) );
  NAND4_X1 U8323 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n5033)
         );
  AOI22_X1 U8324 ( .A1(n25572), .A2(\xmem_data[112][4] ), .B1(n25519), .B2(
        \xmem_data[113][4] ), .ZN(n5026) );
  AOI22_X1 U8325 ( .A1(n22677), .A2(\xmem_data[114][4] ), .B1(n25635), .B2(
        \xmem_data[115][4] ), .ZN(n5025) );
  AOI22_X1 U8326 ( .A1(n25520), .A2(\xmem_data[116][4] ), .B1(n20730), .B2(
        \xmem_data[117][4] ), .ZN(n5024) );
  AOI22_X1 U8327 ( .A1(n30515), .A2(\xmem_data[118][4] ), .B1(n25521), .B2(
        \xmem_data[119][4] ), .ZN(n5023) );
  NAND4_X1 U8328 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n5032)
         );
  AOI22_X1 U8329 ( .A1(n30955), .A2(\xmem_data[120][4] ), .B1(n23724), .B2(
        \xmem_data[121][4] ), .ZN(n5030) );
  AOI22_X1 U8330 ( .A1(n14975), .A2(\xmem_data[122][4] ), .B1(n25526), .B2(
        \xmem_data[123][4] ), .ZN(n5029) );
  AOI22_X1 U8331 ( .A1(n25527), .A2(\xmem_data[124][4] ), .B1(n13127), .B2(
        \xmem_data[125][4] ), .ZN(n5028) );
  AOI22_X1 U8332 ( .A1(n25528), .A2(\xmem_data[126][4] ), .B1(n29124), .B2(
        \xmem_data[127][4] ), .ZN(n5027) );
  NAND4_X1 U8333 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5031)
         );
  OR4_X1 U8334 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5035) );
  AOI22_X1 U8335 ( .A1(n5036), .A2(n25558), .B1(n5035), .B2(n25560), .ZN(n5059) );
  AOI22_X1 U8336 ( .A1(n25561), .A2(\xmem_data[32][4] ), .B1(n28039), .B2(
        \xmem_data[33][4] ), .ZN(n5040) );
  AOI22_X1 U8337 ( .A1(n25687), .A2(\xmem_data[34][4] ), .B1(n27439), .B2(
        \xmem_data[35][4] ), .ZN(n5039) );
  AOI22_X1 U8338 ( .A1(n3217), .A2(\xmem_data[36][4] ), .B1(n24563), .B2(
        \xmem_data[37][4] ), .ZN(n5038) );
  AOI22_X1 U8339 ( .A1(n25562), .A2(\xmem_data[38][4] ), .B1(n3342), .B2(
        \xmem_data[39][4] ), .ZN(n5037) );
  NAND4_X1 U8340 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n5056)
         );
  AOI22_X1 U8341 ( .A1(n25486), .A2(\xmem_data[40][4] ), .B1(n30698), .B2(
        \xmem_data[41][4] ), .ZN(n5044) );
  AOI22_X1 U8342 ( .A1(n25450), .A2(\xmem_data[42][4] ), .B1(n27910), .B2(
        \xmem_data[43][4] ), .ZN(n5043) );
  AOI22_X1 U8343 ( .A1(n29180), .A2(\xmem_data[44][4] ), .B1(n24157), .B2(
        \xmem_data[45][4] ), .ZN(n5042) );
  AOI22_X1 U8344 ( .A1(n21075), .A2(\xmem_data[46][4] ), .B1(n25567), .B2(
        \xmem_data[47][4] ), .ZN(n5041) );
  NAND4_X1 U8345 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n5055)
         );
  AOI22_X1 U8346 ( .A1(n28052), .A2(\xmem_data[48][4] ), .B1(n27455), .B2(
        \xmem_data[49][4] ), .ZN(n5048) );
  AOI22_X1 U8347 ( .A1(n25574), .A2(\xmem_data[50][4] ), .B1(n25573), .B2(
        \xmem_data[51][4] ), .ZN(n5047) );
  AOI22_X1 U8348 ( .A1(n25398), .A2(\xmem_data[52][4] ), .B1(n28687), .B2(
        \xmem_data[53][4] ), .ZN(n5046) );
  AOI22_X1 U8349 ( .A1(n25576), .A2(\xmem_data[54][4] ), .B1(n25575), .B2(
        \xmem_data[55][4] ), .ZN(n5045) );
  NAND4_X1 U8350 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n5054)
         );
  AOI22_X1 U8351 ( .A1(n29281), .A2(\xmem_data[56][4] ), .B1(n30600), .B2(
        \xmem_data[57][4] ), .ZN(n5052) );
  AOI22_X1 U8352 ( .A1(n25583), .A2(\xmem_data[58][4] ), .B1(n25582), .B2(
        \xmem_data[59][4] ), .ZN(n5051) );
  AOI22_X1 U8353 ( .A1(n14981), .A2(\xmem_data[60][4] ), .B1(n25584), .B2(
        \xmem_data[61][4] ), .ZN(n5050) );
  AOI22_X1 U8354 ( .A1(n21059), .A2(\xmem_data[62][4] ), .B1(n20710), .B2(
        \xmem_data[63][4] ), .ZN(n5049) );
  NAND4_X1 U8355 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5053)
         );
  OR4_X1 U8356 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n5057) );
  NAND2_X1 U8357 ( .A1(n5057), .A2(n25593), .ZN(n5058) );
  BUF_X1 U8358 ( .A(n14981), .Z(n20488) );
  AOI22_X1 U8359 ( .A1(n20488), .A2(\xmem_data[0][5] ), .B1(n20985), .B2(
        \xmem_data[1][5] ), .ZN(n5065) );
  AOI22_X1 U8360 ( .A1(n20769), .A2(\xmem_data[2][5] ), .B1(n30588), .B2(
        \xmem_data[3][5] ), .ZN(n5064) );
  BUF_X1 U8361 ( .A(n28947), .Z(n20489) );
  AOI22_X1 U8362 ( .A1(n20489), .A2(\xmem_data[4][5] ), .B1(n3318), .B2(
        \xmem_data[5][5] ), .ZN(n5063) );
  AND2_X1 U8363 ( .A1(n25360), .A2(\xmem_data[6][5] ), .ZN(n5061) );
  AOI21_X1 U8364 ( .B1(n28318), .B2(\xmem_data[7][5] ), .A(n5061), .ZN(n5062)
         );
  NAND4_X1 U8365 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5089)
         );
  AOI22_X1 U8366 ( .A1(n28493), .A2(\xmem_data[27][5] ), .B1(
        \xmem_data[26][5] ), .B2(n13481), .ZN(n5066) );
  INV_X1 U8367 ( .A(n5066), .ZN(n5071) );
  BUF_X1 U8368 ( .A(n14882), .Z(n20506) );
  AOI22_X1 U8369 ( .A1(n24222), .A2(\xmem_data[28][5] ), .B1(n3337), .B2(
        \xmem_data[29][5] ), .ZN(n5069) );
  BUF_X1 U8370 ( .A(n14912), .Z(n20505) );
  AOI22_X1 U8371 ( .A1(n20505), .A2(\xmem_data[24][5] ), .B1(n23802), .B2(
        \xmem_data[25][5] ), .ZN(n5068) );
  BUF_X1 U8372 ( .A(n14914), .Z(n20507) );
  AOI22_X1 U8373 ( .A1(n20507), .A2(\xmem_data[30][5] ), .B1(n20552), .B2(
        \xmem_data[31][5] ), .ZN(n5067) );
  NOR2_X1 U8374 ( .A1(n5071), .A2(n5070), .ZN(n5087) );
  AOI22_X1 U8375 ( .A1(n20806), .A2(\xmem_data[12][5] ), .B1(n21074), .B2(
        \xmem_data[13][5] ), .ZN(n5072) );
  INV_X1 U8376 ( .A(n5072), .ZN(n5076) );
  AOI22_X1 U8377 ( .A1(n20500), .A2(\xmem_data[10][5] ), .B1(n20994), .B2(
        \xmem_data[11][5] ), .ZN(n5074) );
  NAND2_X1 U8378 ( .A1(n20809), .A2(\xmem_data[15][5] ), .ZN(n5073) );
  NAND2_X1 U8379 ( .A1(n5074), .A2(n5073), .ZN(n5075) );
  NOR2_X1 U8380 ( .A1(n5076), .A2(n5075), .ZN(n5086) );
  AOI22_X1 U8381 ( .A1(n3222), .A2(\xmem_data[8][5] ), .B1(n29627), .B2(
        \xmem_data[9][5] ), .ZN(n5085) );
  AOI22_X1 U8382 ( .A1(n29188), .A2(\xmem_data[22][5] ), .B1(n24593), .B2(
        \xmem_data[23][5] ), .ZN(n5077) );
  INV_X1 U8383 ( .A(n5077), .ZN(n5083) );
  AOI22_X1 U8384 ( .A1(n25606), .A2(\xmem_data[20][5] ), .B1(n30892), .B2(
        \xmem_data[21][5] ), .ZN(n5079) );
  BUF_X1 U8385 ( .A(n10977), .Z(n20495) );
  AOI22_X1 U8386 ( .A1(n24555), .A2(\xmem_data[18][5] ), .B1(n27537), .B2(
        \xmem_data[19][5] ), .ZN(n5078) );
  NAND2_X1 U8387 ( .A1(n5079), .A2(n5078), .ZN(n5082) );
  AOI22_X1 U8388 ( .A1(n30854), .A2(\xmem_data[16][5] ), .B1(n25424), .B2(
        \xmem_data[17][5] ), .ZN(n5080) );
  INV_X1 U8389 ( .A(n5080), .ZN(n5081) );
  NOR3_X1 U8390 ( .A1(n5083), .A2(n5082), .A3(n5081), .ZN(n5084) );
  NAND4_X1 U8391 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5088)
         );
  AOI21_X1 U8392 ( .B1(n5090), .B2(n6990), .A(n10589), .ZN(n5091) );
  INV_X1 U8393 ( .A(n5091), .ZN(n5092) );
  AOI22_X1 U8394 ( .A1(n37191), .A2(n5092), .B1(n5091), .B2(n4499), .ZN(n5159)
         );
  NAND2_X1 U8395 ( .A1(load_xaddr_val[5]), .A2(n5092), .ZN(n5093) );
  XOR2_X1 U8396 ( .A(n39040), .B(n5093), .Z(n5136) );
  NOR2_X1 U8397 ( .A1(n5159), .A2(n5136), .ZN(n20515) );
  OAI21_X1 U8398 ( .B1(n3967), .B2(n3499), .A(n20515), .ZN(n5164) );
  BUF_X1 U8399 ( .A(n13420), .Z(n20567) );
  AOI22_X1 U8400 ( .A1(n20488), .A2(\xmem_data[96][5] ), .B1(n20567), .B2(
        \xmem_data[97][5] ), .ZN(n5097) );
  AOI22_X1 U8401 ( .A1(n24524), .A2(\xmem_data[98][5] ), .B1(n20827), .B2(
        \xmem_data[99][5] ), .ZN(n5096) );
  AOI22_X1 U8402 ( .A1(n22752), .A2(\xmem_data[100][5] ), .B1(n28718), .B2(
        \xmem_data[101][5] ), .ZN(n5095) );
  BUF_X1 U8403 ( .A(n13468), .Z(n20568) );
  AOI22_X1 U8404 ( .A1(n20568), .A2(\xmem_data[102][5] ), .B1(n24694), .B2(
        \xmem_data[103][5] ), .ZN(n5094) );
  NAND4_X1 U8405 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n5113)
         );
  AOI22_X1 U8406 ( .A1(n3222), .A2(\xmem_data[104][5] ), .B1(n24696), .B2(
        \xmem_data[105][5] ), .ZN(n5101) );
  BUF_X1 U8407 ( .A(n14989), .Z(n20558) );
  AOI22_X1 U8408 ( .A1(n20558), .A2(\xmem_data[106][5] ), .B1(n3340), .B2(
        \xmem_data[107][5] ), .ZN(n5100) );
  BUF_X1 U8409 ( .A(n14927), .Z(n20559) );
  AOI22_X1 U8410 ( .A1(n20559), .A2(\xmem_data[108][5] ), .B1(n27905), .B2(
        \xmem_data[109][5] ), .ZN(n5099) );
  AOI22_X1 U8411 ( .A1(n25450), .A2(\xmem_data[110][5] ), .B1(n24554), .B2(
        \xmem_data[111][5] ), .ZN(n5098) );
  NAND4_X1 U8412 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n5112)
         );
  BUF_X1 U8413 ( .A(n14997), .Z(n20545) );
  AOI22_X1 U8414 ( .A1(n20546), .A2(\xmem_data[112][5] ), .B1(n20545), .B2(
        \xmem_data[113][5] ), .ZN(n5105) );
  BUF_X1 U8415 ( .A(n10977), .Z(n20541) );
  AOI22_X1 U8416 ( .A1(n24516), .A2(\xmem_data[114][5] ), .B1(n25710), .B2(
        \xmem_data[115][5] ), .ZN(n5104) );
  BUF_X1 U8417 ( .A(n14898), .Z(n20544) );
  AOI22_X1 U8418 ( .A1(n20544), .A2(\xmem_data[116][5] ), .B1(n29770), .B2(
        \xmem_data[117][5] ), .ZN(n5103) );
  BUF_X1 U8419 ( .A(n13149), .Z(n20542) );
  AOI22_X1 U8420 ( .A1(n20543), .A2(\xmem_data[118][5] ), .B1(n20542), .B2(
        \xmem_data[119][5] ), .ZN(n5102) );
  NAND4_X1 U8421 ( .A1(n5105), .A2(n5104), .A3(n5103), .A4(n5102), .ZN(n5111)
         );
  AOI22_X1 U8422 ( .A1(n24219), .A2(\xmem_data[120][5] ), .B1(n23722), .B2(
        \xmem_data[121][5] ), .ZN(n5109) );
  AOI22_X1 U8423 ( .A1(n31254), .A2(\xmem_data[122][5] ), .B1(n29100), .B2(
        \xmem_data[123][5] ), .ZN(n5108) );
  BUF_X1 U8424 ( .A(n14973), .Z(n20551) );
  AOI22_X1 U8425 ( .A1(n20551), .A2(\xmem_data[124][5] ), .B1(n3269), .B2(
        \xmem_data[125][5] ), .ZN(n5107) );
  BUF_X1 U8426 ( .A(n14883), .Z(n20553) );
  BUF_X1 U8427 ( .A(n13486), .Z(n20552) );
  AOI22_X1 U8428 ( .A1(n20553), .A2(\xmem_data[126][5] ), .B1(n20552), .B2(
        \xmem_data[127][5] ), .ZN(n5106) );
  NAND4_X1 U8429 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5110)
         );
  OR4_X1 U8430 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n5138) );
  AND2_X1 U8431 ( .A1(n5159), .A2(n5136), .ZN(n20538) );
  BUF_X1 U8432 ( .A(n13127), .Z(n20577) );
  AND2_X1 U8433 ( .A1(n25359), .A2(\xmem_data[64][5] ), .ZN(n5114) );
  AOI21_X1 U8434 ( .B1(n20577), .B2(\xmem_data[65][5] ), .A(n5114), .ZN(n5119)
         );
  BUF_X1 U8435 ( .A(n13487), .Z(n20579) );
  AOI22_X1 U8436 ( .A1(n20579), .A2(\xmem_data[66][5] ), .B1(n27436), .B2(
        \xmem_data[67][5] ), .ZN(n5118) );
  BUF_X1 U8437 ( .A(n28974), .Z(n20578) );
  AOI22_X1 U8438 ( .A1(n20578), .A2(\xmem_data[68][5] ), .B1(n24693), .B2(
        \xmem_data[69][5] ), .ZN(n5117) );
  BUF_X1 U8439 ( .A(n29064), .Z(n20518) );
  AND2_X1 U8440 ( .A1(n25360), .A2(\xmem_data[70][5] ), .ZN(n5115) );
  AOI21_X1 U8441 ( .B1(n20518), .B2(\xmem_data[71][5] ), .A(n5115), .ZN(n5116)
         );
  NAND4_X1 U8442 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n5116), .ZN(n5135)
         );
  BUF_X1 U8443 ( .A(n10999), .Z(n20588) );
  BUF_X1 U8444 ( .A(n14997), .Z(n20587) );
  AOI22_X1 U8445 ( .A1(n20588), .A2(\xmem_data[80][5] ), .B1(n20587), .B2(
        \xmem_data[81][5] ), .ZN(n5123) );
  AOI22_X1 U8446 ( .A1(n30552), .A2(\xmem_data[82][5] ), .B1(n28298), .B2(
        \xmem_data[83][5] ), .ZN(n5122) );
  BUF_X1 U8447 ( .A(n14935), .Z(n20584) );
  AOI22_X1 U8448 ( .A1(n20584), .A2(\xmem_data[84][5] ), .B1(n20776), .B2(
        \xmem_data[85][5] ), .ZN(n5121) );
  AOI22_X1 U8449 ( .A1(n20586), .A2(\xmem_data[86][5] ), .B1(n20585), .B2(
        \xmem_data[87][5] ), .ZN(n5120) );
  NAND4_X1 U8450 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n5134)
         );
  AOI22_X1 U8451 ( .A1(n29316), .A2(\xmem_data[88][5] ), .B1(n23802), .B2(
        \xmem_data[89][5] ), .ZN(n5127) );
  AOI22_X1 U8452 ( .A1(n25367), .A2(\xmem_data[90][5] ), .B1(n17002), .B2(
        \xmem_data[91][5] ), .ZN(n5126) );
  AOI22_X1 U8453 ( .A1(n20551), .A2(\xmem_data[92][5] ), .B1(n20950), .B2(
        \xmem_data[93][5] ), .ZN(n5125) );
  AOI22_X1 U8454 ( .A1(n28098), .A2(\xmem_data[94][5] ), .B1(n29325), .B2(
        \xmem_data[95][5] ), .ZN(n5124) );
  NAND4_X1 U8455 ( .A1(n5127), .A2(n5126), .A3(n5125), .A4(n5124), .ZN(n5133)
         );
  AOI22_X1 U8456 ( .A1(n3217), .A2(\xmem_data[72][5] ), .B1(n20805), .B2(
        \xmem_data[73][5] ), .ZN(n5131) );
  BUF_X1 U8457 ( .A(n13469), .Z(n20598) );
  AOI22_X1 U8458 ( .A1(n20598), .A2(\xmem_data[74][5] ), .B1(n24534), .B2(
        \xmem_data[75][5] ), .ZN(n5130) );
  AOI22_X1 U8459 ( .A1(n29104), .A2(\xmem_data[76][5] ), .B1(n28308), .B2(
        \xmem_data[77][5] ), .ZN(n5129) );
  AOI22_X1 U8460 ( .A1(n27446), .A2(\xmem_data[78][5] ), .B1(n31321), .B2(
        \xmem_data[79][5] ), .ZN(n5128) );
  NAND4_X1 U8461 ( .A1(n5131), .A2(n5130), .A3(n5129), .A4(n5128), .ZN(n5132)
         );
  OR4_X1 U8462 ( .A1(n5135), .A2(n5134), .A3(n5133), .A4(n5132), .ZN(n5137) );
  INV_X1 U8463 ( .A(n5136), .ZN(n5160) );
  NOR2_X1 U8464 ( .A1(n5159), .A2(n5160), .ZN(n20573) );
  AOI22_X1 U8465 ( .A1(n5138), .A2(n20538), .B1(n5137), .B2(n20573), .ZN(n5163) );
  AOI22_X1 U8466 ( .A1(n25406), .A2(\xmem_data[32][5] ), .B1(n20577), .B2(
        \xmem_data[33][5] ), .ZN(n5142) );
  AOI22_X1 U8467 ( .A1(n20579), .A2(\xmem_data[34][5] ), .B1(n21061), .B2(
        \xmem_data[35][5] ), .ZN(n5141) );
  AOI22_X1 U8468 ( .A1(n20578), .A2(\xmem_data[36][5] ), .B1(n28245), .B2(
        \xmem_data[37][5] ), .ZN(n5140) );
  BUF_X1 U8469 ( .A(n29064), .Z(n20576) );
  AOI22_X1 U8470 ( .A1(n28501), .A2(\xmem_data[38][5] ), .B1(n20576), .B2(
        \xmem_data[39][5] ), .ZN(n5139) );
  NAND4_X1 U8471 ( .A1(n5142), .A2(n5141), .A3(n5140), .A4(n5139), .ZN(n5158)
         );
  AOI22_X1 U8472 ( .A1(n3221), .A2(\xmem_data[40][5] ), .B1(n27708), .B2(
        \xmem_data[41][5] ), .ZN(n5146) );
  AOI22_X1 U8473 ( .A1(n20598), .A2(\xmem_data[42][5] ), .B1(n20807), .B2(
        \xmem_data[43][5] ), .ZN(n5145) );
  AOI22_X1 U8474 ( .A1(n31275), .A2(\xmem_data[44][5] ), .B1(n29567), .B2(
        \xmem_data[45][5] ), .ZN(n5144) );
  AOI22_X1 U8475 ( .A1(n25450), .A2(\xmem_data[46][5] ), .B1(n27910), .B2(
        \xmem_data[47][5] ), .ZN(n5143) );
  NAND4_X1 U8476 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n5157)
         );
  AOI22_X1 U8477 ( .A1(n20588), .A2(\xmem_data[48][5] ), .B1(n20587), .B2(
        \xmem_data[49][5] ), .ZN(n5150) );
  AOI22_X1 U8478 ( .A1(n22740), .A2(\xmem_data[50][5] ), .B1(n17041), .B2(
        \xmem_data[51][5] ), .ZN(n5149) );
  AOI22_X1 U8479 ( .A1(n20584), .A2(\xmem_data[52][5] ), .B1(n29237), .B2(
        \xmem_data[53][5] ), .ZN(n5148) );
  AOI22_X1 U8480 ( .A1(n20586), .A2(\xmem_data[54][5] ), .B1(n20585), .B2(
        \xmem_data[55][5] ), .ZN(n5147) );
  NAND4_X1 U8481 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n5156)
         );
  AOI22_X1 U8482 ( .A1(n31270), .A2(\xmem_data[56][5] ), .B1(n29239), .B2(
        \xmem_data[57][5] ), .ZN(n5154) );
  AOI22_X1 U8483 ( .A1(n27460), .A2(\xmem_data[58][5] ), .B1(n20593), .B2(
        \xmem_data[59][5] ), .ZN(n5153) );
  AOI22_X1 U8484 ( .A1(n21051), .A2(\xmem_data[60][5] ), .B1(n29816), .B2(
        \xmem_data[61][5] ), .ZN(n5152) );
  AOI22_X1 U8485 ( .A1(n31314), .A2(\xmem_data[62][5] ), .B1(n31316), .B2(
        \xmem_data[63][5] ), .ZN(n5151) );
  NAND4_X1 U8486 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n5155)
         );
  OR4_X1 U8487 ( .A1(n5158), .A2(n5157), .A3(n5156), .A4(n5155), .ZN(n5161) );
  NAND2_X1 U8488 ( .A1(n5161), .A2(n20606), .ZN(n5162) );
  NAND3_X1 U8489 ( .A1(n5164), .A2(n5163), .A3(n5162), .ZN(n31882) );
  XNOR2_X1 U8490 ( .A(n31882), .B(\fmem_data[21][7] ), .ZN(n31661) );
  AOI22_X1 U8491 ( .A1(n20488), .A2(\xmem_data[0][4] ), .B1(n25628), .B2(
        \xmem_data[1][4] ), .ZN(n5165) );
  INV_X1 U8492 ( .A(n5165), .ZN(n5180) );
  NAND2_X1 U8493 ( .A1(n25450), .A2(\xmem_data[14][4] ), .ZN(n5166) );
  AOI22_X1 U8494 ( .A1(n25581), .A2(\xmem_data[28][4] ), .B1(n3301), .B2(
        \xmem_data[29][4] ), .ZN(n5168) );
  AOI22_X1 U8495 ( .A1(n30542), .A2(\xmem_data[22][4] ), .B1(n25434), .B2(
        \xmem_data[23][4] ), .ZN(n5167) );
  AOI22_X1 U8496 ( .A1(n29104), .A2(\xmem_data[12][4] ), .B1(n22668), .B2(
        \xmem_data[13][4] ), .ZN(n5169) );
  INV_X1 U8497 ( .A(n5169), .ZN(n5170) );
  AOI21_X1 U8498 ( .B1(\xmem_data[7][4] ), .B2(n20576), .A(n5170), .ZN(n5177)
         );
  AOI22_X1 U8499 ( .A1(n22701), .A2(\xmem_data[16][4] ), .B1(n25457), .B2(
        \xmem_data[17][4] ), .ZN(n5176) );
  AOI22_X1 U8500 ( .A1(n29271), .A2(\xmem_data[20][4] ), .B1(n27945), .B2(
        \xmem_data[21][4] ), .ZN(n5175) );
  AOI22_X1 U8501 ( .A1(n20507), .A2(\xmem_data[30][4] ), .B1(n27847), .B2(
        \xmem_data[31][4] ), .ZN(n5171) );
  INV_X1 U8502 ( .A(n5171), .ZN(n5173) );
  AND2_X1 U8503 ( .A1(n31347), .A2(\xmem_data[6][4] ), .ZN(n5172) );
  NOR2_X1 U8504 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  NAND4_X1 U8505 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n5178)
         );
  NOR3_X1 U8506 ( .A1(n5180), .A2(n5179), .A3(n5178), .ZN(n5196) );
  AOI22_X1 U8507 ( .A1(n3222), .A2(\xmem_data[8][4] ), .B1(n30964), .B2(
        \xmem_data[9][4] ), .ZN(n5181) );
  INV_X1 U8508 ( .A(n5181), .ZN(n5185) );
  AOI22_X1 U8509 ( .A1(n20500), .A2(\xmem_data[10][4] ), .B1(n28083), .B2(
        \xmem_data[11][4] ), .ZN(n5182) );
  INV_X1 U8510 ( .A(n5182), .ZN(n5184) );
  AND2_X1 U8511 ( .A1(n28050), .A2(\xmem_data[15][4] ), .ZN(n5183) );
  NOR3_X1 U8512 ( .A1(n5185), .A2(n5184), .A3(n5183), .ZN(n5194) );
  AOI22_X1 U8513 ( .A1(n13481), .A2(\xmem_data[26][4] ), .B1(n30956), .B2(
        \xmem_data[27][4] ), .ZN(n5186) );
  INV_X1 U8514 ( .A(n5186), .ZN(n5191) );
  AOI22_X1 U8515 ( .A1(n24159), .A2(\xmem_data[18][4] ), .B1(n20541), .B2(
        \xmem_data[19][4] ), .ZN(n5189) );
  AOI22_X1 U8516 ( .A1(n28329), .A2(\xmem_data[2][4] ), .B1(n21061), .B2(
        \xmem_data[3][4] ), .ZN(n5188) );
  AOI22_X1 U8517 ( .A1(n20505), .A2(\xmem_data[24][4] ), .B1(n22682), .B2(
        \xmem_data[25][4] ), .ZN(n5187) );
  NOR2_X1 U8518 ( .A1(n5191), .A2(n5190), .ZN(n5193) );
  AOI22_X1 U8519 ( .A1(n20489), .A2(\xmem_data[4][4] ), .B1(n28718), .B2(
        \xmem_data[5][4] ), .ZN(n5192) );
  AND3_X1 U8520 ( .A1(n5194), .A2(n5193), .A3(n5192), .ZN(n5195) );
  AOI21_X1 U8521 ( .B1(n5196), .B2(n5195), .A(n3232), .ZN(n5197) );
  INV_X1 U8522 ( .A(n5197), .ZN(n5265) );
  AOI22_X1 U8523 ( .A1(n28292), .A2(\xmem_data[32][4] ), .B1(n20577), .B2(
        \xmem_data[33][4] ), .ZN(n5202) );
  AOI22_X1 U8524 ( .A1(n20579), .A2(\xmem_data[34][4] ), .B1(n28076), .B2(
        \xmem_data[35][4] ), .ZN(n5201) );
  AOI22_X1 U8525 ( .A1(n20578), .A2(\xmem_data[36][4] ), .B1(n3153), .B2(
        \xmem_data[37][4] ), .ZN(n5200) );
  AND2_X1 U8526 ( .A1(n24439), .A2(\xmem_data[38][4] ), .ZN(n5198) );
  AOI21_X1 U8527 ( .B1(n28044), .B2(\xmem_data[39][4] ), .A(n5198), .ZN(n5199)
         );
  NAND4_X1 U8528 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n5219)
         );
  AOI22_X1 U8529 ( .A1(n25398), .A2(\xmem_data[56][4] ), .B1(n28754), .B2(
        \xmem_data[57][4] ), .ZN(n5206) );
  AOI22_X1 U8530 ( .A1(n29238), .A2(\xmem_data[58][4] ), .B1(n25717), .B2(
        \xmem_data[59][4] ), .ZN(n5205) );
  AOI22_X1 U8531 ( .A1(n27856), .A2(\xmem_data[60][4] ), .B1(n3300), .B2(
        \xmem_data[61][4] ), .ZN(n5204) );
  AOI22_X1 U8532 ( .A1(n27525), .A2(\xmem_data[62][4] ), .B1(n24572), .B2(
        \xmem_data[63][4] ), .ZN(n5203) );
  NAND4_X1 U8533 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n5217)
         );
  AOI22_X1 U8534 ( .A1(n20588), .A2(\xmem_data[48][4] ), .B1(n20587), .B2(
        \xmem_data[49][4] ), .ZN(n5210) );
  AOI22_X1 U8535 ( .A1(n17012), .A2(\xmem_data[50][4] ), .B1(n28980), .B2(
        \xmem_data[51][4] ), .ZN(n5209) );
  AOI22_X1 U8536 ( .A1(n20584), .A2(\xmem_data[52][4] ), .B1(n28154), .B2(
        \xmem_data[53][4] ), .ZN(n5208) );
  AOI22_X1 U8537 ( .A1(n20586), .A2(\xmem_data[54][4] ), .B1(n20585), .B2(
        \xmem_data[55][4] ), .ZN(n5207) );
  NAND4_X1 U8538 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n5216)
         );
  AOI22_X1 U8539 ( .A1(n3219), .A2(\xmem_data[40][4] ), .B1(n28733), .B2(
        \xmem_data[41][4] ), .ZN(n5214) );
  AOI22_X1 U8540 ( .A1(n20598), .A2(\xmem_data[42][4] ), .B1(n28475), .B2(
        \xmem_data[43][4] ), .ZN(n5213) );
  AOI22_X1 U8541 ( .A1(n13444), .A2(\xmem_data[44][4] ), .B1(n25451), .B2(
        \xmem_data[45][4] ), .ZN(n5212) );
  AOI22_X1 U8542 ( .A1(n25450), .A2(\xmem_data[46][4] ), .B1(n24450), .B2(
        \xmem_data[47][4] ), .ZN(n5211) );
  NAND4_X1 U8543 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n5215)
         );
  OR3_X1 U8544 ( .A1(n5217), .A2(n5216), .A3(n5215), .ZN(n5218) );
  OAI21_X1 U8545 ( .B1(n5219), .B2(n5218), .A(n20606), .ZN(n5264) );
  AOI22_X1 U8546 ( .A1(n20488), .A2(\xmem_data[96][4] ), .B1(n20567), .B2(
        \xmem_data[97][4] ), .ZN(n5223) );
  AOI22_X1 U8547 ( .A1(n30498), .A2(\xmem_data[98][4] ), .B1(n17030), .B2(
        \xmem_data[99][4] ), .ZN(n5222) );
  AOI22_X1 U8548 ( .A1(n25357), .A2(\xmem_data[100][4] ), .B1(n23754), .B2(
        \xmem_data[101][4] ), .ZN(n5221) );
  AOI22_X1 U8549 ( .A1(n20568), .A2(\xmem_data[102][4] ), .B1(n20576), .B2(
        \xmem_data[103][4] ), .ZN(n5220) );
  NAND4_X1 U8550 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n5240)
         );
  AOI22_X1 U8551 ( .A1(n29048), .A2(\xmem_data[120][4] ), .B1(n30950), .B2(
        \xmem_data[121][4] ), .ZN(n5227) );
  AOI22_X1 U8552 ( .A1(n25435), .A2(\xmem_data[122][4] ), .B1(n3178), .B2(
        \xmem_data[123][4] ), .ZN(n5226) );
  AOI22_X1 U8553 ( .A1(n20551), .A2(\xmem_data[124][4] ), .B1(n30645), .B2(
        \xmem_data[125][4] ), .ZN(n5225) );
  AOI22_X1 U8554 ( .A1(n20553), .A2(\xmem_data[126][4] ), .B1(n20552), .B2(
        \xmem_data[127][4] ), .ZN(n5224) );
  NAND4_X1 U8555 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n5238)
         );
  AOI22_X1 U8556 ( .A1(n20546), .A2(\xmem_data[112][4] ), .B1(n20545), .B2(
        \xmem_data[113][4] ), .ZN(n5231) );
  AOI22_X1 U8557 ( .A1(n23761), .A2(\xmem_data[114][4] ), .B1(n30891), .B2(
        \xmem_data[115][4] ), .ZN(n5230) );
  AOI22_X1 U8558 ( .A1(n20544), .A2(\xmem_data[116][4] ), .B1(n28091), .B2(
        \xmem_data[117][4] ), .ZN(n5229) );
  AOI22_X1 U8559 ( .A1(n20543), .A2(\xmem_data[118][4] ), .B1(n20542), .B2(
        \xmem_data[119][4] ), .ZN(n5228) );
  NAND4_X1 U8560 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n5237)
         );
  AOI22_X1 U8561 ( .A1(n3218), .A2(\xmem_data[104][4] ), .B1(n29256), .B2(
        \xmem_data[105][4] ), .ZN(n5235) );
  AOI22_X1 U8562 ( .A1(n20558), .A2(\xmem_data[106][4] ), .B1(n24534), .B2(
        \xmem_data[107][4] ), .ZN(n5234) );
  AOI22_X1 U8563 ( .A1(n20559), .A2(\xmem_data[108][4] ), .B1(n24702), .B2(
        \xmem_data[109][4] ), .ZN(n5233) );
  AOI22_X1 U8564 ( .A1(n30877), .A2(\xmem_data[110][4] ), .B1(n30607), .B2(
        \xmem_data[111][4] ), .ZN(n5232) );
  NAND4_X1 U8565 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n5236)
         );
  OR3_X1 U8566 ( .A1(n5238), .A2(n5237), .A3(n5236), .ZN(n5239) );
  OAI21_X1 U8567 ( .B1(n5240), .B2(n5239), .A(n20538), .ZN(n5263) );
  AOI22_X1 U8568 ( .A1(n14981), .A2(\xmem_data[64][4] ), .B1(n20577), .B2(
        \xmem_data[65][4] ), .ZN(n5244) );
  AOI22_X1 U8569 ( .A1(n20579), .A2(\xmem_data[66][4] ), .B1(n29057), .B2(
        \xmem_data[67][4] ), .ZN(n5243) );
  AOI22_X1 U8570 ( .A1(n20578), .A2(\xmem_data[68][4] ), .B1(n30864), .B2(
        \xmem_data[69][4] ), .ZN(n5242) );
  AOI22_X1 U8571 ( .A1(n29253), .A2(\xmem_data[70][4] ), .B1(n27439), .B2(
        \xmem_data[71][4] ), .ZN(n5241) );
  NAND4_X1 U8572 ( .A1(n5244), .A2(n5243), .A3(n5242), .A4(n5241), .ZN(n5261)
         );
  AOI22_X1 U8573 ( .A1(n20588), .A2(\xmem_data[80][4] ), .B1(n20587), .B2(
        \xmem_data[81][4] ), .ZN(n5248) );
  AOI22_X1 U8574 ( .A1(n29232), .A2(\xmem_data[82][4] ), .B1(n27537), .B2(
        \xmem_data[83][4] ), .ZN(n5247) );
  AOI22_X1 U8575 ( .A1(n20584), .A2(\xmem_data[84][4] ), .B1(n30543), .B2(
        \xmem_data[85][4] ), .ZN(n5246) );
  AOI22_X1 U8576 ( .A1(n20586), .A2(\xmem_data[86][4] ), .B1(n20585), .B2(
        \xmem_data[87][4] ), .ZN(n5245) );
  NAND4_X1 U8577 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n5259)
         );
  AOI22_X1 U8578 ( .A1(n16989), .A2(\xmem_data[88][4] ), .B1(n29410), .B2(
        \xmem_data[89][4] ), .ZN(n5252) );
  AOI22_X1 U8579 ( .A1(n28097), .A2(\xmem_data[90][4] ), .B1(n24548), .B2(
        \xmem_data[91][4] ), .ZN(n5251) );
  AOI22_X1 U8580 ( .A1(n28462), .A2(\xmem_data[92][4] ), .B1(n30686), .B2(
        \xmem_data[93][4] ), .ZN(n5250) );
  AOI22_X1 U8581 ( .A1(n27365), .A2(\xmem_data[94][4] ), .B1(n24685), .B2(
        \xmem_data[95][4] ), .ZN(n5249) );
  NAND4_X1 U8582 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n5258)
         );
  AOI22_X1 U8583 ( .A1(n3222), .A2(\xmem_data[72][4] ), .B1(n30593), .B2(
        \xmem_data[73][4] ), .ZN(n5256) );
  AOI22_X1 U8584 ( .A1(n20598), .A2(\xmem_data[74][4] ), .B1(n3340), .B2(
        \xmem_data[75][4] ), .ZN(n5255) );
  AOI22_X1 U8585 ( .A1(n28509), .A2(\xmem_data[76][4] ), .B1(n28344), .B2(
        \xmem_data[77][4] ), .ZN(n5254) );
  AOI22_X1 U8586 ( .A1(n25514), .A2(\xmem_data[78][4] ), .B1(n25707), .B2(
        \xmem_data[79][4] ), .ZN(n5253) );
  NAND4_X1 U8587 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n5257)
         );
  OR3_X1 U8588 ( .A1(n5259), .A2(n5258), .A3(n5257), .ZN(n5260) );
  OAI21_X1 U8589 ( .B1(n5261), .B2(n5260), .A(n20573), .ZN(n5262) );
  XNOR2_X1 U8590 ( .A(n31489), .B(\fmem_data[21][7] ), .ZN(n25747) );
  XOR2_X1 U8591 ( .A(\fmem_data[21][6] ), .B(\fmem_data[21][7] ), .Z(n5266) );
  OAI22_X1 U8592 ( .A1(n31661), .A2(n35508), .B1(n25747), .B2(n35507), .ZN(
        n35093) );
  AOI22_X1 U8593 ( .A1(n20993), .A2(\xmem_data[96][5] ), .B1(n3140), .B2(
        \xmem_data[97][5] ), .ZN(n5270) );
  BUF_X1 U8594 ( .A(n25604), .Z(n28972) );
  AOI22_X1 U8595 ( .A1(n25450), .A2(\xmem_data[98][5] ), .B1(n28972), .B2(
        \xmem_data[99][5] ), .ZN(n5269) );
  AOI22_X1 U8596 ( .A1(n3358), .A2(\xmem_data[100][5] ), .B1(n20799), .B2(
        \xmem_data[101][5] ), .ZN(n5268) );
  AOI22_X1 U8597 ( .A1(n21075), .A2(\xmem_data[102][5] ), .B1(n20541), .B2(
        \xmem_data[103][5] ), .ZN(n5267) );
  NAND4_X1 U8598 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n5286)
         );
  BUF_X1 U8599 ( .A(n14935), .Z(n29009) );
  BUF_X1 U8600 ( .A(n3464), .Z(n29008) );
  AOI22_X1 U8601 ( .A1(n29009), .A2(\xmem_data[104][5] ), .B1(n29008), .B2(
        \xmem_data[105][5] ), .ZN(n5274) );
  BUF_X1 U8602 ( .A(n14937), .Z(n29010) );
  AOI22_X1 U8603 ( .A1(n3212), .A2(\xmem_data[106][5] ), .B1(n29010), .B2(
        \xmem_data[107][5] ), .ZN(n5273) );
  BUF_X1 U8604 ( .A(n14971), .Z(n29012) );
  AOI22_X1 U8605 ( .A1(n17043), .A2(\xmem_data[108][5] ), .B1(n29012), .B2(
        \xmem_data[109][5] ), .ZN(n5272) );
  AOI22_X1 U8606 ( .A1(n29238), .A2(\xmem_data[110][5] ), .B1(n28428), .B2(
        \xmem_data[111][5] ), .ZN(n5271) );
  NAND4_X1 U8607 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n5285)
         );
  BUF_X1 U8608 ( .A(n14974), .Z(n28955) );
  AOI22_X1 U8609 ( .A1(n25581), .A2(\xmem_data[112][5] ), .B1(n28955), .B2(
        \xmem_data[113][5] ), .ZN(n5278) );
  AOI22_X1 U8610 ( .A1(n28098), .A2(\xmem_data[114][5] ), .B1(n20782), .B2(
        \xmem_data[115][5] ), .ZN(n5277) );
  BUF_X1 U8611 ( .A(n14981), .Z(n29017) );
  AOI22_X1 U8612 ( .A1(n29017), .A2(\xmem_data[116][5] ), .B1(n31308), .B2(
        \xmem_data[117][5] ), .ZN(n5276) );
  AOI22_X1 U8613 ( .A1(n31344), .A2(\xmem_data[118][5] ), .B1(n21061), .B2(
        \xmem_data[119][5] ), .ZN(n5275) );
  NAND4_X1 U8614 ( .A1(n5278), .A2(n5277), .A3(n5276), .A4(n5275), .ZN(n5284)
         );
  BUF_X1 U8615 ( .A(n28974), .Z(n12471) );
  AOI22_X1 U8616 ( .A1(n12471), .A2(\xmem_data[120][5] ), .B1(n30864), .B2(
        \xmem_data[121][5] ), .ZN(n5282) );
  AOI22_X1 U8617 ( .A1(n25360), .A2(\xmem_data[122][5] ), .B1(n29064), .B2(
        \xmem_data[123][5] ), .ZN(n5281) );
  BUF_X1 U8618 ( .A(n14988), .Z(n29026) );
  AOI22_X1 U8619 ( .A1(n3217), .A2(\xmem_data[124][5] ), .B1(n29026), .B2(
        \xmem_data[125][5] ), .ZN(n5280) );
  BUF_X1 U8620 ( .A(n14989), .Z(n29028) );
  BUF_X1 U8621 ( .A(n14990), .Z(n29027) );
  AOI22_X1 U8622 ( .A1(n29028), .A2(\xmem_data[126][5] ), .B1(n29027), .B2(
        \xmem_data[127][5] ), .ZN(n5279) );
  NAND4_X1 U8623 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n5283)
         );
  OR4_X1 U8624 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n5312) );
  INV_X1 U8625 ( .A(n10589), .ZN(n13432) );
  AOI21_X1 U8626 ( .B1(n13132), .B2(n39035), .A(n13432), .ZN(n5288) );
  INV_X1 U8627 ( .A(n5288), .ZN(n5287) );
  AOI22_X1 U8628 ( .A1(n37191), .A2(n5288), .B1(n5287), .B2(n4499), .ZN(n5360)
         );
  AND2_X1 U8629 ( .A1(n5360), .A2(n5359), .ZN(n28968) );
  BUF_X1 U8630 ( .A(n14973), .Z(n29055) );
  BUF_X1 U8631 ( .A(n14974), .Z(n29054) );
  AOI22_X1 U8632 ( .A1(n29055), .A2(\xmem_data[80][5] ), .B1(n29054), .B2(
        \xmem_data[81][5] ), .ZN(n5294) );
  AOI22_X1 U8633 ( .A1(n20949), .A2(\xmem_data[82][5] ), .B1(n24685), .B2(
        \xmem_data[83][5] ), .ZN(n5293) );
  AND2_X1 U8634 ( .A1(n25527), .A2(\xmem_data[84][5] ), .ZN(n5290) );
  AOI21_X1 U8635 ( .B1(n29657), .B2(\xmem_data[85][5] ), .A(n5290), .ZN(n5292)
         );
  BUF_X1 U8636 ( .A(n31263), .Z(n29057) );
  AOI22_X1 U8637 ( .A1(n16999), .A2(\xmem_data[86][5] ), .B1(n29057), .B2(
        \xmem_data[87][5] ), .ZN(n5291) );
  NAND4_X1 U8638 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n5310)
         );
  BUF_X1 U8639 ( .A(n14898), .Z(n29046) );
  AOI22_X1 U8640 ( .A1(n29046), .A2(\xmem_data[72][5] ), .B1(n24458), .B2(
        \xmem_data[73][5] ), .ZN(n5298) );
  AOI22_X1 U8641 ( .A1(n3212), .A2(\xmem_data[74][5] ), .B1(n24509), .B2(
        \xmem_data[75][5] ), .ZN(n5297) );
  BUF_X1 U8642 ( .A(n14971), .Z(n29047) );
  AOI22_X1 U8643 ( .A1(n29048), .A2(\xmem_data[76][5] ), .B1(n29047), .B2(
        \xmem_data[77][5] ), .ZN(n5296) );
  BUF_X1 U8644 ( .A(n13481), .Z(n29049) );
  AOI22_X1 U8645 ( .A1(n29049), .A2(\xmem_data[78][5] ), .B1(n28428), .B2(
        \xmem_data[79][5] ), .ZN(n5295) );
  NAND4_X1 U8646 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n5309)
         );
  AOI22_X1 U8647 ( .A1(n12471), .A2(\xmem_data[88][5] ), .B1(n3382), .B2(
        \xmem_data[89][5] ), .ZN(n5302) );
  AOI22_X1 U8648 ( .A1(n31347), .A2(\xmem_data[90][5] ), .B1(n29064), .B2(
        \xmem_data[91][5] ), .ZN(n5301) );
  BUF_X1 U8649 ( .A(n14988), .Z(n29065) );
  AOI22_X1 U8650 ( .A1(n3219), .A2(\xmem_data[92][5] ), .B1(n29065), .B2(
        \xmem_data[93][5] ), .ZN(n5300) );
  AOI22_X1 U8651 ( .A1(n23739), .A2(\xmem_data[94][5] ), .B1(n25617), .B2(
        \xmem_data[95][5] ), .ZN(n5299) );
  NAND4_X1 U8652 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), .ZN(n5308)
         );
  BUF_X1 U8653 ( .A(n14991), .Z(n28952) );
  AOI22_X1 U8654 ( .A1(n13444), .A2(\xmem_data[64][5] ), .B1(n28952), .B2(
        \xmem_data[65][5] ), .ZN(n5306) );
  AOI22_X1 U8655 ( .A1(n28510), .A2(\xmem_data[66][5] ), .B1(n24638), .B2(
        \xmem_data[67][5] ), .ZN(n5305) );
  AOI22_X1 U8656 ( .A1(n22739), .A2(\xmem_data[68][5] ), .B1(n22738), .B2(
        \xmem_data[69][5] ), .ZN(n5304) );
  AOI22_X1 U8657 ( .A1(n13168), .A2(\xmem_data[70][5] ), .B1(n24131), .B2(
        \xmem_data[71][5] ), .ZN(n5303) );
  NAND4_X1 U8658 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), .ZN(n5307)
         );
  OR4_X1 U8659 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n5311) );
  INV_X1 U8660 ( .A(n5359), .ZN(n5336) );
  AOI22_X1 U8661 ( .A1(n5312), .A2(n28968), .B1(n5311), .B2(n29041), .ZN(n5364) );
  AOI22_X1 U8662 ( .A1(n22759), .A2(\xmem_data[32][5] ), .B1(n28952), .B2(
        \xmem_data[33][5] ), .ZN(n5316) );
  AOI22_X1 U8663 ( .A1(n28007), .A2(\xmem_data[34][5] ), .B1(n20809), .B2(
        \xmem_data[35][5] ), .ZN(n5315) );
  AOI22_X1 U8664 ( .A1(n13475), .A2(\xmem_data[36][5] ), .B1(n25708), .B2(
        \xmem_data[37][5] ), .ZN(n5314) );
  AOI22_X1 U8665 ( .A1(n28515), .A2(\xmem_data[38][5] ), .B1(n25425), .B2(
        \xmem_data[39][5] ), .ZN(n5313) );
  NAND4_X1 U8666 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n5335)
         );
  AOI22_X1 U8667 ( .A1(n29046), .A2(\xmem_data[40][5] ), .B1(n28154), .B2(
        \xmem_data[41][5] ), .ZN(n5320) );
  AOI22_X1 U8668 ( .A1(n25460), .A2(\xmem_data[42][5] ), .B1(n25573), .B2(
        \xmem_data[43][5] ), .ZN(n5319) );
  AOI22_X1 U8669 ( .A1(n29048), .A2(\xmem_data[44][5] ), .B1(n29047), .B2(
        \xmem_data[45][5] ), .ZN(n5318) );
  AOI22_X1 U8670 ( .A1(n29049), .A2(\xmem_data[46][5] ), .B1(n30899), .B2(
        \xmem_data[47][5] ), .ZN(n5317) );
  NAND4_X1 U8671 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n5334)
         );
  AOI22_X1 U8672 ( .A1(n25406), .A2(\xmem_data[52][5] ), .B1(n28241), .B2(
        \xmem_data[53][5] ), .ZN(n5327) );
  AOI22_X1 U8673 ( .A1(n10456), .A2(\xmem_data[54][5] ), .B1(n29057), .B2(
        \xmem_data[55][5] ), .ZN(n5322) );
  AOI22_X1 U8674 ( .A1(n20949), .A2(\xmem_data[50][5] ), .B1(n30525), .B2(
        \xmem_data[51][5] ), .ZN(n5321) );
  NAND2_X1 U8675 ( .A1(n5322), .A2(n5321), .ZN(n5325) );
  AOI22_X1 U8676 ( .A1(n29055), .A2(\xmem_data[48][5] ), .B1(n29054), .B2(
        \xmem_data[49][5] ), .ZN(n5323) );
  INV_X1 U8677 ( .A(n5323), .ZN(n5324) );
  NOR2_X1 U8678 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  NAND2_X1 U8679 ( .A1(n5327), .A2(n5326), .ZN(n5333) );
  BUF_X1 U8680 ( .A(n28974), .Z(n21309) );
  AOI22_X1 U8681 ( .A1(n21309), .A2(\xmem_data[56][5] ), .B1(n3412), .B2(
        \xmem_data[57][5] ), .ZN(n5331) );
  AOI22_X1 U8682 ( .A1(n29253), .A2(\xmem_data[58][5] ), .B1(n29064), .B2(
        \xmem_data[59][5] ), .ZN(n5330) );
  AOI22_X1 U8683 ( .A1(n3220), .A2(\xmem_data[60][5] ), .B1(n29065), .B2(
        \xmem_data[61][5] ), .ZN(n5329) );
  AOI22_X1 U8684 ( .A1(n31367), .A2(\xmem_data[62][5] ), .B1(n25416), .B2(
        \xmem_data[63][5] ), .ZN(n5328) );
  NAND4_X1 U8685 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .ZN(n5332)
         );
  OR4_X1 U8686 ( .A1(n5335), .A2(n5334), .A3(n5333), .A4(n5332), .ZN(n5337) );
  AND2_X1 U8687 ( .A1(n5336), .A2(n5360), .ZN(n29078) );
  NAND2_X1 U8688 ( .A1(n5337), .A2(n29078), .ZN(n5363) );
  AOI22_X1 U8689 ( .A1(n3256), .A2(\xmem_data[0][5] ), .B1(n3126), .B2(
        \xmem_data[1][5] ), .ZN(n5341) );
  AOI22_X1 U8690 ( .A1(n3231), .A2(\xmem_data[2][5] ), .B1(n28972), .B2(
        \xmem_data[3][5] ), .ZN(n5340) );
  AOI22_X1 U8691 ( .A1(n28373), .A2(\xmem_data[4][5] ), .B1(n29451), .B2(
        \xmem_data[5][5] ), .ZN(n5339) );
  AOI22_X1 U8692 ( .A1(n24448), .A2(\xmem_data[6][5] ), .B1(n30891), .B2(
        \xmem_data[7][5] ), .ZN(n5338) );
  NAND4_X1 U8693 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n5358)
         );
  AOI22_X1 U8694 ( .A1(n25671), .A2(\xmem_data[8][5] ), .B1(n20776), .B2(
        \xmem_data[9][5] ), .ZN(n5345) );
  BUF_X1 U8695 ( .A(n14936), .Z(n28993) );
  AOI22_X1 U8696 ( .A1(n28993), .A2(\xmem_data[10][5] ), .B1(n29317), .B2(
        \xmem_data[11][5] ), .ZN(n5344) );
  BUF_X1 U8697 ( .A(n14971), .Z(n28994) );
  AOI22_X1 U8698 ( .A1(n31329), .A2(\xmem_data[12][5] ), .B1(n28994), .B2(
        \xmem_data[13][5] ), .ZN(n5343) );
  AOI22_X1 U8699 ( .A1(n30515), .A2(\xmem_data[14][5] ), .B1(n28493), .B2(
        \xmem_data[15][5] ), .ZN(n5342) );
  NAND4_X1 U8700 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n5357)
         );
  AOI22_X1 U8701 ( .A1(n3372), .A2(\xmem_data[16][5] ), .B1(n30269), .B2(
        \xmem_data[17][5] ), .ZN(n5350) );
  BUF_X1 U8702 ( .A(n14914), .Z(n28983) );
  AOI22_X1 U8703 ( .A1(n28983), .A2(\xmem_data[18][5] ), .B1(n24606), .B2(
        \xmem_data[19][5] ), .ZN(n5349) );
  BUF_X1 U8704 ( .A(n14919), .Z(n28979) );
  AND2_X1 U8705 ( .A1(n28979), .A2(\xmem_data[20][5] ), .ZN(n5346) );
  AOI21_X1 U8706 ( .B1(n20567), .B2(\xmem_data[21][5] ), .A(n5346), .ZN(n5348)
         );
  AOI22_X1 U8707 ( .A1(n24122), .A2(\xmem_data[22][5] ), .B1(n30588), .B2(
        \xmem_data[23][5] ), .ZN(n5347) );
  NAND4_X1 U8708 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n5356)
         );
  BUF_X1 U8709 ( .A(n28973), .Z(n21308) );
  AOI22_X1 U8710 ( .A1(n12471), .A2(\xmem_data[24][5] ), .B1(n21308), .B2(
        \xmem_data[25][5] ), .ZN(n5354) );
  AOI22_X1 U8711 ( .A1(n25485), .A2(\xmem_data[26][5] ), .B1(n29064), .B2(
        \xmem_data[27][5] ), .ZN(n5353) );
  AOI22_X1 U8712 ( .A1(n3218), .A2(\xmem_data[28][5] ), .B1(n29494), .B2(
        \xmem_data[29][5] ), .ZN(n5352) );
  AOI22_X1 U8713 ( .A1(n20500), .A2(\xmem_data[30][5] ), .B1(n24565), .B2(
        \xmem_data[31][5] ), .ZN(n5351) );
  NAND4_X1 U8714 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n5355)
         );
  OR4_X1 U8715 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n5361) );
  NAND2_X1 U8716 ( .A1(n5361), .A2(n29002), .ZN(n5362) );
  AOI22_X1 U8717 ( .A1(n12471), .A2(\xmem_data[120][4] ), .B1(n21308), .B2(
        \xmem_data[121][4] ), .ZN(n5368) );
  AOI22_X1 U8718 ( .A1(n24439), .A2(\xmem_data[122][4] ), .B1(n28364), .B2(
        \xmem_data[123][4] ), .ZN(n5367) );
  AOI22_X1 U8719 ( .A1(n3220), .A2(\xmem_data[124][4] ), .B1(n29026), .B2(
        \xmem_data[125][4] ), .ZN(n5366) );
  AOI22_X1 U8720 ( .A1(n29028), .A2(\xmem_data[126][4] ), .B1(n29027), .B2(
        \xmem_data[127][4] ), .ZN(n5365) );
  NAND4_X1 U8721 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n5379)
         );
  AOI22_X1 U8722 ( .A1(n27994), .A2(\xmem_data[96][4] ), .B1(n28952), .B2(
        \xmem_data[97][4] ), .ZN(n5372) );
  AOI22_X1 U8723 ( .A1(n28007), .A2(\xmem_data[98][4] ), .B1(n27447), .B2(
        \xmem_data[99][4] ), .ZN(n5371) );
  AOI22_X1 U8724 ( .A1(n29307), .A2(\xmem_data[100][4] ), .B1(n27514), .B2(
        \xmem_data[101][4] ), .ZN(n5370) );
  AOI22_X1 U8725 ( .A1(n24159), .A2(\xmem_data[102][4] ), .B1(n20495), .B2(
        \xmem_data[103][4] ), .ZN(n5369) );
  NAND4_X1 U8726 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n5378)
         );
  AOI22_X1 U8727 ( .A1(n29009), .A2(\xmem_data[104][4] ), .B1(n29008), .B2(
        \xmem_data[105][4] ), .ZN(n5376) );
  AOI22_X1 U8728 ( .A1(n3213), .A2(\xmem_data[106][4] ), .B1(n29010), .B2(
        \xmem_data[107][4] ), .ZN(n5375) );
  AOI22_X1 U8729 ( .A1(n24459), .A2(\xmem_data[108][4] ), .B1(n29012), .B2(
        \xmem_data[109][4] ), .ZN(n5374) );
  AOI22_X1 U8730 ( .A1(n27523), .A2(\xmem_data[110][4] ), .B1(n17002), .B2(
        \xmem_data[111][4] ), .ZN(n5373) );
  NAND4_X1 U8731 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n5377)
         );
  AOI22_X1 U8732 ( .A1(n20506), .A2(\xmem_data[112][4] ), .B1(n28955), .B2(
        \xmem_data[113][4] ), .ZN(n5383) );
  AOI22_X1 U8733 ( .A1(n29245), .A2(\xmem_data[114][4] ), .B1(n24685), .B2(
        \xmem_data[115][4] ), .ZN(n5382) );
  AOI22_X1 U8734 ( .A1(n29017), .A2(\xmem_data[116][4] ), .B1(n30901), .B2(
        \xmem_data[117][4] ), .ZN(n5381) );
  AOI22_X1 U8735 ( .A1(n20769), .A2(\xmem_data[118][4] ), .B1(n28354), .B2(
        \xmem_data[119][4] ), .ZN(n5380) );
  NAND4_X1 U8736 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n5384)
         );
  AOI22_X1 U8737 ( .A1(n29055), .A2(\xmem_data[80][4] ), .B1(n29054), .B2(
        \xmem_data[81][4] ), .ZN(n5390) );
  AOI22_X1 U8738 ( .A1(n24622), .A2(\xmem_data[82][4] ), .B1(n3209), .B2(
        \xmem_data[83][4] ), .ZN(n5389) );
  AND2_X1 U8739 ( .A1(n29136), .A2(\xmem_data[84][4] ), .ZN(n5386) );
  AOI21_X1 U8740 ( .B1(n17051), .B2(\xmem_data[85][4] ), .A(n5386), .ZN(n5388)
         );
  AOI22_X1 U8741 ( .A1(n20707), .A2(\xmem_data[86][4] ), .B1(n29057), .B2(
        \xmem_data[87][4] ), .ZN(n5387) );
  NAND4_X1 U8742 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n5406)
         );
  AOI22_X1 U8743 ( .A1(n29046), .A2(\xmem_data[72][4] ), .B1(n17018), .B2(
        \xmem_data[73][4] ), .ZN(n5394) );
  AOI22_X1 U8744 ( .A1(n31269), .A2(\xmem_data[74][4] ), .B1(n24708), .B2(
        \xmem_data[75][4] ), .ZN(n5393) );
  AOI22_X1 U8745 ( .A1(n29048), .A2(\xmem_data[76][4] ), .B1(n29047), .B2(
        \xmem_data[77][4] ), .ZN(n5392) );
  AOI22_X1 U8746 ( .A1(n29049), .A2(\xmem_data[78][4] ), .B1(n24647), .B2(
        \xmem_data[79][4] ), .ZN(n5391) );
  NAND4_X1 U8747 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n5405)
         );
  AOI22_X1 U8748 ( .A1(n25629), .A2(\xmem_data[88][4] ), .B1(n3228), .B2(
        \xmem_data[89][4] ), .ZN(n5398) );
  AOI22_X1 U8749 ( .A1(n22753), .A2(\xmem_data[90][4] ), .B1(n29064), .B2(
        \xmem_data[91][4] ), .ZN(n5397) );
  AOI22_X1 U8750 ( .A1(n3219), .A2(\xmem_data[92][4] ), .B1(n29065), .B2(
        \xmem_data[93][4] ), .ZN(n5396) );
  AOI22_X1 U8751 ( .A1(n23739), .A2(\xmem_data[94][4] ), .B1(n20994), .B2(
        \xmem_data[95][4] ), .ZN(n5395) );
  NAND4_X1 U8752 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n5404)
         );
  AOI22_X1 U8753 ( .A1(n28372), .A2(\xmem_data[64][4] ), .B1(n30698), .B2(
        \xmem_data[65][4] ), .ZN(n5402) );
  AOI22_X1 U8754 ( .A1(n28343), .A2(\xmem_data[66][4] ), .B1(n28972), .B2(
        \xmem_data[67][4] ), .ZN(n5401) );
  AOI22_X1 U8755 ( .A1(n24158), .A2(\xmem_data[68][4] ), .B1(n28089), .B2(
        \xmem_data[69][4] ), .ZN(n5400) );
  AOI22_X1 U8756 ( .A1(n24212), .A2(\xmem_data[70][4] ), .B1(n25459), .B2(
        \xmem_data[71][4] ), .ZN(n5399) );
  NAND4_X1 U8757 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5403)
         );
  AOI22_X1 U8758 ( .A1(n29055), .A2(\xmem_data[48][4] ), .B1(n29054), .B2(
        \xmem_data[49][4] ), .ZN(n5412) );
  AOI22_X1 U8759 ( .A1(n14975), .A2(\xmem_data[50][4] ), .B1(n29325), .B2(
        \xmem_data[51][4] ), .ZN(n5411) );
  AND2_X1 U8760 ( .A1(n25359), .A2(\xmem_data[52][4] ), .ZN(n5408) );
  AOI21_X1 U8761 ( .B1(n27568), .B2(\xmem_data[53][4] ), .A(n5408), .ZN(n5410)
         );
  AOI22_X1 U8762 ( .A1(n24468), .A2(\xmem_data[54][4] ), .B1(n29057), .B2(
        \xmem_data[55][4] ), .ZN(n5409) );
  NAND4_X1 U8763 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n5428)
         );
  AOI22_X1 U8764 ( .A1(n29046), .A2(\xmem_data[40][4] ), .B1(n28091), .B2(
        \xmem_data[41][4] ), .ZN(n5416) );
  AOI22_X1 U8765 ( .A1(n28993), .A2(\xmem_data[42][4] ), .B1(n29010), .B2(
        \xmem_data[43][4] ), .ZN(n5415) );
  AOI22_X1 U8766 ( .A1(n29048), .A2(\xmem_data[44][4] ), .B1(n29047), .B2(
        \xmem_data[45][4] ), .ZN(n5414) );
  AOI22_X1 U8767 ( .A1(n29049), .A2(\xmem_data[46][4] ), .B1(n25521), .B2(
        \xmem_data[47][4] ), .ZN(n5413) );
  NAND4_X1 U8768 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n5427)
         );
  AOI22_X1 U8769 ( .A1(n12471), .A2(\xmem_data[56][4] ), .B1(n3305), .B2(
        \xmem_data[57][4] ), .ZN(n5420) );
  AOI22_X1 U8770 ( .A1(n28501), .A2(\xmem_data[58][4] ), .B1(n28364), .B2(
        \xmem_data[59][4] ), .ZN(n5419) );
  AOI22_X1 U8771 ( .A1(n3217), .A2(\xmem_data[60][4] ), .B1(n29065), .B2(
        \xmem_data[61][4] ), .ZN(n5418) );
  AOI22_X1 U8772 ( .A1(n23739), .A2(\xmem_data[62][4] ), .B1(n20994), .B2(
        \xmem_data[63][4] ), .ZN(n5417) );
  NAND4_X1 U8773 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n5426)
         );
  AOI22_X1 U8774 ( .A1(n27550), .A2(\xmem_data[32][4] ), .B1(n21074), .B2(
        \xmem_data[33][4] ), .ZN(n5424) );
  BUF_X1 U8775 ( .A(n13474), .Z(n29045) );
  AOI22_X1 U8776 ( .A1(n29045), .A2(\xmem_data[34][4] ), .B1(n27447), .B2(
        \xmem_data[35][4] ), .ZN(n5423) );
  AOI22_X1 U8777 ( .A1(n20546), .A2(\xmem_data[36][4] ), .B1(n25457), .B2(
        \xmem_data[37][4] ), .ZN(n5422) );
  AOI22_X1 U8778 ( .A1(n27535), .A2(\xmem_data[38][4] ), .B1(n28298), .B2(
        \xmem_data[39][4] ), .ZN(n5421) );
  NAND4_X1 U8779 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n5425)
         );
  AOI22_X1 U8780 ( .A1(n29281), .A2(\xmem_data[16][4] ), .B1(n17004), .B2(
        \xmem_data[17][4] ), .ZN(n5433) );
  AOI22_X1 U8781 ( .A1(n28983), .A2(\xmem_data[18][4] ), .B1(n29325), .B2(
        \xmem_data[19][4] ), .ZN(n5432) );
  AOI22_X1 U8782 ( .A1(n28979), .A2(\xmem_data[20][4] ), .B1(n27717), .B2(
        \xmem_data[21][4] ), .ZN(n5431) );
  AOI22_X1 U8783 ( .A1(n29248), .A2(\xmem_data[22][4] ), .B1(n20953), .B2(
        \xmem_data[23][4] ), .ZN(n5430) );
  NAND4_X1 U8784 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n5450)
         );
  AOI22_X1 U8785 ( .A1(n21309), .A2(\xmem_data[24][4] ), .B1(n3383), .B2(
        \xmem_data[25][4] ), .ZN(n5437) );
  AOI22_X1 U8786 ( .A1(n30589), .A2(\xmem_data[26][4] ), .B1(n29064), .B2(
        \xmem_data[27][4] ), .ZN(n5436) );
  AOI22_X1 U8787 ( .A1(n3219), .A2(\xmem_data[28][4] ), .B1(n24632), .B2(
        \xmem_data[29][4] ), .ZN(n5435) );
  AOI22_X1 U8788 ( .A1(n31367), .A2(\xmem_data[30][4] ), .B1(n3340), .B2(
        \xmem_data[31][4] ), .ZN(n5434) );
  NAND4_X1 U8789 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n5448)
         );
  AOI22_X1 U8790 ( .A1(n25616), .A2(\xmem_data[0][4] ), .B1(n3374), .B2(
        \xmem_data[1][4] ), .ZN(n5441) );
  AOI22_X1 U8791 ( .A1(n25514), .A2(\xmem_data[2][4] ), .B1(n24554), .B2(
        \xmem_data[3][4] ), .ZN(n5440) );
  AOI22_X1 U8792 ( .A1(n22739), .A2(\xmem_data[4][4] ), .B1(n28051), .B2(
        \xmem_data[5][4] ), .ZN(n5439) );
  AOI22_X1 U8793 ( .A1(n24212), .A2(\xmem_data[6][4] ), .B1(n25710), .B2(
        \xmem_data[7][4] ), .ZN(n5438) );
  NAND4_X1 U8794 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n5447)
         );
  AOI22_X1 U8795 ( .A1(n25382), .A2(\xmem_data[8][4] ), .B1(n17018), .B2(
        \xmem_data[9][4] ), .ZN(n5445) );
  AOI22_X1 U8796 ( .A1(n28993), .A2(\xmem_data[10][4] ), .B1(n21007), .B2(
        \xmem_data[11][4] ), .ZN(n5444) );
  AOI22_X1 U8797 ( .A1(n25520), .A2(\xmem_data[12][4] ), .B1(n28994), .B2(
        \xmem_data[13][4] ), .ZN(n5443) );
  AOI22_X1 U8798 ( .A1(n30616), .A2(\xmem_data[14][4] ), .B1(n28061), .B2(
        \xmem_data[15][4] ), .ZN(n5442) );
  NAND4_X1 U8799 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n5446)
         );
  XNOR2_X1 U8800 ( .A(n32617), .B(\fmem_data[9][7] ), .ZN(n31977) );
  XOR2_X1 U8801 ( .A(\fmem_data[9][6] ), .B(\fmem_data[9][7] ), .Z(n5455) );
  OAI22_X1 U8802 ( .A1(n35022), .A2(n35726), .B1(n31977), .B2(n35725), .ZN(
        n35092) );
  AND2_X1 U8803 ( .A1(n24439), .A2(\xmem_data[86][5] ), .ZN(n5456) );
  AOI21_X1 U8804 ( .B1(n25730), .B2(\xmem_data[87][5] ), .A(n5456), .ZN(n5457)
         );
  INV_X1 U8805 ( .A(n5457), .ZN(n5465) );
  AOI22_X1 U8806 ( .A1(n22702), .A2(\xmem_data[66][5] ), .B1(n28980), .B2(
        \xmem_data[67][5] ), .ZN(n5459) );
  AOI22_X1 U8807 ( .A1(n22701), .A2(\xmem_data[64][5] ), .B1(n22738), .B2(
        \xmem_data[65][5] ), .ZN(n5458) );
  NAND2_X1 U8808 ( .A1(n5459), .A2(n5458), .ZN(n5464) );
  AOI22_X1 U8809 ( .A1(n24457), .A2(\xmem_data[70][5] ), .B1(n29317), .B2(
        \xmem_data[71][5] ), .ZN(n5462) );
  AOI22_X1 U8810 ( .A1(n22703), .A2(\xmem_data[68][5] ), .B1(n31328), .B2(
        \xmem_data[69][5] ), .ZN(n5461) );
  AOI22_X1 U8811 ( .A1(n22727), .A2(\xmem_data[82][5] ), .B1(n30909), .B2(
        \xmem_data[83][5] ), .ZN(n5460) );
  NOR3_X1 U8812 ( .A1(n5465), .A2(n5464), .A3(n5463), .ZN(n5466) );
  INV_X1 U8813 ( .A(n22663), .ZN(n5520) );
  NOR2_X1 U8814 ( .A1(n5466), .A2(n5520), .ZN(n5506) );
  AOI22_X1 U8815 ( .A1(n22701), .A2(\xmem_data[32][5] ), .B1(n25708), .B2(
        \xmem_data[33][5] ), .ZN(n5470) );
  AOI22_X1 U8816 ( .A1(n22702), .A2(\xmem_data[34][5] ), .B1(n31268), .B2(
        \xmem_data[35][5] ), .ZN(n5469) );
  AOI22_X1 U8817 ( .A1(n22703), .A2(\xmem_data[36][5] ), .B1(n30666), .B2(
        \xmem_data[37][5] ), .ZN(n5468) );
  AOI22_X1 U8818 ( .A1(n28299), .A2(\xmem_data[38][5] ), .B1(n25573), .B2(
        \xmem_data[39][5] ), .ZN(n5467) );
  NAND4_X1 U8819 ( .A1(n5470), .A2(n5469), .A3(n5468), .A4(n5467), .ZN(n5474)
         );
  NAND2_X1 U8820 ( .A1(n28772), .A2(\xmem_data[49][5] ), .ZN(n5472) );
  NAND2_X1 U8821 ( .A1(n27526), .A2(\xmem_data[48][5] ), .ZN(n5471) );
  NAND2_X1 U8822 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NOR2_X1 U8823 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  INV_X1 U8824 ( .A(n22735), .ZN(n5535) );
  NOR2_X1 U8825 ( .A1(n5475), .A2(n5535), .ZN(n5505) );
  AOI22_X1 U8826 ( .A1(n27943), .A2(\xmem_data[96][5] ), .B1(n24556), .B2(
        \xmem_data[97][5] ), .ZN(n5479) );
  AOI22_X1 U8827 ( .A1(n22675), .A2(\xmem_data[98][5] ), .B1(n28298), .B2(
        \xmem_data[99][5] ), .ZN(n5478) );
  AOI22_X1 U8828 ( .A1(n22674), .A2(\xmem_data[100][5] ), .B1(n17018), .B2(
        \xmem_data[101][5] ), .ZN(n5477) );
  AOI22_X1 U8829 ( .A1(n22677), .A2(\xmem_data[102][5] ), .B1(n22676), .B2(
        \xmem_data[103][5] ), .ZN(n5476) );
  NAND4_X1 U8830 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n5483)
         );
  NAND2_X1 U8831 ( .A1(n29725), .A2(\xmem_data[113][5] ), .ZN(n5481) );
  NAND2_X1 U8832 ( .A1(n29017), .A2(\xmem_data[112][5] ), .ZN(n5480) );
  NAND2_X1 U8833 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NOR2_X1 U8834 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  INV_X1 U8835 ( .A(n22698), .ZN(n5533) );
  NOR2_X1 U8836 ( .A1(n5484), .A2(n5533), .ZN(n5504) );
  AOI22_X1 U8837 ( .A1(n3219), .A2(\xmem_data[56][5] ), .B1(n22708), .B2(
        \xmem_data[57][5] ), .ZN(n5488) );
  AOI22_X1 U8838 ( .A1(n22710), .A2(\xmem_data[58][5] ), .B1(n22709), .B2(
        \xmem_data[59][5] ), .ZN(n5487) );
  AOI22_X1 U8839 ( .A1(n22711), .A2(\xmem_data[60][5] ), .B1(n29231), .B2(
        \xmem_data[61][5] ), .ZN(n5486) );
  AOI22_X1 U8840 ( .A1(n27547), .A2(\xmem_data[62][5] ), .B1(n22712), .B2(
        \xmem_data[63][5] ), .ZN(n5485) );
  NAND4_X1 U8841 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n5492)
         );
  AOI22_X1 U8842 ( .A1(n22729), .A2(\xmem_data[52][5] ), .B1(n22728), .B2(
        \xmem_data[53][5] ), .ZN(n5490) );
  AOI22_X1 U8843 ( .A1(n22727), .A2(\xmem_data[50][5] ), .B1(n20986), .B2(
        \xmem_data[51][5] ), .ZN(n5489) );
  NAND2_X1 U8844 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NOR2_X1 U8845 ( .A1(n5492), .A2(n5491), .ZN(n5502) );
  AOI22_X1 U8846 ( .A1(n3221), .A2(\xmem_data[120][5] ), .B1(n25448), .B2(
        \xmem_data[121][5] ), .ZN(n5496) );
  AOI22_X1 U8847 ( .A1(n22667), .A2(\xmem_data[122][5] ), .B1(n22666), .B2(
        \xmem_data[123][5] ), .ZN(n5495) );
  AOI22_X1 U8848 ( .A1(n22669), .A2(\xmem_data[124][5] ), .B1(n22668), .B2(
        \xmem_data[125][5] ), .ZN(n5494) );
  AOI22_X1 U8849 ( .A1(n28045), .A2(\xmem_data[126][5] ), .B1(n28374), .B2(
        \xmem_data[127][5] ), .ZN(n5493) );
  NAND4_X1 U8850 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n5500)
         );
  AOI22_X1 U8851 ( .A1(n30861), .A2(\xmem_data[116][5] ), .B1(n3412), .B2(
        \xmem_data[117][5] ), .ZN(n5498) );
  AOI22_X1 U8852 ( .A1(n25388), .A2(\xmem_data[114][5] ), .B1(n25630), .B2(
        \xmem_data[115][5] ), .ZN(n5497) );
  NAND2_X1 U8853 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NOR2_X1 U8854 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  OAI22_X1 U8855 ( .A1(n5502), .A2(n5535), .B1(n5501), .B2(n5533), .ZN(n5503)
         );
  NOR4_X1 U8856 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n5568)
         );
  AOI22_X1 U8857 ( .A1(n3220), .A2(\xmem_data[88][5] ), .B1(n22708), .B2(
        \xmem_data[89][5] ), .ZN(n5510) );
  AOI22_X1 U8858 ( .A1(n22710), .A2(\xmem_data[90][5] ), .B1(n22709), .B2(
        \xmem_data[91][5] ), .ZN(n5509) );
  AOI22_X1 U8859 ( .A1(n22711), .A2(\xmem_data[92][5] ), .B1(n3282), .B2(
        \xmem_data[93][5] ), .ZN(n5508) );
  AOI22_X1 U8860 ( .A1(n28045), .A2(\xmem_data[94][5] ), .B1(n22712), .B2(
        \xmem_data[95][5] ), .ZN(n5507) );
  NAND4_X1 U8861 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .ZN(n5513)
         );
  AOI22_X1 U8862 ( .A1(n22729), .A2(\xmem_data[84][5] ), .B1(n22728), .B2(
        \xmem_data[85][5] ), .ZN(n5511) );
  INV_X1 U8863 ( .A(n5511), .ZN(n5512) );
  NOR2_X1 U8864 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NOR2_X1 U8865 ( .A1(n5514), .A2(n5520), .ZN(n5539) );
  AOI22_X1 U8866 ( .A1(n22718), .A2(\xmem_data[72][5] ), .B1(n22717), .B2(
        \xmem_data[73][5] ), .ZN(n5518) );
  AOI22_X1 U8867 ( .A1(n29049), .A2(\xmem_data[74][5] ), .B1(n30899), .B2(
        \xmem_data[75][5] ), .ZN(n5517) );
  AOI22_X1 U8868 ( .A1(n20943), .A2(\xmem_data[76][5] ), .B1(n3328), .B2(
        \xmem_data[77][5] ), .ZN(n5516) );
  AOI22_X1 U8869 ( .A1(n24223), .A2(\xmem_data[78][5] ), .B1(n22719), .B2(
        \xmem_data[79][5] ), .ZN(n5515) );
  AOI22_X1 U8870 ( .A1(n29253), .A2(\xmem_data[118][5] ), .B1(n25692), .B2(
        \xmem_data[119][5] ), .ZN(n5519) );
  OAI22_X1 U8871 ( .A1(n3751), .A2(n5520), .B1(n5519), .B2(n5533), .ZN(n5538)
         );
  AOI22_X1 U8872 ( .A1(n28501), .A2(\xmem_data[54][5] ), .B1(n27902), .B2(
        \xmem_data[55][5] ), .ZN(n5522) );
  AOI22_X1 U8873 ( .A1(n29017), .A2(\xmem_data[80][5] ), .B1(n14982), .B2(
        \xmem_data[81][5] ), .ZN(n5521) );
  OAI22_X1 U8874 ( .A1(n5522), .A2(n5535), .B1(n5521), .B2(n5520), .ZN(n5537)
         );
  AOI22_X1 U8875 ( .A1(n22718), .A2(\xmem_data[40][5] ), .B1(n22717), .B2(
        \xmem_data[41][5] ), .ZN(n5526) );
  AOI22_X1 U8876 ( .A1(n30871), .A2(\xmem_data[42][5] ), .B1(n24615), .B2(
        \xmem_data[43][5] ), .ZN(n5525) );
  AOI22_X1 U8877 ( .A1(n28291), .A2(\xmem_data[44][5] ), .B1(n3329), .B2(
        \xmem_data[45][5] ), .ZN(n5524) );
  AOI22_X1 U8878 ( .A1(n23779), .A2(\xmem_data[46][5] ), .B1(n22719), .B2(
        \xmem_data[47][5] ), .ZN(n5523) );
  AOI22_X1 U8879 ( .A1(n25435), .A2(\xmem_data[106][5] ), .B1(n22683), .B2(
        \xmem_data[107][5] ), .ZN(n5527) );
  INV_X1 U8880 ( .A(n5527), .ZN(n5532) );
  AOI22_X1 U8881 ( .A1(n28327), .A2(\xmem_data[108][5] ), .B1(n21056), .B2(
        \xmem_data[109][5] ), .ZN(n5530) );
  AOI22_X1 U8882 ( .A1(n22685), .A2(\xmem_data[110][5] ), .B1(n22684), .B2(
        \xmem_data[111][5] ), .ZN(n5529) );
  AOI22_X1 U8883 ( .A1(n17043), .A2(\xmem_data[104][5] ), .B1(n22682), .B2(
        \xmem_data[105][5] ), .ZN(n5528) );
  NOR2_X1 U8884 ( .A1(n5532), .A2(n5531), .ZN(n5534) );
  OAI22_X1 U8885 ( .A1(n3743), .A2(n5535), .B1(n5534), .B2(n5533), .ZN(n5536)
         );
  NOR4_X1 U8886 ( .A1(n5539), .A2(n5538), .A3(n5537), .A4(n5536), .ZN(n5567)
         );
  AOI22_X1 U8887 ( .A1(n3219), .A2(\xmem_data[24][5] ), .B1(n29789), .B2(
        \xmem_data[25][5] ), .ZN(n5544) );
  AOI22_X1 U8888 ( .A1(n22759), .A2(\xmem_data[28][5] ), .B1(n23742), .B2(
        \xmem_data[29][5] ), .ZN(n5540) );
  AOI22_X1 U8889 ( .A1(n20558), .A2(\xmem_data[26][5] ), .B1(n22758), .B2(
        \xmem_data[27][5] ), .ZN(n5542) );
  NAND2_X1 U8890 ( .A1(n27447), .A2(\xmem_data[31][5] ), .ZN(n5541) );
  NAND2_X1 U8891 ( .A1(n5544), .A2(n5543), .ZN(n5550) );
  AOI22_X1 U8892 ( .A1(n22739), .A2(\xmem_data[0][5] ), .B1(n22738), .B2(
        \xmem_data[1][5] ), .ZN(n5548) );
  AOI22_X1 U8893 ( .A1(n22740), .A2(\xmem_data[2][5] ), .B1(n20541), .B2(
        \xmem_data[3][5] ), .ZN(n5547) );
  AOI22_X1 U8894 ( .A1(n22741), .A2(\xmem_data[4][5] ), .B1(n3158), .B2(
        \xmem_data[5][5] ), .ZN(n5546) );
  AOI22_X1 U8895 ( .A1(n22742), .A2(\xmem_data[6][5] ), .B1(n25434), .B2(
        \xmem_data[7][5] ), .ZN(n5545) );
  NAND4_X1 U8896 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n5549)
         );
  OR2_X1 U8897 ( .A1(n5550), .A2(n5549), .ZN(n5563) );
  AND2_X1 U8898 ( .A1(n22751), .A2(\xmem_data[16][5] ), .ZN(n5551) );
  AOI21_X1 U8899 ( .B1(n29820), .B2(\xmem_data[17][5] ), .A(n5551), .ZN(n5555)
         );
  AOI22_X1 U8900 ( .A1(n24468), .A2(\xmem_data[18][5] ), .B1(n24607), .B2(
        \xmem_data[19][5] ), .ZN(n5554) );
  AOI22_X1 U8901 ( .A1(n22752), .A2(\xmem_data[20][5] ), .B1(n28039), .B2(
        \xmem_data[21][5] ), .ZN(n5553) );
  AOI22_X1 U8902 ( .A1(n22753), .A2(\xmem_data[22][5] ), .B1(n29064), .B2(
        \xmem_data[23][5] ), .ZN(n5552) );
  NAND4_X1 U8903 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n5561)
         );
  AOI22_X1 U8904 ( .A1(n24219), .A2(\xmem_data[8][5] ), .B1(n27825), .B2(
        \xmem_data[9][5] ), .ZN(n5559) );
  AOI22_X1 U8905 ( .A1(n30871), .A2(\xmem_data[10][5] ), .B1(n28428), .B2(
        \xmem_data[11][5] ), .ZN(n5558) );
  AOI22_X1 U8906 ( .A1(n20506), .A2(\xmem_data[12][5] ), .B1(n20817), .B2(
        \xmem_data[13][5] ), .ZN(n5557) );
  AOI22_X1 U8907 ( .A1(n31362), .A2(\xmem_data[14][5] ), .B1(n29325), .B2(
        \xmem_data[15][5] ), .ZN(n5556) );
  NAND4_X1 U8908 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n5560)
         );
  OR2_X1 U8909 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  OR2_X1 U8910 ( .A1(n5563), .A2(n5562), .ZN(n5565) );
  INV_X1 U8911 ( .A(n22768), .ZN(n22022) );
  NOR2_X1 U8912 ( .A1(n22022), .A2(n39023), .ZN(n5564) );
  AOI21_X1 U8913 ( .B1(n5565), .B2(n22768), .A(n3882), .ZN(n5566) );
  AOI22_X1 U8914 ( .A1(n22718), .A2(\xmem_data[72][4] ), .B1(n22717), .B2(
        \xmem_data[73][4] ), .ZN(n5572) );
  AOI22_X1 U8915 ( .A1(n29280), .A2(\xmem_data[74][4] ), .B1(n25632), .B2(
        \xmem_data[75][4] ), .ZN(n5571) );
  AOI22_X1 U8916 ( .A1(n23778), .A2(\xmem_data[76][4] ), .B1(n3337), .B2(
        \xmem_data[77][4] ), .ZN(n5570) );
  AOI22_X1 U8917 ( .A1(n28098), .A2(\xmem_data[78][4] ), .B1(n22719), .B2(
        \xmem_data[79][4] ), .ZN(n5569) );
  NAND4_X1 U8918 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(n5576)
         );
  AND2_X1 U8919 ( .A1(n20568), .A2(\xmem_data[86][4] ), .ZN(n5573) );
  AOI21_X1 U8920 ( .B1(n23734), .B2(\xmem_data[87][4] ), .A(n5573), .ZN(n5574)
         );
  INV_X1 U8921 ( .A(n5574), .ZN(n5575) );
  AOI22_X1 U8922 ( .A1(n22703), .A2(\xmem_data[68][4] ), .B1(n3465), .B2(
        \xmem_data[69][4] ), .ZN(n5580) );
  AOI22_X1 U8923 ( .A1(n22702), .A2(\xmem_data[66][4] ), .B1(n30891), .B2(
        \xmem_data[67][4] ), .ZN(n5579) );
  AOI22_X1 U8924 ( .A1(n22701), .A2(\xmem_data[64][4] ), .B1(n28309), .B2(
        \xmem_data[65][4] ), .ZN(n5578) );
  AOI22_X1 U8925 ( .A1(n24457), .A2(\xmem_data[70][4] ), .B1(n20585), .B2(
        \xmem_data[71][4] ), .ZN(n5577) );
  NAND4_X1 U8926 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n5583)
         );
  AOI22_X1 U8927 ( .A1(n22729), .A2(\xmem_data[84][4] ), .B1(n22728), .B2(
        \xmem_data[85][4] ), .ZN(n5581) );
  INV_X1 U8928 ( .A(n5581), .ZN(n5582) );
  NOR2_X1 U8929 ( .A1(n5583), .A2(n5582), .ZN(n5593) );
  AOI22_X1 U8930 ( .A1(n3218), .A2(\xmem_data[88][4] ), .B1(n22708), .B2(
        \xmem_data[89][4] ), .ZN(n5587) );
  AOI22_X1 U8931 ( .A1(n22710), .A2(\xmem_data[90][4] ), .B1(n22709), .B2(
        \xmem_data[91][4] ), .ZN(n5586) );
  AOI22_X1 U8932 ( .A1(n22711), .A2(\xmem_data[92][4] ), .B1(n3375), .B2(
        \xmem_data[93][4] ), .ZN(n5585) );
  AOI22_X1 U8933 ( .A1(n13474), .A2(\xmem_data[94][4] ), .B1(n22712), .B2(
        \xmem_data[95][4] ), .ZN(n5584) );
  NAND4_X1 U8934 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n5590)
         );
  AOI22_X1 U8935 ( .A1(n22727), .A2(\xmem_data[82][4] ), .B1(n28038), .B2(
        \xmem_data[83][4] ), .ZN(n5588) );
  INV_X1 U8936 ( .A(n5588), .ZN(n5589) );
  NOR2_X1 U8937 ( .A1(n5590), .A2(n5589), .ZN(n5592) );
  AOI22_X1 U8938 ( .A1(n29017), .A2(\xmem_data[80][4] ), .B1(n29820), .B2(
        \xmem_data[81][4] ), .ZN(n5591) );
  NAND3_X1 U8939 ( .A1(n5593), .A2(n5592), .A3(n5591), .ZN(n5594) );
  OAI21_X1 U8940 ( .B1(n3983), .B2(n5594), .A(n22663), .ZN(n5666) );
  AOI22_X1 U8941 ( .A1(n31355), .A2(\xmem_data[104][4] ), .B1(n22682), .B2(
        \xmem_data[105][4] ), .ZN(n5598) );
  AOI22_X1 U8942 ( .A1(n24221), .A2(\xmem_data[106][4] ), .B1(n22683), .B2(
        \xmem_data[107][4] ), .ZN(n5597) );
  AOI22_X1 U8943 ( .A1(n25364), .A2(\xmem_data[108][4] ), .B1(n20950), .B2(
        \xmem_data[109][4] ), .ZN(n5596) );
  AOI22_X1 U8944 ( .A1(n22685), .A2(\xmem_data[110][4] ), .B1(n22684), .B2(
        \xmem_data[111][4] ), .ZN(n5595) );
  NAND4_X1 U8945 ( .A1(n5598), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n5602)
         );
  AND2_X1 U8946 ( .A1(n25485), .A2(\xmem_data[118][4] ), .ZN(n5599) );
  AOI21_X1 U8947 ( .B1(n24443), .B2(\xmem_data[119][4] ), .A(n5599), .ZN(n5600) );
  INV_X1 U8948 ( .A(n5600), .ZN(n5601) );
  AOI22_X1 U8949 ( .A1(n27943), .A2(\xmem_data[96][4] ), .B1(n24640), .B2(
        \xmem_data[97][4] ), .ZN(n5606) );
  AOI22_X1 U8950 ( .A1(n22675), .A2(\xmem_data[98][4] ), .B1(n25425), .B2(
        \xmem_data[99][4] ), .ZN(n5605) );
  AOI22_X1 U8951 ( .A1(n22674), .A2(\xmem_data[100][4] ), .B1(n29437), .B2(
        \xmem_data[101][4] ), .ZN(n5604) );
  AOI22_X1 U8952 ( .A1(n22677), .A2(\xmem_data[102][4] ), .B1(n22676), .B2(
        \xmem_data[103][4] ), .ZN(n5603) );
  NAND4_X1 U8953 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n5609)
         );
  AOI22_X1 U8954 ( .A1(n20578), .A2(\xmem_data[116][4] ), .B1(n3413), .B2(
        \xmem_data[117][4] ), .ZN(n5607) );
  INV_X1 U8955 ( .A(n5607), .ZN(n5608) );
  NOR2_X1 U8956 ( .A1(n5609), .A2(n5608), .ZN(n5619) );
  AOI22_X1 U8957 ( .A1(n3221), .A2(\xmem_data[120][4] ), .B1(n25414), .B2(
        \xmem_data[121][4] ), .ZN(n5613) );
  AOI22_X1 U8958 ( .A1(n22667), .A2(\xmem_data[122][4] ), .B1(n22666), .B2(
        \xmem_data[123][4] ), .ZN(n5612) );
  AOI22_X1 U8959 ( .A1(n22669), .A2(\xmem_data[124][4] ), .B1(n22668), .B2(
        \xmem_data[125][4] ), .ZN(n5611) );
  AOI22_X1 U8960 ( .A1(n27446), .A2(\xmem_data[126][4] ), .B1(n28374), .B2(
        \xmem_data[127][4] ), .ZN(n5610) );
  NAND4_X1 U8961 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5616)
         );
  AOI22_X1 U8962 ( .A1(n29326), .A2(\xmem_data[114][4] ), .B1(n25358), .B2(
        \xmem_data[115][4] ), .ZN(n5614) );
  INV_X1 U8963 ( .A(n5614), .ZN(n5615) );
  NOR2_X1 U8964 ( .A1(n5616), .A2(n5615), .ZN(n5618) );
  AOI22_X1 U8965 ( .A1(n23725), .A2(\xmem_data[112][4] ), .B1(n20567), .B2(
        \xmem_data[113][4] ), .ZN(n5617) );
  OAI21_X1 U8966 ( .B1(n3984), .B2(n5620), .A(n22698), .ZN(n5665) );
  AOI22_X1 U8967 ( .A1(n22718), .A2(\xmem_data[40][4] ), .B1(n22717), .B2(
        \xmem_data[41][4] ), .ZN(n5624) );
  AOI22_X1 U8968 ( .A1(n31360), .A2(\xmem_data[42][4] ), .B1(n30899), .B2(
        \xmem_data[43][4] ), .ZN(n5623) );
  AOI22_X1 U8969 ( .A1(n30898), .A2(\xmem_data[44][4] ), .B1(n23780), .B2(
        \xmem_data[45][4] ), .ZN(n5622) );
  AOI22_X1 U8970 ( .A1(n24622), .A2(\xmem_data[46][4] ), .B1(n22719), .B2(
        \xmem_data[47][4] ), .ZN(n5621) );
  AOI22_X1 U8971 ( .A1(n25527), .A2(\xmem_data[48][4] ), .B1(n20577), .B2(
        \xmem_data[49][4] ), .ZN(n5626) );
  AOI22_X1 U8972 ( .A1(n31347), .A2(\xmem_data[54][4] ), .B1(n25354), .B2(
        \xmem_data[55][4] ), .ZN(n5625) );
  AOI22_X1 U8973 ( .A1(n22701), .A2(\xmem_data[32][4] ), .B1(n28089), .B2(
        \xmem_data[33][4] ), .ZN(n5630) );
  AOI22_X1 U8974 ( .A1(n22702), .A2(\xmem_data[34][4] ), .B1(n3175), .B2(
        \xmem_data[35][4] ), .ZN(n5629) );
  AOI22_X1 U8975 ( .A1(n22703), .A2(\xmem_data[36][4] ), .B1(n29315), .B2(
        \xmem_data[37][4] ), .ZN(n5628) );
  AOI22_X1 U8976 ( .A1(n31269), .A2(\xmem_data[38][4] ), .B1(n13149), .B2(
        \xmem_data[39][4] ), .ZN(n5627) );
  AOI22_X1 U8977 ( .A1(n22727), .A2(\xmem_data[50][4] ), .B1(n30588), .B2(
        \xmem_data[51][4] ), .ZN(n5636) );
  AOI22_X1 U8978 ( .A1(n3218), .A2(\xmem_data[56][4] ), .B1(n22708), .B2(
        \xmem_data[57][4] ), .ZN(n5634) );
  AOI22_X1 U8979 ( .A1(n22710), .A2(\xmem_data[58][4] ), .B1(n22709), .B2(
        \xmem_data[59][4] ), .ZN(n5633) );
  AOI22_X1 U8980 ( .A1(n22711), .A2(\xmem_data[60][4] ), .B1(n21074), .B2(
        \xmem_data[61][4] ), .ZN(n5632) );
  AOI22_X1 U8981 ( .A1(n25450), .A2(\xmem_data[62][4] ), .B1(n22712), .B2(
        \xmem_data[63][4] ), .ZN(n5631) );
  AOI22_X1 U8982 ( .A1(n22729), .A2(\xmem_data[52][4] ), .B1(n22728), .B2(
        \xmem_data[53][4] ), .ZN(n5635) );
  NAND4_X1 U8983 ( .A1(n3845), .A2(n5636), .A3(n3527), .A4(n5635), .ZN(n5637)
         );
  OAI21_X1 U8984 ( .B1(n5638), .B2(n5637), .A(n22735), .ZN(n5664) );
  AOI22_X1 U8985 ( .A1(n28510), .A2(\xmem_data[30][4] ), .B1(n23813), .B2(
        \xmem_data[31][4] ), .ZN(n5639) );
  INV_X1 U8986 ( .A(n5639), .ZN(n5645) );
  AOI22_X1 U8987 ( .A1(n22751), .A2(\xmem_data[16][4] ), .B1(n28192), .B2(
        \xmem_data[17][4] ), .ZN(n5640) );
  INV_X1 U8988 ( .A(n5640), .ZN(n5644) );
  AOI22_X1 U8989 ( .A1(n27567), .A2(\xmem_data[18][4] ), .B1(n25358), .B2(
        \xmem_data[19][4] ), .ZN(n5642) );
  AOI22_X1 U8990 ( .A1(n22753), .A2(\xmem_data[22][4] ), .B1(n29064), .B2(
        \xmem_data[23][4] ), .ZN(n5641) );
  NAND2_X1 U8991 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  NOR3_X1 U8992 ( .A1(n5645), .A2(n5644), .A3(n5643), .ZN(n5661) );
  AOI22_X1 U8993 ( .A1(n24707), .A2(\xmem_data[8][4] ), .B1(n28687), .B2(
        \xmem_data[9][4] ), .ZN(n5649) );
  AOI22_X1 U8994 ( .A1(n29238), .A2(\xmem_data[10][4] ), .B1(n28428), .B2(
        \xmem_data[11][4] ), .ZN(n5648) );
  AOI22_X1 U8995 ( .A1(n28327), .A2(\xmem_data[12][4] ), .B1(n23780), .B2(
        \xmem_data[13][4] ), .ZN(n5647) );
  AOI22_X1 U8996 ( .A1(n28495), .A2(\xmem_data[14][4] ), .B1(n29325), .B2(
        \xmem_data[15][4] ), .ZN(n5646) );
  AOI22_X1 U8997 ( .A1(n22759), .A2(\xmem_data[28][4] ), .B1(n3344), .B2(
        \xmem_data[29][4] ), .ZN(n5652) );
  AOI22_X1 U8998 ( .A1(n30963), .A2(\xmem_data[26][4] ), .B1(n22758), .B2(
        \xmem_data[27][4] ), .ZN(n5651) );
  AOI22_X1 U8999 ( .A1(n3217), .A2(\xmem_data[24][4] ), .B1(n27831), .B2(
        \xmem_data[25][4] ), .ZN(n5650) );
  NAND3_X1 U9000 ( .A1(n5652), .A2(n5651), .A3(n5650), .ZN(n5655) );
  AOI22_X1 U9001 ( .A1(n22752), .A2(\xmem_data[20][4] ), .B1(n24630), .B2(
        \xmem_data[21][4] ), .ZN(n5653) );
  INV_X1 U9002 ( .A(n5653), .ZN(n5654) );
  NOR2_X1 U9003 ( .A1(n5655), .A2(n5654), .ZN(n5660) );
  AOI22_X1 U9004 ( .A1(n22739), .A2(\xmem_data[0][4] ), .B1(n22738), .B2(
        \xmem_data[1][4] ), .ZN(n5659) );
  AOI22_X1 U9005 ( .A1(n22740), .A2(\xmem_data[2][4] ), .B1(n25459), .B2(
        \xmem_data[3][4] ), .ZN(n5658) );
  AOI22_X1 U9006 ( .A1(n22741), .A2(\xmem_data[4][4] ), .B1(n29315), .B2(
        \xmem_data[5][4] ), .ZN(n5657) );
  AOI22_X1 U9007 ( .A1(n22742), .A2(\xmem_data[6][4] ), .B1(n30949), .B2(
        \xmem_data[7][4] ), .ZN(n5656) );
  NAND4_X1 U9008 ( .A1(n5661), .A2(n3790), .A3(n5660), .A4(n3500), .ZN(n5662)
         );
  NAND2_X1 U9009 ( .A1(n5662), .A2(n22768), .ZN(n5663) );
  XNOR2_X1 U9010 ( .A(n31233), .B(\fmem_data[5][7] ), .ZN(n23920) );
  XOR2_X1 U9011 ( .A(\fmem_data[5][6] ), .B(\fmem_data[5][7] ), .Z(n5667) );
  XOR2_X1 U9012 ( .A(\fmem_data[28][3] ), .B(\fmem_data[28][2] ), .Z(n5668) );
  BUF_X1 U9013 ( .A(n13435), .Z(n20775) );
  AOI22_X1 U9014 ( .A1(n25457), .A2(\xmem_data[24][7] ), .B1(n20775), .B2(
        \xmem_data[25][7] ), .ZN(n5672) );
  AOI22_X1 U9015 ( .A1(n29023), .A2(\xmem_data[26][7] ), .B1(n25709), .B2(
        \xmem_data[27][7] ), .ZN(n5671) );
  BUF_X1 U9016 ( .A(n29187), .Z(n20776) );
  AOI22_X1 U9017 ( .A1(n28752), .A2(\xmem_data[28][7] ), .B1(n24457), .B2(
        \xmem_data[29][7] ), .ZN(n5670) );
  AOI22_X1 U9018 ( .A1(n20585), .A2(\xmem_data[30][7] ), .B1(n24546), .B2(
        \xmem_data[31][7] ), .ZN(n5669) );
  AND4_X1 U9019 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n5680)
         );
  BUF_X1 U9020 ( .A(n13469), .Z(n20787) );
  AOI22_X1 U9021 ( .A1(n23740), .A2(\xmem_data[16][7] ), .B1(n20787), .B2(
        \xmem_data[17][7] ), .ZN(n5673) );
  INV_X1 U9022 ( .A(n5673), .ZN(n5678) );
  AOI22_X1 U9023 ( .A1(n28083), .A2(\xmem_data[18][7] ), .B1(n30550), .B2(
        \xmem_data[19][7] ), .ZN(n5676) );
  AOI22_X1 U9024 ( .A1(n25422), .A2(\xmem_data[22][7] ), .B1(n3357), .B2(
        \xmem_data[23][7] ), .ZN(n5675) );
  NAND2_X1 U9025 ( .A1(n25417), .A2(\xmem_data[20][7] ), .ZN(n5674) );
  NAND3_X1 U9026 ( .A1(n5676), .A2(n5675), .A3(n5674), .ZN(n5677) );
  NOR2_X1 U9027 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  NAND2_X1 U9028 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  NOR2_X1 U9029 ( .A1(n5681), .A2(n3874), .ZN(n5694) );
  AOI22_X1 U9030 ( .A1(n30950), .A2(\xmem_data[0][7] ), .B1(n29318), .B2(
        \xmem_data[1][7] ), .ZN(n5685) );
  AOI22_X1 U9031 ( .A1(n29100), .A2(\xmem_data[2][7] ), .B1(n27951), .B2(
        \xmem_data[3][7] ), .ZN(n5684) );
  BUF_X1 U9032 ( .A(n14914), .Z(n20781) );
  AOI22_X1 U9033 ( .A1(n3271), .A2(\xmem_data[4][7] ), .B1(n20781), .B2(
        \xmem_data[5][7] ), .ZN(n5683) );
  AOI22_X1 U9034 ( .A1(n20782), .A2(\xmem_data[6][7] ), .B1(n28979), .B2(
        \xmem_data[7][7] ), .ZN(n5682) );
  BUF_X1 U9035 ( .A(n13420), .Z(n20770) );
  AOI22_X1 U9036 ( .A1(n20770), .A2(\xmem_data[8][7] ), .B1(n20769), .B2(
        \xmem_data[9][7] ), .ZN(n5689) );
  AOI22_X1 U9037 ( .A1(n25354), .A2(\xmem_data[14][7] ), .B1(n3217), .B2(
        \xmem_data[15][7] ), .ZN(n5688) );
  AOI22_X1 U9038 ( .A1(n30588), .A2(\xmem_data[10][7] ), .B1(n27958), .B2(
        \xmem_data[11][7] ), .ZN(n5687) );
  AOI22_X1 U9039 ( .A1(n3434), .A2(\xmem_data[12][7] ), .B1(n25687), .B2(
        \xmem_data[13][7] ), .ZN(n5686) );
  NAND4_X1 U9040 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n5690)
         );
  NOR2_X1 U9041 ( .A1(n3978), .A2(n5690), .ZN(n5693) );
  INV_X1 U9042 ( .A(n5692), .ZN(n8227) );
  AOI22_X1 U9043 ( .A1(load_xaddr_val[5]), .A2(n8227), .B1(n5692), .B2(n39041), 
        .ZN(n5759) );
  AOI21_X1 U9044 ( .B1(load_xaddr_val[6]), .B2(n4499), .A(n20311), .ZN(n14909)
         );
  AOI22_X1 U9045 ( .A1(n5692), .A2(n39040), .B1(n14909), .B2(n8227), .ZN(n5737) );
  NOR2_X1 U9046 ( .A1(n5759), .A2(n5737), .ZN(n20795) );
  INV_X1 U9047 ( .A(n20795), .ZN(n20188) );
  AOI21_X1 U9048 ( .B1(n5694), .B2(n5693), .A(n20188), .ZN(n5695) );
  INV_X1 U9049 ( .A(n5695), .ZN(n5765) );
  BUF_X1 U9050 ( .A(n14971), .Z(n20815) );
  BUF_X1 U9051 ( .A(n13452), .Z(n20814) );
  AOI22_X1 U9052 ( .A1(n20815), .A2(\xmem_data[64][7] ), .B1(n20814), .B2(
        \xmem_data[65][7] ), .ZN(n5699) );
  BUF_X1 U9053 ( .A(n14882), .Z(n20816) );
  AOI22_X1 U9054 ( .A1(n17002), .A2(\xmem_data[66][7] ), .B1(n28327), .B2(
        \xmem_data[67][7] ), .ZN(n5698) );
  BUF_X1 U9055 ( .A(n14974), .Z(n20817) );
  AOI22_X1 U9056 ( .A1(n20817), .A2(\xmem_data[68][7] ), .B1(n14883), .B2(
        \xmem_data[69][7] ), .ZN(n5697) );
  BUF_X1 U9057 ( .A(n13486), .Z(n20818) );
  AOI22_X1 U9058 ( .A1(n20818), .A2(\xmem_data[70][7] ), .B1(n23725), .B2(
        \xmem_data[71][7] ), .ZN(n5696) );
  NAND4_X1 U9059 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n5715)
         );
  BUF_X1 U9060 ( .A(n13420), .Z(n20826) );
  AOI22_X1 U9061 ( .A1(n20826), .A2(\xmem_data[72][7] ), .B1(n30524), .B2(
        \xmem_data[73][7] ), .ZN(n5703) );
  BUF_X1 U9062 ( .A(n31263), .Z(n20827) );
  AOI22_X1 U9063 ( .A1(n20827), .A2(\xmem_data[74][7] ), .B1(n31262), .B2(
        \xmem_data[75][7] ), .ZN(n5702) );
  BUF_X1 U9064 ( .A(n28973), .Z(n20828) );
  AOI22_X1 U9065 ( .A1(n20828), .A2(\xmem_data[76][7] ), .B1(n31347), .B2(
        \xmem_data[77][7] ), .ZN(n5701) );
  AOI22_X1 U9066 ( .A1(n28503), .A2(\xmem_data[78][7] ), .B1(n3218), .B2(
        \xmem_data[79][7] ), .ZN(n5700) );
  NAND4_X1 U9067 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n5714)
         );
  BUF_X1 U9068 ( .A(n14988), .Z(n20805) );
  AOI22_X1 U9069 ( .A1(n20805), .A2(\xmem_data[80][7] ), .B1(n20787), .B2(
        \xmem_data[81][7] ), .ZN(n5707) );
  BUF_X1 U9070 ( .A(n14926), .Z(n20807) );
  BUF_X1 U9071 ( .A(n14927), .Z(n20806) );
  AOI22_X1 U9072 ( .A1(n20807), .A2(\xmem_data[82][7] ), .B1(n20806), .B2(
        \xmem_data[83][7] ), .ZN(n5706) );
  BUF_X1 U9073 ( .A(n14991), .Z(n20808) );
  AOI22_X1 U9074 ( .A1(n20808), .A2(\xmem_data[84][7] ), .B1(n25514), .B2(
        \xmem_data[85][7] ), .ZN(n5705) );
  BUF_X1 U9075 ( .A(n31276), .Z(n20809) );
  AOI22_X1 U9076 ( .A1(n20809), .A2(\xmem_data[86][7] ), .B1(n20546), .B2(
        \xmem_data[87][7] ), .ZN(n5704) );
  NAND4_X1 U9077 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n5713)
         );
  BUF_X1 U9078 ( .A(n14997), .Z(n20799) );
  AOI22_X1 U9079 ( .A1(n20799), .A2(\xmem_data[88][7] ), .B1(n27513), .B2(
        \xmem_data[89][7] ), .ZN(n5711) );
  BUF_X1 U9080 ( .A(n14935), .Z(n20798) );
  AOI22_X1 U9081 ( .A1(n30514), .A2(\xmem_data[90][7] ), .B1(n20798), .B2(
        \xmem_data[91][7] ), .ZN(n5710) );
  AOI22_X1 U9082 ( .A1(n24458), .A2(\xmem_data[92][7] ), .B1(n30542), .B2(
        \xmem_data[93][7] ), .ZN(n5709) );
  BUF_X1 U9083 ( .A(n14937), .Z(n20800) );
  AOI22_X1 U9084 ( .A1(n20800), .A2(\xmem_data[94][7] ), .B1(n25398), .B2(
        \xmem_data[95][7] ), .ZN(n5708) );
  NAND4_X1 U9085 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n5712)
         );
  OR4_X1 U9086 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n5716) );
  INV_X1 U9087 ( .A(n5737), .ZN(n5760) );
  NAND2_X1 U9088 ( .A1(n5716), .A2(n20833), .ZN(n5764) );
  BUF_X1 U9089 ( .A(n14971), .Z(n20730) );
  AOI22_X1 U9090 ( .A1(n20730), .A2(\xmem_data[96][7] ), .B1(n25435), .B2(
        \xmem_data[97][7] ), .ZN(n5720) );
  BUF_X1 U9091 ( .A(n14881), .Z(n20731) );
  AOI22_X1 U9092 ( .A1(n20731), .A2(\xmem_data[98][7] ), .B1(n28327), .B2(
        \xmem_data[99][7] ), .ZN(n5719) );
  BUF_X1 U9093 ( .A(n14974), .Z(n20732) );
  AOI22_X1 U9094 ( .A1(n20732), .A2(\xmem_data[100][7] ), .B1(n28062), .B2(
        \xmem_data[101][7] ), .ZN(n5718) );
  BUF_X1 U9095 ( .A(n14981), .Z(n20733) );
  AOI22_X1 U9096 ( .A1(n20734), .A2(\xmem_data[102][7] ), .B1(n20733), .B2(
        \xmem_data[103][7] ), .ZN(n5717) );
  NAND4_X1 U9097 ( .A1(n5720), .A2(n5719), .A3(n5718), .A4(n5717), .ZN(n5736)
         );
  BUF_X1 U9098 ( .A(n13420), .Z(n20708) );
  BUF_X1 U9099 ( .A(n10456), .Z(n20707) );
  AOI22_X1 U9100 ( .A1(n20708), .A2(\xmem_data[104][7] ), .B1(n20707), .B2(
        \xmem_data[105][7] ), .ZN(n5724) );
  BUF_X1 U9101 ( .A(n31263), .Z(n20710) );
  BUF_X1 U9102 ( .A(n28947), .Z(n20709) );
  AOI22_X1 U9103 ( .A1(n20710), .A2(\xmem_data[106][7] ), .B1(n20709), .B2(
        \xmem_data[107][7] ), .ZN(n5723) );
  BUF_X1 U9104 ( .A(n13468), .Z(n20711) );
  AOI22_X1 U9105 ( .A1(n3382), .A2(\xmem_data[108][7] ), .B1(n20711), .B2(
        \xmem_data[109][7] ), .ZN(n5722) );
  AOI22_X1 U9106 ( .A1(n20518), .A2(\xmem_data[110][7] ), .B1(n3217), .B2(
        \xmem_data[111][7] ), .ZN(n5721) );
  NAND4_X1 U9107 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n5735)
         );
  BUF_X1 U9108 ( .A(n14988), .Z(n20724) );
  AOI22_X1 U9109 ( .A1(n20724), .A2(\xmem_data[112][7] ), .B1(n20723), .B2(
        \xmem_data[113][7] ), .ZN(n5728) );
  AOI22_X1 U9110 ( .A1(n20725), .A2(\xmem_data[114][7] ), .B1(n27550), .B2(
        \xmem_data[115][7] ), .ZN(n5727) );
  AOI22_X1 U9111 ( .A1(n29706), .A2(\xmem_data[116][7] ), .B1(n25450), .B2(
        \xmem_data[117][7] ), .ZN(n5726) );
  AOI22_X1 U9112 ( .A1(n27447), .A2(\xmem_data[118][7] ), .B1(n27863), .B2(
        \xmem_data[119][7] ), .ZN(n5725) );
  NAND4_X1 U9113 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n5734)
         );
  BUF_X1 U9114 ( .A(n14997), .Z(n20716) );
  AOI22_X1 U9115 ( .A1(n20716), .A2(\xmem_data[120][7] ), .B1(n24212), .B2(
        \xmem_data[121][7] ), .ZN(n5732) );
  BUF_X1 U9116 ( .A(n14935), .Z(n20717) );
  AOI22_X1 U9117 ( .A1(n28980), .A2(\xmem_data[122][7] ), .B1(n20717), .B2(
        \xmem_data[123][7] ), .ZN(n5731) );
  BUF_X1 U9118 ( .A(n29187), .Z(n20718) );
  AOI22_X1 U9119 ( .A1(n23795), .A2(\xmem_data[124][7] ), .B1(n30542), .B2(
        \xmem_data[125][7] ), .ZN(n5730) );
  AOI22_X1 U9120 ( .A1(n21007), .A2(\xmem_data[126][7] ), .B1(n28427), .B2(
        \xmem_data[127][7] ), .ZN(n5729) );
  NAND4_X1 U9121 ( .A1(n5732), .A2(n5731), .A3(n5730), .A4(n5729), .ZN(n5733)
         );
  OR4_X1 U9122 ( .A1(n5736), .A2(n5735), .A3(n5734), .A4(n5733), .ZN(n5738) );
  AND2_X1 U9123 ( .A1(n5759), .A2(n5737), .ZN(n20742) );
  NAND2_X1 U9124 ( .A1(n5738), .A2(n20742), .ZN(n5763) );
  AOI22_X1 U9125 ( .A1(n20815), .A2(\xmem_data[32][7] ), .B1(n20814), .B2(
        \xmem_data[33][7] ), .ZN(n5742) );
  AOI22_X1 U9126 ( .A1(n27462), .A2(\xmem_data[34][7] ), .B1(n27951), .B2(
        \xmem_data[35][7] ), .ZN(n5741) );
  AOI22_X1 U9127 ( .A1(n20817), .A2(\xmem_data[36][7] ), .B1(n24521), .B2(
        \xmem_data[37][7] ), .ZN(n5740) );
  AOI22_X1 U9128 ( .A1(n20818), .A2(\xmem_data[38][7] ), .B1(n27526), .B2(
        \xmem_data[39][7] ), .ZN(n5739) );
  NAND4_X1 U9129 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n5758)
         );
  AOI22_X1 U9130 ( .A1(n20826), .A2(\xmem_data[40][7] ), .B1(n30524), .B2(
        \xmem_data[41][7] ), .ZN(n5746) );
  AOI22_X1 U9131 ( .A1(n20827), .A2(\xmem_data[42][7] ), .B1(n30861), .B2(
        \xmem_data[43][7] ), .ZN(n5745) );
  AOI22_X1 U9132 ( .A1(n20828), .A2(\xmem_data[44][7] ), .B1(n22753), .B2(
        \xmem_data[45][7] ), .ZN(n5744) );
  AOI22_X1 U9133 ( .A1(n25413), .A2(\xmem_data[46][7] ), .B1(n3220), .B2(
        \xmem_data[47][7] ), .ZN(n5743) );
  NAND4_X1 U9134 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n5757)
         );
  AOI22_X1 U9135 ( .A1(n20805), .A2(\xmem_data[48][7] ), .B1(n20598), .B2(
        \xmem_data[49][7] ), .ZN(n5750) );
  AOI22_X1 U9136 ( .A1(n20807), .A2(\xmem_data[50][7] ), .B1(n20806), .B2(
        \xmem_data[51][7] ), .ZN(n5749) );
  AOI22_X1 U9137 ( .A1(n20808), .A2(\xmem_data[52][7] ), .B1(n3231), .B2(
        \xmem_data[53][7] ), .ZN(n5748) );
  AOI22_X1 U9138 ( .A1(n20809), .A2(\xmem_data[54][7] ), .B1(n25481), .B2(
        \xmem_data[55][7] ), .ZN(n5747) );
  NAND4_X1 U9139 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n5756)
         );
  AOI22_X1 U9140 ( .A1(n20799), .A2(\xmem_data[56][7] ), .B1(n22675), .B2(
        \xmem_data[57][7] ), .ZN(n5754) );
  AOI22_X1 U9141 ( .A1(n28334), .A2(\xmem_data[58][7] ), .B1(n20798), .B2(
        \xmem_data[59][7] ), .ZN(n5753) );
  AOI22_X1 U9142 ( .A1(n25519), .A2(\xmem_data[60][7] ), .B1(n27516), .B2(
        \xmem_data[61][7] ), .ZN(n5752) );
  AOI22_X1 U9143 ( .A1(n20800), .A2(\xmem_data[62][7] ), .B1(n16989), .B2(
        \xmem_data[63][7] ), .ZN(n5751) );
  NAND4_X1 U9144 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n5755)
         );
  OR4_X1 U9145 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n5761) );
  NAND2_X1 U9146 ( .A1(n5761), .A2(n20765), .ZN(n5762) );
  NAND4_X1 U9147 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n35399)
         );
  XNOR2_X1 U9148 ( .A(n35399), .B(\fmem_data[28][3] ), .ZN(n30379) );
  INV_X1 U9149 ( .A(n5766), .ZN(n11341) );
  INV_X1 U9150 ( .A(n5767), .ZN(n5768) );
  AOI22_X1 U9151 ( .A1(n37191), .A2(n5768), .B1(n5767), .B2(n4499), .ZN(n5862)
         );
  NAND2_X1 U9152 ( .A1(n37191), .A2(n5768), .ZN(n5769) );
  XOR2_X1 U9153 ( .A(n39040), .B(n5769), .Z(n5838) );
  BUF_X1 U9154 ( .A(n14988), .Z(n31368) );
  BUF_X1 U9155 ( .A(n14925), .Z(n31367) );
  AOI22_X1 U9156 ( .A1(n31368), .A2(\xmem_data[96][3] ), .B1(n31367), .B2(
        \xmem_data[97][3] ), .ZN(n5773) );
  AOI22_X1 U9157 ( .A1(n27904), .A2(\xmem_data[98][3] ), .B1(n22669), .B2(
        \xmem_data[99][3] ), .ZN(n5772) );
  AOI22_X1 U9158 ( .A1(n3126), .A2(\xmem_data[100][3] ), .B1(n29103), .B2(
        \xmem_data[101][3] ), .ZN(n5771) );
  AOI22_X1 U9159 ( .A1(n28972), .A2(\xmem_data[102][3] ), .B1(n3358), .B2(
        \xmem_data[103][3] ), .ZN(n5770) );
  NAND4_X1 U9160 ( .A1(n5773), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n5789)
         );
  BUF_X1 U9161 ( .A(n14997), .Z(n31353) );
  AOI22_X1 U9162 ( .A1(n31353), .A2(\xmem_data[104][3] ), .B1(n24159), .B2(
        \xmem_data[105][3] ), .ZN(n5777) );
  AOI22_X1 U9163 ( .A1(n3176), .A2(\xmem_data[106][3] ), .B1(n29309), .B2(
        \xmem_data[107][3] ), .ZN(n5776) );
  BUF_X1 U9164 ( .A(n3464), .Z(n31354) );
  AOI22_X1 U9165 ( .A1(n30948), .A2(\xmem_data[108][3] ), .B1(n20586), .B2(
        \xmem_data[109][3] ), .ZN(n5775) );
  BUF_X1 U9166 ( .A(n13415), .Z(n31355) );
  AOI22_X1 U9167 ( .A1(n31330), .A2(\xmem_data[110][3] ), .B1(n31355), .B2(
        \xmem_data[111][3] ), .ZN(n5774) );
  NAND4_X1 U9168 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n5788)
         );
  BUF_X1 U9169 ( .A(n13452), .Z(n31360) );
  AOI22_X1 U9170 ( .A1(n30872), .A2(\xmem_data[112][3] ), .B1(n31360), .B2(
        \xmem_data[113][3] ), .ZN(n5781) );
  BUF_X1 U9171 ( .A(n14973), .Z(n31361) );
  AOI22_X1 U9172 ( .A1(n30557), .A2(\xmem_data[114][3] ), .B1(n31361), .B2(
        \xmem_data[115][3] ), .ZN(n5780) );
  BUF_X1 U9173 ( .A(n14914), .Z(n31362) );
  AOI22_X1 U9174 ( .A1(n29379), .A2(\xmem_data[116][3] ), .B1(n31362), .B2(
        \xmem_data[117][3] ), .ZN(n5779) );
  AOI22_X1 U9175 ( .A1(n27847), .A2(\xmem_data[118][3] ), .B1(n22751), .B2(
        \xmem_data[119][3] ), .ZN(n5778) );
  NAND4_X1 U9176 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n5787)
         );
  BUF_X1 U9177 ( .A(n13420), .Z(n31345) );
  BUF_X1 U9178 ( .A(n13487), .Z(n31344) );
  AOI22_X1 U9179 ( .A1(n31345), .A2(\xmem_data[120][3] ), .B1(n31344), .B2(
        \xmem_data[121][3] ), .ZN(n5785) );
  BUF_X1 U9180 ( .A(n28947), .Z(n31346) );
  AOI22_X1 U9181 ( .A1(n21061), .A2(\xmem_data[122][3] ), .B1(n31346), .B2(
        \xmem_data[123][3] ), .ZN(n5784) );
  AOI22_X1 U9182 ( .A1(n28677), .A2(\xmem_data[124][3] ), .B1(n31347), .B2(
        \xmem_data[125][3] ), .ZN(n5783) );
  BUF_X1 U9183 ( .A(n29064), .Z(n31348) );
  AOI22_X1 U9184 ( .A1(n31348), .A2(\xmem_data[126][3] ), .B1(n3222), .B2(
        \xmem_data[127][3] ), .ZN(n5782) );
  NAND4_X1 U9185 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5786)
         );
  OR4_X1 U9186 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n5812) );
  INV_X1 U9187 ( .A(n5838), .ZN(n5863) );
  NOR2_X1 U9188 ( .A1(n5862), .A2(n5863), .ZN(n31342) );
  AOI22_X1 U9189 ( .A1(n31368), .A2(\xmem_data[64][3] ), .B1(n31367), .B2(
        \xmem_data[65][3] ), .ZN(n5793) );
  AOI22_X1 U9190 ( .A1(n29289), .A2(\xmem_data[66][3] ), .B1(n21068), .B2(
        \xmem_data[67][3] ), .ZN(n5792) );
  AOI22_X1 U9191 ( .A1(n29762), .A2(\xmem_data[68][3] ), .B1(n25450), .B2(
        \xmem_data[69][3] ), .ZN(n5791) );
  AOI22_X1 U9192 ( .A1(n27508), .A2(\xmem_data[70][3] ), .B1(n3357), .B2(
        \xmem_data[71][3] ), .ZN(n5790) );
  NAND4_X1 U9193 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n5810)
         );
  AOI22_X1 U9194 ( .A1(n31353), .A2(\xmem_data[72][3] ), .B1(n25423), .B2(
        \xmem_data[73][3] ), .ZN(n5797) );
  AOI22_X1 U9195 ( .A1(n28980), .A2(\xmem_data[74][3] ), .B1(n29271), .B2(
        \xmem_data[75][3] ), .ZN(n5796) );
  AOI22_X1 U9196 ( .A1(n21005), .A2(\xmem_data[76][3] ), .B1(n20543), .B2(
        \xmem_data[77][3] ), .ZN(n5795) );
  AOI22_X1 U9197 ( .A1(n25573), .A2(\xmem_data[78][3] ), .B1(n31355), .B2(
        \xmem_data[79][3] ), .ZN(n5794) );
  NAND4_X1 U9198 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n5809)
         );
  AOI22_X1 U9199 ( .A1(n14971), .A2(\xmem_data[80][3] ), .B1(n31360), .B2(
        \xmem_data[81][3] ), .ZN(n5801) );
  AOI22_X1 U9200 ( .A1(n28428), .A2(\xmem_data[82][3] ), .B1(n31361), .B2(
        \xmem_data[83][3] ), .ZN(n5800) );
  AOI22_X1 U9201 ( .A1(n17004), .A2(\xmem_data[84][3] ), .B1(n31362), .B2(
        \xmem_data[85][3] ), .ZN(n5799) );
  AOI22_X1 U9202 ( .A1(n22684), .A2(\xmem_data[86][3] ), .B1(n17003), .B2(
        \xmem_data[87][3] ), .ZN(n5798) );
  NAND4_X1 U9203 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n5808)
         );
  AOI22_X1 U9204 ( .A1(n31345), .A2(\xmem_data[88][3] ), .B1(n31344), .B2(
        \xmem_data[89][3] ), .ZN(n5806) );
  AOI22_X1 U9205 ( .A1(n17056), .A2(\xmem_data[90][3] ), .B1(n31346), .B2(
        \xmem_data[91][3] ), .ZN(n5805) );
  AOI22_X1 U9206 ( .A1(n25725), .A2(\xmem_data[92][3] ), .B1(n31347), .B2(
        \xmem_data[93][3] ), .ZN(n5804) );
  AND2_X1 U9207 ( .A1(n3221), .A2(\xmem_data[95][3] ), .ZN(n5802) );
  AOI21_X1 U9208 ( .B1(n31348), .B2(\xmem_data[94][3] ), .A(n5802), .ZN(n5803)
         );
  NAND4_X1 U9209 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n5807)
         );
  OR4_X1 U9210 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n5811) );
  AOI22_X1 U9211 ( .A1(n31376), .A2(n5812), .B1(n31342), .B2(n5811), .ZN(n5867) );
  AOI22_X1 U9212 ( .A1(n3335), .A2(\xmem_data[28][3] ), .B1(n3247), .B2(
        \xmem_data[29][3] ), .ZN(n5814) );
  BUF_X1 U9213 ( .A(n13457), .Z(n31261) );
  AOI22_X1 U9214 ( .A1(n28470), .A2(\xmem_data[30][3] ), .B1(n3219), .B2(
        \xmem_data[31][3] ), .ZN(n5821) );
  BUF_X1 U9215 ( .A(n28947), .Z(n31262) );
  AOI22_X1 U9216 ( .A1(n3380), .A2(\xmem_data[26][3] ), .B1(n31262), .B2(
        \xmem_data[27][3] ), .ZN(n5820) );
  BUF_X1 U9217 ( .A(n14971), .Z(n31255) );
  BUF_X1 U9218 ( .A(n13452), .Z(n31254) );
  AOI22_X1 U9219 ( .A1(n31255), .A2(\xmem_data[16][3] ), .B1(n31254), .B2(
        \xmem_data[17][3] ), .ZN(n5819) );
  AOI22_X1 U9220 ( .A1(n17002), .A2(\xmem_data[18][3] ), .B1(n25364), .B2(
        \xmem_data[19][3] ), .ZN(n5818) );
  AOI22_X1 U9221 ( .A1(n23724), .A2(\xmem_data[20][3] ), .B1(n29245), .B2(
        \xmem_data[21][3] ), .ZN(n5817) );
  BUF_X1 U9222 ( .A(n14919), .Z(n31256) );
  AOI22_X1 U9223 ( .A1(n21058), .A2(\xmem_data[22][3] ), .B1(n31256), .B2(
        \xmem_data[23][3] ), .ZN(n5816) );
  NAND4_X1 U9224 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n3755), .ZN(n5837)
         );
  AOI22_X1 U9225 ( .A1(n27708), .A2(\xmem_data[0][3] ), .B1(n20787), .B2(
        \xmem_data[1][3] ), .ZN(n5829) );
  BUF_X1 U9226 ( .A(n14927), .Z(n31275) );
  AOI22_X1 U9227 ( .A1(n30883), .A2(\xmem_data[2][3] ), .B1(n31275), .B2(
        \xmem_data[3][3] ), .ZN(n5823) );
  INV_X1 U9228 ( .A(n5823), .ZN(n5827) );
  AOI22_X1 U9229 ( .A1(n31276), .A2(\xmem_data[6][3] ), .B1(n28415), .B2(
        \xmem_data[7][3] ), .ZN(n5825) );
  NAND2_X1 U9230 ( .A1(n29157), .A2(\xmem_data[4][3] ), .ZN(n5824) );
  NAND2_X1 U9231 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  NOR2_X1 U9232 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND2_X1 U9233 ( .A1(n5829), .A2(n5828), .ZN(n5835) );
  AOI22_X1 U9234 ( .A1(n27944), .A2(\xmem_data[8][3] ), .B1(n20958), .B2(
        \xmem_data[9][3] ), .ZN(n5833) );
  AOI22_X1 U9235 ( .A1(n31268), .A2(\xmem_data[10][3] ), .B1(n22703), .B2(
        \xmem_data[11][3] ), .ZN(n5832) );
  BUF_X1 U9236 ( .A(n14936), .Z(n31269) );
  AOI22_X1 U9237 ( .A1(n3465), .A2(\xmem_data[12][3] ), .B1(n31269), .B2(
        \xmem_data[13][3] ), .ZN(n5831) );
  BUF_X1 U9238 ( .A(n14912), .Z(n31270) );
  AOI22_X1 U9239 ( .A1(n22676), .A2(\xmem_data[14][3] ), .B1(n31270), .B2(
        \xmem_data[15][3] ), .ZN(n5830) );
  NAND4_X1 U9240 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n5834)
         );
  OR2_X1 U9241 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NOR2_X1 U9242 ( .A1(n5837), .A2(n5836), .ZN(n5840) );
  BUF_X1 U9243 ( .A(n14928), .Z(n31252) );
  NAND2_X1 U9244 ( .A1(n28510), .A2(\xmem_data[5][3] ), .ZN(n5839) );
  NOR2_X1 U9245 ( .A1(n5862), .A2(n5838), .ZN(n31284) );
  INV_X1 U9246 ( .A(n31284), .ZN(n31041) );
  AOI21_X1 U9247 ( .B1(n5840), .B2(n5839), .A(n31041), .ZN(n5841) );
  INV_X1 U9248 ( .A(n5841), .ZN(n5866) );
  AOI22_X1 U9249 ( .A1(n21067), .A2(\xmem_data[32][3] ), .B1(n23739), .B2(
        \xmem_data[33][3] ), .ZN(n5845) );
  AOI22_X1 U9250 ( .A1(n30606), .A2(\xmem_data[34][3] ), .B1(n28372), .B2(
        \xmem_data[35][3] ), .ZN(n5844) );
  AOI22_X1 U9251 ( .A1(n3375), .A2(\xmem_data[36][3] ), .B1(n29045), .B2(
        \xmem_data[37][3] ), .ZN(n5843) );
  BUF_X1 U9252 ( .A(n25604), .Z(n31321) );
  AOI22_X1 U9253 ( .A1(n31321), .A2(\xmem_data[38][3] ), .B1(n20546), .B2(
        \xmem_data[39][3] ), .ZN(n5842) );
  NAND4_X1 U9254 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n5861)
         );
  BUF_X1 U9255 ( .A(n14997), .Z(n31327) );
  BUF_X1 U9256 ( .A(n13435), .Z(n31326) );
  AOI22_X1 U9257 ( .A1(n31327), .A2(\xmem_data[40][3] ), .B1(n31326), .B2(
        \xmem_data[41][3] ), .ZN(n5849) );
  AOI22_X1 U9258 ( .A1(n20495), .A2(\xmem_data[42][3] ), .B1(n29271), .B2(
        \xmem_data[43][3] ), .ZN(n5848) );
  BUF_X1 U9259 ( .A(n3464), .Z(n31328) );
  AOI22_X1 U9260 ( .A1(n31328), .A2(\xmem_data[44][3] ), .B1(n27516), .B2(
        \xmem_data[45][3] ), .ZN(n5847) );
  BUF_X1 U9261 ( .A(n14937), .Z(n31330) );
  BUF_X1 U9262 ( .A(n13415), .Z(n31329) );
  AOI22_X1 U9263 ( .A1(n31330), .A2(\xmem_data[46][3] ), .B1(n31329), .B2(
        \xmem_data[47][3] ), .ZN(n5846) );
  NAND4_X1 U9264 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n5860)
         );
  AOI22_X1 U9265 ( .A1(n29410), .A2(\xmem_data[48][3] ), .B1(n30515), .B2(
        \xmem_data[49][3] ), .ZN(n5853) );
  AOI22_X1 U9266 ( .A1(n27974), .A2(\xmem_data[50][3] ), .B1(n25581), .B2(
        \xmem_data[51][3] ), .ZN(n5852) );
  BUF_X1 U9267 ( .A(n14974), .Z(n31315) );
  BUF_X1 U9268 ( .A(n14914), .Z(n31314) );
  AOI22_X1 U9269 ( .A1(n31315), .A2(\xmem_data[52][3] ), .B1(n31314), .B2(
        \xmem_data[53][3] ), .ZN(n5851) );
  BUF_X1 U9270 ( .A(n13486), .Z(n31316) );
  AOI22_X1 U9271 ( .A1(n31316), .A2(\xmem_data[54][3] ), .B1(n17003), .B2(
        \xmem_data[55][3] ), .ZN(n5850) );
  NAND4_X1 U9272 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n5859)
         );
  BUF_X1 U9273 ( .A(n13127), .Z(n31308) );
  AOI22_X1 U9274 ( .A1(n31308), .A2(\xmem_data[56][3] ), .B1(n28329), .B2(
        \xmem_data[57][3] ), .ZN(n5857) );
  BUF_X1 U9275 ( .A(n28974), .Z(n31309) );
  AOI22_X1 U9276 ( .A1(n20986), .A2(\xmem_data[58][3] ), .B1(n31309), .B2(
        \xmem_data[59][3] ), .ZN(n5856) );
  AOI22_X1 U9277 ( .A1(n3449), .A2(\xmem_data[60][3] ), .B1(n14875), .B2(
        \xmem_data[61][3] ), .ZN(n5855) );
  AOI22_X1 U9278 ( .A1(n30503), .A2(\xmem_data[62][3] ), .B1(n3222), .B2(
        \xmem_data[63][3] ), .ZN(n5854) );
  NAND4_X1 U9279 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n5858)
         );
  OR4_X1 U9280 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n5864) );
  AND2_X1 U9281 ( .A1(n5863), .A2(n5862), .ZN(n31340) );
  NAND2_X1 U9282 ( .A1(n5864), .A2(n31340), .ZN(n5865) );
  XOR2_X1 U9283 ( .A(\fmem_data[12][6] ), .B(\fmem_data[12][7] ), .Z(n5868) );
  AOI22_X1 U9284 ( .A1(n27831), .A2(\xmem_data[32][4] ), .B1(n25562), .B2(
        \xmem_data[33][4] ), .ZN(n5872) );
  AOI22_X1 U9285 ( .A1(n20807), .A2(\xmem_data[34][4] ), .B1(n13444), .B2(
        \xmem_data[35][4] ), .ZN(n5871) );
  AOI22_X1 U9286 ( .A1(n3345), .A2(\xmem_data[36][4] ), .B1(n28307), .B2(
        \xmem_data[37][4] ), .ZN(n5870) );
  AOI22_X1 U9287 ( .A1(n31321), .A2(\xmem_data[38][4] ), .B1(n3358), .B2(
        \xmem_data[39][4] ), .ZN(n5869) );
  NAND4_X1 U9288 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n5888)
         );
  AOI22_X1 U9289 ( .A1(n31327), .A2(\xmem_data[40][4] ), .B1(n31326), .B2(
        \xmem_data[41][4] ), .ZN(n5876) );
  AOI22_X1 U9290 ( .A1(n28334), .A2(\xmem_data[42][4] ), .B1(n25606), .B2(
        \xmem_data[43][4] ), .ZN(n5875) );
  AOI22_X1 U9291 ( .A1(n31328), .A2(\xmem_data[44][4] ), .B1(n22677), .B2(
        \xmem_data[45][4] ), .ZN(n5874) );
  AOI22_X1 U9292 ( .A1(n31330), .A2(\xmem_data[46][4] ), .B1(n31329), .B2(
        \xmem_data[47][4] ), .ZN(n5873) );
  NAND4_X1 U9293 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n5887)
         );
  AOI22_X1 U9294 ( .A1(n29439), .A2(\xmem_data[48][4] ), .B1(n24460), .B2(
        \xmem_data[49][4] ), .ZN(n5880) );
  AOI22_X1 U9295 ( .A1(n28493), .A2(\xmem_data[50][4] ), .B1(n3372), .B2(
        \xmem_data[51][4] ), .ZN(n5879) );
  AOI22_X1 U9296 ( .A1(n31315), .A2(\xmem_data[52][4] ), .B1(n31314), .B2(
        \xmem_data[53][4] ), .ZN(n5878) );
  AOI22_X1 U9297 ( .A1(n31316), .A2(\xmem_data[54][4] ), .B1(n17049), .B2(
        \xmem_data[55][4] ), .ZN(n5877) );
  NAND4_X1 U9298 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n5886)
         );
  AOI22_X1 U9299 ( .A1(n31308), .A2(\xmem_data[56][4] ), .B1(n31261), .B2(
        \xmem_data[57][4] ), .ZN(n5884) );
  AOI22_X1 U9300 ( .A1(n27436), .A2(\xmem_data[58][4] ), .B1(n31309), .B2(
        \xmem_data[59][4] ), .ZN(n5883) );
  AOI22_X1 U9301 ( .A1(n28718), .A2(\xmem_data[60][4] ), .B1(n28501), .B2(
        \xmem_data[61][4] ), .ZN(n5882) );
  AOI22_X1 U9302 ( .A1(n28355), .A2(\xmem_data[62][4] ), .B1(n3217), .B2(
        \xmem_data[63][4] ), .ZN(n5881) );
  NAND4_X1 U9303 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n5885)
         );
  OR4_X1 U9304 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n5889) );
  AND2_X1 U9305 ( .A1(n5889), .A2(n31340), .ZN(n5959) );
  AOI22_X1 U9306 ( .A1(n31353), .A2(\xmem_data[104][4] ), .B1(n20958), .B2(
        \xmem_data[105][4] ), .ZN(n5893) );
  AOI22_X1 U9307 ( .A1(n16986), .A2(\xmem_data[106][4] ), .B1(n20798), .B2(
        \xmem_data[107][4] ), .ZN(n5892) );
  AOI22_X1 U9308 ( .A1(n27455), .A2(\xmem_data[108][4] ), .B1(n29188), .B2(
        \xmem_data[109][4] ), .ZN(n5891) );
  AOI22_X1 U9309 ( .A1(n28337), .A2(\xmem_data[110][4] ), .B1(n31355), .B2(
        \xmem_data[111][4] ), .ZN(n5890) );
  NAND4_X1 U9310 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n5904)
         );
  AOI22_X1 U9311 ( .A1(n29239), .A2(\xmem_data[112][4] ), .B1(n31360), .B2(
        \xmem_data[113][4] ), .ZN(n5897) );
  AOI22_X1 U9312 ( .A1(n25575), .A2(\xmem_data[114][4] ), .B1(n31361), .B2(
        \xmem_data[115][4] ), .ZN(n5896) );
  AOI22_X1 U9313 ( .A1(n3307), .A2(\xmem_data[116][4] ), .B1(n31362), .B2(
        \xmem_data[117][4] ), .ZN(n5895) );
  AOI22_X1 U9314 ( .A1(n3172), .A2(\xmem_data[118][4] ), .B1(n27463), .B2(
        \xmem_data[119][4] ), .ZN(n5894) );
  NAND4_X1 U9315 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n5903)
         );
  AOI22_X1 U9316 ( .A1(n31368), .A2(\xmem_data[96][4] ), .B1(n31367), .B2(
        \xmem_data[97][4] ), .ZN(n5901) );
  AOI22_X1 U9317 ( .A1(n20725), .A2(\xmem_data[98][4] ), .B1(n22669), .B2(
        \xmem_data[99][4] ), .ZN(n5900) );
  AOI22_X1 U9318 ( .A1(n29706), .A2(\xmem_data[100][4] ), .B1(n29103), .B2(
        \xmem_data[101][4] ), .ZN(n5899) );
  AOI22_X1 U9319 ( .A1(n25422), .A2(\xmem_data[102][4] ), .B1(n3357), .B2(
        \xmem_data[103][4] ), .ZN(n5898) );
  NAND4_X1 U9320 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5902)
         );
  OR3_X1 U9321 ( .A1(n5904), .A2(n5903), .A3(n5902), .ZN(n5911) );
  AOI22_X1 U9322 ( .A1(n31345), .A2(\xmem_data[120][4] ), .B1(n31344), .B2(
        \xmem_data[121][4] ), .ZN(n5909) );
  AOI22_X1 U9323 ( .A1(n27925), .A2(\xmem_data[122][4] ), .B1(n31346), .B2(
        \xmem_data[123][4] ), .ZN(n5908) );
  AOI22_X1 U9324 ( .A1(n28164), .A2(\xmem_data[124][4] ), .B1(n31347), .B2(
        \xmem_data[125][4] ), .ZN(n5907) );
  AND2_X1 U9325 ( .A1(n3217), .A2(\xmem_data[127][4] ), .ZN(n5905) );
  AOI21_X1 U9326 ( .B1(n31348), .B2(\xmem_data[126][4] ), .A(n5905), .ZN(n5906) );
  NAND4_X1 U9327 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n5910)
         );
  AOI22_X1 U9328 ( .A1(n24607), .A2(\xmem_data[90][4] ), .B1(n31309), .B2(
        \xmem_data[91][4] ), .ZN(n5915) );
  AOI22_X1 U9329 ( .A1(n31308), .A2(\xmem_data[88][4] ), .B1(n20951), .B2(
        \xmem_data[89][4] ), .ZN(n5914) );
  AOI22_X1 U9330 ( .A1(n3333), .A2(\xmem_data[92][4] ), .B1(n20568), .B2(
        \xmem_data[93][4] ), .ZN(n5913) );
  AOI22_X1 U9331 ( .A1(n27439), .A2(\xmem_data[94][4] ), .B1(n3221), .B2(
        \xmem_data[95][4] ), .ZN(n5912) );
  NAND4_X1 U9332 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n5932)
         );
  AOI22_X1 U9333 ( .A1(n23777), .A2(\xmem_data[80][4] ), .B1(n30616), .B2(
        \xmem_data[81][4] ), .ZN(n5919) );
  AOI22_X1 U9334 ( .A1(n24190), .A2(\xmem_data[82][4] ), .B1(n28060), .B2(
        \xmem_data[83][4] ), .ZN(n5918) );
  AOI22_X1 U9335 ( .A1(n31315), .A2(\xmem_data[84][4] ), .B1(n31314), .B2(
        \xmem_data[85][4] ), .ZN(n5917) );
  AOI22_X1 U9336 ( .A1(n31316), .A2(\xmem_data[86][4] ), .B1(n28500), .B2(
        \xmem_data[87][4] ), .ZN(n5916) );
  NAND4_X1 U9337 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n5930)
         );
  AOI22_X1 U9338 ( .A1(n28367), .A2(\xmem_data[64][4] ), .B1(n24207), .B2(
        \xmem_data[65][4] ), .ZN(n5923) );
  AOI22_X1 U9339 ( .A1(n23741), .A2(\xmem_data[66][4] ), .B1(n3255), .B2(
        \xmem_data[67][4] ), .ZN(n5922) );
  AOI22_X1 U9340 ( .A1(n30698), .A2(\xmem_data[68][4] ), .B1(n29103), .B2(
        \xmem_data[69][4] ), .ZN(n5921) );
  AOI22_X1 U9341 ( .A1(n31321), .A2(\xmem_data[70][4] ), .B1(n13475), .B2(
        \xmem_data[71][4] ), .ZN(n5920) );
  NAND4_X1 U9342 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n5929)
         );
  AOI22_X1 U9343 ( .A1(n31327), .A2(\xmem_data[72][4] ), .B1(n31326), .B2(
        \xmem_data[73][4] ), .ZN(n5927) );
  AOI22_X1 U9344 ( .A1(n28980), .A2(\xmem_data[74][4] ), .B1(n27536), .B2(
        \xmem_data[75][4] ), .ZN(n5926) );
  AOI22_X1 U9345 ( .A1(n31328), .A2(\xmem_data[76][4] ), .B1(n15000), .B2(
        \xmem_data[77][4] ), .ZN(n5925) );
  AOI22_X1 U9346 ( .A1(n31330), .A2(\xmem_data[78][4] ), .B1(n31329), .B2(
        \xmem_data[79][4] ), .ZN(n5924) );
  NAND4_X1 U9347 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n5928)
         );
  AOI22_X1 U9348 ( .A1(n29725), .A2(\xmem_data[24][4] ), .B1(n31261), .B2(
        \xmem_data[25][4] ), .ZN(n5936) );
  AOI22_X1 U9349 ( .A1(n3380), .A2(\xmem_data[26][4] ), .B1(n31262), .B2(
        \xmem_data[27][4] ), .ZN(n5935) );
  AOI22_X1 U9350 ( .A1(n28164), .A2(\xmem_data[28][4] ), .B1(n25442), .B2(
        \xmem_data[29][4] ), .ZN(n5934) );
  AOI22_X1 U9351 ( .A1(n28318), .A2(\xmem_data[30][4] ), .B1(n3218), .B2(
        \xmem_data[31][4] ), .ZN(n5933) );
  NAND4_X1 U9352 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n5954)
         );
  AOI22_X1 U9353 ( .A1(n29403), .A2(\xmem_data[8][4] ), .B1(n24212), .B2(
        \xmem_data[9][4] ), .ZN(n5940) );
  AOI22_X1 U9354 ( .A1(n31268), .A2(\xmem_data[10][4] ), .B1(n25382), .B2(
        \xmem_data[11][4] ), .ZN(n5939) );
  AOI22_X1 U9355 ( .A1(n29437), .A2(\xmem_data[12][4] ), .B1(n31269), .B2(
        \xmem_data[13][4] ), .ZN(n5938) );
  AOI22_X1 U9356 ( .A1(n25573), .A2(\xmem_data[14][4] ), .B1(n31270), .B2(
        \xmem_data[15][4] ), .ZN(n5937) );
  NAND4_X1 U9357 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n5952)
         );
  AOI22_X1 U9358 ( .A1(n31255), .A2(\xmem_data[16][4] ), .B1(n31254), .B2(
        \xmem_data[17][4] ), .ZN(n5944) );
  AOI22_X1 U9359 ( .A1(n22683), .A2(\xmem_data[18][4] ), .B1(n20506), .B2(
        \xmem_data[19][4] ), .ZN(n5943) );
  AOI22_X1 U9360 ( .A1(n28202), .A2(\xmem_data[20][4] ), .B1(n24622), .B2(
        \xmem_data[21][4] ), .ZN(n5942) );
  AOI22_X1 U9361 ( .A1(n24572), .A2(\xmem_data[22][4] ), .B1(n31256), .B2(
        \xmem_data[23][4] ), .ZN(n5941) );
  NAND4_X1 U9362 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5951)
         );
  AOI22_X1 U9363 ( .A1(n27396), .A2(\xmem_data[4][4] ), .B1(n28343), .B2(
        \xmem_data[5][4] ), .ZN(n5945) );
  INV_X1 U9364 ( .A(n5945), .ZN(n5950) );
  AOI22_X1 U9365 ( .A1(n24438), .A2(\xmem_data[2][4] ), .B1(n31275), .B2(
        \xmem_data[3][4] ), .ZN(n5948) );
  AOI22_X1 U9366 ( .A1(n31276), .A2(\xmem_data[6][4] ), .B1(n3358), .B2(
        \xmem_data[7][4] ), .ZN(n5947) );
  AOI22_X1 U9367 ( .A1(n24632), .A2(\xmem_data[0][4] ), .B1(n20500), .B2(
        \xmem_data[1][4] ), .ZN(n5946) );
  NAND3_X1 U9368 ( .A1(n5948), .A2(n5947), .A3(n5946), .ZN(n5949) );
  NAND3_X1 U9369 ( .A1(n5957), .A2(n5956), .A3(n5955), .ZN(n5958) );
  NAND2_X1 U9370 ( .A1(n24657), .A2(\xmem_data[6][5] ), .ZN(n5984) );
  BUF_X1 U9371 ( .A(n14988), .Z(n24139) );
  AOI22_X1 U9372 ( .A1(n3222), .A2(\xmem_data[0][5] ), .B1(n24139), .B2(
        \xmem_data[1][5] ), .ZN(n5960) );
  INV_X1 U9373 ( .A(n5960), .ZN(n5967) );
  BUF_X1 U9374 ( .A(n13435), .Z(n24132) );
  BUF_X1 U9375 ( .A(n10977), .Z(n24131) );
  AOI22_X1 U9376 ( .A1(n24132), .A2(\xmem_data[10][5] ), .B1(n30891), .B2(
        \xmem_data[11][5] ), .ZN(n5961) );
  INV_X1 U9377 ( .A(n5961), .ZN(n5966) );
  BUF_X1 U9378 ( .A(n14927), .Z(n24140) );
  AOI22_X1 U9379 ( .A1(n24140), .A2(\xmem_data[4][5] ), .B1(n3146), .B2(
        \xmem_data[5][5] ), .ZN(n5964) );
  BUF_X1 U9380 ( .A(n14926), .Z(n24141) );
  AOI22_X1 U9381 ( .A1(n25562), .A2(\xmem_data[2][5] ), .B1(n24141), .B2(
        \xmem_data[3][5] ), .ZN(n5963) );
  NAND2_X1 U9382 ( .A1(n23813), .A2(\xmem_data[7][5] ), .ZN(n5962) );
  NAND3_X1 U9383 ( .A1(n5964), .A2(n5963), .A3(n5962), .ZN(n5965) );
  NOR3_X1 U9384 ( .A1(n5967), .A2(n5966), .A3(n5965), .ZN(n5983) );
  BUF_X1 U9385 ( .A(n14971), .Z(n24115) );
  AOI22_X1 U9386 ( .A1(n31270), .A2(\xmem_data[16][5] ), .B1(n24115), .B2(
        \xmem_data[17][5] ), .ZN(n5971) );
  BUF_X1 U9387 ( .A(n13452), .Z(n24116) );
  AOI22_X1 U9388 ( .A1(n24116), .A2(\xmem_data[18][5] ), .B1(n30899), .B2(
        \xmem_data[19][5] ), .ZN(n5970) );
  BUF_X1 U9389 ( .A(n14973), .Z(n24117) );
  AOI22_X1 U9390 ( .A1(n24117), .A2(\xmem_data[20][5] ), .B1(n28226), .B2(
        \xmem_data[21][5] ), .ZN(n5969) );
  AOI22_X1 U9391 ( .A1(n29245), .A2(\xmem_data[22][5] ), .B1(n24606), .B2(
        \xmem_data[23][5] ), .ZN(n5968) );
  NAND4_X1 U9392 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n5977)
         );
  AOI22_X1 U9393 ( .A1(n17003), .A2(\xmem_data[24][5] ), .B1(n21060), .B2(
        \xmem_data[25][5] ), .ZN(n5975) );
  BUF_X1 U9394 ( .A(n13457), .Z(n24122) );
  AOI22_X1 U9395 ( .A1(n24122), .A2(\xmem_data[26][5] ), .B1(n20827), .B2(
        \xmem_data[27][5] ), .ZN(n5974) );
  AOI22_X1 U9396 ( .A1(n31346), .A2(\xmem_data[28][5] ), .B1(n28677), .B2(
        \xmem_data[29][5] ), .ZN(n5973) );
  AOI22_X1 U9397 ( .A1(n30589), .A2(\xmem_data[30][5] ), .B1(n25508), .B2(
        \xmem_data[31][5] ), .ZN(n5972) );
  NAND4_X1 U9398 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n5976)
         );
  NOR2_X1 U9399 ( .A1(n5977), .A2(n5976), .ZN(n5982) );
  BUF_X1 U9400 ( .A(n10999), .Z(n24130) );
  AOI22_X1 U9401 ( .A1(n24130), .A2(\xmem_data[8][5] ), .B1(n28743), .B2(
        \xmem_data[9][5] ), .ZN(n5980) );
  BUF_X1 U9402 ( .A(n14936), .Z(n24134) );
  BUF_X1 U9403 ( .A(n14937), .Z(n24133) );
  AOI22_X1 U9404 ( .A1(n24134), .A2(\xmem_data[14][5] ), .B1(n24133), .B2(
        \xmem_data[15][5] ), .ZN(n5979) );
  AOI22_X1 U9405 ( .A1(n20584), .A2(\xmem_data[12][5] ), .B1(n28231), .B2(
        \xmem_data[13][5] ), .ZN(n5978) );
  AND3_X1 U9406 ( .A1(n5980), .A2(n5979), .A3(n5978), .ZN(n5981) );
  NAND4_X1 U9407 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n5988)
         );
  OAI21_X1 U9408 ( .B1(n6172), .B2(n5985), .A(n10589), .ZN(n5986) );
  NOR2_X1 U9409 ( .A1(n39041), .A2(n5986), .ZN(n5987) );
  AOI21_X1 U9410 ( .B1(n4499), .B2(n5986), .A(n5987), .ZN(n6067) );
  OAI22_X1 U9411 ( .A1(n5987), .A2(n39040), .B1(n20978), .B2(n5986), .ZN(n6035) );
  NOR2_X1 U9412 ( .A1(n6067), .A2(n6035), .ZN(n17389) );
  NAND2_X1 U9413 ( .A1(n5988), .A2(n17389), .ZN(n6074) );
  AOI22_X1 U9414 ( .A1(n28500), .A2(\xmem_data[56][5] ), .B1(n29298), .B2(
        \xmem_data[57][5] ), .ZN(n5993) );
  AOI22_X1 U9415 ( .A1(n29125), .A2(\xmem_data[58][5] ), .B1(n28354), .B2(
        \xmem_data[59][5] ), .ZN(n5992) );
  AOI22_X1 U9416 ( .A1(n28317), .A2(\xmem_data[60][5] ), .B1(n16980), .B2(
        \xmem_data[61][5] ), .ZN(n5991) );
  AND2_X1 U9417 ( .A1(n30863), .A2(\xmem_data[62][5] ), .ZN(n5989) );
  AOI21_X1 U9418 ( .B1(n28503), .B2(\xmem_data[63][5] ), .A(n5989), .ZN(n5990)
         );
  NAND4_X1 U9419 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n6010)
         );
  AOI22_X1 U9420 ( .A1(n27943), .A2(\xmem_data[40][5] ), .B1(n23792), .B2(
        \xmem_data[41][5] ), .ZN(n5997) );
  AOI22_X1 U9421 ( .A1(n24212), .A2(\xmem_data[42][5] ), .B1(n29310), .B2(
        \xmem_data[43][5] ), .ZN(n5996) );
  BUF_X1 U9422 ( .A(n29187), .Z(n24213) );
  AOI22_X1 U9423 ( .A1(n22703), .A2(\xmem_data[44][5] ), .B1(n27818), .B2(
        \xmem_data[45][5] ), .ZN(n5995) );
  BUF_X1 U9424 ( .A(n13149), .Z(n24214) );
  AOI22_X1 U9425 ( .A1(n3213), .A2(\xmem_data[46][5] ), .B1(n24214), .B2(
        \xmem_data[47][5] ), .ZN(n5994) );
  NAND4_X1 U9426 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n6008)
         );
  BUF_X1 U9427 ( .A(n13415), .Z(n24219) );
  AOI22_X1 U9428 ( .A1(n24219), .A2(\xmem_data[48][5] ), .B1(n20942), .B2(
        \xmem_data[49][5] ), .ZN(n6001) );
  BUF_X1 U9429 ( .A(n13452), .Z(n24221) );
  AOI22_X1 U9430 ( .A1(n24221), .A2(\xmem_data[50][5] ), .B1(n30557), .B2(
        \xmem_data[51][5] ), .ZN(n6000) );
  BUF_X1 U9431 ( .A(n14973), .Z(n24222) );
  AOI22_X1 U9432 ( .A1(n24222), .A2(\xmem_data[52][5] ), .B1(n29246), .B2(
        \xmem_data[53][5] ), .ZN(n5999) );
  BUF_X1 U9433 ( .A(n14883), .Z(n24223) );
  AOI22_X1 U9434 ( .A1(n24223), .A2(\xmem_data[54][5] ), .B1(n25526), .B2(
        \xmem_data[55][5] ), .ZN(n5998) );
  NAND4_X1 U9435 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6007)
         );
  AOI22_X1 U9436 ( .A1(n3220), .A2(\xmem_data[32][5] ), .B1(n29698), .B2(
        \xmem_data[33][5] ), .ZN(n6005) );
  BUF_X1 U9437 ( .A(n14989), .Z(n24207) );
  AOI22_X1 U9438 ( .A1(n24207), .A2(\xmem_data[34][5] ), .B1(n29289), .B2(
        \xmem_data[35][5] ), .ZN(n6004) );
  AOI22_X1 U9439 ( .A1(n30550), .A2(\xmem_data[36][5] ), .B1(n29157), .B2(
        \xmem_data[37][5] ), .ZN(n6003) );
  AOI22_X1 U9440 ( .A1(n25450), .A2(\xmem_data[38][5] ), .B1(n25604), .B2(
        \xmem_data[39][5] ), .ZN(n6002) );
  NAND4_X1 U9441 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n6006)
         );
  OR3_X1 U9442 ( .A1(n6008), .A2(n6007), .A3(n6006), .ZN(n6009) );
  OR2_X1 U9443 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  INV_X1 U9444 ( .A(n6035), .ZN(n6066) );
  AND2_X1 U9445 ( .A1(n6066), .A2(n6067), .ZN(n24236) );
  AOI22_X1 U9446 ( .A1(n24564), .A2(\xmem_data[100][5] ), .B1(n29762), .B2(
        \xmem_data[101][5] ), .ZN(n6014) );
  AOI22_X1 U9447 ( .A1(n20598), .A2(\xmem_data[98][5] ), .B1(n24438), .B2(
        \xmem_data[99][5] ), .ZN(n6013) );
  AOI22_X1 U9448 ( .A1(n3221), .A2(\xmem_data[96][5] ), .B1(n29494), .B2(
        \xmem_data[97][5] ), .ZN(n6012) );
  NAND3_X1 U9449 ( .A1(n6014), .A2(n6013), .A3(n6012), .ZN(n6018) );
  BUF_X1 U9450 ( .A(n10999), .Z(n24158) );
  BUF_X1 U9451 ( .A(n14997), .Z(n24157) );
  AOI22_X1 U9452 ( .A1(n24158), .A2(\xmem_data[104][5] ), .B1(n24157), .B2(
        \xmem_data[105][5] ), .ZN(n6016) );
  AOI22_X1 U9453 ( .A1(n24160), .A2(\xmem_data[108][5] ), .B1(n17018), .B2(
        \xmem_data[109][5] ), .ZN(n6015) );
  NAND2_X1 U9454 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NOR2_X1 U9455 ( .A1(n6018), .A2(n6017), .ZN(n6026) );
  AOI22_X1 U9456 ( .A1(n31329), .A2(\xmem_data[112][5] ), .B1(n20942), .B2(
        \xmem_data[113][5] ), .ZN(n6022) );
  BUF_X1 U9457 ( .A(n13452), .Z(n24165) );
  AOI22_X1 U9458 ( .A1(n24165), .A2(\xmem_data[114][5] ), .B1(n24190), .B2(
        \xmem_data[115][5] ), .ZN(n6021) );
  AOI22_X1 U9459 ( .A1(n21051), .A2(\xmem_data[116][5] ), .B1(n29297), .B2(
        \xmem_data[117][5] ), .ZN(n6020) );
  BUF_X1 U9460 ( .A(n14914), .Z(n24167) );
  BUF_X1 U9461 ( .A(n13486), .Z(n24166) );
  AOI22_X1 U9462 ( .A1(n24167), .A2(\xmem_data[118][5] ), .B1(n24166), .B2(
        \xmem_data[119][5] ), .ZN(n6019) );
  AND2_X1 U9463 ( .A1(n28337), .A2(\xmem_data[111][5] ), .ZN(n6023) );
  AOI21_X1 U9464 ( .B1(n23716), .B2(\xmem_data[110][5] ), .A(n6023), .ZN(n6025) );
  BUF_X1 U9465 ( .A(n13435), .Z(n24159) );
  AOI22_X1 U9466 ( .A1(n24159), .A2(\xmem_data[106][5] ), .B1(n25567), .B2(
        \xmem_data[107][5] ), .ZN(n6024) );
  NAND4_X1 U9467 ( .A1(n6026), .A2(n3806), .A3(n6025), .A4(n6024), .ZN(n6034)
         );
  BUF_X1 U9468 ( .A(n13468), .Z(n24172) );
  AND2_X1 U9469 ( .A1(n24172), .A2(\xmem_data[126][5] ), .ZN(n6027) );
  AOI21_X1 U9470 ( .B1(n30962), .B2(\xmem_data[127][5] ), .A(n6027), .ZN(n6032) );
  AND2_X1 U9471 ( .A1(n28979), .A2(\xmem_data[120][5] ), .ZN(n6028) );
  AOI21_X1 U9472 ( .B1(n20577), .B2(\xmem_data[121][5] ), .A(n6028), .ZN(n6031) );
  AOI22_X1 U9473 ( .A1(n25561), .A2(\xmem_data[124][5] ), .B1(n22728), .B2(
        \xmem_data[125][5] ), .ZN(n6030) );
  AOI22_X1 U9474 ( .A1(n24624), .A2(\xmem_data[122][5] ), .B1(n17056), .B2(
        \xmem_data[123][5] ), .ZN(n6029) );
  NAND4_X1 U9475 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n6033)
         );
  NOR2_X1 U9476 ( .A1(n6034), .A2(n6033), .ZN(n6038) );
  AOI22_X1 U9477 ( .A1(n25450), .A2(\xmem_data[102][5] ), .B1(n28374), .B2(
        \xmem_data[103][5] ), .ZN(n6037) );
  AND2_X1 U9478 ( .A1(n6067), .A2(n6035), .ZN(n24205) );
  INV_X1 U9479 ( .A(n24205), .ZN(n6036) );
  AOI21_X1 U9480 ( .B1(n6038), .B2(n6037), .A(n6036), .ZN(n6039) );
  INV_X1 U9481 ( .A(n6039), .ZN(n6073) );
  AND2_X1 U9482 ( .A1(n23731), .A2(\xmem_data[94][5] ), .ZN(n6040) );
  AOI21_X1 U9483 ( .B1(n28082), .B2(\xmem_data[95][5] ), .A(n6040), .ZN(n6041)
         );
  INV_X1 U9484 ( .A(n6041), .ZN(n6048) );
  AOI22_X1 U9485 ( .A1(n31262), .A2(\xmem_data[92][5] ), .B1(n3245), .B2(
        \xmem_data[93][5] ), .ZN(n6043) );
  AOI22_X1 U9486 ( .A1(n25388), .A2(\xmem_data[90][5] ), .B1(n30588), .B2(
        \xmem_data[91][5] ), .ZN(n6042) );
  NAND2_X1 U9487 ( .A1(n6043), .A2(n6042), .ZN(n6047) );
  AND2_X1 U9488 ( .A1(n20733), .A2(\xmem_data[88][5] ), .ZN(n6044) );
  AOI21_X1 U9489 ( .B1(n20708), .B2(\xmem_data[89][5] ), .A(n6044), .ZN(n6045)
         );
  INV_X1 U9490 ( .A(n6045), .ZN(n6046) );
  NOR3_X1 U9491 ( .A1(n6048), .A2(n6047), .A3(n6046), .ZN(n6070) );
  AOI22_X1 U9492 ( .A1(n31252), .A2(\xmem_data[70][5] ), .B1(n25604), .B2(
        \xmem_data[71][5] ), .ZN(n6049) );
  INV_X1 U9493 ( .A(n6049), .ZN(n6059) );
  AOI22_X1 U9494 ( .A1(n24219), .A2(\xmem_data[80][5] ), .B1(n23722), .B2(
        \xmem_data[81][5] ), .ZN(n6053) );
  AOI22_X1 U9495 ( .A1(n24221), .A2(\xmem_data[82][5] ), .B1(n3326), .B2(
        \xmem_data[83][5] ), .ZN(n6052) );
  AOI22_X1 U9496 ( .A1(n24222), .A2(\xmem_data[84][5] ), .B1(n31315), .B2(
        \xmem_data[85][5] ), .ZN(n6051) );
  AOI22_X1 U9497 ( .A1(n24223), .A2(\xmem_data[86][5] ), .B1(n22719), .B2(
        \xmem_data[87][5] ), .ZN(n6050) );
  NAND4_X1 U9498 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n6058)
         );
  AOI22_X1 U9499 ( .A1(n13444), .A2(\xmem_data[68][5] ), .B1(n16973), .B2(
        \xmem_data[69][5] ), .ZN(n6056) );
  AOI22_X1 U9500 ( .A1(n24207), .A2(\xmem_data[66][5] ), .B1(n3322), .B2(
        \xmem_data[67][5] ), .ZN(n6055) );
  AOI22_X1 U9501 ( .A1(n3221), .A2(\xmem_data[64][5] ), .B1(n25414), .B2(
        \xmem_data[65][5] ), .ZN(n6054) );
  NAND3_X1 U9502 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n6057) );
  OR3_X1 U9503 ( .A1(n6059), .A2(n6058), .A3(n6057), .ZN(n6065) );
  AOI22_X1 U9504 ( .A1(n25481), .A2(\xmem_data[72][5] ), .B1(n23762), .B2(
        \xmem_data[73][5] ), .ZN(n6063) );
  AOI22_X1 U9505 ( .A1(n24212), .A2(\xmem_data[74][5] ), .B1(n13476), .B2(
        \xmem_data[75][5] ), .ZN(n6062) );
  AOI22_X1 U9506 ( .A1(n14999), .A2(\xmem_data[76][5] ), .B1(n3466), .B2(
        \xmem_data[77][5] ), .ZN(n6061) );
  AOI22_X1 U9507 ( .A1(n25460), .A2(\xmem_data[78][5] ), .B1(n24214), .B2(
        \xmem_data[79][5] ), .ZN(n6060) );
  NAND4_X1 U9508 ( .A1(n6063), .A2(n6062), .A3(n6061), .A4(n6060), .ZN(n6064)
         );
  NOR2_X1 U9509 ( .A1(n6065), .A2(n6064), .ZN(n6069) );
  INV_X1 U9510 ( .A(n24204), .ZN(n6068) );
  AOI21_X1 U9511 ( .B1(n6070), .B2(n6069), .A(n6068), .ZN(n6071) );
  INV_X1 U9512 ( .A(n6071), .ZN(n6072) );
  XNOR2_X1 U9513 ( .A(n31668), .B(\fmem_data[13][5] ), .ZN(n24726) );
  XOR2_X1 U9514 ( .A(\fmem_data[13][5] ), .B(\fmem_data[13][4] ), .Z(n6075) );
  AOI22_X1 U9515 ( .A1(n25514), .A2(\xmem_data[6][6] ), .B1(n23813), .B2(
        \xmem_data[7][6] ), .ZN(n6076) );
  INV_X1 U9516 ( .A(n6076), .ZN(n6098) );
  AOI22_X1 U9517 ( .A1(n24130), .A2(\xmem_data[8][6] ), .B1(n30663), .B2(
        \xmem_data[9][6] ), .ZN(n6080) );
  AOI22_X1 U9518 ( .A1(n24132), .A2(\xmem_data[10][6] ), .B1(n25710), .B2(
        \xmem_data[11][6] ), .ZN(n6079) );
  AOI22_X1 U9519 ( .A1(n25572), .A2(\xmem_data[12][6] ), .B1(n28154), .B2(
        \xmem_data[13][6] ), .ZN(n6078) );
  AOI22_X1 U9520 ( .A1(n24134), .A2(\xmem_data[14][6] ), .B1(n24133), .B2(
        \xmem_data[15][6] ), .ZN(n6077) );
  NAND4_X1 U9521 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n6097)
         );
  AOI22_X1 U9522 ( .A1(n3220), .A2(\xmem_data[0][6] ), .B1(n24139), .B2(
        \xmem_data[1][6] ), .ZN(n6083) );
  AOI22_X1 U9523 ( .A1(n24140), .A2(\xmem_data[4][6] ), .B1(n30295), .B2(
        \xmem_data[5][6] ), .ZN(n6082) );
  AOI22_X1 U9524 ( .A1(n24695), .A2(\xmem_data[2][6] ), .B1(n24141), .B2(
        \xmem_data[3][6] ), .ZN(n6081) );
  NAND3_X1 U9525 ( .A1(n6083), .A2(n6082), .A3(n6081), .ZN(n6096) );
  AOI22_X1 U9526 ( .A1(n30589), .A2(\xmem_data[30][6] ), .B1(n28318), .B2(
        \xmem_data[31][6] ), .ZN(n6094) );
  AOI22_X1 U9527 ( .A1(n27958), .A2(\xmem_data[28][6] ), .B1(n3433), .B2(
        \xmem_data[29][6] ), .ZN(n6084) );
  INV_X1 U9528 ( .A(n6084), .ZN(n6087) );
  AOI22_X1 U9529 ( .A1(n24122), .A2(\xmem_data[26][6] ), .B1(n29057), .B2(
        \xmem_data[27][6] ), .ZN(n6085) );
  INV_X1 U9530 ( .A(n6085), .ZN(n6086) );
  NOR2_X1 U9531 ( .A1(n6087), .A2(n6086), .ZN(n6093) );
  AOI22_X1 U9532 ( .A1(n28492), .A2(\xmem_data[16][6] ), .B1(n24115), .B2(
        \xmem_data[17][6] ), .ZN(n6091) );
  AOI22_X1 U9533 ( .A1(n24116), .A2(\xmem_data[18][6] ), .B1(n25717), .B2(
        \xmem_data[19][6] ), .ZN(n6090) );
  AOI22_X1 U9534 ( .A1(n24117), .A2(\xmem_data[20][6] ), .B1(n30645), .B2(
        \xmem_data[21][6] ), .ZN(n6089) );
  AOI22_X1 U9535 ( .A1(n28098), .A2(\xmem_data[22][6] ), .B1(n24606), .B2(
        \xmem_data[23][6] ), .ZN(n6088) );
  AOI22_X1 U9536 ( .A1(n28468), .A2(\xmem_data[24][6] ), .B1(n27717), .B2(
        \xmem_data[25][6] ), .ZN(n6092) );
  NAND4_X1 U9537 ( .A1(n6094), .A2(n6093), .A3(n3796), .A4(n6092), .ZN(n6095)
         );
  NOR4_X1 U9538 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n6166)
         );
  AOI22_X1 U9539 ( .A1(n3220), .A2(\xmem_data[32][6] ), .B1(n29698), .B2(
        \xmem_data[33][6] ), .ZN(n6102) );
  AOI22_X1 U9540 ( .A1(n24207), .A2(\xmem_data[34][6] ), .B1(n21069), .B2(
        \xmem_data[35][6] ), .ZN(n6101) );
  AOI22_X1 U9541 ( .A1(n14890), .A2(\xmem_data[36][6] ), .B1(n29157), .B2(
        \xmem_data[37][6] ), .ZN(n6100) );
  AOI22_X1 U9542 ( .A1(n28007), .A2(\xmem_data[38][6] ), .B1(n25604), .B2(
        \xmem_data[39][6] ), .ZN(n6099) );
  NAND4_X1 U9543 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n6118)
         );
  AOI22_X1 U9544 ( .A1(n20982), .A2(\xmem_data[40][6] ), .B1(n29179), .B2(
        \xmem_data[41][6] ), .ZN(n6106) );
  AOI22_X1 U9545 ( .A1(n24212), .A2(\xmem_data[42][6] ), .B1(n28334), .B2(
        \xmem_data[43][6] ), .ZN(n6105) );
  AOI22_X1 U9546 ( .A1(n20717), .A2(\xmem_data[44][6] ), .B1(n30666), .B2(
        \xmem_data[45][6] ), .ZN(n6104) );
  AOI22_X1 U9547 ( .A1(n28993), .A2(\xmem_data[46][6] ), .B1(n24214), .B2(
        \xmem_data[47][6] ), .ZN(n6103) );
  NAND4_X1 U9548 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n6117)
         );
  AOI22_X1 U9549 ( .A1(n24219), .A2(\xmem_data[48][6] ), .B1(n20730), .B2(
        \xmem_data[49][6] ), .ZN(n6110) );
  AOI22_X1 U9550 ( .A1(n24221), .A2(\xmem_data[50][6] ), .B1(n24548), .B2(
        \xmem_data[51][6] ), .ZN(n6109) );
  AOI22_X1 U9551 ( .A1(n24222), .A2(\xmem_data[52][6] ), .B1(n30311), .B2(
        \xmem_data[53][6] ), .ZN(n6108) );
  AOI22_X1 U9552 ( .A1(n24223), .A2(\xmem_data[54][6] ), .B1(n3171), .B2(
        \xmem_data[55][6] ), .ZN(n6107) );
  NAND4_X1 U9553 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6116)
         );
  AOI22_X1 U9554 ( .A1(n21057), .A2(\xmem_data[56][6] ), .B1(n25628), .B2(
        \xmem_data[57][6] ), .ZN(n6114) );
  AOI22_X1 U9555 ( .A1(n20707), .A2(\xmem_data[58][6] ), .B1(n28038), .B2(
        \xmem_data[59][6] ), .ZN(n6113) );
  AOI22_X1 U9556 ( .A1(n20709), .A2(\xmem_data[60][6] ), .B1(n3413), .B2(
        \xmem_data[61][6] ), .ZN(n6112) );
  AOI22_X1 U9557 ( .A1(n27501), .A2(\xmem_data[62][6] ), .B1(n25413), .B2(
        \xmem_data[63][6] ), .ZN(n6111) );
  NAND4_X1 U9558 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n6115)
         );
  OR4_X1 U9559 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n6119) );
  NAND2_X1 U9560 ( .A1(n6119), .A2(n24236), .ZN(n6165) );
  AOI22_X1 U9561 ( .A1(n3221), .A2(\xmem_data[64][6] ), .B1(n24563), .B2(
        \xmem_data[65][6] ), .ZN(n6123) );
  AOI22_X1 U9562 ( .A1(n24207), .A2(\xmem_data[66][6] ), .B1(n22666), .B2(
        \xmem_data[67][6] ), .ZN(n6122) );
  AOI22_X1 U9563 ( .A1(n17061), .A2(\xmem_data[68][6] ), .B1(n28084), .B2(
        \xmem_data[69][6] ), .ZN(n6121) );
  AOI22_X1 U9564 ( .A1(n24657), .A2(\xmem_data[70][6] ), .B1(n25604), .B2(
        \xmem_data[71][6] ), .ZN(n6120) );
  NAND4_X1 U9565 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n6140)
         );
  AOI22_X1 U9566 ( .A1(n28415), .A2(\xmem_data[72][6] ), .B1(n20587), .B2(
        \xmem_data[73][6] ), .ZN(n6127) );
  AOI22_X1 U9567 ( .A1(n24212), .A2(\xmem_data[74][6] ), .B1(n28334), .B2(
        \xmem_data[75][6] ), .ZN(n6126) );
  AOI22_X1 U9568 ( .A1(n27912), .A2(\xmem_data[76][6] ), .B1(n27945), .B2(
        \xmem_data[77][6] ), .ZN(n6125) );
  AOI22_X1 U9569 ( .A1(n23716), .A2(\xmem_data[78][6] ), .B1(n24214), .B2(
        \xmem_data[79][6] ), .ZN(n6124) );
  NAND4_X1 U9570 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n6139)
         );
  AOI22_X1 U9571 ( .A1(n24219), .A2(\xmem_data[80][6] ), .B1(n30309), .B2(
        \xmem_data[81][6] ), .ZN(n6131) );
  AOI22_X1 U9572 ( .A1(n24221), .A2(\xmem_data[82][6] ), .B1(n17002), .B2(
        \xmem_data[83][6] ), .ZN(n6130) );
  AOI22_X1 U9573 ( .A1(n24222), .A2(\xmem_data[84][6] ), .B1(n29816), .B2(
        \xmem_data[85][6] ), .ZN(n6129) );
  AOI22_X1 U9574 ( .A1(n24223), .A2(\xmem_data[86][6] ), .B1(n25582), .B2(
        \xmem_data[87][6] ), .ZN(n6128) );
  NAND4_X1 U9575 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n6138)
         );
  AOI22_X1 U9576 ( .A1(n28500), .A2(\xmem_data[88][6] ), .B1(n29298), .B2(
        \xmem_data[89][6] ), .ZN(n6136) );
  AOI22_X1 U9577 ( .A1(n30524), .A2(\xmem_data[90][6] ), .B1(n24607), .B2(
        \xmem_data[91][6] ), .ZN(n6135) );
  AOI22_X1 U9578 ( .A1(n24470), .A2(\xmem_data[92][6] ), .B1(n3229), .B2(
        \xmem_data[93][6] ), .ZN(n6134) );
  AND2_X1 U9579 ( .A1(n24439), .A2(\xmem_data[94][6] ), .ZN(n6132) );
  AOI21_X1 U9580 ( .B1(n28355), .B2(\xmem_data[95][6] ), .A(n6132), .ZN(n6133)
         );
  NAND4_X1 U9581 ( .A1(n6136), .A2(n6135), .A3(n6134), .A4(n6133), .ZN(n6137)
         );
  OR4_X1 U9582 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n6163) );
  AOI22_X1 U9583 ( .A1(n29086), .A2(\xmem_data[120][6] ), .B1(n27717), .B2(
        \xmem_data[121][6] ), .ZN(n6145) );
  AOI22_X1 U9584 ( .A1(n22727), .A2(\xmem_data[122][6] ), .B1(n27436), .B2(
        \xmem_data[123][6] ), .ZN(n6144) );
  AOI22_X1 U9585 ( .A1(n27563), .A2(\xmem_data[124][6] ), .B1(n28718), .B2(
        \xmem_data[125][6] ), .ZN(n6143) );
  AND2_X1 U9586 ( .A1(n24172), .A2(\xmem_data[126][6] ), .ZN(n6141) );
  AOI21_X1 U9587 ( .B1(n27502), .B2(\xmem_data[127][6] ), .A(n6141), .ZN(n6142) );
  NAND4_X1 U9588 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n6161)
         );
  AOI22_X1 U9589 ( .A1(n24158), .A2(\xmem_data[104][6] ), .B1(n24157), .B2(
        \xmem_data[105][6] ), .ZN(n6149) );
  AOI22_X1 U9590 ( .A1(n24159), .A2(\xmem_data[106][6] ), .B1(n30514), .B2(
        \xmem_data[107][6] ), .ZN(n6148) );
  AOI22_X1 U9591 ( .A1(n24160), .A2(\xmem_data[108][6] ), .B1(n30303), .B2(
        \xmem_data[109][6] ), .ZN(n6147) );
  AOI22_X1 U9592 ( .A1(n24457), .A2(\xmem_data[110][6] ), .B1(n14937), .B2(
        \xmem_data[111][6] ), .ZN(n6146) );
  NAND4_X1 U9593 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n6160)
         );
  AOI22_X1 U9594 ( .A1(n20940), .A2(\xmem_data[112][6] ), .B1(n25400), .B2(
        \xmem_data[113][6] ), .ZN(n6153) );
  AOI22_X1 U9595 ( .A1(n24165), .A2(\xmem_data[114][6] ), .B1(n24220), .B2(
        \xmem_data[115][6] ), .ZN(n6152) );
  AOI22_X1 U9596 ( .A1(n28494), .A2(\xmem_data[116][6] ), .B1(n20732), .B2(
        \xmem_data[117][6] ), .ZN(n6151) );
  AOI22_X1 U9597 ( .A1(n24167), .A2(\xmem_data[118][6] ), .B1(n24166), .B2(
        \xmem_data[119][6] ), .ZN(n6150) );
  NAND4_X1 U9598 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n6159)
         );
  AOI22_X1 U9599 ( .A1(n3222), .A2(\xmem_data[96][6] ), .B1(n30964), .B2(
        \xmem_data[97][6] ), .ZN(n6157) );
  AOI22_X1 U9600 ( .A1(n27507), .A2(\xmem_data[98][6] ), .B1(n20807), .B2(
        \xmem_data[99][6] ), .ZN(n6156) );
  AOI22_X1 U9601 ( .A1(n13444), .A2(\xmem_data[100][6] ), .B1(n3282), .B2(
        \xmem_data[101][6] ), .ZN(n6155) );
  AOI22_X1 U9602 ( .A1(n28045), .A2(\xmem_data[102][6] ), .B1(n28374), .B2(
        \xmem_data[103][6] ), .ZN(n6154) );
  NAND4_X1 U9603 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n6158)
         );
  OR4_X1 U9604 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n6162) );
  AOI22_X1 U9605 ( .A1(n6163), .A2(n24204), .B1(n6162), .B2(n24205), .ZN(n6164) );
  XNOR2_X1 U9606 ( .A(n31669), .B(\fmem_data[13][5] ), .ZN(n33102) );
  INV_X1 U9607 ( .A(n6990), .ZN(n6486) );
  NAND3_X1 U9608 ( .A1(n6486), .A2(n6485), .A3(n39052), .ZN(n6181) );
  NAND2_X1 U9609 ( .A1(n6181), .A2(n10589), .ZN(n6180) );
  INV_X1 U9610 ( .A(n6180), .ZN(n6167) );
  AOI22_X1 U9611 ( .A1(n37191), .A2(n6167), .B1(n6180), .B2(n39041), .ZN(n6278) );
  NAND2_X1 U9612 ( .A1(n37191), .A2(n6167), .ZN(n6168) );
  XOR2_X1 U9613 ( .A(n39040), .B(n6168), .Z(n6255) );
  AND2_X1 U9614 ( .A1(n6278), .A2(n6255), .ZN(n30287) );
  NOR2_X2 U9615 ( .A1(n6171), .A2(n6586), .ZN(n7215) );
  AOI21_X1 U9616 ( .B1(n7215), .B2(n6990), .A(n10589), .ZN(n7599) );
  NOR2_X1 U9617 ( .A1(n7599), .A2(n6169), .ZN(n6188) );
  INV_X1 U9618 ( .A(n6990), .ZN(n8418) );
  NAND2_X1 U9619 ( .A1(n39035), .A2(n3402), .ZN(n6170) );
  OAI21_X2 U9620 ( .B1(n7215), .B2(n8418), .A(n3944), .ZN(n6196) );
  INV_X1 U9621 ( .A(n6196), .ZN(n6190) );
  NAND2_X2 U9622 ( .A1(n3394), .A2(n6190), .ZN(n8010) );
  INV_X1 U9623 ( .A(n6183), .ZN(n6175) );
  NOR2_X1 U9624 ( .A1(n6172), .A2(n6171), .ZN(n6178) );
  NAND2_X2 U9625 ( .A1(n6175), .A2(n6177), .ZN(n11358) );
  NOR2_X2 U9626 ( .A1(n8010), .A2(n11358), .ZN(n11489) );
  AND2_X1 U9627 ( .A1(n6178), .A2(n3248), .ZN(n6174) );
  NAND2_X2 U9628 ( .A1(n6175), .A2(n6174), .ZN(n11359) );
  NOR2_X1 U9629 ( .A1(n11359), .A2(n8010), .ZN(n6999) );
  BUF_X2 U9630 ( .A(n6999), .Z(n10861) );
  BUF_X2 U9631 ( .A(n10861), .Z(n26616) );
  AOI22_X1 U9632 ( .A1(n29788), .A2(\xmem_data[96][5] ), .B1(n29672), .B2(
        \xmem_data[97][5] ), .ZN(n6187) );
  INV_X1 U9633 ( .A(n6178), .ZN(n11343) );
  NOR2_X2 U9634 ( .A1(n8010), .A2(n3377), .ZN(n11451) );
  BUF_X2 U9635 ( .A(n11451), .Z(n30279) );
  BUF_X1 U9636 ( .A(n14988), .Z(n30278) );
  AOI22_X1 U9637 ( .A1(n30279), .A2(\xmem_data[98][5] ), .B1(n30278), .B2(
        \xmem_data[99][5] ), .ZN(n6186) );
  NAND2_X1 U9638 ( .A1(n8020), .A2(n7421), .ZN(n6189) );
  NAND2_X2 U9639 ( .A1(n6183), .A2(n6177), .ZN(n11361) );
  NOR2_X2 U9640 ( .A1(n3447), .A2(n11361), .ZN(n11484) );
  NOR2_X2 U9641 ( .A1(n3447), .A2(n3246), .ZN(n11780) );
  AOI22_X1 U9642 ( .A1(n30280), .A2(\xmem_data[100][5] ), .B1(n29556), .B2(
        \xmem_data[101][5] ), .ZN(n6185) );
  NAND2_X1 U9643 ( .A1(n6180), .A2(n6179), .ZN(n8216) );
  INV_X1 U9644 ( .A(n8216), .ZN(n6201) );
  INV_X1 U9645 ( .A(n6201), .ZN(n8210) );
  OR2_X1 U9646 ( .A1(n6992), .A2(n39035), .ZN(n6182) );
  NAND2_X2 U9647 ( .A1(n6182), .A2(n6181), .ZN(n11357) );
  BUF_X1 U9648 ( .A(n6183), .Z(n11342) );
  NOR2_X1 U9649 ( .A1(n8211), .A2(n7645), .ZN(n6234) );
  BUF_X1 U9650 ( .A(n6234), .Z(n30282) );
  BUF_X1 U9651 ( .A(n14991), .Z(n30281) );
  AOI22_X1 U9652 ( .A1(n30282), .A2(\xmem_data[102][5] ), .B1(n3138), .B2(
        \xmem_data[103][5] ), .ZN(n6184) );
  NAND4_X1 U9653 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n6210)
         );
  NOR2_X2 U9654 ( .A1(n3446), .A2(n11358), .ZN(n11436) );
  BUF_X1 U9655 ( .A(n11436), .Z(n30248) );
  NOR2_X2 U9656 ( .A1(n3446), .A2(n11359), .ZN(n11437) );
  AOI22_X1 U9657 ( .A1(n30633), .A2(\xmem_data[104][5] ), .B1(n29589), .B2(
        \xmem_data[105][5] ), .ZN(n6195) );
  NAND2_X1 U9658 ( .A1(n11357), .A2(n8210), .ZN(n6191) );
  AOI22_X1 U9659 ( .A1(n30171), .A2(\xmem_data[106][5] ), .B1(n24157), .B2(
        \xmem_data[107][5] ), .ZN(n6194) );
  OR2_X2 U9660 ( .A1(n6188), .A2(n6196), .ZN(n8000) );
  NOR2_X2 U9661 ( .A1(n8000), .A2(n11361), .ZN(n11439) );
  BUF_X1 U9662 ( .A(n11439), .Z(n30250) );
  NAND2_X1 U9663 ( .A1(n3395), .A2(n3443), .ZN(n7408) );
  BUF_X1 U9664 ( .A(n8700), .Z(n30301) );
  AOI22_X1 U9665 ( .A1(n30745), .A2(\xmem_data[108][5] ), .B1(n29739), .B2(
        \xmem_data[109][5] ), .ZN(n6193) );
  NOR2_X1 U9666 ( .A1(n7206), .A2(n6191), .ZN(n6281) );
  AOI22_X1 U9667 ( .A1(n30251), .A2(\xmem_data[110][5] ), .B1(n25607), .B2(
        \xmem_data[111][5] ), .ZN(n6192) );
  NAND4_X1 U9668 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n6209)
         );
  AOI22_X1 U9669 ( .A1(n3167), .A2(\xmem_data[112][5] ), .B1(n3186), .B2(
        \xmem_data[113][5] ), .ZN(n6200) );
  NOR2_X2 U9670 ( .A1(n3378), .A2(n8000), .ZN(n15549) );
  BUF_X1 U9671 ( .A(n15549), .Z(n28689) );
  AOI22_X1 U9672 ( .A1(n28689), .A2(\xmem_data[114][5] ), .B1(n29012), .B2(
        \xmem_data[115][5] ), .ZN(n6199) );
  NAND3_X2 U9673 ( .A1(n8020), .A2(n7421), .A3(n6196), .ZN(n8005) );
  NOR2_X2 U9674 ( .A1(n8005), .A2(n11361), .ZN(n10802) );
  BUF_X1 U9675 ( .A(n10802), .Z(n30063) );
  NOR2_X2 U9676 ( .A1(n8005), .A2(n3457), .ZN(n18518) );
  BUF_X2 U9677 ( .A(n18518), .Z(n30170) );
  AOI22_X1 U9678 ( .A1(n29488), .A2(\xmem_data[116][5] ), .B1(n29487), .B2(
        \xmem_data[117][5] ), .ZN(n6198) );
  INV_X1 U9679 ( .A(n8216), .ZN(n8204) );
  NOR2_X1 U9680 ( .A1(n7010), .A2(n8199), .ZN(n6239) );
  BUF_X2 U9681 ( .A(n6239), .Z(n30270) );
  BUF_X1 U9682 ( .A(n14974), .Z(n30269) );
  AOI22_X1 U9683 ( .A1(n30270), .A2(\xmem_data[118][5] ), .B1(n30269), .B2(
        \xmem_data[119][5] ), .ZN(n6197) );
  NAND4_X1 U9684 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n6208)
         );
  NOR2_X1 U9685 ( .A1(n11358), .A2(n6202), .ZN(n6246) );
  AOI22_X1 U9686 ( .A1(n3211), .A2(\xmem_data[120][5] ), .B1(n30256), .B2(
        \xmem_data[121][5] ), .ZN(n6206) );
  NOR2_X1 U9687 ( .A1(n3377), .A2(n6202), .ZN(n6309) );
  BUF_X1 U9688 ( .A(n6309), .Z(n30048) );
  BUF_X1 U9689 ( .A(n13127), .Z(n30257) );
  AOI22_X1 U9690 ( .A1(n30048), .A2(\xmem_data[122][5] ), .B1(n30257), .B2(
        \xmem_data[123][5] ), .ZN(n6205) );
  NOR2_X1 U9691 ( .A1(n11361), .A2(n6202), .ZN(n6244) );
  BUF_X1 U9692 ( .A(n6244), .Z(n30260) );
  AOI22_X1 U9693 ( .A1(n30260), .A2(\xmem_data[124][5] ), .B1(n3420), .B2(
        \xmem_data[125][5] ), .ZN(n6204) );
  NOR2_X1 U9694 ( .A1(n11370), .A2(n6202), .ZN(n6245) );
  AOI22_X1 U9695 ( .A1(n30200), .A2(\xmem_data[126][5] ), .B1(n3434), .B2(
        \xmem_data[127][5] ), .ZN(n6203) );
  NAND4_X1 U9696 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n6207)
         );
  OR4_X1 U9697 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n6232) );
  INV_X1 U9698 ( .A(n6255), .ZN(n6279) );
  NOR2_X2 U9699 ( .A1(n6278), .A2(n6279), .ZN(n30188) );
  BUF_X1 U9700 ( .A(n11489), .Z(n30291) );
  BUF_X2 U9701 ( .A(n10861), .Z(n29697) );
  AOI22_X1 U9702 ( .A1(n28734), .A2(\xmem_data[64][5] ), .B1(n29697), .B2(
        \xmem_data[65][5] ), .ZN(n6214) );
  AOI22_X1 U9703 ( .A1(n28138), .A2(\xmem_data[66][5] ), .B1(n30278), .B2(
        \xmem_data[67][5] ), .ZN(n6213) );
  BUF_X1 U9704 ( .A(n11484), .Z(n30294) );
  AOI22_X1 U9705 ( .A1(n30294), .A2(\xmem_data[68][5] ), .B1(n29708), .B2(
        \xmem_data[69][5] ), .ZN(n6212) );
  AOI22_X1 U9706 ( .A1(n30219), .A2(\xmem_data[70][5] ), .B1(n30295), .B2(
        \xmem_data[71][5] ), .ZN(n6211) );
  NAND4_X1 U9707 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6230)
         );
  AOI22_X1 U9708 ( .A1(n29481), .A2(\xmem_data[72][5] ), .B1(n3369), .B2(
        \xmem_data[73][5] ), .ZN(n6218) );
  BUF_X1 U9709 ( .A(n14997), .Z(n30083) );
  AOI22_X1 U9710 ( .A1(n30192), .A2(\xmem_data[74][5] ), .B1(n30083), .B2(
        \xmem_data[75][5] ), .ZN(n6217) );
  BUF_X1 U9711 ( .A(n11439), .Z(n30302) );
  AOI22_X1 U9712 ( .A1(n27754), .A2(\xmem_data[76][5] ), .B1(n30090), .B2(
        \xmem_data[77][5] ), .ZN(n6216) );
  BUF_X1 U9713 ( .A(n29187), .Z(n30303) );
  AOI22_X1 U9714 ( .A1(n30304), .A2(\xmem_data[78][5] ), .B1(n30666), .B2(
        \xmem_data[79][5] ), .ZN(n6215) );
  NAND4_X1 U9715 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n6229)
         );
  AOI22_X1 U9716 ( .A1(n3164), .A2(\xmem_data[80][5] ), .B1(n3191), .B2(
        \xmem_data[81][5] ), .ZN(n6222) );
  BUF_X1 U9717 ( .A(n15549), .Z(n23901) );
  BUF_X1 U9718 ( .A(n14971), .Z(n30309) );
  AOI22_X1 U9719 ( .A1(n23901), .A2(\xmem_data[82][5] ), .B1(n30309), .B2(
        \xmem_data[83][5] ), .ZN(n6221) );
  BUF_X1 U9720 ( .A(n10802), .Z(n30717) );
  BUF_X4 U9721 ( .A(n18518), .Z(n29640) );
  AOI22_X1 U9722 ( .A1(n30717), .A2(\xmem_data[84][5] ), .B1(n30644), .B2(
        \xmem_data[85][5] ), .ZN(n6220) );
  BUF_X1 U9723 ( .A(n14974), .Z(n30311) );
  AOI22_X1 U9724 ( .A1(n30270), .A2(\xmem_data[86][5] ), .B1(n30311), .B2(
        \xmem_data[87][5] ), .ZN(n6219) );
  NAND4_X1 U9725 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(n6228)
         );
  AOI22_X1 U9726 ( .A1(n3210), .A2(\xmem_data[88][5] ), .B1(n3193), .B2(
        \xmem_data[89][5] ), .ZN(n6226) );
  AOI22_X1 U9727 ( .A1(n30258), .A2(\xmem_data[90][5] ), .B1(n20952), .B2(
        \xmem_data[91][5] ), .ZN(n6225) );
  BUF_X1 U9728 ( .A(n6244), .Z(n30318) );
  AOI22_X1 U9729 ( .A1(n30318), .A2(\xmem_data[92][5] ), .B1(n30317), .B2(
        \xmem_data[93][5] ), .ZN(n6224) );
  BUF_X1 U9730 ( .A(n6245), .Z(n30320) );
  BUF_X1 U9731 ( .A(n28973), .Z(n30319) );
  AOI22_X1 U9732 ( .A1(n30320), .A2(\xmem_data[94][5] ), .B1(n3153), .B2(
        \xmem_data[95][5] ), .ZN(n6223) );
  NAND4_X1 U9733 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6223), .ZN(n6227)
         );
  OR4_X1 U9734 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n6231) );
  AOI22_X1 U9735 ( .A1(n30287), .A2(n6232), .B1(n30188), .B2(n6231), .ZN(n6293) );
  BUF_X1 U9736 ( .A(n11780), .Z(n30217) );
  AOI22_X1 U9737 ( .A1(n30280), .A2(\xmem_data[4][5] ), .B1(n29556), .B2(
        \xmem_data[5][5] ), .ZN(n6233) );
  INV_X1 U9738 ( .A(n6233), .ZN(n6238) );
  BUF_X1 U9739 ( .A(n11451), .Z(n30215) );
  AOI22_X1 U9740 ( .A1(n28138), .A2(\xmem_data[2][5] ), .B1(n29565), .B2(
        \xmem_data[3][5] ), .ZN(n6236) );
  BUF_X1 U9741 ( .A(n14991), .Z(n30218) );
  AOI22_X1 U9742 ( .A1(n30219), .A2(\xmem_data[6][5] ), .B1(n3131), .B2(
        \xmem_data[7][5] ), .ZN(n6235) );
  NAND2_X1 U9743 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  NOR2_X1 U9744 ( .A1(n6238), .A2(n6237), .ZN(n6257) );
  AOI22_X1 U9745 ( .A1(n3162), .A2(\xmem_data[16][5] ), .B1(n11426), .B2(
        \xmem_data[17][5] ), .ZN(n6243) );
  BUF_X1 U9746 ( .A(n15549), .Z(n26812) );
  AOI22_X1 U9747 ( .A1(n26812), .A2(\xmem_data[18][5] ), .B1(n30309), .B2(
        \xmem_data[19][5] ), .ZN(n6242) );
  BUF_X2 U9748 ( .A(n18518), .Z(n30644) );
  AOI22_X1 U9749 ( .A1(n30076), .A2(\xmem_data[20][5] ), .B1(n29487), .B2(
        \xmem_data[21][5] ), .ZN(n6241) );
  BUF_X1 U9750 ( .A(n6239), .Z(n30205) );
  AOI22_X1 U9751 ( .A1(n30205), .A2(\xmem_data[22][5] ), .B1(n3308), .B2(
        \xmem_data[23][5] ), .ZN(n6240) );
  NAND4_X1 U9752 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n6254)
         );
  BUF_X1 U9753 ( .A(n6244), .Z(n30199) );
  AOI22_X1 U9754 ( .A1(n30199), .A2(\xmem_data[28][5] ), .B1(n30317), .B2(
        \xmem_data[29][5] ), .ZN(n6252) );
  AOI22_X1 U9755 ( .A1(n30320), .A2(\xmem_data[30][5] ), .B1(n3149), .B2(
        \xmem_data[31][5] ), .ZN(n6251) );
  AOI22_X1 U9756 ( .A1(n3211), .A2(\xmem_data[24][5] ), .B1(n3193), .B2(
        \xmem_data[25][5] ), .ZN(n6249) );
  AOI22_X1 U9757 ( .A1(n30048), .A2(\xmem_data[26][5] ), .B1(n29657), .B2(
        \xmem_data[27][5] ), .ZN(n6248) );
  AND2_X1 U9758 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND3_X1 U9759 ( .A1(n6252), .A2(n6251), .A3(n6250), .ZN(n6253) );
  NOR2_X1 U9760 ( .A1(n6254), .A2(n6253), .ZN(n6256) );
  NOR2_X2 U9761 ( .A1(n6278), .A2(n6255), .ZN(n30228) );
  AOI21_X1 U9762 ( .B1(n6257), .B2(n6256), .A(n30229), .ZN(n6291) );
  BUF_X1 U9763 ( .A(n10861), .Z(n30695) );
  AOI22_X1 U9764 ( .A1(n27710), .A2(\xmem_data[32][5] ), .B1(n30290), .B2(
        \xmem_data[33][5] ), .ZN(n6261) );
  AOI22_X1 U9765 ( .A1(n3392), .A2(\xmem_data[34][5] ), .B1(n30292), .B2(
        \xmem_data[35][5] ), .ZN(n6260) );
  AOI22_X1 U9766 ( .A1(n30294), .A2(\xmem_data[36][5] ), .B1(n29798), .B2(
        \xmem_data[37][5] ), .ZN(n6259) );
  AOI22_X1 U9767 ( .A1(n30219), .A2(\xmem_data[38][5] ), .B1(n30295), .B2(
        \xmem_data[39][5] ), .ZN(n6258) );
  AND4_X1 U9768 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n6277)
         );
  AOI22_X1 U9769 ( .A1(n29647), .A2(\xmem_data[40][5] ), .B1(n29482), .B2(
        \xmem_data[41][5] ), .ZN(n6265) );
  AOI22_X1 U9770 ( .A1(n30171), .A2(\xmem_data[42][5] ), .B1(n30083), .B2(
        \xmem_data[43][5] ), .ZN(n6264) );
  BUF_X1 U9771 ( .A(n8700), .Z(n27728) );
  AOI22_X1 U9772 ( .A1(n29395), .A2(\xmem_data[44][5] ), .B1(n29592), .B2(
        \xmem_data[45][5] ), .ZN(n6263) );
  AOI22_X1 U9773 ( .A1(n30304), .A2(\xmem_data[46][5] ), .B1(n29315), .B2(
        \xmem_data[47][5] ), .ZN(n6262) );
  AND4_X1 U9774 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n6276)
         );
  AOI22_X1 U9775 ( .A1(n3165), .A2(\xmem_data[48][5] ), .B1(n3184), .B2(
        \xmem_data[49][5] ), .ZN(n6269) );
  AOI22_X1 U9776 ( .A1(n30075), .A2(\xmem_data[50][5] ), .B1(n30309), .B2(
        \xmem_data[51][5] ), .ZN(n6268) );
  AOI22_X1 U9777 ( .A1(n27713), .A2(\xmem_data[52][5] ), .B1(n29721), .B2(
        \xmem_data[53][5] ), .ZN(n6267) );
  AOI22_X1 U9778 ( .A1(n30205), .A2(\xmem_data[54][5] ), .B1(n30311), .B2(
        \xmem_data[55][5] ), .ZN(n6266) );
  AND4_X1 U9779 ( .A1(n6269), .A2(n6268), .A3(n6267), .A4(n6266), .ZN(n6275)
         );
  AOI22_X1 U9780 ( .A1(n3211), .A2(\xmem_data[56][5] ), .B1(n3193), .B2(
        \xmem_data[57][5] ), .ZN(n6273) );
  AOI22_X1 U9781 ( .A1(n30258), .A2(\xmem_data[58][5] ), .B1(n17051), .B2(
        \xmem_data[59][5] ), .ZN(n6272) );
  AOI22_X1 U9782 ( .A1(n30318), .A2(\xmem_data[60][5] ), .B1(n30317), .B2(
        \xmem_data[61][5] ), .ZN(n6271) );
  AOI22_X1 U9783 ( .A1(n30320), .A2(\xmem_data[62][5] ), .B1(n3153), .B2(
        \xmem_data[63][5] ), .ZN(n6270) );
  AND4_X1 U9784 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n6274)
         );
  NAND4_X1 U9785 ( .A1(n6277), .A2(n6276), .A3(n6275), .A4(n6274), .ZN(n6280)
         );
  AND2_X1 U9786 ( .A1(n6279), .A2(n6278), .ZN(n30329) );
  BUF_X1 U9787 ( .A(n11436), .Z(n30191) );
  BUF_X1 U9788 ( .A(n11437), .Z(n30190) );
  AOI22_X1 U9789 ( .A1(n29647), .A2(\xmem_data[8][5] ), .B1(n29589), .B2(
        \xmem_data[9][5] ), .ZN(n6285) );
  AOI22_X1 U9790 ( .A1(n30171), .A2(\xmem_data[10][5] ), .B1(n30083), .B2(
        \xmem_data[11][5] ), .ZN(n6284) );
  BUF_X1 U9791 ( .A(n8700), .Z(n28778) );
  AOI22_X1 U9792 ( .A1(n29604), .A2(\xmem_data[12][5] ), .B1(n29739), .B2(
        \xmem_data[13][5] ), .ZN(n6283) );
  AOI22_X1 U9793 ( .A1(n30304), .A2(\xmem_data[14][5] ), .B1(n27517), .B2(
        \xmem_data[15][5] ), .ZN(n6282) );
  AND4_X1 U9794 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n6289)
         );
  BUF_X1 U9795 ( .A(n11489), .Z(n30223) );
  AOI22_X1 U9796 ( .A1(n30223), .A2(\xmem_data[0][5] ), .B1(n29697), .B2(
        \xmem_data[1][5] ), .ZN(n6286) );
  INV_X1 U9797 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U9798 ( .A1(n6287), .A2(n30228), .ZN(n6288) );
  OAI21_X1 U9799 ( .B1(n30229), .B2(n6289), .A(n6288), .ZN(n6290) );
  NOR3_X1 U9800 ( .A1(n6291), .A2(n3834), .A3(n6290), .ZN(n6292) );
  NAND2_X1 U9801 ( .A1(n6293), .A2(n6292), .ZN(n32211) );
  BUF_X2 U9802 ( .A(n15549), .Z(n30715) );
  AND2_X1 U9803 ( .A1(n29639), .A2(\xmem_data[115][4] ), .ZN(n6294) );
  AOI21_X1 U9804 ( .B1(n30715), .B2(\xmem_data[114][4] ), .A(n6294), .ZN(n6298) );
  AOI22_X1 U9805 ( .A1(n3166), .A2(\xmem_data[112][4] ), .B1(n3182), .B2(
        \xmem_data[113][4] ), .ZN(n6297) );
  AOI22_X1 U9806 ( .A1(n30063), .A2(\xmem_data[116][4] ), .B1(n30765), .B2(
        \xmem_data[117][4] ), .ZN(n6296) );
  AOI22_X1 U9807 ( .A1(n30270), .A2(\xmem_data[118][4] ), .B1(n30269), .B2(
        \xmem_data[119][4] ), .ZN(n6295) );
  NAND4_X1 U9808 ( .A1(n6298), .A2(n6297), .A3(n6296), .A4(n6295), .ZN(n6304)
         );
  BUF_X1 U9809 ( .A(n15549), .Z(n27031) );
  AOI22_X1 U9810 ( .A1(n27031), .A2(\xmem_data[50][4] ), .B1(n30309), .B2(
        \xmem_data[51][4] ), .ZN(n6302) );
  BUF_X1 U9811 ( .A(n10802), .Z(n29722) );
  BUF_X2 U9812 ( .A(n18518), .Z(n30716) );
  AOI22_X1 U9813 ( .A1(n30198), .A2(\xmem_data[52][4] ), .B1(n30644), .B2(
        \xmem_data[53][4] ), .ZN(n6301) );
  AOI22_X1 U9814 ( .A1(n3167), .A2(\xmem_data[48][4] ), .B1(n3190), .B2(
        \xmem_data[49][4] ), .ZN(n6300) );
  AOI22_X1 U9815 ( .A1(n30270), .A2(\xmem_data[54][4] ), .B1(n30311), .B2(
        \xmem_data[55][4] ), .ZN(n6299) );
  NAND4_X1 U9816 ( .A1(n6302), .A2(n6301), .A3(n6300), .A4(n6299), .ZN(n6303)
         );
  AOI22_X1 U9817 ( .A1(n30287), .A2(n6304), .B1(n6303), .B2(n30329), .ZN(n6337) );
  AOI22_X1 U9818 ( .A1(n30633), .A2(\xmem_data[8][4] ), .B1(n30662), .B2(
        \xmem_data[9][4] ), .ZN(n6308) );
  AOI22_X1 U9819 ( .A1(n30192), .A2(\xmem_data[10][4] ), .B1(n29308), .B2(
        \xmem_data[11][4] ), .ZN(n6307) );
  BUF_X1 U9820 ( .A(n8700), .Z(n30193) );
  AOI22_X1 U9821 ( .A1(n29436), .A2(\xmem_data[12][4] ), .B1(n30301), .B2(
        \xmem_data[13][4] ), .ZN(n6306) );
  AOI22_X1 U9822 ( .A1(n30304), .A2(\xmem_data[14][4] ), .B1(n28231), .B2(
        \xmem_data[15][4] ), .ZN(n6305) );
  NAND4_X1 U9823 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6323)
         );
  AOI22_X1 U9824 ( .A1(n3211), .A2(\xmem_data[24][4] ), .B1(n3192), .B2(
        \xmem_data[25][4] ), .ZN(n6313) );
  AOI22_X1 U9825 ( .A1(n30258), .A2(\xmem_data[26][4] ), .B1(n23753), .B2(
        \xmem_data[27][4] ), .ZN(n6312) );
  AOI22_X1 U9826 ( .A1(n30199), .A2(\xmem_data[28][4] ), .B1(n3420), .B2(
        \xmem_data[29][4] ), .ZN(n6311) );
  AOI22_X1 U9827 ( .A1(n30320), .A2(\xmem_data[30][4] ), .B1(n28164), .B2(
        \xmem_data[31][4] ), .ZN(n6310) );
  NAND4_X1 U9828 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n6310), .ZN(n6314)
         );
  NAND2_X1 U9829 ( .A1(n6314), .A2(n30228), .ZN(n6321) );
  AOI22_X1 U9830 ( .A1(n3210), .A2(\xmem_data[120][4] ), .B1(n30256), .B2(
        \xmem_data[121][4] ), .ZN(n6318) );
  AOI22_X1 U9831 ( .A1(n30258), .A2(\xmem_data[122][4] ), .B1(n30257), .B2(
        \xmem_data[123][4] ), .ZN(n6317) );
  AOI22_X1 U9832 ( .A1(n30260), .A2(\xmem_data[124][4] ), .B1(n3420), .B2(
        \xmem_data[125][4] ), .ZN(n6316) );
  AOI22_X1 U9833 ( .A1(n30200), .A2(\xmem_data[126][4] ), .B1(n3412), .B2(
        \xmem_data[127][4] ), .ZN(n6315) );
  NAND4_X1 U9834 ( .A1(n6318), .A2(n6317), .A3(n6316), .A4(n6315), .ZN(n6319)
         );
  NAND2_X1 U9835 ( .A1(n6319), .A2(n30287), .ZN(n6320) );
  NAND2_X1 U9836 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  AOI21_X1 U9837 ( .B1(n6323), .B2(n30228), .A(n6322), .ZN(n6336) );
  AOI22_X1 U9838 ( .A1(n29390), .A2(\xmem_data[40][4] ), .B1(n29646), .B2(
        \xmem_data[41][4] ), .ZN(n6327) );
  AOI22_X1 U9839 ( .A1(n30171), .A2(\xmem_data[42][4] ), .B1(n30083), .B2(
        \xmem_data[43][4] ), .ZN(n6326) );
  AOI22_X1 U9840 ( .A1(n30635), .A2(\xmem_data[44][4] ), .B1(n27728), .B2(
        \xmem_data[45][4] ), .ZN(n6325) );
  AOI22_X1 U9841 ( .A1(n30304), .A2(\xmem_data[46][4] ), .B1(n28091), .B2(
        \xmem_data[47][4] ), .ZN(n6324) );
  NAND4_X1 U9842 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n6328)
         );
  NAND2_X1 U9843 ( .A1(n6328), .A2(n30329), .ZN(n6335) );
  AOI22_X1 U9844 ( .A1(n29590), .A2(\xmem_data[72][4] ), .B1(n30662), .B2(
        \xmem_data[73][4] ), .ZN(n6332) );
  AOI22_X1 U9845 ( .A1(n30171), .A2(\xmem_data[74][4] ), .B1(n30083), .B2(
        \xmem_data[75][4] ), .ZN(n6331) );
  BUF_X1 U9846 ( .A(n8700), .Z(n30237) );
  AOI22_X1 U9847 ( .A1(n29604), .A2(\xmem_data[76][4] ), .B1(n30090), .B2(
        \xmem_data[77][4] ), .ZN(n6330) );
  AOI22_X1 U9848 ( .A1(n30304), .A2(\xmem_data[78][4] ), .B1(n29605), .B2(
        \xmem_data[79][4] ), .ZN(n6329) );
  NAND4_X1 U9849 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n6333)
         );
  NAND2_X1 U9850 ( .A1(n6333), .A2(n30188), .ZN(n6334) );
  NAND4_X1 U9851 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n6392)
         );
  AOI22_X1 U9852 ( .A1(n3211), .A2(\xmem_data[56][4] ), .B1(n3193), .B2(
        \xmem_data[57][4] ), .ZN(n6342) );
  AOI22_X1 U9853 ( .A1(n30258), .A2(\xmem_data[58][4] ), .B1(n20826), .B2(
        \xmem_data[59][4] ), .ZN(n6341) );
  AOI22_X1 U9854 ( .A1(n30200), .A2(\xmem_data[62][4] ), .B1(n3153), .B2(
        \xmem_data[63][4] ), .ZN(n6339) );
  NAND4_X1 U9855 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n6348)
         );
  BUF_X2 U9856 ( .A(n10861), .Z(n29672) );
  AOI22_X1 U9857 ( .A1(n30291), .A2(\xmem_data[96][4] ), .B1(n30106), .B2(
        \xmem_data[97][4] ), .ZN(n6346) );
  BUF_X1 U9858 ( .A(n14988), .Z(n30292) );
  AOI22_X1 U9859 ( .A1(n28700), .A2(\xmem_data[98][4] ), .B1(n30292), .B2(
        \xmem_data[99][4] ), .ZN(n6345) );
  AOI22_X1 U9860 ( .A1(n30280), .A2(\xmem_data[100][4] ), .B1(n30293), .B2(
        \xmem_data[101][4] ), .ZN(n6344) );
  AOI22_X1 U9861 ( .A1(n30282), .A2(\xmem_data[102][4] ), .B1(n3137), .B2(
        \xmem_data[103][4] ), .ZN(n6343) );
  NAND4_X1 U9862 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n6347)
         );
  AOI22_X1 U9863 ( .A1(n30329), .A2(n6348), .B1(n6347), .B2(n30287), .ZN(n6372) );
  AOI22_X1 U9864 ( .A1(n3392), .A2(\xmem_data[34][4] ), .B1(n29832), .B2(
        \xmem_data[35][4] ), .ZN(n6352) );
  AOI22_X1 U9865 ( .A1(n27710), .A2(\xmem_data[32][4] ), .B1(n30707), .B2(
        \xmem_data[33][4] ), .ZN(n6351) );
  AOI22_X1 U9866 ( .A1(n30294), .A2(\xmem_data[36][4] ), .B1(n28786), .B2(
        \xmem_data[37][4] ), .ZN(n6350) );
  AOI22_X1 U9867 ( .A1(n30219), .A2(\xmem_data[38][4] ), .B1(n30295), .B2(
        \xmem_data[39][4] ), .ZN(n6349) );
  NAND4_X1 U9868 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n6353)
         );
  NAND2_X1 U9869 ( .A1(n6353), .A2(n30329), .ZN(n6371) );
  AOI22_X1 U9870 ( .A1(n3167), .A2(\xmem_data[80][4] ), .B1(n3186), .B2(
        \xmem_data[81][4] ), .ZN(n6357) );
  AOI22_X1 U9871 ( .A1(n30075), .A2(\xmem_data[82][4] ), .B1(n30309), .B2(
        \xmem_data[83][4] ), .ZN(n6356) );
  BUF_X1 U9872 ( .A(n10802), .Z(n29547) );
  AOI22_X1 U9873 ( .A1(n29547), .A2(\xmem_data[84][4] ), .B1(n29640), .B2(
        \xmem_data[85][4] ), .ZN(n6355) );
  AOI22_X1 U9874 ( .A1(n30205), .A2(\xmem_data[86][4] ), .B1(n30311), .B2(
        \xmem_data[87][4] ), .ZN(n6354) );
  NAND4_X1 U9875 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n6363)
         );
  AOI22_X1 U9876 ( .A1(n29716), .A2(\xmem_data[18][4] ), .B1(n29639), .B2(
        \xmem_data[19][4] ), .ZN(n6361) );
  AOI22_X1 U9877 ( .A1(n3168), .A2(\xmem_data[16][4] ), .B1(n3188), .B2(
        \xmem_data[17][4] ), .ZN(n6360) );
  BUF_X4 U9878 ( .A(n18518), .Z(n30266) );
  AOI22_X1 U9879 ( .A1(n27713), .A2(\xmem_data[20][4] ), .B1(n29640), .B2(
        \xmem_data[21][4] ), .ZN(n6359) );
  AOI22_X1 U9880 ( .A1(n30205), .A2(\xmem_data[22][4] ), .B1(n28955), .B2(
        \xmem_data[23][4] ), .ZN(n6358) );
  NAND4_X1 U9881 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n6362)
         );
  AOI22_X1 U9882 ( .A1(n6363), .A2(n30188), .B1(n6362), .B2(n30228), .ZN(n6370) );
  AOI22_X1 U9883 ( .A1(n29590), .A2(\xmem_data[104][4] ), .B1(n30190), .B2(
        \xmem_data[105][4] ), .ZN(n6367) );
  AOI22_X1 U9884 ( .A1(n3214), .A2(\xmem_data[106][4] ), .B1(n29403), .B2(
        \xmem_data[107][4] ), .ZN(n6366) );
  AOI22_X1 U9885 ( .A1(n30665), .A2(\xmem_data[108][4] ), .B1(n28684), .B2(
        \xmem_data[109][4] ), .ZN(n6365) );
  AOI22_X1 U9886 ( .A1(n30251), .A2(\xmem_data[110][4] ), .B1(n30666), .B2(
        \xmem_data[111][4] ), .ZN(n6364) );
  NAND4_X1 U9887 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .ZN(n6368)
         );
  NAND2_X1 U9888 ( .A1(n6368), .A2(n30287), .ZN(n6369) );
  NAND4_X1 U9889 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n6391)
         );
  AOI22_X1 U9890 ( .A1(n28207), .A2(\xmem_data[66][4] ), .B1(n29627), .B2(
        \xmem_data[67][4] ), .ZN(n6376) );
  BUF_X2 U9891 ( .A(n10861), .Z(n27013) );
  AOI22_X1 U9892 ( .A1(n27710), .A2(\xmem_data[64][4] ), .B1(n26616), .B2(
        \xmem_data[65][4] ), .ZN(n6375) );
  AOI22_X1 U9893 ( .A1(n30294), .A2(\xmem_data[68][4] ), .B1(n29708), .B2(
        \xmem_data[69][4] ), .ZN(n6374) );
  AOI22_X1 U9894 ( .A1(n30219), .A2(\xmem_data[70][4] ), .B1(n30295), .B2(
        \xmem_data[71][4] ), .ZN(n6373) );
  NAND4_X1 U9895 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n6382)
         );
  AOI22_X1 U9896 ( .A1(n3210), .A2(\xmem_data[88][4] ), .B1(n3193), .B2(
        \xmem_data[89][4] ), .ZN(n6380) );
  AOI22_X1 U9897 ( .A1(n6309), .A2(\xmem_data[90][4] ), .B1(n29383), .B2(
        \xmem_data[91][4] ), .ZN(n6379) );
  AOI22_X1 U9898 ( .A1(n30318), .A2(\xmem_data[92][4] ), .B1(n30317), .B2(
        \xmem_data[93][4] ), .ZN(n6378) );
  AOI22_X1 U9899 ( .A1(n30200), .A2(\xmem_data[94][4] ), .B1(n3153), .B2(
        \xmem_data[95][4] ), .ZN(n6377) );
  NAND4_X1 U9900 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n6381)
         );
  OAI21_X1 U9901 ( .B1(n6382), .B2(n6381), .A(n30188), .ZN(n6389) );
  BUF_X1 U9902 ( .A(n10861), .Z(n30106) );
  AOI22_X1 U9903 ( .A1(n28136), .A2(\xmem_data[0][4] ), .B1(n29753), .B2(
        \xmem_data[1][4] ), .ZN(n6386) );
  AOI22_X1 U9904 ( .A1(n29628), .A2(\xmem_data[2][4] ), .B1(n30292), .B2(
        \xmem_data[3][4] ), .ZN(n6385) );
  AOI22_X1 U9905 ( .A1(n28740), .A2(\xmem_data[4][4] ), .B1(n28786), .B2(
        \xmem_data[5][4] ), .ZN(n6384) );
  AOI22_X1 U9906 ( .A1(n30219), .A2(\xmem_data[6][4] ), .B1(n3132), .B2(
        \xmem_data[7][4] ), .ZN(n6383) );
  NAND4_X1 U9907 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n6387)
         );
  NAND2_X1 U9908 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  XOR2_X1 U9909 ( .A(\fmem_data[15][6] ), .B(\fmem_data[15][7] ), .Z(n6393) );
  OAI22_X1 U9910 ( .A1(n35031), .A2(n35697), .B1(n33235), .B2(n35696), .ZN(
        n35094) );
  XNOR2_X1 U9911 ( .A(n35096), .B(n35094), .ZN(n6989) );
  AOI22_X1 U9912 ( .A1(n31345), .A2(\xmem_data[120][7] ), .B1(n31344), .B2(
        \xmem_data[121][7] ), .ZN(n6397) );
  AOI22_X1 U9913 ( .A1(n27925), .A2(\xmem_data[122][7] ), .B1(n31346), .B2(
        \xmem_data[123][7] ), .ZN(n6396) );
  AOI22_X1 U9914 ( .A1(n3434), .A2(\xmem_data[124][7] ), .B1(n31347), .B2(
        \xmem_data[125][7] ), .ZN(n6395) );
  AOI22_X1 U9915 ( .A1(n31348), .A2(\xmem_data[126][7] ), .B1(n3217), .B2(
        \xmem_data[127][7] ), .ZN(n6394) );
  NAND4_X1 U9916 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n6414)
         );
  AOI22_X1 U9917 ( .A1(n31353), .A2(\xmem_data[104][7] ), .B1(n22702), .B2(
        \xmem_data[105][7] ), .ZN(n6401) );
  AOI22_X1 U9918 ( .A1(n25710), .A2(\xmem_data[106][7] ), .B1(n30513), .B2(
        \xmem_data[107][7] ), .ZN(n6400) );
  AOI22_X1 U9919 ( .A1(n17018), .A2(\xmem_data[108][7] ), .B1(n29188), .B2(
        \xmem_data[109][7] ), .ZN(n6399) );
  AOI22_X1 U9920 ( .A1(n24133), .A2(\xmem_data[110][7] ), .B1(n31355), .B2(
        \xmem_data[111][7] ), .ZN(n6398) );
  NAND4_X1 U9921 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n6412)
         );
  AOI22_X1 U9922 ( .A1(n28687), .A2(\xmem_data[112][7] ), .B1(n31360), .B2(
        \xmem_data[113][7] ), .ZN(n6405) );
  AOI22_X1 U9923 ( .A1(n27952), .A2(\xmem_data[114][7] ), .B1(n31361), .B2(
        \xmem_data[115][7] ), .ZN(n6404) );
  AOI22_X1 U9924 ( .A1(n28202), .A2(\xmem_data[116][7] ), .B1(n31362), .B2(
        \xmem_data[117][7] ), .ZN(n6403) );
  AOI22_X1 U9925 ( .A1(n31316), .A2(\xmem_data[118][7] ), .B1(n27526), .B2(
        \xmem_data[119][7] ), .ZN(n6402) );
  NAND4_X1 U9926 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n6411)
         );
  AOI22_X1 U9927 ( .A1(n31368), .A2(\xmem_data[96][7] ), .B1(n31367), .B2(
        \xmem_data[97][7] ), .ZN(n6409) );
  AOI22_X1 U9928 ( .A1(n20725), .A2(\xmem_data[98][7] ), .B1(n25415), .B2(
        \xmem_data[99][7] ), .ZN(n6408) );
  AOI22_X1 U9929 ( .A1(n20808), .A2(\xmem_data[100][7] ), .B1(n15011), .B2(
        \xmem_data[101][7] ), .ZN(n6407) );
  AOI22_X1 U9930 ( .A1(n25422), .A2(\xmem_data[102][7] ), .B1(n3358), .B2(
        \xmem_data[103][7] ), .ZN(n6406) );
  NAND4_X1 U9931 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n6410)
         );
  OR3_X1 U9932 ( .A1(n6412), .A2(n6411), .A3(n6410), .ZN(n6413) );
  OAI21_X1 U9933 ( .B1(n6414), .B2(n6413), .A(n31376), .ZN(n6437) );
  AOI22_X1 U9934 ( .A1(n31308), .A2(\xmem_data[88][7] ), .B1(n30524), .B2(
        \xmem_data[89][7] ), .ZN(n6418) );
  AOI22_X1 U9935 ( .A1(n17056), .A2(\xmem_data[90][7] ), .B1(n31309), .B2(
        \xmem_data[91][7] ), .ZN(n6417) );
  AOI22_X1 U9936 ( .A1(n3348), .A2(\xmem_data[92][7] ), .B1(n24172), .B2(
        \xmem_data[93][7] ), .ZN(n6416) );
  AOI22_X1 U9937 ( .A1(n20991), .A2(\xmem_data[94][7] ), .B1(n3220), .B2(
        \xmem_data[95][7] ), .ZN(n6415) );
  NAND4_X1 U9938 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n6435)
         );
  AOI22_X1 U9939 ( .A1(n31327), .A2(\xmem_data[72][7] ), .B1(n31326), .B2(
        \xmem_data[73][7] ), .ZN(n6422) );
  AOI22_X1 U9940 ( .A1(n30891), .A2(\xmem_data[74][7] ), .B1(n28517), .B2(
        \xmem_data[75][7] ), .ZN(n6421) );
  AOI22_X1 U9941 ( .A1(n31328), .A2(\xmem_data[76][7] ), .B1(n30615), .B2(
        \xmem_data[77][7] ), .ZN(n6420) );
  AOI22_X1 U9942 ( .A1(n31330), .A2(\xmem_data[78][7] ), .B1(n31329), .B2(
        \xmem_data[79][7] ), .ZN(n6419) );
  NAND4_X1 U9943 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6419), .ZN(n6433)
         );
  AOI22_X1 U9944 ( .A1(n16990), .A2(\xmem_data[80][7] ), .B1(n27523), .B2(
        \xmem_data[81][7] ), .ZN(n6426) );
  AOI22_X1 U9945 ( .A1(n21010), .A2(\xmem_data[82][7] ), .B1(n25581), .B2(
        \xmem_data[83][7] ), .ZN(n6425) );
  AOI22_X1 U9946 ( .A1(n31315), .A2(\xmem_data[84][7] ), .B1(n31314), .B2(
        \xmem_data[85][7] ), .ZN(n6424) );
  AOI22_X1 U9947 ( .A1(n31316), .A2(\xmem_data[86][7] ), .B1(n28500), .B2(
        \xmem_data[87][7] ), .ZN(n6423) );
  NAND4_X1 U9948 ( .A1(n6426), .A2(n6425), .A3(n6424), .A4(n6423), .ZN(n6432)
         );
  AOI22_X1 U9949 ( .A1(n23770), .A2(\xmem_data[64][7] ), .B1(n29255), .B2(
        \xmem_data[65][7] ), .ZN(n6430) );
  AOI22_X1 U9950 ( .A1(n28475), .A2(\xmem_data[66][7] ), .B1(n13444), .B2(
        \xmem_data[67][7] ), .ZN(n6429) );
  AOI22_X1 U9951 ( .A1(n29157), .A2(\xmem_data[68][7] ), .B1(n24553), .B2(
        \xmem_data[69][7] ), .ZN(n6428) );
  AOI22_X1 U9952 ( .A1(n31321), .A2(\xmem_data[70][7] ), .B1(n13475), .B2(
        \xmem_data[71][7] ), .ZN(n6427) );
  NAND4_X1 U9953 ( .A1(n6430), .A2(n6429), .A3(n6428), .A4(n6427), .ZN(n6431)
         );
  OR3_X1 U9954 ( .A1(n6433), .A2(n6432), .A3(n6431), .ZN(n6434) );
  OAI21_X1 U9955 ( .B1(n6435), .B2(n6434), .A(n31342), .ZN(n6436) );
  NAND2_X1 U9956 ( .A1(n6437), .A2(n6436), .ZN(n6481) );
  AOI22_X1 U9957 ( .A1(n20808), .A2(\xmem_data[4][7] ), .B1(n23771), .B2(
        \xmem_data[5][7] ), .ZN(n6438) );
  AOI22_X1 U9958 ( .A1(n27911), .A2(\xmem_data[8][7] ), .B1(n20775), .B2(
        \xmem_data[9][7] ), .ZN(n6441) );
  AOI22_X1 U9959 ( .A1(n24214), .A2(\xmem_data[14][7] ), .B1(n31270), .B2(
        \xmem_data[15][7] ), .ZN(n6440) );
  AOI22_X1 U9960 ( .A1(n31269), .A2(\xmem_data[13][7] ), .B1(
        \xmem_data[12][7] ), .B2(n24545), .ZN(n6439) );
  AOI22_X1 U9961 ( .A1(n31255), .A2(\xmem_data[16][7] ), .B1(n31254), .B2(
        \xmem_data[17][7] ), .ZN(n6445) );
  AOI22_X1 U9962 ( .A1(n20593), .A2(\xmem_data[18][7] ), .B1(n20506), .B2(
        \xmem_data[19][7] ), .ZN(n6444) );
  AOI22_X1 U9963 ( .A1(n3330), .A2(\xmem_data[20][7] ), .B1(n29245), .B2(
        \xmem_data[21][7] ), .ZN(n6443) );
  AOI22_X1 U9964 ( .A1(n22719), .A2(\xmem_data[22][7] ), .B1(n31256), .B2(
        \xmem_data[23][7] ), .ZN(n6442) );
  AOI22_X1 U9965 ( .A1(n3341), .A2(\xmem_data[2][7] ), .B1(n31275), .B2(
        \xmem_data[3][7] ), .ZN(n6448) );
  AOI22_X1 U9966 ( .A1(n31276), .A2(\xmem_data[6][7] ), .B1(n3358), .B2(
        \xmem_data[7][7] ), .ZN(n6447) );
  AOI22_X1 U9967 ( .A1(n30964), .A2(\xmem_data[0][7] ), .B1(n20500), .B2(
        \xmem_data[1][7] ), .ZN(n6446) );
  AOI22_X1 U9968 ( .A1(n31268), .A2(\xmem_data[10][7] ), .B1(n25382), .B2(
        \xmem_data[11][7] ), .ZN(n6449) );
  NAND4_X1 U9969 ( .A1(n6450), .A2(n3480), .A3(n3949), .A4(n6449), .ZN(n6456)
         );
  AOI22_X1 U9970 ( .A1(n27498), .A2(\xmem_data[24][7] ), .B1(n31261), .B2(
        \xmem_data[25][7] ), .ZN(n6454) );
  AOI22_X1 U9971 ( .A1(n3380), .A2(\xmem_data[26][7] ), .B1(n31262), .B2(
        \xmem_data[27][7] ), .ZN(n6453) );
  AOI22_X1 U9972 ( .A1(n3144), .A2(\xmem_data[28][7] ), .B1(n30589), .B2(
        \xmem_data[29][7] ), .ZN(n6452) );
  AOI22_X1 U9973 ( .A1(n24443), .A2(\xmem_data[30][7] ), .B1(n3220), .B2(
        \xmem_data[31][7] ), .ZN(n6451) );
  NAND4_X1 U9974 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n6451), .ZN(n6455)
         );
  OAI21_X1 U9975 ( .B1(n6456), .B2(n6455), .A(n31284), .ZN(n6457) );
  AOI22_X1 U9976 ( .A1(n24563), .A2(\xmem_data[32][7] ), .B1(n25562), .B2(
        \xmem_data[33][7] ), .ZN(n6461) );
  AOI22_X1 U9977 ( .A1(n28475), .A2(\xmem_data[34][7] ), .B1(n28342), .B2(
        \xmem_data[35][7] ), .ZN(n6460) );
  AOI22_X1 U9978 ( .A1(n16973), .A2(\xmem_data[36][7] ), .B1(n29103), .B2(
        \xmem_data[37][7] ), .ZN(n6459) );
  AOI22_X1 U9979 ( .A1(n31321), .A2(\xmem_data[38][7] ), .B1(n13475), .B2(
        \xmem_data[39][7] ), .ZN(n6458) );
  NAND4_X1 U9980 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6477)
         );
  AOI22_X1 U9981 ( .A1(n31327), .A2(\xmem_data[40][7] ), .B1(n31326), .B2(
        \xmem_data[41][7] ), .ZN(n6465) );
  AOI22_X1 U9982 ( .A1(n28980), .A2(\xmem_data[42][7] ), .B1(n24597), .B2(
        \xmem_data[43][7] ), .ZN(n6464) );
  AOI22_X1 U9983 ( .A1(n31328), .A2(\xmem_data[44][7] ), .B1(n29188), .B2(
        \xmem_data[45][7] ), .ZN(n6463) );
  AOI22_X1 U9984 ( .A1(n31330), .A2(\xmem_data[46][7] ), .B1(n31329), .B2(
        \xmem_data[47][7] ), .ZN(n6462) );
  NAND4_X1 U9985 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n6476)
         );
  AOI22_X1 U9986 ( .A1(n23802), .A2(\xmem_data[48][7] ), .B1(n24592), .B2(
        \xmem_data[49][7] ), .ZN(n6469) );
  AOI22_X1 U9987 ( .A1(n28428), .A2(\xmem_data[50][7] ), .B1(n28429), .B2(
        \xmem_data[51][7] ), .ZN(n6468) );
  AOI22_X1 U9988 ( .A1(n31315), .A2(\xmem_data[52][7] ), .B1(n31314), .B2(
        \xmem_data[53][7] ), .ZN(n6467) );
  AOI22_X1 U9989 ( .A1(n31316), .A2(\xmem_data[54][7] ), .B1(n28500), .B2(
        \xmem_data[55][7] ), .ZN(n6466) );
  NAND4_X1 U9990 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n6475)
         );
  AOI22_X1 U9991 ( .A1(n31308), .A2(\xmem_data[56][7] ), .B1(n20769), .B2(
        \xmem_data[57][7] ), .ZN(n6473) );
  AOI22_X1 U9992 ( .A1(n17056), .A2(\xmem_data[58][7] ), .B1(n31309), .B2(
        \xmem_data[59][7] ), .ZN(n6472) );
  AOI22_X1 U9993 ( .A1(n21308), .A2(\xmem_data[60][7] ), .B1(n28501), .B2(
        \xmem_data[61][7] ), .ZN(n6471) );
  AOI22_X1 U9994 ( .A1(n31348), .A2(\xmem_data[62][7] ), .B1(n3222), .B2(
        \xmem_data[63][7] ), .ZN(n6470) );
  NAND4_X1 U9995 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6474)
         );
  OR4_X1 U9996 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n6478) );
  AND2_X1 U9997 ( .A1(n6478), .A2(n31340), .ZN(n6479) );
  XNOR2_X1 U9998 ( .A(n35122), .B(\fmem_data[12][3] ), .ZN(n25603) );
  XOR2_X1 U9999 ( .A(\fmem_data[12][3] ), .B(\fmem_data[12][2] ), .Z(n6482) );
  AND2_X1 U10000 ( .A1(n33582), .A2(n34340), .ZN(n6483) );
  OR2_X1 U10001 ( .A1(n25603), .A2(n6483), .ZN(n33239) );
  XOR2_X1 U10002 ( .A(\fmem_data[14][3] ), .B(\fmem_data[14][2] ), .Z(n6484)
         );
  XOR2_X1 U10003 ( .A(n39040), .B(n6489), .Z(n6578) );
  INV_X1 U10004 ( .A(n6578), .ZN(n6554) );
  INV_X1 U10005 ( .A(n6489), .ZN(n6490) );
  AOI21_X1 U10006 ( .B1(n39041), .B2(n6491), .A(n6490), .ZN(n6579) );
  AND2_X1 U10007 ( .A1(n6554), .A2(n6579), .ZN(n27968) );
  AOI22_X1 U10008 ( .A1(n31348), .A2(\xmem_data[32][7] ), .B1(n3218), .B2(
        \xmem_data[33][7] ), .ZN(n6495) );
  AOI22_X1 U10009 ( .A1(n20805), .A2(\xmem_data[34][7] ), .B1(n24695), .B2(
        \xmem_data[35][7] ), .ZN(n6494) );
  AOI22_X1 U10010 ( .A1(n27938), .A2(\xmem_data[36][7] ), .B1(n3256), .B2(
        \xmem_data[37][7] ), .ZN(n6493) );
  AOI22_X1 U10011 ( .A1(n30295), .A2(\xmem_data[38][7] ), .B1(n28343), .B2(
        \xmem_data[39][7] ), .ZN(n6492) );
  NAND4_X1 U10012 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6511)
         );
  AOI22_X1 U10013 ( .A1(n24606), .A2(\xmem_data[56][7] ), .B1(n17003), .B2(
        \xmem_data[57][7] ), .ZN(n6499) );
  BUF_X1 U10014 ( .A(n13457), .Z(n27957) );
  AOI22_X1 U10015 ( .A1(n28467), .A2(\xmem_data[58][7] ), .B1(n27957), .B2(
        \xmem_data[59][7] ), .ZN(n6498) );
  BUF_X1 U10016 ( .A(n31263), .Z(n27959) );
  BUF_X1 U10017 ( .A(n28947), .Z(n27958) );
  AOI22_X1 U10018 ( .A1(n27959), .A2(\xmem_data[60][7] ), .B1(n27958), .B2(
        \xmem_data[61][7] ), .ZN(n6497) );
  AOI22_X1 U10019 ( .A1(n23732), .A2(\xmem_data[62][7] ), .B1(n31347), .B2(
        \xmem_data[63][7] ), .ZN(n6496) );
  NAND4_X1 U10020 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6510)
         );
  AOI22_X1 U10021 ( .A1(n20809), .A2(\xmem_data[40][7] ), .B1(n24590), .B2(
        \xmem_data[41][7] ), .ZN(n6503) );
  BUF_X1 U10022 ( .A(n14997), .Z(n27944) );
  AOI22_X1 U10023 ( .A1(n27944), .A2(\xmem_data[42][7] ), .B1(n24212), .B2(
        \xmem_data[43][7] ), .ZN(n6502) );
  AOI22_X1 U10024 ( .A1(n31268), .A2(\xmem_data[44][7] ), .B1(n29009), .B2(
        \xmem_data[45][7] ), .ZN(n6501) );
  BUF_X1 U10025 ( .A(n29187), .Z(n27945) );
  AOI22_X1 U10026 ( .A1(n29237), .A2(\xmem_data[46][7] ), .B1(n27516), .B2(
        \xmem_data[47][7] ), .ZN(n6500) );
  NAND4_X1 U10027 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n6509)
         );
  AOI22_X1 U10028 ( .A1(n21007), .A2(\xmem_data[48][7] ), .B1(n22718), .B2(
        \xmem_data[49][7] ), .ZN(n6507) );
  BUF_X1 U10029 ( .A(n13452), .Z(n27950) );
  AOI22_X1 U10030 ( .A1(n29319), .A2(\xmem_data[50][7] ), .B1(n27950), .B2(
        \xmem_data[51][7] ), .ZN(n6506) );
  BUF_X1 U10031 ( .A(n14881), .Z(n27952) );
  BUF_X1 U10032 ( .A(n14973), .Z(n27951) );
  AOI22_X1 U10033 ( .A1(n27952), .A2(\xmem_data[52][7] ), .B1(n27951), .B2(
        \xmem_data[53][7] ), .ZN(n6505) );
  AOI22_X1 U10034 ( .A1(n24571), .A2(\xmem_data[54][7] ), .B1(n28062), .B2(
        \xmem_data[55][7] ), .ZN(n6504) );
  NAND4_X1 U10035 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .ZN(n6508)
         );
  OR4_X1 U10036 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(n6533)
         );
  BUF_X1 U10037 ( .A(n29064), .Z(n27902) );
  AOI22_X1 U10038 ( .A1(n27902), .A2(\xmem_data[96][7] ), .B1(n3217), .B2(
        \xmem_data[97][7] ), .ZN(n6515) );
  AOI22_X1 U10039 ( .A1(n17033), .A2(\xmem_data[98][7] ), .B1(n30963), .B2(
        \xmem_data[99][7] ), .ZN(n6514) );
  BUF_X1 U10040 ( .A(n14926), .Z(n27904) );
  BUF_X1 U10041 ( .A(n14927), .Z(n27903) );
  AOI22_X1 U10042 ( .A1(n27904), .A2(\xmem_data[100][7] ), .B1(n27903), .B2(
        \xmem_data[101][7] ), .ZN(n6513) );
  BUF_X1 U10043 ( .A(n14991), .Z(n27905) );
  AOI22_X1 U10044 ( .A1(n27905), .A2(\xmem_data[102][7] ), .B1(n25514), .B2(
        \xmem_data[103][7] ), .ZN(n6512) );
  NAND4_X1 U10045 ( .A1(n6515), .A2(n6514), .A3(n6513), .A4(n6512), .ZN(n6531)
         );
  AOI22_X1 U10046 ( .A1(n20818), .A2(\xmem_data[120][7] ), .B1(n30496), .B2(
        \xmem_data[121][7] ), .ZN(n6519) );
  AOI22_X1 U10047 ( .A1(n28467), .A2(\xmem_data[122][7] ), .B1(n20769), .B2(
        \xmem_data[123][7] ), .ZN(n6518) );
  BUF_X1 U10048 ( .A(n31263), .Z(n27925) );
  AOI22_X1 U10049 ( .A1(n27925), .A2(\xmem_data[124][7] ), .B1(n22729), .B2(
        \xmem_data[125][7] ), .ZN(n6517) );
  AOI22_X1 U10050 ( .A1(n3333), .A2(\xmem_data[126][7] ), .B1(n24172), .B2(
        \xmem_data[127][7] ), .ZN(n6516) );
  NAND4_X1 U10051 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n6530)
         );
  BUF_X1 U10052 ( .A(n25604), .Z(n27910) );
  AOI22_X1 U10053 ( .A1(n27910), .A2(\xmem_data[104][7] ), .B1(n3357), .B2(
        \xmem_data[105][7] ), .ZN(n6523) );
  BUF_X1 U10054 ( .A(n14997), .Z(n27911) );
  AOI22_X1 U10055 ( .A1(n27911), .A2(\xmem_data[106][7] ), .B1(n24132), .B2(
        \xmem_data[107][7] ), .ZN(n6522) );
  BUF_X1 U10056 ( .A(n13476), .Z(n27913) );
  BUF_X1 U10057 ( .A(n14935), .Z(n27912) );
  AOI22_X1 U10058 ( .A1(n3176), .A2(\xmem_data[108][7] ), .B1(n27912), .B2(
        \xmem_data[109][7] ), .ZN(n6521) );
  AOI22_X1 U10059 ( .A1(n20939), .A2(\xmem_data[110][7] ), .B1(n25383), .B2(
        \xmem_data[111][7] ), .ZN(n6520) );
  NAND4_X1 U10060 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n6529)
         );
  BUF_X1 U10061 ( .A(n14937), .Z(n27919) );
  BUF_X1 U10062 ( .A(n13415), .Z(n27918) );
  AOI22_X1 U10063 ( .A1(n27919), .A2(\xmem_data[112][7] ), .B1(n27918), .B2(
        \xmem_data[113][7] ), .ZN(n6527) );
  BUF_X1 U10064 ( .A(n13452), .Z(n27920) );
  AOI22_X1 U10065 ( .A1(n30872), .A2(\xmem_data[114][7] ), .B1(n27920), .B2(
        \xmem_data[115][7] ), .ZN(n6526) );
  AOI22_X1 U10066 ( .A1(n20593), .A2(\xmem_data[116][7] ), .B1(n17001), .B2(
        \xmem_data[117][7] ), .ZN(n6525) );
  AOI22_X1 U10067 ( .A1(n28955), .A2(\xmem_data[118][7] ), .B1(n31362), .B2(
        \xmem_data[119][7] ), .ZN(n6524) );
  NAND4_X1 U10068 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n6528)
         );
  AND2_X1 U10069 ( .A1(n6579), .A2(n6578), .ZN(n27937) );
  AOI22_X1 U10070 ( .A1(n24467), .A2(\xmem_data[88][7] ), .B1(n25723), .B2(
        \xmem_data[89][7] ), .ZN(n6537) );
  AOI22_X1 U10071 ( .A1(n27959), .A2(\xmem_data[92][7] ), .B1(n27958), .B2(
        \xmem_data[93][7] ), .ZN(n6536) );
  AOI22_X1 U10072 ( .A1(n27498), .A2(\xmem_data[90][7] ), .B1(n27957), .B2(
        \xmem_data[91][7] ), .ZN(n6535) );
  AOI22_X1 U10073 ( .A1(n3414), .A2(\xmem_data[94][7] ), .B1(n29286), .B2(
        \xmem_data[95][7] ), .ZN(n6534) );
  NAND4_X1 U10074 ( .A1(n6537), .A2(n6536), .A3(n6535), .A4(n6534), .ZN(n6553)
         );
  AOI22_X1 U10075 ( .A1(n25508), .A2(\xmem_data[64][7] ), .B1(n3222), .B2(
        \xmem_data[65][7] ), .ZN(n6541) );
  AOI22_X1 U10076 ( .A1(n30593), .A2(\xmem_data[66][7] ), .B1(n20558), .B2(
        \xmem_data[67][7] ), .ZN(n6540) );
  AOI22_X1 U10077 ( .A1(n27938), .A2(\xmem_data[68][7] ), .B1(n22759), .B2(
        \xmem_data[69][7] ), .ZN(n6539) );
  AOI22_X1 U10078 ( .A1(n22668), .A2(\xmem_data[70][7] ), .B1(n24553), .B2(
        \xmem_data[71][7] ), .ZN(n6538) );
  NAND4_X1 U10079 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6552)
         );
  AOI22_X1 U10080 ( .A1(n13149), .A2(\xmem_data[80][7] ), .B1(n24546), .B2(
        \xmem_data[81][7] ), .ZN(n6545) );
  AOI22_X1 U10081 ( .A1(n23802), .A2(\xmem_data[82][7] ), .B1(n27950), .B2(
        \xmem_data[83][7] ), .ZN(n6544) );
  AOI22_X1 U10082 ( .A1(n27952), .A2(\xmem_data[84][7] ), .B1(n27951), .B2(
        \xmem_data[85][7] ), .ZN(n6543) );
  AOI22_X1 U10083 ( .A1(n24522), .A2(\xmem_data[86][7] ), .B1(n31362), .B2(
        \xmem_data[87][7] ), .ZN(n6542) );
  NAND4_X1 U10084 ( .A1(n6545), .A2(n6544), .A3(n6543), .A4(n6542), .ZN(n6551)
         );
  AOI22_X1 U10085 ( .A1(n20809), .A2(\xmem_data[72][7] ), .B1(n28415), .B2(
        \xmem_data[73][7] ), .ZN(n6549) );
  AOI22_X1 U10086 ( .A1(n27944), .A2(\xmem_data[74][7] ), .B1(n24212), .B2(
        \xmem_data[75][7] ), .ZN(n6548) );
  AOI22_X1 U10087 ( .A1(n3175), .A2(\xmem_data[76][7] ), .B1(n22703), .B2(
        \xmem_data[77][7] ), .ZN(n6547) );
  AOI22_X1 U10088 ( .A1(n29315), .A2(\xmem_data[78][7] ), .B1(n3208), .B2(
        \xmem_data[79][7] ), .ZN(n6546) );
  NAND4_X1 U10089 ( .A1(n6549), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(n6550)
         );
  NOR2_X1 U10090 ( .A1(n6579), .A2(n6554), .ZN(n27935) );
  AOI22_X1 U10091 ( .A1(n28355), .A2(\xmem_data[0][7] ), .B1(n3220), .B2(
        \xmem_data[1][7] ), .ZN(n6558) );
  AOI22_X1 U10092 ( .A1(n25490), .A2(\xmem_data[4][7] ), .B1(n30882), .B2(
        \xmem_data[5][7] ), .ZN(n6557) );
  BUF_X1 U10093 ( .A(n14925), .Z(n27869) );
  AOI22_X1 U10094 ( .A1(n29565), .A2(\xmem_data[2][7] ), .B1(n27869), .B2(
        \xmem_data[3][7] ), .ZN(n6556) );
  NAND3_X1 U10095 ( .A1(n6558), .A2(n6557), .A3(n6556), .ZN(n6574) );
  BUF_X1 U10096 ( .A(n10999), .Z(n27863) );
  AOI22_X1 U10097 ( .A1(n27910), .A2(\xmem_data[8][7] ), .B1(n27863), .B2(
        \xmem_data[9][7] ), .ZN(n6562) );
  AOI22_X1 U10098 ( .A1(n27763), .A2(\xmem_data[10][7] ), .B1(n31326), .B2(
        \xmem_data[11][7] ), .ZN(n6561) );
  AOI22_X1 U10099 ( .A1(n25425), .A2(\xmem_data[12][7] ), .B1(n25382), .B2(
        \xmem_data[13][7] ), .ZN(n6560) );
  BUF_X1 U10100 ( .A(n14936), .Z(n27864) );
  AOI22_X1 U10101 ( .A1(n30666), .A2(\xmem_data[14][7] ), .B1(n27864), .B2(
        \xmem_data[15][7] ), .ZN(n6559) );
  NAND4_X1 U10102 ( .A1(n6562), .A2(n6561), .A3(n6560), .A4(n6559), .ZN(n6573)
         );
  AOI22_X1 U10103 ( .A1(n28096), .A2(\xmem_data[16][7] ), .B1(n24459), .B2(
        \xmem_data[17][7] ), .ZN(n6566) );
  BUF_X1 U10104 ( .A(n14971), .Z(n27855) );
  AOI22_X1 U10105 ( .A1(n27855), .A2(\xmem_data[18][7] ), .B1(n24116), .B2(
        \xmem_data[19][7] ), .ZN(n6565) );
  BUF_X1 U10106 ( .A(n14882), .Z(n27856) );
  AOI22_X1 U10107 ( .A1(n30956), .A2(\xmem_data[20][7] ), .B1(n25679), .B2(
        \xmem_data[21][7] ), .ZN(n6564) );
  AOI22_X1 U10108 ( .A1(n30686), .A2(\xmem_data[22][7] ), .B1(n27975), .B2(
        \xmem_data[23][7] ), .ZN(n6563) );
  NAND4_X1 U10109 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .ZN(n6572)
         );
  BUF_X1 U10110 ( .A(n14976), .Z(n27847) );
  AOI22_X1 U10111 ( .A1(n27847), .A2(\xmem_data[24][7] ), .B1(n28468), .B2(
        \xmem_data[25][7] ), .ZN(n6570) );
  BUF_X1 U10112 ( .A(n13127), .Z(n27852) );
  AOI22_X1 U10113 ( .A1(n27852), .A2(\xmem_data[26][7] ), .B1(n25528), .B2(
        \xmem_data[27][7] ), .ZN(n6569) );
  AOI22_X1 U10114 ( .A1(n20710), .A2(\xmem_data[28][7] ), .B1(n25357), .B2(
        \xmem_data[29][7] ), .ZN(n6568) );
  AOI22_X1 U10115 ( .A1(n3153), .A2(\xmem_data[30][7] ), .B1(n25360), .B2(
        \xmem_data[31][7] ), .ZN(n6567) );
  NAND4_X1 U10116 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n6571)
         );
  OR4_X1 U10117 ( .A1(n6574), .A2(n6573), .A3(n6572), .A4(n6571), .ZN(n6581)
         );
  AND2_X1 U10118 ( .A1(n3345), .A2(\xmem_data[6][7] ), .ZN(n6575) );
  NOR2_X1 U10119 ( .A1(n6579), .A2(n6578), .ZN(n9896) );
  INV_X1 U10120 ( .A(n9896), .ZN(n27877) );
  XNOR2_X1 U10121 ( .A(n35102), .B(\fmem_data[14][3] ), .ZN(n25602) );
  INV_X1 U10122 ( .A(n6585), .ZN(n33240) );
  AOI22_X1 U10123 ( .A1(n24511), .A2(\xmem_data[72][3] ), .B1(n21009), .B2(
        \xmem_data[73][3] ), .ZN(n6594) );
  NOR2_X1 U10124 ( .A1(n6586), .A2(n39010), .ZN(n6621) );
  INV_X1 U10125 ( .A(n6621), .ZN(n8856) );
  AND2_X1 U10126 ( .A1(n8856), .A2(n9417), .ZN(n6587) );
  OR3_X1 U10127 ( .A1(n8409), .A2(n3248), .A3(n6587), .ZN(n6613) );
  AND2_X1 U10128 ( .A1(n10590), .A2(n8409), .ZN(n6588) );
  NOR2_X1 U10129 ( .A1(n10589), .A2(n6588), .ZN(n6816) );
  INV_X1 U10130 ( .A(n10590), .ZN(n6589) );
  OR2_X1 U10131 ( .A1(n6621), .A2(n6990), .ZN(n10069) );
  OR2_X1 U10132 ( .A1(n6612), .A2(n6611), .ZN(n6590) );
  NOR2_X1 U10133 ( .A1(n6613), .A2(n6590), .ZN(n6675) );
  AOI22_X1 U10134 ( .A1(n3271), .A2(\xmem_data[74][3] ), .B1(n3200), .B2(
        \xmem_data[75][3] ), .ZN(n6593) );
  AOI22_X1 U10135 ( .A1(n20552), .A2(\xmem_data[76][3] ), .B1(n25527), .B2(
        \xmem_data[77][3] ), .ZN(n6592) );
  AOI22_X1 U10136 ( .A1(n13420), .A2(\xmem_data[78][3] ), .B1(n20769), .B2(
        \xmem_data[79][3] ), .ZN(n6591) );
  BUF_X1 U10137 ( .A(n28973), .Z(n16980) );
  NAND2_X1 U10138 ( .A1(n6612), .A2(n6611), .ZN(n6595) );
  NOR2_X1 U10139 ( .A1(n6613), .A2(n6595), .ZN(n6680) );
  AOI22_X1 U10140 ( .A1(n16980), .A2(\xmem_data[82][3] ), .B1(n16979), .B2(
        \xmem_data[83][3] ), .ZN(n6596) );
  INV_X1 U10141 ( .A(n6596), .ZN(n6597) );
  AOI21_X1 U10142 ( .B1(n21066), .B2(\xmem_data[84][3] ), .A(n6597), .ZN(n6620) );
  AOI22_X1 U10143 ( .A1(n3342), .A2(\xmem_data[88][3] ), .B1(n30882), .B2(
        \xmem_data[89][3] ), .ZN(n6603) );
  BUF_X1 U10144 ( .A(n14991), .Z(n16973) );
  INV_X1 U10145 ( .A(n6611), .ZN(n6598) );
  NAND2_X1 U10146 ( .A1(n6612), .A2(n6598), .ZN(n6599) );
  NOR2_X1 U10147 ( .A1(n6613), .A2(n6599), .ZN(n6685) );
  BUF_X1 U10148 ( .A(n6685), .Z(n16972) );
  AOI22_X1 U10149 ( .A1(n16973), .A2(\xmem_data[90][3] ), .B1(n16972), .B2(
        \xmem_data[91][3] ), .ZN(n6602) );
  BUF_X1 U10150 ( .A(n25604), .Z(n16974) );
  AOI22_X1 U10151 ( .A1(n16974), .A2(\xmem_data[92][3] ), .B1(n3358), .B2(
        \xmem_data[93][3] ), .ZN(n6601) );
  AOI22_X1 U10152 ( .A1(n25424), .A2(\xmem_data[94][3] ), .B1(n28375), .B2(
        \xmem_data[95][3] ), .ZN(n6600) );
  NAND4_X1 U10153 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6610)
         );
  NAND2_X1 U10154 ( .A1(n3221), .A2(\xmem_data[85][3] ), .ZN(n6605) );
  NAND2_X1 U10155 ( .A1(n17056), .A2(\xmem_data[80][3] ), .ZN(n6604) );
  NAND2_X1 U10156 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  AOI21_X1 U10157 ( .B1(n27563), .B2(\xmem_data[81][3] ), .A(n6606), .ZN(n6608) );
  AOI22_X1 U10158 ( .A1(n25731), .A2(\xmem_data[86][3] ), .B1(n20598), .B2(
        \xmem_data[87][3] ), .ZN(n6607) );
  NAND2_X1 U10159 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  NOR2_X1 U10160 ( .A1(n6610), .A2(n6609), .ZN(n6619) );
  AOI22_X1 U10161 ( .A1(n16986), .A2(\xmem_data[64][3] ), .B1(n24160), .B2(
        \xmem_data[65][3] ), .ZN(n6618) );
  BUF_X1 U10162 ( .A(n3464), .Z(n16988) );
  OR2_X1 U10163 ( .A1(n6612), .A2(n6598), .ZN(n6614) );
  NOR2_X1 U10164 ( .A1(n6614), .A2(n6613), .ZN(n17042) );
  BUF_X1 U10165 ( .A(n17042), .Z(n16987) );
  AOI22_X1 U10166 ( .A1(n16988), .A2(\xmem_data[66][3] ), .B1(n16987), .B2(
        \xmem_data[67][3] ), .ZN(n6617) );
  BUF_X1 U10167 ( .A(n14970), .Z(n16989) );
  AOI22_X1 U10168 ( .A1(n28337), .A2(\xmem_data[68][3] ), .B1(n16989), .B2(
        \xmem_data[69][3] ), .ZN(n6616) );
  BUF_X1 U10169 ( .A(n14971), .Z(n16990) );
  AOI22_X1 U10170 ( .A1(n16990), .A2(\xmem_data[70][3] ), .B1(n28097), .B2(
        \xmem_data[71][3] ), .ZN(n6615) );
  NAND4_X1 U10171 ( .A1(n3509), .A2(n6620), .A3(n6619), .A4(n3846), .ZN(n6624)
         );
  NAND2_X1 U10172 ( .A1(n7216), .A2(n6621), .ZN(n6622) );
  NOR2_X1 U10173 ( .A1(n8856), .A2(n11381), .ZN(n6623) );
  AOI21_X1 U10174 ( .B1(n4499), .B2(n6622), .A(n6623), .ZN(n6695) );
  XOR2_X1 U10175 ( .A(n6623), .B(load_xaddr_val[6]), .Z(n6694) );
  INV_X1 U10176 ( .A(n6694), .ZN(n6669) );
  NAND2_X1 U10177 ( .A1(n6624), .A2(n16966), .ZN(n6700) );
  AOI22_X1 U10178 ( .A1(n27974), .A2(\xmem_data[104][3] ), .B1(n24222), .B2(
        \xmem_data[105][3] ), .ZN(n6628) );
  AOI22_X1 U10179 ( .A1(n3270), .A2(\xmem_data[106][3] ), .B1(n3200), .B2(
        \xmem_data[107][3] ), .ZN(n6627) );
  AOI22_X1 U10180 ( .A1(n29151), .A2(\xmem_data[108][3] ), .B1(n23781), .B2(
        \xmem_data[109][3] ), .ZN(n6626) );
  AOI22_X1 U10181 ( .A1(n31308), .A2(\xmem_data[110][3] ), .B1(n25388), .B2(
        \xmem_data[111][3] ), .ZN(n6625) );
  AOI22_X1 U10182 ( .A1(n16980), .A2(\xmem_data[114][3] ), .B1(n16979), .B2(
        \xmem_data[115][3] ), .ZN(n6629) );
  INV_X1 U10183 ( .A(n6629), .ZN(n6630) );
  AOI21_X1 U10184 ( .B1(n28364), .B2(\xmem_data[116][3] ), .A(n6630), .ZN(
        n6647) );
  AOI22_X1 U10185 ( .A1(n22709), .A2(\xmem_data[120][3] ), .B1(n27903), .B2(
        \xmem_data[121][3] ), .ZN(n6634) );
  AOI22_X1 U10186 ( .A1(n16973), .A2(\xmem_data[122][3] ), .B1(n16972), .B2(
        \xmem_data[123][3] ), .ZN(n6633) );
  AOI22_X1 U10187 ( .A1(n16974), .A2(\xmem_data[124][3] ), .B1(n27943), .B2(
        \xmem_data[125][3] ), .ZN(n6632) );
  AOI22_X1 U10188 ( .A1(n30943), .A2(\xmem_data[126][3] ), .B1(n30552), .B2(
        \xmem_data[127][3] ), .ZN(n6631) );
  NAND4_X1 U10189 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6641)
         );
  NAND2_X1 U10190 ( .A1(n3220), .A2(\xmem_data[117][3] ), .ZN(n6636) );
  NAND2_X1 U10191 ( .A1(n17056), .A2(\xmem_data[112][3] ), .ZN(n6635) );
  NAND2_X1 U10192 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  AOI21_X1 U10193 ( .B1(n25685), .B2(\xmem_data[113][3] ), .A(n6637), .ZN(
        n6639) );
  AOI22_X1 U10194 ( .A1(n24563), .A2(\xmem_data[118][3] ), .B1(n24695), .B2(
        \xmem_data[119][3] ), .ZN(n6638) );
  NAND2_X1 U10195 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  NOR2_X1 U10196 ( .A1(n6641), .A2(n6640), .ZN(n6646) );
  AOI22_X1 U10197 ( .A1(n16986), .A2(\xmem_data[96][3] ), .B1(n28090), .B2(
        \xmem_data[97][3] ), .ZN(n6645) );
  AOI22_X1 U10198 ( .A1(n16988), .A2(\xmem_data[98][3] ), .B1(n16987), .B2(
        \xmem_data[99][3] ), .ZN(n6644) );
  AOI22_X1 U10199 ( .A1(n13149), .A2(\xmem_data[100][3] ), .B1(n16989), .B2(
        \xmem_data[101][3] ), .ZN(n6643) );
  AOI22_X1 U10200 ( .A1(n16990), .A2(\xmem_data[102][3] ), .B1(n23801), .B2(
        \xmem_data[103][3] ), .ZN(n6642) );
  NAND4_X1 U10201 ( .A1(n3510), .A2(n6647), .A3(n6646), .A4(n3847), .ZN(n6648)
         );
  AND2_X1 U10202 ( .A1(n6695), .A2(n6694), .ZN(n16997) );
  NAND2_X1 U10203 ( .A1(n6648), .A2(n16997), .ZN(n6699) );
  AOI22_X1 U10204 ( .A1(n31268), .A2(\xmem_data[32][3] ), .B1(n23793), .B2(
        \xmem_data[33][3] ), .ZN(n6652) );
  BUF_X1 U10205 ( .A(n3464), .Z(n17018) );
  AOI22_X1 U10206 ( .A1(n29396), .A2(\xmem_data[34][3] ), .B1(n3202), .B2(
        \xmem_data[35][3] ), .ZN(n6651) );
  BUF_X1 U10207 ( .A(n14937), .Z(n17020) );
  AOI22_X1 U10208 ( .A1(n17020), .A2(\xmem_data[36][3] ), .B1(n29048), .B2(
        \xmem_data[37][3] ), .ZN(n6650) );
  BUF_X1 U10209 ( .A(n14971), .Z(n17021) );
  AOI22_X1 U10210 ( .A1(n17021), .A2(\xmem_data[38][3] ), .B1(n20941), .B2(
        \xmem_data[39][3] ), .ZN(n6649) );
  NAND4_X1 U10211 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6668)
         );
  BUF_X1 U10212 ( .A(n3324), .Z(n17002) );
  BUF_X1 U10213 ( .A(n14973), .Z(n17001) );
  AOI22_X1 U10214 ( .A1(n24615), .A2(\xmem_data[40][3] ), .B1(n17001), .B2(
        \xmem_data[41][3] ), .ZN(n6656) );
  BUF_X1 U10215 ( .A(n14974), .Z(n17004) );
  AOI22_X1 U10216 ( .A1(n17004), .A2(\xmem_data[42][3] ), .B1(n3199), .B2(
        \xmem_data[43][3] ), .ZN(n6655) );
  BUF_X1 U10217 ( .A(n14981), .Z(n17003) );
  AOI22_X1 U10218 ( .A1(n27847), .A2(\xmem_data[44][3] ), .B1(n17003), .B2(
        \xmem_data[45][3] ), .ZN(n6654) );
  BUF_X1 U10219 ( .A(n13457), .Z(n16999) );
  AOI22_X1 U10220 ( .A1(n20952), .A2(\xmem_data[46][3] ), .B1(n16999), .B2(
        \xmem_data[47][3] ), .ZN(n6653) );
  NAND4_X1 U10221 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6667)
         );
  BUF_X1 U10222 ( .A(n31263), .Z(n17030) );
  AOI22_X1 U10223 ( .A1(n17030), .A2(\xmem_data[48][3] ), .B1(n22729), .B2(
        \xmem_data[49][3] ), .ZN(n6660) );
  BUF_X1 U10224 ( .A(n6680), .Z(n17031) );
  AOI22_X1 U10225 ( .A1(n3388), .A2(\xmem_data[50][3] ), .B1(n17031), .B2(
        \xmem_data[51][3] ), .ZN(n6659) );
  AOI22_X1 U10226 ( .A1(n31348), .A2(\xmem_data[52][3] ), .B1(n3219), .B2(
        \xmem_data[53][3] ), .ZN(n6658) );
  BUF_X1 U10227 ( .A(n14988), .Z(n17033) );
  AOI22_X1 U10228 ( .A1(n17033), .A2(\xmem_data[54][3] ), .B1(n22710), .B2(
        \xmem_data[55][3] ), .ZN(n6657) );
  NAND4_X1 U10229 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6666)
         );
  BUF_X1 U10230 ( .A(n14990), .Z(n17010) );
  AOI22_X1 U10231 ( .A1(n17010), .A2(\xmem_data[56][3] ), .B1(n21068), .B2(
        \xmem_data[57][3] ), .ZN(n6664) );
  BUF_X1 U10232 ( .A(n6685), .Z(n17011) );
  AOI22_X1 U10233 ( .A1(n29762), .A2(\xmem_data[58][3] ), .B1(n17011), .B2(
        \xmem_data[59][3] ), .ZN(n6663) );
  AOI22_X1 U10234 ( .A1(n28050), .A2(\xmem_data[60][3] ), .B1(n22739), .B2(
        \xmem_data[61][3] ), .ZN(n6662) );
  BUF_X1 U10235 ( .A(n14997), .Z(n17013) );
  BUF_X1 U10236 ( .A(n13435), .Z(n17012) );
  AOI22_X1 U10237 ( .A1(n17013), .A2(\xmem_data[62][3] ), .B1(n17012), .B2(
        \xmem_data[63][3] ), .ZN(n6661) );
  NAND4_X1 U10238 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6665)
         );
  OR4_X1 U10239 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6670)
         );
  AND2_X1 U10240 ( .A1(n6669), .A2(n6695), .ZN(n17038) );
  NAND2_X1 U10241 ( .A1(n6670), .A2(n17038), .ZN(n6698) );
  AOI22_X1 U10242 ( .A1(n17041), .A2(\xmem_data[0][3] ), .B1(n29271), .B2(
        \xmem_data[1][3] ), .ZN(n6674) );
  AOI22_X1 U10243 ( .A1(n28752), .A2(\xmem_data[2][3] ), .B1(n17019), .B2(
        \xmem_data[3][3] ), .ZN(n6673) );
  BUF_X1 U10244 ( .A(n13415), .Z(n17043) );
  AOI22_X1 U10245 ( .A1(n27919), .A2(\xmem_data[4][3] ), .B1(n17043), .B2(
        \xmem_data[5][3] ), .ZN(n6672) );
  BUF_X1 U10246 ( .A(n14971), .Z(n17044) );
  AOI22_X1 U10247 ( .A1(n17044), .A2(\xmem_data[6][3] ), .B1(n29318), .B2(
        \xmem_data[7][3] ), .ZN(n6671) );
  NAND4_X1 U10248 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6693)
         );
  AOI22_X1 U10249 ( .A1(n22683), .A2(\xmem_data[8][3] ), .B1(n29089), .B2(
        \xmem_data[9][3] ), .ZN(n6679) );
  AOI22_X1 U10250 ( .A1(n25401), .A2(\xmem_data[10][3] ), .B1(n3200), .B2(
        \xmem_data[11][3] ), .ZN(n6678) );
  BUF_X1 U10251 ( .A(n14919), .Z(n17049) );
  AOI22_X1 U10252 ( .A1(n24685), .A2(\xmem_data[12][3] ), .B1(n17049), .B2(
        \xmem_data[13][3] ), .ZN(n6677) );
  BUF_X1 U10253 ( .A(n13127), .Z(n17051) );
  BUF_X1 U10254 ( .A(n13457), .Z(n17050) );
  AOI22_X1 U10255 ( .A1(n17051), .A2(\xmem_data[14][3] ), .B1(n17050), .B2(
        \xmem_data[15][3] ), .ZN(n6676) );
  NAND4_X1 U10256 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6692)
         );
  BUF_X1 U10257 ( .A(n31263), .Z(n17056) );
  AOI22_X1 U10258 ( .A1(n17056), .A2(\xmem_data[16][3] ), .B1(n24470), .B2(
        \xmem_data[17][3] ), .ZN(n6684) );
  AOI22_X1 U10259 ( .A1(n3317), .A2(\xmem_data[18][3] ), .B1(n16979), .B2(
        \xmem_data[19][3] ), .ZN(n6683) );
  AOI22_X1 U10260 ( .A1(n30906), .A2(\xmem_data[20][3] ), .B1(n3219), .B2(
        \xmem_data[21][3] ), .ZN(n6682) );
  AOI22_X1 U10261 ( .A1(n23770), .A2(\xmem_data[22][3] ), .B1(n25509), .B2(
        \xmem_data[23][3] ), .ZN(n6681) );
  NAND4_X1 U10262 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6691)
         );
  BUF_X1 U10263 ( .A(n14927), .Z(n17061) );
  AOI22_X1 U10264 ( .A1(n29027), .A2(\xmem_data[24][3] ), .B1(n17061), .B2(
        \xmem_data[25][3] ), .ZN(n6689) );
  BUF_X1 U10265 ( .A(n14991), .Z(n17063) );
  BUF_X1 U10266 ( .A(n6685), .Z(n17062) );
  AOI22_X1 U10267 ( .A1(n17063), .A2(\xmem_data[26][3] ), .B1(n17062), .B2(
        \xmem_data[27][3] ), .ZN(n6688) );
  AOI22_X1 U10268 ( .A1(n25422), .A2(\xmem_data[28][3] ), .B1(n20588), .B2(
        \xmem_data[29][3] ), .ZN(n6687) );
  BUF_X1 U10269 ( .A(n14997), .Z(n17064) );
  AOI22_X1 U10270 ( .A1(n17064), .A2(\xmem_data[30][3] ), .B1(n28515), .B2(
        \xmem_data[31][3] ), .ZN(n6686) );
  NAND4_X1 U10271 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6690)
         );
  OR4_X1 U10272 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6696)
         );
  NOR2_X1 U10273 ( .A1(n6695), .A2(n6694), .ZN(n17073) );
  NAND2_X1 U10274 ( .A1(n6696), .A2(n17073), .ZN(n6697) );
  NAND4_X1 U10275 ( .A1(n6699), .A2(n6700), .A3(n6698), .A4(n6697), .ZN(n32165) );
  XNOR2_X1 U10276 ( .A(n32165), .B(\fmem_data[2][7] ), .ZN(n32019) );
  XOR2_X1 U10277 ( .A(\fmem_data[2][6] ), .B(\fmem_data[2][7] ), .Z(n6701) );
  AOI22_X1 U10278 ( .A1(n17041), .A2(\xmem_data[32][4] ), .B1(n23793), .B2(
        \xmem_data[33][4] ), .ZN(n6705) );
  AOI22_X1 U10279 ( .A1(n16988), .A2(\xmem_data[34][4] ), .B1(n16987), .B2(
        \xmem_data[35][4] ), .ZN(n6704) );
  AOI22_X1 U10280 ( .A1(n17020), .A2(\xmem_data[36][4] ), .B1(n25398), .B2(
        \xmem_data[37][4] ), .ZN(n6703) );
  AOI22_X1 U10281 ( .A1(n17021), .A2(\xmem_data[38][4] ), .B1(n30616), .B2(
        \xmem_data[39][4] ), .ZN(n6702) );
  NAND4_X1 U10282 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6721)
         );
  AOI22_X1 U10283 ( .A1(n17002), .A2(\xmem_data[40][4] ), .B1(n17001), .B2(
        \xmem_data[41][4] ), .ZN(n6709) );
  AOI22_X1 U10284 ( .A1(n17004), .A2(\xmem_data[42][4] ), .B1(n3201), .B2(
        \xmem_data[43][4] ), .ZN(n6708) );
  AOI22_X1 U10285 ( .A1(n24572), .A2(\xmem_data[44][4] ), .B1(n17003), .B2(
        \xmem_data[45][4] ), .ZN(n6707) );
  AOI22_X1 U10286 ( .A1(n20985), .A2(\xmem_data[46][4] ), .B1(n16999), .B2(
        \xmem_data[47][4] ), .ZN(n6706) );
  NAND4_X1 U10287 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n6720)
         );
  AOI22_X1 U10288 ( .A1(n17030), .A2(\xmem_data[48][4] ), .B1(n28037), .B2(
        \xmem_data[49][4] ), .ZN(n6713) );
  AOI22_X1 U10289 ( .A1(n3387), .A2(\xmem_data[50][4] ), .B1(n17031), .B2(
        \xmem_data[51][4] ), .ZN(n6712) );
  AOI22_X1 U10290 ( .A1(n28364), .A2(\xmem_data[52][4] ), .B1(n3222), .B2(
        \xmem_data[53][4] ), .ZN(n6711) );
  AOI22_X1 U10291 ( .A1(n17033), .A2(\xmem_data[54][4] ), .B1(n25562), .B2(
        \xmem_data[55][4] ), .ZN(n6710) );
  NAND4_X1 U10292 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6719)
         );
  AOI22_X1 U10293 ( .A1(n17010), .A2(\xmem_data[56][4] ), .B1(n27994), .B2(
        \xmem_data[57][4] ), .ZN(n6717) );
  AOI22_X1 U10294 ( .A1(n28308), .A2(\xmem_data[58][4] ), .B1(n17011), .B2(
        \xmem_data[59][4] ), .ZN(n6716) );
  AOI22_X1 U10295 ( .A1(n25422), .A2(\xmem_data[60][4] ), .B1(n24590), .B2(
        \xmem_data[61][4] ), .ZN(n6715) );
  AOI22_X1 U10296 ( .A1(n17013), .A2(\xmem_data[62][4] ), .B1(n17012), .B2(
        \xmem_data[63][4] ), .ZN(n6714) );
  NAND4_X1 U10297 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6718)
         );
  OR4_X1 U10298 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6743)
         );
  AOI22_X1 U10299 ( .A1(n17041), .A2(\xmem_data[0][4] ), .B1(n20544), .B2(
        \xmem_data[1][4] ), .ZN(n6725) );
  AOI22_X1 U10300 ( .A1(n29605), .A2(\xmem_data[2][4] ), .B1(n3202), .B2(
        \xmem_data[3][4] ), .ZN(n6724) );
  AOI22_X1 U10301 ( .A1(n21007), .A2(\xmem_data[4][4] ), .B1(n17043), .B2(
        \xmem_data[5][4] ), .ZN(n6723) );
  AOI22_X1 U10302 ( .A1(n17044), .A2(\xmem_data[6][4] ), .B1(n31254), .B2(
        \xmem_data[7][4] ), .ZN(n6722) );
  NAND4_X1 U10303 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6741)
         );
  AOI22_X1 U10304 ( .A1(n28385), .A2(\xmem_data[8][4] ), .B1(n28327), .B2(
        \xmem_data[9][4] ), .ZN(n6729) );
  AOI22_X1 U10305 ( .A1(n31315), .A2(\xmem_data[10][4] ), .B1(n3200), .B2(
        \xmem_data[11][4] ), .ZN(n6728) );
  AOI22_X1 U10306 ( .A1(n3171), .A2(\xmem_data[12][4] ), .B1(n17049), .B2(
        \xmem_data[13][4] ), .ZN(n6727) );
  AOI22_X1 U10307 ( .A1(n17051), .A2(\xmem_data[14][4] ), .B1(n17050), .B2(
        \xmem_data[15][4] ), .ZN(n6726) );
  NAND4_X1 U10308 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6740)
         );
  AOI22_X1 U10309 ( .A1(n31348), .A2(\xmem_data[20][4] ), .B1(n3222), .B2(
        \xmem_data[21][4] ), .ZN(n6733) );
  AOI22_X1 U10310 ( .A1(n3334), .A2(\xmem_data[18][4] ), .B1(n16979), .B2(
        \xmem_data[19][4] ), .ZN(n6732) );
  AOI22_X1 U10311 ( .A1(n17056), .A2(\xmem_data[16][4] ), .B1(n29328), .B2(
        \xmem_data[17][4] ), .ZN(n6731) );
  AOI22_X1 U10312 ( .A1(n20805), .A2(\xmem_data[22][4] ), .B1(n20723), .B2(
        \xmem_data[23][4] ), .ZN(n6730) );
  NAND4_X1 U10313 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6739)
         );
  AOI22_X1 U10314 ( .A1(n27938), .A2(\xmem_data[24][4] ), .B1(n17061), .B2(
        \xmem_data[25][4] ), .ZN(n6737) );
  AOI22_X1 U10315 ( .A1(n17063), .A2(\xmem_data[26][4] ), .B1(n17062), .B2(
        \xmem_data[27][4] ), .ZN(n6736) );
  AOI22_X1 U10316 ( .A1(n25422), .A2(\xmem_data[28][4] ), .B1(n28415), .B2(
        \xmem_data[29][4] ), .ZN(n6735) );
  AOI22_X1 U10317 ( .A1(n17064), .A2(\xmem_data[30][4] ), .B1(n23761), .B2(
        \xmem_data[31][4] ), .ZN(n6734) );
  NAND4_X1 U10318 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n6738)
         );
  OR4_X1 U10319 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6742)
         );
  AOI22_X1 U10320 ( .A1(n17038), .A2(n6743), .B1(n17073), .B2(n6742), .ZN(
        n6796) );
  AOI22_X1 U10321 ( .A1(n16980), .A2(\xmem_data[114][4] ), .B1(n16979), .B2(
        \xmem_data[115][4] ), .ZN(n6744) );
  INV_X1 U10322 ( .A(n6744), .ZN(n6745) );
  AOI21_X1 U10323 ( .B1(n28355), .B2(\xmem_data[116][4] ), .A(n6745), .ZN(
        n6771) );
  NAND2_X1 U10324 ( .A1(n3220), .A2(\xmem_data[117][4] ), .ZN(n6747) );
  NAND2_X1 U10325 ( .A1(n25724), .A2(\xmem_data[112][4] ), .ZN(n6746) );
  NAND2_X1 U10326 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  AOI21_X1 U10327 ( .B1(n24470), .B2(\xmem_data[113][4] ), .A(n6748), .ZN(
        n6750) );
  AOI22_X1 U10328 ( .A1(n30754), .A2(\xmem_data[110][4] ), .B1(n28329), .B2(
        \xmem_data[111][4] ), .ZN(n6749) );
  NAND2_X1 U10329 ( .A1(n6750), .A2(n6749), .ZN(n6760) );
  AOI22_X1 U10330 ( .A1(n16986), .A2(\xmem_data[96][4] ), .B1(n24160), .B2(
        \xmem_data[97][4] ), .ZN(n6752) );
  AOI22_X1 U10331 ( .A1(n17033), .A2(\xmem_data[118][4] ), .B1(n28319), .B2(
        \xmem_data[119][4] ), .ZN(n6751) );
  NAND2_X1 U10332 ( .A1(n6752), .A2(n6751), .ZN(n6758) );
  AOI22_X1 U10333 ( .A1(n16990), .A2(\xmem_data[102][4] ), .B1(n25367), .B2(
        \xmem_data[103][4] ), .ZN(n6756) );
  AOI22_X1 U10334 ( .A1(n3171), .A2(\xmem_data[108][4] ), .B1(n11008), .B2(
        \xmem_data[109][4] ), .ZN(n6755) );
  AOI22_X1 U10335 ( .A1(n20585), .A2(\xmem_data[100][4] ), .B1(n16989), .B2(
        \xmem_data[101][4] ), .ZN(n6754) );
  AOI22_X1 U10336 ( .A1(n3270), .A2(\xmem_data[106][4] ), .B1(n3200), .B2(
        \xmem_data[107][4] ), .ZN(n6753) );
  NAND4_X1 U10337 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6757)
         );
  OR2_X1 U10338 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NOR2_X1 U10339 ( .A1(n6760), .A2(n6759), .ZN(n6770) );
  AOI22_X1 U10340 ( .A1(n30606), .A2(\xmem_data[120][4] ), .B1(n28509), .B2(
        \xmem_data[121][4] ), .ZN(n6764) );
  AOI22_X1 U10341 ( .A1(n16973), .A2(\xmem_data[122][4] ), .B1(n16972), .B2(
        \xmem_data[123][4] ), .ZN(n6763) );
  AOI22_X1 U10342 ( .A1(n16974), .A2(\xmem_data[124][4] ), .B1(n24590), .B2(
        \xmem_data[125][4] ), .ZN(n6762) );
  AOI22_X1 U10343 ( .A1(n29451), .A2(\xmem_data[126][4] ), .B1(n24639), .B2(
        \xmem_data[127][4] ), .ZN(n6761) );
  AOI22_X1 U10344 ( .A1(n16988), .A2(\xmem_data[98][4] ), .B1(n16987), .B2(
        \xmem_data[99][4] ), .ZN(n6765) );
  INV_X1 U10345 ( .A(n6765), .ZN(n6768) );
  AOI22_X1 U10346 ( .A1(n27462), .A2(\xmem_data[104][4] ), .B1(n25679), .B2(
        \xmem_data[105][4] ), .ZN(n6766) );
  INV_X1 U10347 ( .A(n6766), .ZN(n6767) );
  NOR2_X1 U10348 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  NAND4_X1 U10349 ( .A1(n6771), .A2(n6770), .A3(n3793), .A4(n6769), .ZN(n6772)
         );
  NAND2_X1 U10350 ( .A1(n6772), .A2(n16997), .ZN(n6795) );
  AOI22_X1 U10351 ( .A1(n16986), .A2(\xmem_data[64][4] ), .B1(n29309), .B2(
        \xmem_data[65][4] ), .ZN(n6776) );
  AOI22_X1 U10352 ( .A1(n3465), .A2(\xmem_data[66][4] ), .B1(n17019), .B2(
        \xmem_data[67][4] ), .ZN(n6775) );
  AOI22_X1 U10353 ( .A1(n17020), .A2(\xmem_data[68][4] ), .B1(n27918), .B2(
        \xmem_data[69][4] ), .ZN(n6774) );
  AOI22_X1 U10354 ( .A1(n17021), .A2(\xmem_data[70][4] ), .B1(n24592), .B2(
        \xmem_data[71][4] ), .ZN(n6773) );
  NAND4_X1 U10355 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6792)
         );
  AOI22_X1 U10356 ( .A1(n24190), .A2(\xmem_data[72][4] ), .B1(n17001), .B2(
        \xmem_data[73][4] ), .ZN(n6780) );
  AOI22_X1 U10357 ( .A1(n17004), .A2(\xmem_data[74][4] ), .B1(n3200), .B2(
        \xmem_data[75][4] ), .ZN(n6779) );
  AOI22_X1 U10358 ( .A1(n20782), .A2(\xmem_data[76][4] ), .B1(n17003), .B2(
        \xmem_data[77][4] ), .ZN(n6778) );
  AOI22_X1 U10359 ( .A1(n29725), .A2(\xmem_data[78][4] ), .B1(n16999), .B2(
        \xmem_data[79][4] ), .ZN(n6777) );
  NAND4_X1 U10360 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6791)
         );
  AOI22_X1 U10361 ( .A1(n17030), .A2(\xmem_data[80][4] ), .B1(n28366), .B2(
        \xmem_data[81][4] ), .ZN(n6784) );
  AOI22_X1 U10362 ( .A1(n3387), .A2(\xmem_data[82][4] ), .B1(n17031), .B2(
        \xmem_data[83][4] ), .ZN(n6783) );
  AOI22_X1 U10363 ( .A1(n24694), .A2(\xmem_data[84][4] ), .B1(n3221), .B2(
        \xmem_data[85][4] ), .ZN(n6782) );
  AOI22_X1 U10364 ( .A1(n17033), .A2(\xmem_data[86][4] ), .B1(n20723), .B2(
        \xmem_data[87][4] ), .ZN(n6781) );
  NAND4_X1 U10365 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(n6790)
         );
  AOI22_X1 U10366 ( .A1(n17010), .A2(\xmem_data[88][4] ), .B1(n31275), .B2(
        \xmem_data[89][4] ), .ZN(n6788) );
  AOI22_X1 U10367 ( .A1(n25417), .A2(\xmem_data[90][4] ), .B1(n17011), .B2(
        \xmem_data[91][4] ), .ZN(n6787) );
  AOI22_X1 U10368 ( .A1(n30885), .A2(\xmem_data[92][4] ), .B1(n29180), .B2(
        \xmem_data[93][4] ), .ZN(n6786) );
  AOI22_X1 U10369 ( .A1(n17013), .A2(\xmem_data[94][4] ), .B1(n17012), .B2(
        \xmem_data[95][4] ), .ZN(n6785) );
  NAND4_X1 U10370 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6789)
         );
  OR4_X1 U10371 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6793)
         );
  NAND2_X1 U10372 ( .A1(n6793), .A2(n16966), .ZN(n6794) );
  XNOR2_X1 U10373 ( .A(n31221), .B(\fmem_data[2][7] ), .ZN(n33324) );
  OAI22_X1 U10374 ( .A1(n32019), .A2(n35721), .B1(n33324), .B2(n35722), .ZN(
        n33320) );
  BUF_X1 U10375 ( .A(n14973), .Z(n28291) );
  AOI22_X1 U10376 ( .A1(n27974), .A2(\xmem_data[120][5] ), .B1(n28291), .B2(
        \xmem_data[121][5] ), .ZN(n6800) );
  AOI22_X1 U10377 ( .A1(n31315), .A2(\xmem_data[122][5] ), .B1(n20949), .B2(
        \xmem_data[123][5] ), .ZN(n6799) );
  BUF_X1 U10378 ( .A(n13486), .Z(n28293) );
  BUF_X1 U10379 ( .A(n14981), .Z(n28292) );
  AOI22_X1 U10380 ( .A1(n28293), .A2(\xmem_data[124][5] ), .B1(n28292), .B2(
        \xmem_data[125][5] ), .ZN(n6798) );
  AOI22_X1 U10381 ( .A1(n29298), .A2(\xmem_data[126][5] ), .B1(n24468), .B2(
        \xmem_data[127][5] ), .ZN(n6797) );
  NAND4_X1 U10382 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6811)
         );
  AOI22_X1 U10383 ( .A1(n28298), .A2(\xmem_data[112][5] ), .B1(n24160), .B2(
        \xmem_data[113][5] ), .ZN(n6804) );
  BUF_X1 U10384 ( .A(n3464), .Z(n28300) );
  BUF_X1 U10385 ( .A(n14936), .Z(n28299) );
  AOI22_X1 U10386 ( .A1(n30303), .A2(\xmem_data[114][5] ), .B1(n28299), .B2(
        \xmem_data[115][5] ), .ZN(n6803) );
  AOI22_X1 U10387 ( .A1(n20585), .A2(\xmem_data[116][5] ), .B1(n31329), .B2(
        \xmem_data[117][5] ), .ZN(n6802) );
  BUF_X1 U10388 ( .A(n14971), .Z(n28302) );
  BUF_X1 U10389 ( .A(n13481), .Z(n28301) );
  AOI22_X1 U10390 ( .A1(n28302), .A2(\xmem_data[118][5] ), .B1(n28301), .B2(
        \xmem_data[119][5] ), .ZN(n6801) );
  NAND4_X1 U10391 ( .A1(n6804), .A2(n6803), .A3(n6802), .A4(n6801), .ZN(n6810)
         );
  AOI22_X1 U10392 ( .A1(n3322), .A2(\xmem_data[104][5] ), .B1(n30882), .B2(
        \xmem_data[105][5] ), .ZN(n6808) );
  BUF_X1 U10393 ( .A(n14991), .Z(n28308) );
  BUF_X1 U10394 ( .A(n13474), .Z(n28307) );
  AOI22_X1 U10395 ( .A1(n28308), .A2(\xmem_data[106][5] ), .B1(n28307), .B2(
        \xmem_data[107][5] ), .ZN(n6807) );
  AOI22_X1 U10396 ( .A1(n25707), .A2(\xmem_data[108][5] ), .B1(n25456), .B2(
        \xmem_data[109][5] ), .ZN(n6806) );
  BUF_X1 U10397 ( .A(n14997), .Z(n28309) );
  AOI22_X1 U10398 ( .A1(n28309), .A2(\xmem_data[110][5] ), .B1(n25423), .B2(
        \xmem_data[111][5] ), .ZN(n6805) );
  NAND4_X1 U10399 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6809)
         );
  OR3_X1 U10400 ( .A1(n6811), .A2(n6810), .A3(n6809), .ZN(n6820) );
  BUF_X1 U10401 ( .A(n29064), .Z(n28318) );
  AOI22_X1 U10402 ( .A1(n28318), .A2(\xmem_data[100][5] ), .B1(n3217), .B2(
        \xmem_data[101][5] ), .ZN(n6815) );
  AOI22_X1 U10403 ( .A1(n3245), .A2(\xmem_data[98][5] ), .B1(n28501), .B2(
        \xmem_data[99][5] ), .ZN(n6814) );
  AOI22_X1 U10404 ( .A1(n27564), .A2(\xmem_data[96][5] ), .B1(n28317), .B2(
        \xmem_data[97][5] ), .ZN(n6813) );
  BUF_X1 U10405 ( .A(n14989), .Z(n28319) );
  AOI22_X1 U10406 ( .A1(n25693), .A2(\xmem_data[102][5] ), .B1(n28319), .B2(
        \xmem_data[103][5] ), .ZN(n6812) );
  NAND4_X1 U10407 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6819)
         );
  INV_X1 U10408 ( .A(n6816), .ZN(n6817) );
  AOI22_X1 U10409 ( .A1(n37191), .A2(n6817), .B1(n6816), .B2(n39041), .ZN(
        n6890) );
  NAND2_X1 U10410 ( .A1(load_xaddr_val[5]), .A2(n6817), .ZN(n6818) );
  XOR2_X1 U10411 ( .A(n39040), .B(n6818), .Z(n6889) );
  AND2_X1 U10412 ( .A1(n6890), .A2(n6889), .ZN(n28288) );
  OAI21_X1 U10413 ( .B1(n6820), .B2(n6819), .A(n28288), .ZN(n6895) );
  BUF_X1 U10414 ( .A(n14882), .Z(n28327) );
  AOI22_X1 U10415 ( .A1(n27952), .A2(\xmem_data[56][5] ), .B1(n29281), .B2(
        \xmem_data[57][5] ), .ZN(n6824) );
  AOI22_X1 U10416 ( .A1(n25718), .A2(\xmem_data[58][5] ), .B1(n28098), .B2(
        \xmem_data[59][5] ), .ZN(n6823) );
  BUF_X1 U10417 ( .A(n14919), .Z(n28328) );
  AOI22_X1 U10418 ( .A1(n3179), .A2(\xmem_data[60][5] ), .B1(n28328), .B2(
        \xmem_data[61][5] ), .ZN(n6822) );
  BUF_X1 U10419 ( .A(n10456), .Z(n28329) );
  AOI22_X1 U10420 ( .A1(n30674), .A2(\xmem_data[62][5] ), .B1(n28329), .B2(
        \xmem_data[63][5] ), .ZN(n6821) );
  NAND4_X1 U10421 ( .A1(n6824), .A2(n6823), .A3(n6822), .A4(n6821), .ZN(n6835)
         );
  AOI22_X1 U10422 ( .A1(n28334), .A2(\xmem_data[48][5] ), .B1(n25709), .B2(
        \xmem_data[49][5] ), .ZN(n6828) );
  BUF_X1 U10423 ( .A(n3464), .Z(n28336) );
  BUF_X1 U10424 ( .A(n14936), .Z(n28335) );
  AOI22_X1 U10425 ( .A1(n28336), .A2(\xmem_data[50][5] ), .B1(n28335), .B2(
        \xmem_data[51][5] ), .ZN(n6827) );
  BUF_X1 U10426 ( .A(n14937), .Z(n28337) );
  AOI22_X1 U10427 ( .A1(n28337), .A2(\xmem_data[52][5] ), .B1(n27518), .B2(
        \xmem_data[53][5] ), .ZN(n6826) );
  AOI22_X1 U10428 ( .A1(n20730), .A2(\xmem_data[54][5] ), .B1(n30545), .B2(
        \xmem_data[55][5] ), .ZN(n6825) );
  NAND4_X1 U10429 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n6825), .ZN(n6834)
         );
  BUF_X1 U10430 ( .A(n14927), .Z(n28342) );
  AOI22_X1 U10431 ( .A1(n21069), .A2(\xmem_data[40][5] ), .B1(n28342), .B2(
        \xmem_data[41][5] ), .ZN(n6832) );
  BUF_X1 U10432 ( .A(n14991), .Z(n28344) );
  BUF_X1 U10433 ( .A(n14928), .Z(n28343) );
  AOI22_X1 U10434 ( .A1(n28344), .A2(\xmem_data[42][5] ), .B1(n28007), .B2(
        \xmem_data[43][5] ), .ZN(n6831) );
  AOI22_X1 U10435 ( .A1(n27910), .A2(\xmem_data[44][5] ), .B1(n30884), .B2(
        \xmem_data[45][5] ), .ZN(n6830) );
  BUF_X1 U10436 ( .A(n14997), .Z(n28346) );
  BUF_X1 U10437 ( .A(n14934), .Z(n28345) );
  AOI22_X1 U10438 ( .A1(n28346), .A2(\xmem_data[46][5] ), .B1(n28345), .B2(
        \xmem_data[47][5] ), .ZN(n6829) );
  NAND4_X1 U10439 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6833)
         );
  OR3_X1 U10440 ( .A1(n6835), .A2(n6834), .A3(n6833), .ZN(n6842) );
  BUF_X1 U10441 ( .A(n29064), .Z(n28355) );
  AND2_X1 U10442 ( .A1(n3219), .A2(\xmem_data[37][5] ), .ZN(n6836) );
  AOI21_X1 U10443 ( .B1(n28355), .B2(\xmem_data[36][5] ), .A(n6836), .ZN(n6840) );
  AOI22_X1 U10444 ( .A1(n28718), .A2(\xmem_data[34][5] ), .B1(n27501), .B2(
        \xmem_data[35][5] ), .ZN(n6839) );
  BUF_X1 U10445 ( .A(n31263), .Z(n28354) );
  AOI22_X1 U10446 ( .A1(n28354), .A2(\xmem_data[32][5] ), .B1(n21309), .B2(
        \xmem_data[33][5] ), .ZN(n6838) );
  BUF_X1 U10447 ( .A(n14989), .Z(n28356) );
  AOI22_X1 U10448 ( .A1(n25612), .A2(\xmem_data[38][5] ), .B1(n28356), .B2(
        \xmem_data[39][5] ), .ZN(n6837) );
  NAND4_X1 U10449 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6841)
         );
  INV_X1 U10450 ( .A(n6889), .ZN(n6867) );
  AND2_X1 U10451 ( .A1(n6867), .A2(n6890), .ZN(n28361) );
  OAI21_X1 U10452 ( .B1(n6842), .B2(n6841), .A(n28361), .ZN(n6894) );
  AND2_X1 U10453 ( .A1(n3217), .A2(\xmem_data[69][5] ), .ZN(n6843) );
  AOI21_X1 U10454 ( .B1(n28355), .B2(\xmem_data[68][5] ), .A(n6843), .ZN(n6850) );
  AOI22_X1 U10455 ( .A1(n28354), .A2(\xmem_data[64][5] ), .B1(n28037), .B2(
        \xmem_data[65][5] ), .ZN(n6849) );
  AOI22_X1 U10456 ( .A1(n24139), .A2(\xmem_data[70][5] ), .B1(n28356), .B2(
        \xmem_data[71][5] ), .ZN(n6844) );
  INV_X1 U10457 ( .A(n6844), .ZN(n6847) );
  AOI22_X1 U10458 ( .A1(n3424), .A2(\xmem_data[66][5] ), .B1(n28501), .B2(
        \xmem_data[67][5] ), .ZN(n6845) );
  INV_X1 U10459 ( .A(n6845), .ZN(n6846) );
  NOR2_X1 U10460 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  NAND3_X1 U10461 ( .A1(n6850), .A2(n6849), .A3(n6848), .ZN(n6866) );
  AOI22_X1 U10462 ( .A1(n28334), .A2(\xmem_data[80][5] ), .B1(n23793), .B2(
        \xmem_data[81][5] ), .ZN(n6854) );
  AOI22_X1 U10463 ( .A1(n28336), .A2(\xmem_data[82][5] ), .B1(n28335), .B2(
        \xmem_data[83][5] ), .ZN(n6853) );
  AOI22_X1 U10464 ( .A1(n28337), .A2(\xmem_data[84][5] ), .B1(n16989), .B2(
        \xmem_data[85][5] ), .ZN(n6852) );
  AOI22_X1 U10465 ( .A1(n20815), .A2(\xmem_data[86][5] ), .B1(n29049), .B2(
        \xmem_data[87][5] ), .ZN(n6851) );
  NAND4_X1 U10466 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6865)
         );
  AOI22_X1 U10467 ( .A1(n20807), .A2(\xmem_data[72][5] ), .B1(n28342), .B2(
        \xmem_data[73][5] ), .ZN(n6858) );
  AOI22_X1 U10468 ( .A1(n28344), .A2(\xmem_data[74][5] ), .B1(n30877), .B2(
        \xmem_data[75][5] ), .ZN(n6857) );
  AOI22_X1 U10469 ( .A1(n31321), .A2(\xmem_data[76][5] ), .B1(n20546), .B2(
        \xmem_data[77][5] ), .ZN(n6856) );
  AOI22_X1 U10470 ( .A1(n28346), .A2(\xmem_data[78][5] ), .B1(n28345), .B2(
        \xmem_data[79][5] ), .ZN(n6855) );
  NAND4_X1 U10471 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6864)
         );
  AOI22_X1 U10472 ( .A1(n25632), .A2(\xmem_data[88][5] ), .B1(n25581), .B2(
        \xmem_data[89][5] ), .ZN(n6862) );
  AOI22_X1 U10473 ( .A1(n20817), .A2(\xmem_data[90][5] ), .B1(n24167), .B2(
        \xmem_data[91][5] ), .ZN(n6861) );
  AOI22_X1 U10474 ( .A1(n3179), .A2(\xmem_data[92][5] ), .B1(n28328), .B2(
        \xmem_data[93][5] ), .ZN(n6860) );
  AOI22_X1 U10475 ( .A1(n21060), .A2(\xmem_data[94][5] ), .B1(n28329), .B2(
        \xmem_data[95][5] ), .ZN(n6859) );
  NAND4_X1 U10476 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6863)
         );
  OR4_X1 U10477 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6868)
         );
  NAND2_X1 U10478 ( .A1(n6868), .A2(n28324), .ZN(n6893) );
  BUF_X1 U10479 ( .A(n28974), .Z(n28366) );
  AOI22_X1 U10480 ( .A1(n27436), .A2(\xmem_data[0][5] ), .B1(n28366), .B2(
        \xmem_data[1][5] ), .ZN(n6872) );
  AOI22_X1 U10481 ( .A1(n3306), .A2(\xmem_data[2][5] ), .B1(n29253), .B2(
        \xmem_data[3][5] ), .ZN(n6871) );
  BUF_X1 U10482 ( .A(n29064), .Z(n28364) );
  AOI22_X1 U10483 ( .A1(n28364), .A2(\xmem_data[4][5] ), .B1(n3220), .B2(
        \xmem_data[5][5] ), .ZN(n6870) );
  BUF_X1 U10484 ( .A(n14988), .Z(n28367) );
  AOI22_X1 U10485 ( .A1(n28367), .A2(\xmem_data[6][5] ), .B1(n27444), .B2(
        \xmem_data[7][5] ), .ZN(n6869) );
  NAND4_X1 U10486 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6888)
         );
  BUF_X1 U10487 ( .A(n4158), .Z(n28385) );
  AOI22_X1 U10488 ( .A1(n28385), .A2(\xmem_data[24][5] ), .B1(n25581), .B2(
        \xmem_data[25][5] ), .ZN(n6876) );
  AOI22_X1 U10489 ( .A1(n3338), .A2(\xmem_data[26][5] ), .B1(n30599), .B2(
        \xmem_data[27][5] ), .ZN(n6875) );
  AOI22_X1 U10490 ( .A1(n24685), .A2(\xmem_data[28][5] ), .B1(n27981), .B2(
        \xmem_data[29][5] ), .ZN(n6874) );
  AOI22_X1 U10491 ( .A1(n23730), .A2(\xmem_data[30][5] ), .B1(n27957), .B2(
        \xmem_data[31][5] ), .ZN(n6873) );
  NAND4_X1 U10492 ( .A1(n6876), .A2(n6875), .A3(n6874), .A4(n6873), .ZN(n6887)
         );
  AOI22_X1 U10493 ( .A1(n31268), .A2(\xmem_data[16][5] ), .B1(n28090), .B2(
        \xmem_data[17][5] ), .ZN(n6880) );
  AOI22_X1 U10494 ( .A1(n24458), .A2(\xmem_data[18][5] ), .B1(n29279), .B2(
        \xmem_data[19][5] ), .ZN(n6879) );
  AOI22_X1 U10495 ( .A1(n20585), .A2(\xmem_data[20][5] ), .B1(n24459), .B2(
        \xmem_data[21][5] ), .ZN(n6878) );
  BUF_X1 U10496 ( .A(n14913), .Z(n28380) );
  AOI22_X1 U10497 ( .A1(n30872), .A2(\xmem_data[22][5] ), .B1(n28380), .B2(
        \xmem_data[23][5] ), .ZN(n6877) );
  NAND4_X1 U10498 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6886)
         );
  BUF_X1 U10499 ( .A(n14890), .Z(n28372) );
  AOI22_X1 U10500 ( .A1(n24438), .A2(\xmem_data[8][5] ), .B1(n28372), .B2(
        \xmem_data[9][5] ), .ZN(n6884) );
  AOI22_X1 U10501 ( .A1(n25417), .A2(\xmem_data[10][5] ), .B1(n3231), .B2(
        \xmem_data[11][5] ), .ZN(n6883) );
  BUF_X1 U10502 ( .A(n14933), .Z(n28373) );
  AOI22_X1 U10503 ( .A1(n28374), .A2(\xmem_data[12][5] ), .B1(n3358), .B2(
        \xmem_data[13][5] ), .ZN(n6882) );
  BUF_X1 U10504 ( .A(n13435), .Z(n28375) );
  AOI22_X1 U10505 ( .A1(n20545), .A2(\xmem_data[14][5] ), .B1(n28375), .B2(
        \xmem_data[15][5] ), .ZN(n6881) );
  NAND4_X1 U10506 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6885)
         );
  OR4_X1 U10507 ( .A1(n6888), .A2(n6887), .A3(n6886), .A4(n6885), .ZN(n6891)
         );
  NAND2_X1 U10508 ( .A1(n6891), .A2(n28395), .ZN(n6892) );
  NAND4_X1 U10509 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n32145) );
  XNOR2_X1 U10510 ( .A(n32145), .B(\fmem_data[18][5] ), .ZN(n33034) );
  XOR2_X1 U10511 ( .A(\fmem_data[18][4] ), .B(\fmem_data[18][5] ), .Z(n6896)
         );
  AOI22_X1 U10512 ( .A1(n27974), .A2(\xmem_data[56][6] ), .B1(n25679), .B2(
        \xmem_data[57][6] ), .ZN(n6900) );
  AOI22_X1 U10513 ( .A1(n28955), .A2(\xmem_data[58][6] ), .B1(n14975), .B2(
        \xmem_data[59][6] ), .ZN(n6899) );
  AOI22_X1 U10514 ( .A1(n3179), .A2(\xmem_data[60][6] ), .B1(n28328), .B2(
        \xmem_data[61][6] ), .ZN(n6898) );
  AOI22_X1 U10515 ( .A1(n21060), .A2(\xmem_data[62][6] ), .B1(n28329), .B2(
        \xmem_data[63][6] ), .ZN(n6897) );
  NAND4_X1 U10516 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6911)
         );
  AOI22_X1 U10517 ( .A1(n28334), .A2(\xmem_data[48][6] ), .B1(n29309), .B2(
        \xmem_data[49][6] ), .ZN(n6904) );
  AOI22_X1 U10518 ( .A1(n28336), .A2(\xmem_data[50][6] ), .B1(n28335), .B2(
        \xmem_data[51][6] ), .ZN(n6903) );
  AOI22_X1 U10519 ( .A1(n28337), .A2(\xmem_data[52][6] ), .B1(n29048), .B2(
        \xmem_data[53][6] ), .ZN(n6902) );
  AOI22_X1 U10520 ( .A1(n16990), .A2(\xmem_data[54][6] ), .B1(n28301), .B2(
        \xmem_data[55][6] ), .ZN(n6901) );
  NAND4_X1 U10521 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6910)
         );
  AOI22_X1 U10522 ( .A1(n24697), .A2(\xmem_data[40][6] ), .B1(n28342), .B2(
        \xmem_data[41][6] ), .ZN(n6908) );
  AOI22_X1 U10523 ( .A1(n28344), .A2(\xmem_data[42][6] ), .B1(n28007), .B2(
        \xmem_data[43][6] ), .ZN(n6907) );
  AOI22_X1 U10524 ( .A1(n25670), .A2(\xmem_data[44][6] ), .B1(n20546), .B2(
        \xmem_data[45][6] ), .ZN(n6906) );
  AOI22_X1 U10525 ( .A1(n28346), .A2(\xmem_data[46][6] ), .B1(n28345), .B2(
        \xmem_data[47][6] ), .ZN(n6905) );
  NAND4_X1 U10526 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), .ZN(n6909)
         );
  OR3_X1 U10527 ( .A1(n6911), .A2(n6910), .A3(n6909), .ZN(n6918) );
  AND2_X1 U10528 ( .A1(n3218), .A2(\xmem_data[37][6] ), .ZN(n6912) );
  AOI21_X1 U10529 ( .B1(n28355), .B2(\xmem_data[36][6] ), .A(n6912), .ZN(n6916) );
  AOI22_X1 U10530 ( .A1(n25443), .A2(\xmem_data[34][6] ), .B1(n29253), .B2(
        \xmem_data[35][6] ), .ZN(n6915) );
  AOI22_X1 U10531 ( .A1(n28354), .A2(\xmem_data[32][6] ), .B1(n28366), .B2(
        \xmem_data[33][6] ), .ZN(n6914) );
  AOI22_X1 U10532 ( .A1(n17033), .A2(\xmem_data[38][6] ), .B1(n28356), .B2(
        \xmem_data[39][6] ), .ZN(n6913) );
  NAND4_X1 U10533 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n6917)
         );
  OAI21_X1 U10534 ( .B1(n6918), .B2(n6917), .A(n28361), .ZN(n6985) );
  AOI22_X1 U10535 ( .A1(n25717), .A2(\xmem_data[88][6] ), .B1(n21009), .B2(
        \xmem_data[89][6] ), .ZN(n6922) );
  AOI22_X1 U10536 ( .A1(n30600), .A2(\xmem_data[90][6] ), .B1(n27365), .B2(
        \xmem_data[91][6] ), .ZN(n6921) );
  AOI22_X1 U10537 ( .A1(n3179), .A2(\xmem_data[92][6] ), .B1(n28328), .B2(
        \xmem_data[93][6] ), .ZN(n6920) );
  AOI22_X1 U10538 ( .A1(n24687), .A2(\xmem_data[94][6] ), .B1(n28329), .B2(
        \xmem_data[95][6] ), .ZN(n6919) );
  NAND4_X1 U10539 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n6933)
         );
  AOI22_X1 U10540 ( .A1(n28334), .A2(\xmem_data[80][6] ), .B1(n29009), .B2(
        \xmem_data[81][6] ), .ZN(n6926) );
  AOI22_X1 U10541 ( .A1(n28336), .A2(\xmem_data[82][6] ), .B1(n28335), .B2(
        \xmem_data[83][6] ), .ZN(n6925) );
  AOI22_X1 U10542 ( .A1(n28337), .A2(\xmem_data[84][6] ), .B1(n29316), .B2(
        \xmem_data[85][6] ), .ZN(n6924) );
  AOI22_X1 U10543 ( .A1(n29012), .A2(\xmem_data[86][6] ), .B1(n23776), .B2(
        \xmem_data[87][6] ), .ZN(n6923) );
  NAND4_X1 U10544 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6932)
         );
  AOI22_X1 U10545 ( .A1(n3340), .A2(\xmem_data[72][6] ), .B1(n28342), .B2(
        \xmem_data[73][6] ), .ZN(n6930) );
  AOI22_X1 U10546 ( .A1(n28344), .A2(\xmem_data[74][6] ), .B1(n25450), .B2(
        \xmem_data[75][6] ), .ZN(n6929) );
  AOI22_X1 U10547 ( .A1(n25422), .A2(\xmem_data[76][6] ), .B1(n27943), .B2(
        \xmem_data[77][6] ), .ZN(n6928) );
  AOI22_X1 U10548 ( .A1(n28346), .A2(\xmem_data[78][6] ), .B1(n28345), .B2(
        \xmem_data[79][6] ), .ZN(n6927) );
  NAND4_X1 U10549 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6931)
         );
  OR3_X1 U10550 ( .A1(n6933), .A2(n6932), .A3(n6931), .ZN(n6939) );
  AOI22_X1 U10551 ( .A1(n28355), .A2(\xmem_data[68][6] ), .B1(n3220), .B2(
        \xmem_data[69][6] ), .ZN(n6937) );
  AOI22_X1 U10552 ( .A1(n3434), .A2(\xmem_data[66][6] ), .B1(n25442), .B2(
        \xmem_data[67][6] ), .ZN(n6936) );
  AOI22_X1 U10553 ( .A1(n28354), .A2(\xmem_data[64][6] ), .B1(n25357), .B2(
        \xmem_data[65][6] ), .ZN(n6935) );
  AOI22_X1 U10554 ( .A1(n25448), .A2(\xmem_data[70][6] ), .B1(n28356), .B2(
        \xmem_data[71][6] ), .ZN(n6934) );
  NAND4_X1 U10555 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6938)
         );
  OAI21_X1 U10556 ( .B1(n6939), .B2(n6938), .A(n28324), .ZN(n6984) );
  AOI22_X1 U10557 ( .A1(n28318), .A2(\xmem_data[100][6] ), .B1(n3220), .B2(
        \xmem_data[101][6] ), .ZN(n6943) );
  AOI22_X1 U10558 ( .A1(n3424), .A2(\xmem_data[98][6] ), .B1(n22753), .B2(
        \xmem_data[99][6] ), .ZN(n6942) );
  AOI22_X1 U10559 ( .A1(n25441), .A2(\xmem_data[96][6] ), .B1(n28317), .B2(
        \xmem_data[97][6] ), .ZN(n6941) );
  AOI22_X1 U10560 ( .A1(n29256), .A2(\xmem_data[102][6] ), .B1(n28319), .B2(
        \xmem_data[103][6] ), .ZN(n6940) );
  NAND4_X1 U10561 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n6960)
         );
  AOI22_X1 U10562 ( .A1(n28428), .A2(\xmem_data[120][6] ), .B1(n28291), .B2(
        \xmem_data[121][6] ), .ZN(n6947) );
  AOI22_X1 U10563 ( .A1(n25401), .A2(\xmem_data[122][6] ), .B1(n31362), .B2(
        \xmem_data[123][6] ), .ZN(n6946) );
  AOI22_X1 U10564 ( .A1(n28293), .A2(\xmem_data[124][6] ), .B1(n28292), .B2(
        \xmem_data[125][6] ), .ZN(n6945) );
  AOI22_X1 U10565 ( .A1(n20826), .A2(\xmem_data[126][6] ), .B1(n25388), .B2(
        \xmem_data[127][6] ), .ZN(n6944) );
  NAND4_X1 U10566 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n6958)
         );
  AOI22_X1 U10567 ( .A1(n28298), .A2(\xmem_data[112][6] ), .B1(n25382), .B2(
        \xmem_data[113][6] ), .ZN(n6951) );
  AOI22_X1 U10568 ( .A1(n3120), .A2(\xmem_data[114][6] ), .B1(n28299), .B2(
        \xmem_data[115][6] ), .ZN(n6950) );
  AOI22_X1 U10569 ( .A1(n25573), .A2(\xmem_data[116][6] ), .B1(n22718), .B2(
        \xmem_data[117][6] ), .ZN(n6949) );
  AOI22_X1 U10570 ( .A1(n28302), .A2(\xmem_data[118][6] ), .B1(n28301), .B2(
        \xmem_data[119][6] ), .ZN(n6948) );
  NAND4_X1 U10571 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6957)
         );
  AOI22_X1 U10572 ( .A1(n29257), .A2(\xmem_data[104][6] ), .B1(n25616), .B2(
        \xmem_data[105][6] ), .ZN(n6955) );
  AOI22_X1 U10573 ( .A1(n28308), .A2(\xmem_data[106][6] ), .B1(n28307), .B2(
        \xmem_data[107][6] ), .ZN(n6954) );
  AOI22_X1 U10574 ( .A1(n16974), .A2(\xmem_data[108][6] ), .B1(n30884), .B2(
        \xmem_data[109][6] ), .ZN(n6953) );
  AOI22_X1 U10575 ( .A1(n28309), .A2(\xmem_data[110][6] ), .B1(n23761), .B2(
        \xmem_data[111][6] ), .ZN(n6952) );
  NAND4_X1 U10576 ( .A1(n6955), .A2(n6954), .A3(n6953), .A4(n6952), .ZN(n6956)
         );
  OR3_X1 U10577 ( .A1(n6958), .A2(n6957), .A3(n6956), .ZN(n6959) );
  OAI21_X1 U10578 ( .B1(n6960), .B2(n6959), .A(n28288), .ZN(n6983) );
  AOI22_X1 U10579 ( .A1(n30588), .A2(\xmem_data[0][6] ), .B1(n28366), .B2(
        \xmem_data[1][6] ), .ZN(n6964) );
  AOI22_X1 U10580 ( .A1(n3306), .A2(\xmem_data[2][6] ), .B1(n14875), .B2(
        \xmem_data[3][6] ), .ZN(n6963) );
  AOI22_X1 U10581 ( .A1(n28364), .A2(\xmem_data[4][6] ), .B1(n3221), .B2(
        \xmem_data[5][6] ), .ZN(n6962) );
  AOI22_X1 U10582 ( .A1(n28367), .A2(\xmem_data[6][6] ), .B1(n20787), .B2(
        \xmem_data[7][6] ), .ZN(n6961) );
  NAND4_X1 U10583 ( .A1(n6964), .A2(n6963), .A3(n6962), .A4(n6961), .ZN(n6980)
         );
  AOI22_X1 U10584 ( .A1(n28385), .A2(\xmem_data[24][6] ), .B1(n28327), .B2(
        \xmem_data[25][6] ), .ZN(n6968) );
  AOI22_X1 U10585 ( .A1(n25718), .A2(\xmem_data[26][6] ), .B1(n20983), .B2(
        \xmem_data[27][6] ), .ZN(n6967) );
  AOI22_X1 U10586 ( .A1(n24606), .A2(\xmem_data[28][6] ), .B1(n27526), .B2(
        \xmem_data[29][6] ), .ZN(n6966) );
  AOI22_X1 U10587 ( .A1(n21060), .A2(\xmem_data[30][6] ), .B1(n29248), .B2(
        \xmem_data[31][6] ), .ZN(n6965) );
  NAND4_X1 U10588 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n6979)
         );
  AOI22_X1 U10589 ( .A1(n28980), .A2(\xmem_data[16][6] ), .B1(n30613), .B2(
        \xmem_data[17][6] ), .ZN(n6972) );
  AOI22_X1 U10590 ( .A1(n30746), .A2(\xmem_data[18][6] ), .B1(n3207), .B2(
        \xmem_data[19][6] ), .ZN(n6971) );
  AOI22_X1 U10591 ( .A1(n24509), .A2(\xmem_data[20][6] ), .B1(n28492), .B2(
        \xmem_data[21][6] ), .ZN(n6970) );
  AOI22_X1 U10592 ( .A1(n27855), .A2(\xmem_data[22][6] ), .B1(n28380), .B2(
        \xmem_data[23][6] ), .ZN(n6969) );
  NAND4_X1 U10593 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n6978)
         );
  AOI22_X1 U10594 ( .A1(n22709), .A2(\xmem_data[8][6] ), .B1(n28372), .B2(
        \xmem_data[9][6] ), .ZN(n6976) );
  AOI22_X1 U10595 ( .A1(n28308), .A2(\xmem_data[10][6] ), .B1(n29306), .B2(
        \xmem_data[11][6] ), .ZN(n6975) );
  AOI22_X1 U10596 ( .A1(n28374), .A2(\xmem_data[12][6] ), .B1(n28373), .B2(
        \xmem_data[13][6] ), .ZN(n6974) );
  AOI22_X1 U10597 ( .A1(n29179), .A2(\xmem_data[14][6] ), .B1(n28375), .B2(
        \xmem_data[15][6] ), .ZN(n6973) );
  NAND4_X1 U10598 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), .ZN(n6977)
         );
  OR4_X1 U10599 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n6981)
         );
  NAND2_X1 U10600 ( .A1(n6981), .A2(n28395), .ZN(n6982) );
  NAND4_X1 U10601 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n31672) );
  XNOR2_X1 U10602 ( .A(n3356), .B(\fmem_data[18][5] ), .ZN(n31821) );
  OAI22_X1 U10603 ( .A1(n33034), .A2(n35007), .B1(n31821), .B2(n35006), .ZN(
        n33319) );
  INV_X1 U10604 ( .A(n33319), .ZN(n6986) );
  XNOR2_X1 U10605 ( .A(n33320), .B(n6986), .ZN(n33241) );
  OAI21_X1 U10606 ( .B1(n33239), .B2(n33240), .A(n33241), .ZN(n6988) );
  NAND2_X1 U10607 ( .A1(n33240), .A2(n33239), .ZN(n6987) );
  NAND2_X1 U10608 ( .A1(n6988), .A2(n6987), .ZN(n35095) );
  XNOR2_X1 U10609 ( .A(n6989), .B(n35095), .ZN(n35159) );
  OAI21_X1 U10610 ( .B1(n6992), .B2(n8418), .A(n13432), .ZN(n6993) );
  XOR2_X1 U10611 ( .A(n39040), .B(n6991), .Z(n7068) );
  INV_X1 U10612 ( .A(n7068), .ZN(n7090) );
  MUX2_X1 U10613 ( .A(load_xaddr_val[5]), .B(n39041), .S(n6993), .Z(n7091) );
  INV_X1 U10614 ( .A(n6992), .ZN(n11380) );
  NAND2_X1 U10615 ( .A1(n11380), .A2(n7216), .ZN(n11382) );
  AND2_X2 U10616 ( .A1(n11382), .A2(n6993), .ZN(n11368) );
  NAND2_X1 U10617 ( .A1(n11368), .A2(n11357), .ZN(n6994) );
  NOR2_X1 U10618 ( .A1(n11358), .A2(n6994), .ZN(n7041) );
  BUF_X1 U10619 ( .A(n7041), .Z(n30753) );
  NOR2_X1 U10620 ( .A1(n6994), .A2(n11359), .ZN(n7042) );
  BUF_X1 U10621 ( .A(n7042), .Z(n30752) );
  AOI22_X1 U10622 ( .A1(n30753), .A2(\xmem_data[32][7] ), .B1(n30752), .B2(
        \xmem_data[33][7] ), .ZN(n6998) );
  NOR2_X1 U10623 ( .A1(n6994), .A2(n3377), .ZN(n7043) );
  BUF_X1 U10624 ( .A(n7043), .Z(n30755) );
  BUF_X1 U10625 ( .A(n13127), .Z(n30754) );
  AOI22_X1 U10626 ( .A1(n30755), .A2(\xmem_data[34][7] ), .B1(n30754), .B2(
        \xmem_data[35][7] ), .ZN(n6997) );
  NOR2_X1 U10627 ( .A1(n6994), .A2(n11361), .ZN(n7044) );
  BUF_X1 U10628 ( .A(n7044), .Z(n30757) );
  NOR2_X1 U10629 ( .A1(n6994), .A2(n3246), .ZN(n7045) );
  BUF_X1 U10630 ( .A(n7045), .Z(n30756) );
  AOI22_X1 U10631 ( .A1(n30757), .A2(\xmem_data[36][7] ), .B1(n30756), .B2(
        \xmem_data[37][7] ), .ZN(n6996) );
  NOR2_X1 U10632 ( .A1(n6994), .A2(n7645), .ZN(n7046) );
  BUF_X1 U10633 ( .A(n7046), .Z(n30759) );
  BUF_X1 U10634 ( .A(n28973), .Z(n30758) );
  AOI22_X1 U10635 ( .A1(n30759), .A2(\xmem_data[38][7] ), .B1(n3144), .B2(
        \xmem_data[39][7] ), .ZN(n6995) );
  NAND4_X1 U10636 ( .A1(n6998), .A2(n6997), .A3(n6996), .A4(n6995), .ZN(n7018)
         );
  BUF_X1 U10637 ( .A(n6999), .Z(n7903) );
  BUF_X1 U10638 ( .A(n8293), .Z(n30222) );
  AOI22_X1 U10639 ( .A1(n27710), .A2(\xmem_data[40][7] ), .B1(n30222), .B2(
        \xmem_data[41][7] ), .ZN(n7004) );
  AOI22_X1 U10640 ( .A1(n27740), .A2(\xmem_data[42][7] ), .B1(n29832), .B2(
        \xmem_data[43][7] ), .ZN(n7003) );
  BUF_X1 U10641 ( .A(n11484), .Z(n30777) );
  BUF_X1 U10642 ( .A(n11780), .Z(n30776) );
  AOI22_X1 U10643 ( .A1(n30777), .A2(\xmem_data[44][7] ), .B1(n29556), .B2(
        \xmem_data[45][7] ), .ZN(n7002) );
  NAND2_X1 U10644 ( .A1(n11350), .A2(n11368), .ZN(n7000) );
  NOR2_X1 U10645 ( .A1(n7645), .A2(n7000), .ZN(n26491) );
  AOI22_X1 U10646 ( .A1(n3224), .A2(\xmem_data[46][7] ), .B1(n30698), .B2(
        \xmem_data[47][7] ), .ZN(n7001) );
  NAND4_X1 U10647 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n7017)
         );
  BUF_X2 U10648 ( .A(n11436), .Z(n30633) );
  AOI22_X1 U10649 ( .A1(n29446), .A2(\xmem_data[48][7] ), .B1(n30730), .B2(
        \xmem_data[49][7] ), .ZN(n7009) );
  INV_X1 U10650 ( .A(n11357), .ZN(n7005) );
  NOR2_X1 U10651 ( .A1(n3378), .A2(n11344), .ZN(n26543) );
  BUF_X1 U10652 ( .A(n14997), .Z(n30744) );
  AOI22_X1 U10653 ( .A1(n30664), .A2(\xmem_data[50][7] ), .B1(n30744), .B2(
        \xmem_data[51][7] ), .ZN(n7008) );
  BUF_X1 U10654 ( .A(n11439), .Z(n30635) );
  BUF_X1 U10655 ( .A(n8700), .Z(n28110) );
  AOI22_X1 U10656 ( .A1(n27754), .A2(\xmem_data[52][7] ), .B1(n28110), .B2(
        \xmem_data[53][7] ), .ZN(n7007) );
  NOR2_X1 U10657 ( .A1(n7645), .A2(n11344), .ZN(n7055) );
  BUF_X1 U10658 ( .A(n7055), .Z(n30747) );
  BUF_X1 U10659 ( .A(n29187), .Z(n30746) );
  AOI22_X1 U10660 ( .A1(n30747), .A2(\xmem_data[54][7] ), .B1(n28231), .B2(
        \xmem_data[55][7] ), .ZN(n7006) );
  NAND4_X1 U10661 ( .A1(n7009), .A2(n7008), .A3(n7007), .A4(n7006), .ZN(n7016)
         );
  AOI22_X1 U10662 ( .A1(n3165), .A2(\xmem_data[56][7] ), .B1(n3190), .B2(
        \xmem_data[57][7] ), .ZN(n7014) );
  BUF_X1 U10663 ( .A(n15549), .Z(n29810) );
  AOI22_X1 U10664 ( .A1(n29810), .A2(\xmem_data[58][7] ), .B1(n24710), .B2(
        \xmem_data[59][7] ), .ZN(n7013) );
  BUF_X2 U10665 ( .A(n18518), .Z(n29721) );
  AOI22_X1 U10666 ( .A1(n29363), .A2(\xmem_data[60][7] ), .B1(n29721), .B2(
        \xmem_data[61][7] ), .ZN(n7012) );
  INV_X1 U10667 ( .A(n11368), .ZN(n11349) );
  NOR2_X1 U10668 ( .A1(n7645), .A2(n11351), .ZN(n7077) );
  BUF_X1 U10669 ( .A(n7077), .Z(n30646) );
  BUF_X1 U10670 ( .A(n14974), .Z(n30645) );
  AOI22_X1 U10671 ( .A1(n30646), .A2(\xmem_data[62][7] ), .B1(n30645), .B2(
        \xmem_data[63][7] ), .ZN(n7011) );
  NAND4_X1 U10672 ( .A1(n7014), .A2(n7013), .A3(n7012), .A4(n7011), .ZN(n7015)
         );
  NOR2_X2 U10673 ( .A1(n7091), .A2(n7068), .ZN(n30741) );
  AOI22_X1 U10674 ( .A1(n7041), .A2(\xmem_data[0][7] ), .B1(n30672), .B2(
        \xmem_data[1][7] ), .ZN(n7022) );
  BUF_X1 U10675 ( .A(n7043), .Z(n30722) );
  AOI22_X1 U10676 ( .A1(n30722), .A2(\xmem_data[2][7] ), .B1(n20567), .B2(
        \xmem_data[3][7] ), .ZN(n7021) );
  BUF_X1 U10677 ( .A(n7044), .Z(n30724) );
  BUF_X1 U10678 ( .A(n7045), .Z(n30723) );
  AOI22_X1 U10679 ( .A1(n30724), .A2(\xmem_data[4][7] ), .B1(n30723), .B2(
        \xmem_data[5][7] ), .ZN(n7020) );
  BUF_X1 U10680 ( .A(n7046), .Z(n30725) );
  AOI22_X1 U10681 ( .A1(n30725), .A2(\xmem_data[6][7] ), .B1(n3413), .B2(
        \xmem_data[7][7] ), .ZN(n7019) );
  NAND4_X1 U10682 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n7038)
         );
  BUF_X1 U10683 ( .A(n11489), .Z(n30708) );
  AOI22_X1 U10684 ( .A1(n28136), .A2(\xmem_data[8][7] ), .B1(n30775), .B2(
        \xmem_data[9][7] ), .ZN(n7026) );
  AOI22_X1 U10685 ( .A1(n30279), .A2(\xmem_data[10][7] ), .B1(n27708), .B2(
        \xmem_data[11][7] ), .ZN(n7025) );
  BUF_X1 U10686 ( .A(n11780), .Z(n30709) );
  AOI22_X1 U10687 ( .A1(n28787), .A2(\xmem_data[12][7] ), .B1(n27833), .B2(
        \xmem_data[13][7] ), .ZN(n7024) );
  BUF_X1 U10688 ( .A(n14991), .Z(n30710) );
  AOI22_X1 U10689 ( .A1(n3224), .A2(\xmem_data[14][7] ), .B1(n30710), .B2(
        \xmem_data[15][7] ), .ZN(n7023) );
  NAND4_X1 U10690 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n7023), .ZN(n7037)
         );
  AOI22_X1 U10691 ( .A1(n30633), .A2(\xmem_data[16][7] ), .B1(n28665), .B2(
        \xmem_data[17][7] ), .ZN(n7030) );
  BUF_X1 U10692 ( .A(n26543), .Z(n30731) );
  AOI22_X1 U10693 ( .A1(n30731), .A2(\xmem_data[18][7] ), .B1(n30083), .B2(
        \xmem_data[19][7] ), .ZN(n7029) );
  AOI22_X1 U10694 ( .A1(n29436), .A2(\xmem_data[20][7] ), .B1(n27753), .B2(
        \xmem_data[21][7] ), .ZN(n7028) );
  BUF_X1 U10695 ( .A(n7055), .Z(n30732) );
  AOI22_X1 U10696 ( .A1(n30732), .A2(\xmem_data[22][7] ), .B1(n30666), .B2(
        \xmem_data[23][7] ), .ZN(n7027) );
  NAND4_X1 U10697 ( .A1(n7030), .A2(n7029), .A3(n7028), .A4(n7027), .ZN(n7036)
         );
  AOI22_X1 U10698 ( .A1(n23901), .A2(\xmem_data[26][7] ), .B1(n28147), .B2(
        \xmem_data[27][7] ), .ZN(n7034) );
  AOI22_X1 U10699 ( .A1(n29722), .A2(\xmem_data[28][7] ), .B1(n30716), .B2(
        \xmem_data[29][7] ), .ZN(n7033) );
  AOI22_X1 U10700 ( .A1(n3166), .A2(\xmem_data[24][7] ), .B1(n3185), .B2(
        \xmem_data[25][7] ), .ZN(n7032) );
  AOI22_X1 U10701 ( .A1(n30646), .A2(\xmem_data[30][7] ), .B1(n30645), .B2(
        \xmem_data[31][7] ), .ZN(n7031) );
  NAND4_X1 U10702 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7035)
         );
  OR4_X1 U10703 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .ZN(n7039)
         );
  AOI22_X1 U10704 ( .A1(n30782), .A2(n7040), .B1(n30741), .B2(n7039), .ZN(
        n7095) );
  BUF_X1 U10705 ( .A(n7041), .Z(n30673) );
  BUF_X1 U10706 ( .A(n7042), .Z(n30672) );
  AOI22_X1 U10707 ( .A1(n30673), .A2(\xmem_data[96][7] ), .B1(n30672), .B2(
        \xmem_data[97][7] ), .ZN(n7050) );
  BUF_X1 U10708 ( .A(n7043), .Z(n30675) );
  AOI22_X1 U10709 ( .A1(n30675), .A2(\xmem_data[98][7] ), .B1(n30674), .B2(
        \xmem_data[99][7] ), .ZN(n7049) );
  BUF_X1 U10710 ( .A(n7044), .Z(n30677) );
  BUF_X1 U10711 ( .A(n7045), .Z(n30676) );
  AOI22_X1 U10712 ( .A1(n30677), .A2(\xmem_data[100][7] ), .B1(n30676), .B2(
        \xmem_data[101][7] ), .ZN(n7048) );
  BUF_X1 U10713 ( .A(n7046), .Z(n30678) );
  AOI22_X1 U10714 ( .A1(n30678), .A2(\xmem_data[102][7] ), .B1(n28039), .B2(
        \xmem_data[103][7] ), .ZN(n7047) );
  NAND4_X1 U10715 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n7067)
         );
  BUF_X2 U10716 ( .A(n10861), .Z(n30182) );
  AOI22_X1 U10717 ( .A1(n30223), .A2(\xmem_data[104][7] ), .B1(n26510), .B2(
        \xmem_data[105][7] ), .ZN(n7054) );
  AOI22_X1 U10718 ( .A1(n28138), .A2(\xmem_data[106][7] ), .B1(n28218), .B2(
        \xmem_data[107][7] ), .ZN(n7053) );
  BUF_X1 U10719 ( .A(n11484), .Z(n30697) );
  BUF_X1 U10720 ( .A(n11780), .Z(n30696) );
  AOI22_X1 U10721 ( .A1(n30697), .A2(\xmem_data[108][7] ), .B1(n30217), .B2(
        \xmem_data[109][7] ), .ZN(n7052) );
  BUF_X1 U10722 ( .A(n26491), .Z(n30699) );
  AOI22_X1 U10723 ( .A1(n30699), .A2(\xmem_data[110][7] ), .B1(n30698), .B2(
        \xmem_data[111][7] ), .ZN(n7051) );
  NAND4_X1 U10724 ( .A1(n7054), .A2(n7053), .A3(n7052), .A4(n7051), .ZN(n7066)
         );
  BUF_X1 U10725 ( .A(n11437), .Z(n30662) );
  AOI22_X1 U10726 ( .A1(n29801), .A2(\xmem_data[112][7] ), .B1(n29347), .B2(
        \xmem_data[113][7] ), .ZN(n7059) );
  BUF_X1 U10727 ( .A(n14997), .Z(n30663) );
  AOI22_X1 U10728 ( .A1(n30664), .A2(\xmem_data[114][7] ), .B1(n30663), .B2(
        \xmem_data[115][7] ), .ZN(n7058) );
  BUF_X1 U10729 ( .A(n11439), .Z(n30665) );
  AOI22_X1 U10730 ( .A1(n29395), .A2(\xmem_data[116][7] ), .B1(n27753), .B2(
        \xmem_data[117][7] ), .ZN(n7057) );
  BUF_X1 U10731 ( .A(n7055), .Z(n30667) );
  BUF_X1 U10732 ( .A(n29187), .Z(n30666) );
  AOI22_X1 U10733 ( .A1(n30667), .A2(\xmem_data[118][7] ), .B1(n30543), .B2(
        \xmem_data[119][7] ), .ZN(n7056) );
  NAND4_X1 U10734 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7065)
         );
  AOI22_X1 U10735 ( .A1(n3168), .A2(\xmem_data[120][7] ), .B1(n3186), .B2(
        \xmem_data[121][7] ), .ZN(n7063) );
  AOI22_X1 U10736 ( .A1(n28689), .A2(\xmem_data[122][7] ), .B1(n17021), .B2(
        \xmem_data[123][7] ), .ZN(n7062) );
  AOI22_X1 U10737 ( .A1(n28680), .A2(\xmem_data[124][7] ), .B1(n30170), .B2(
        \xmem_data[125][7] ), .ZN(n7061) );
  BUF_X1 U10738 ( .A(n7077), .Z(n30687) );
  BUF_X1 U10739 ( .A(n14974), .Z(n30686) );
  AOI22_X1 U10740 ( .A1(n30687), .A2(\xmem_data[126][7] ), .B1(n30686), .B2(
        \xmem_data[127][7] ), .ZN(n7060) );
  NAND4_X1 U10741 ( .A1(n7063), .A2(n7062), .A3(n7061), .A4(n7060), .ZN(n7064)
         );
  AND2_X1 U10742 ( .A1(n7091), .A2(n7068), .ZN(n30659) );
  AOI22_X1 U10743 ( .A1(n27740), .A2(\xmem_data[74][7] ), .B1(n27445), .B2(
        \xmem_data[75][7] ), .ZN(n7072) );
  AOI22_X1 U10744 ( .A1(n29626), .A2(\xmem_data[72][7] ), .B1(n29697), .B2(
        \xmem_data[73][7] ), .ZN(n7071) );
  AOI22_X1 U10745 ( .A1(n30777), .A2(\xmem_data[76][7] ), .B1(n28667), .B2(
        \xmem_data[77][7] ), .ZN(n7070) );
  AOI22_X1 U10746 ( .A1(n3224), .A2(\xmem_data[78][7] ), .B1(n3147), .B2(
        \xmem_data[79][7] ), .ZN(n7069) );
  NAND4_X1 U10747 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(n7089)
         );
  BUF_X1 U10748 ( .A(n11436), .Z(n30743) );
  AOI22_X1 U10749 ( .A1(n30248), .A2(\xmem_data[80][7] ), .B1(n29704), .B2(
        \xmem_data[81][7] ), .ZN(n7076) );
  AOI22_X1 U10750 ( .A1(n30664), .A2(\xmem_data[82][7] ), .B1(n30744), .B2(
        \xmem_data[83][7] ), .ZN(n7075) );
  BUF_X1 U10751 ( .A(n11439), .Z(n30745) );
  AOI22_X1 U10752 ( .A1(n28779), .A2(\xmem_data[84][7] ), .B1(n28684), .B2(
        \xmem_data[85][7] ), .ZN(n7074) );
  AOI22_X1 U10753 ( .A1(n30747), .A2(\xmem_data[86][7] ), .B1(n28752), .B2(
        \xmem_data[87][7] ), .ZN(n7073) );
  NAND4_X1 U10754 ( .A1(n7076), .A2(n7075), .A3(n7074), .A4(n7073), .ZN(n7088)
         );
  AOI22_X1 U10755 ( .A1(n3167), .A2(\xmem_data[88][7] ), .B1(n3186), .B2(
        \xmem_data[89][7] ), .ZN(n7081) );
  AOI22_X1 U10756 ( .A1(n28689), .A2(\xmem_data[90][7] ), .B1(n29439), .B2(
        \xmem_data[91][7] ), .ZN(n7080) );
  BUF_X1 U10757 ( .A(n10802), .Z(n29363) );
  BUF_X2 U10758 ( .A(n18518), .Z(n29487) );
  AOI22_X1 U10759 ( .A1(n29815), .A2(\xmem_data[92][7] ), .B1(n29487), .B2(
        \xmem_data[93][7] ), .ZN(n7079) );
  BUF_X1 U10760 ( .A(n7077), .Z(n30767) );
  AOI22_X1 U10761 ( .A1(n30767), .A2(\xmem_data[94][7] ), .B1(n28701), .B2(
        \xmem_data[95][7] ), .ZN(n7078) );
  NAND4_X1 U10762 ( .A1(n7081), .A2(n7080), .A3(n7079), .A4(n7078), .ZN(n7087)
         );
  AOI22_X1 U10763 ( .A1(n30753), .A2(\xmem_data[64][7] ), .B1(n30752), .B2(
        \xmem_data[65][7] ), .ZN(n7085) );
  AOI22_X1 U10764 ( .A1(n30755), .A2(\xmem_data[66][7] ), .B1(n30754), .B2(
        \xmem_data[67][7] ), .ZN(n7084) );
  AOI22_X1 U10765 ( .A1(n30757), .A2(\xmem_data[68][7] ), .B1(n30756), .B2(
        \xmem_data[69][7] ), .ZN(n7083) );
  AOI22_X1 U10766 ( .A1(n30759), .A2(\xmem_data[70][7] ), .B1(n3144), .B2(
        \xmem_data[71][7] ), .ZN(n7082) );
  NAND4_X1 U10767 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n7086)
         );
  OR4_X1 U10768 ( .A1(n7089), .A2(n7088), .A3(n7087), .A4(n7086), .ZN(n7092)
         );
  AOI22_X1 U10769 ( .A1(n7093), .A2(n30659), .B1(n7092), .B2(n30704), .ZN(
        n7094) );
  NAND2_X1 U10770 ( .A1(n7095), .A2(n7094), .ZN(n35258) );
  XNOR2_X1 U10771 ( .A(n3462), .B(\fmem_data[23][3] ), .ZN(n30464) );
  AOI22_X1 U10772 ( .A1(n30291), .A2(\xmem_data[40][6] ), .B1(n29432), .B2(
        \xmem_data[41][6] ), .ZN(n7099) );
  AOI22_X1 U10773 ( .A1(n29628), .A2(\xmem_data[42][6] ), .B1(n30292), .B2(
        \xmem_data[43][6] ), .ZN(n7098) );
  AOI22_X1 U10774 ( .A1(n30777), .A2(\xmem_data[44][6] ), .B1(n28667), .B2(
        \xmem_data[45][6] ), .ZN(n7097) );
  AOI22_X1 U10775 ( .A1(n3224), .A2(\xmem_data[46][6] ), .B1(n3134), .B2(
        \xmem_data[47][6] ), .ZN(n7096) );
  NAND4_X1 U10776 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7100)
         );
  AOI22_X1 U10777 ( .A1(n29788), .A2(\xmem_data[104][6] ), .B1(n30100), .B2(
        \xmem_data[105][6] ), .ZN(n7104) );
  AOI22_X1 U10778 ( .A1(n3392), .A2(\xmem_data[106][6] ), .B1(n24696), .B2(
        \xmem_data[107][6] ), .ZN(n7103) );
  AOI22_X1 U10779 ( .A1(n30697), .A2(\xmem_data[108][6] ), .B1(n29495), .B2(
        \xmem_data[109][6] ), .ZN(n7102) );
  AOI22_X1 U10780 ( .A1(n30699), .A2(\xmem_data[110][6] ), .B1(n30698), .B2(
        \xmem_data[111][6] ), .ZN(n7101) );
  NAND4_X1 U10781 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), .ZN(n7105)
         );
  NAND2_X1 U10782 ( .A1(n7105), .A2(n30659), .ZN(n7106) );
  AOI22_X1 U10783 ( .A1(n29790), .A2(\xmem_data[74][6] ), .B1(n29832), .B2(
        \xmem_data[75][6] ), .ZN(n7111) );
  AOI22_X1 U10784 ( .A1(n30777), .A2(\xmem_data[76][6] ), .B1(n27833), .B2(
        \xmem_data[77][6] ), .ZN(n7110) );
  BUF_X2 U10785 ( .A(n7903), .Z(n29831) );
  AOI22_X1 U10786 ( .A1(n30223), .A2(\xmem_data[72][6] ), .B1(n29831), .B2(
        \xmem_data[73][6] ), .ZN(n7109) );
  AOI22_X1 U10787 ( .A1(n3224), .A2(\xmem_data[78][6] ), .B1(n30698), .B2(
        \xmem_data[79][6] ), .ZN(n7108) );
  NAND4_X1 U10788 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7112)
         );
  AOI22_X1 U10789 ( .A1(n30633), .A2(\xmem_data[16][6] ), .B1(n28738), .B2(
        \xmem_data[17][6] ), .ZN(n7116) );
  AOI22_X1 U10790 ( .A1(n30731), .A2(\xmem_data[18][6] ), .B1(n30663), .B2(
        \xmem_data[19][6] ), .ZN(n7115) );
  BUF_X1 U10791 ( .A(n8700), .Z(n29768) );
  AOI22_X1 U10792 ( .A1(n30665), .A2(\xmem_data[20][6] ), .B1(n29592), .B2(
        \xmem_data[21][6] ), .ZN(n7114) );
  AOI22_X1 U10793 ( .A1(n30732), .A2(\xmem_data[22][6] ), .B1(n28154), .B2(
        \xmem_data[23][6] ), .ZN(n7113) );
  NAND4_X1 U10794 ( .A1(n7116), .A2(n7115), .A3(n7114), .A4(n7113), .ZN(n7122)
         );
  AOI22_X1 U10795 ( .A1(n28689), .A2(\xmem_data[90][6] ), .B1(n22682), .B2(
        \xmem_data[91][6] ), .ZN(n7120) );
  AOI22_X1 U10796 ( .A1(n3161), .A2(\xmem_data[88][6] ), .B1(n3190), .B2(
        \xmem_data[89][6] ), .ZN(n7119) );
  AOI22_X1 U10797 ( .A1(n30198), .A2(\xmem_data[92][6] ), .B1(n30716), .B2(
        \xmem_data[93][6] ), .ZN(n7118) );
  AOI22_X1 U10798 ( .A1(n30767), .A2(\xmem_data[94][6] ), .B1(n3329), .B2(
        \xmem_data[95][6] ), .ZN(n7117) );
  NAND4_X1 U10799 ( .A1(n7120), .A2(n7119), .A3(n7118), .A4(n7117), .ZN(n7121)
         );
  AOI22_X1 U10800 ( .A1(n30741), .A2(n7122), .B1(n7121), .B2(n30704), .ZN(
        n7129) );
  BUF_X1 U10801 ( .A(n15549), .Z(n30764) );
  AOI22_X1 U10802 ( .A1(n30764), .A2(\xmem_data[122][6] ), .B1(n21050), .B2(
        \xmem_data[123][6] ), .ZN(n7126) );
  AOI22_X1 U10803 ( .A1(n3162), .A2(\xmem_data[120][6] ), .B1(n3188), .B2(
        \xmem_data[121][6] ), .ZN(n7125) );
  AOI22_X1 U10804 ( .A1(n30063), .A2(\xmem_data[124][6] ), .B1(n29640), .B2(
        \xmem_data[125][6] ), .ZN(n7124) );
  AOI22_X1 U10805 ( .A1(n30646), .A2(\xmem_data[126][6] ), .B1(n30686), .B2(
        \xmem_data[127][6] ), .ZN(n7123) );
  NAND4_X1 U10806 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .ZN(n7127)
         );
  NAND3_X1 U10807 ( .A1(n7130), .A2(n7129), .A3(n7128), .ZN(n7191) );
  AOI22_X1 U10808 ( .A1(n29390), .A2(\xmem_data[112][6] ), .B1(n29482), .B2(
        \xmem_data[113][6] ), .ZN(n7134) );
  AOI22_X1 U10809 ( .A1(n30664), .A2(\xmem_data[114][6] ), .B1(n30663), .B2(
        \xmem_data[115][6] ), .ZN(n7133) );
  AOI22_X1 U10810 ( .A1(n30635), .A2(\xmem_data[116][6] ), .B1(n30193), .B2(
        \xmem_data[117][6] ), .ZN(n7132) );
  AOI22_X1 U10811 ( .A1(n30667), .A2(\xmem_data[118][6] ), .B1(n20718), .B2(
        \xmem_data[119][6] ), .ZN(n7131) );
  NAND4_X1 U10812 ( .A1(n7134), .A2(n7133), .A3(n7132), .A4(n7131), .ZN(n7135)
         );
  AOI22_X1 U10813 ( .A1(n30753), .A2(\xmem_data[64][6] ), .B1(n30752), .B2(
        \xmem_data[65][6] ), .ZN(n7139) );
  AOI22_X1 U10814 ( .A1(n30755), .A2(\xmem_data[66][6] ), .B1(n30754), .B2(
        \xmem_data[67][6] ), .ZN(n7138) );
  AOI22_X1 U10815 ( .A1(n30757), .A2(\xmem_data[68][6] ), .B1(n30756), .B2(
        \xmem_data[69][6] ), .ZN(n7137) );
  AOI22_X1 U10816 ( .A1(n30759), .A2(\xmem_data[70][6] ), .B1(n3144), .B2(
        \xmem_data[71][6] ), .ZN(n7136) );
  NAND4_X1 U10817 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n7145)
         );
  AOI22_X1 U10818 ( .A1(n7041), .A2(\xmem_data[0][6] ), .B1(n7042), .B2(
        \xmem_data[1][6] ), .ZN(n7143) );
  AOI22_X1 U10819 ( .A1(n30722), .A2(\xmem_data[2][6] ), .B1(n20985), .B2(
        \xmem_data[3][6] ), .ZN(n7142) );
  AOI22_X1 U10820 ( .A1(n30724), .A2(\xmem_data[4][6] ), .B1(n30723), .B2(
        \xmem_data[5][6] ), .ZN(n7141) );
  AOI22_X1 U10821 ( .A1(n30725), .A2(\xmem_data[6][6] ), .B1(n3413), .B2(
        \xmem_data[7][6] ), .ZN(n7140) );
  NAND4_X1 U10822 ( .A1(n7143), .A2(n7142), .A3(n7141), .A4(n7140), .ZN(n7144)
         );
  AOI22_X1 U10823 ( .A1(n7145), .A2(n30704), .B1(n30741), .B2(n7144), .ZN(
        n7163) );
  AOI22_X1 U10824 ( .A1(n30753), .A2(\xmem_data[32][6] ), .B1(n30752), .B2(
        \xmem_data[33][6] ), .ZN(n7149) );
  AOI22_X1 U10825 ( .A1(n30755), .A2(\xmem_data[34][6] ), .B1(n30754), .B2(
        \xmem_data[35][6] ), .ZN(n7148) );
  AOI22_X1 U10826 ( .A1(n30757), .A2(\xmem_data[36][6] ), .B1(n30756), .B2(
        \xmem_data[37][6] ), .ZN(n7147) );
  AOI22_X1 U10827 ( .A1(n30759), .A2(\xmem_data[38][6] ), .B1(n3144), .B2(
        \xmem_data[39][6] ), .ZN(n7146) );
  NAND4_X1 U10828 ( .A1(n7149), .A2(n7148), .A3(n7147), .A4(n7146), .ZN(n7155)
         );
  AOI22_X1 U10829 ( .A1(n30673), .A2(\xmem_data[96][6] ), .B1(n30672), .B2(
        \xmem_data[97][6] ), .ZN(n7153) );
  AOI22_X1 U10830 ( .A1(n30675), .A2(\xmem_data[98][6] ), .B1(n30674), .B2(
        \xmem_data[99][6] ), .ZN(n7152) );
  AOI22_X1 U10831 ( .A1(n30677), .A2(\xmem_data[100][6] ), .B1(n30676), .B2(
        \xmem_data[101][6] ), .ZN(n7151) );
  AOI22_X1 U10832 ( .A1(n30678), .A2(\xmem_data[102][6] ), .B1(n3149), .B2(
        \xmem_data[103][6] ), .ZN(n7150) );
  NAND4_X1 U10833 ( .A1(n7153), .A2(n7152), .A3(n7151), .A4(n7150), .ZN(n7154)
         );
  AOI22_X1 U10834 ( .A1(n3168), .A2(\xmem_data[56][6] ), .B1(n3189), .B2(
        \xmem_data[57][6] ), .ZN(n7159) );
  AOI22_X1 U10835 ( .A1(n29476), .A2(\xmem_data[58][6] ), .B1(n28754), .B2(
        \xmem_data[59][6] ), .ZN(n7158) );
  AOI22_X1 U10836 ( .A1(n28680), .A2(\xmem_data[60][6] ), .B1(n30685), .B2(
        \xmem_data[61][6] ), .ZN(n7157) );
  AOI22_X1 U10837 ( .A1(n30767), .A2(\xmem_data[62][6] ), .B1(n30645), .B2(
        \xmem_data[63][6] ), .ZN(n7156) );
  NAND4_X1 U10838 ( .A1(n7158), .A2(n7157), .A3(n7159), .A4(n7156), .ZN(n7160)
         );
  AOI22_X1 U10839 ( .A1(n29433), .A2(\xmem_data[8][6] ), .B1(n30654), .B2(
        \xmem_data[9][6] ), .ZN(n7168) );
  AOI22_X1 U10840 ( .A1(n30279), .A2(\xmem_data[10][6] ), .B1(n30278), .B2(
        \xmem_data[11][6] ), .ZN(n7167) );
  AOI22_X1 U10841 ( .A1(n29674), .A2(\xmem_data[12][6] ), .B1(n29556), .B2(
        \xmem_data[13][6] ), .ZN(n7166) );
  AOI22_X1 U10842 ( .A1(n3224), .A2(\xmem_data[14][6] ), .B1(n30710), .B2(
        \xmem_data[15][6] ), .ZN(n7165) );
  NAND4_X1 U10843 ( .A1(n7168), .A2(n7167), .A3(n7166), .A4(n7165), .ZN(n7169)
         );
  NAND2_X1 U10844 ( .A1(n7169), .A2(n30741), .ZN(n7188) );
  AOI22_X1 U10845 ( .A1(n29390), .A2(\xmem_data[48][6] ), .B1(n27761), .B2(
        \xmem_data[49][6] ), .ZN(n7173) );
  AOI22_X1 U10846 ( .A1(n30664), .A2(\xmem_data[50][6] ), .B1(n30744), .B2(
        \xmem_data[51][6] ), .ZN(n7172) );
  AOI22_X1 U10847 ( .A1(n27811), .A2(\xmem_data[52][6] ), .B1(n27728), .B2(
        \xmem_data[53][6] ), .ZN(n7171) );
  AOI22_X1 U10848 ( .A1(n30747), .A2(\xmem_data[54][6] ), .B1(n27818), .B2(
        \xmem_data[55][6] ), .ZN(n7170) );
  NAND4_X1 U10849 ( .A1(n7173), .A2(n7172), .A3(n7171), .A4(n7170), .ZN(n7174)
         );
  AOI22_X1 U10850 ( .A1(n29647), .A2(\xmem_data[80][6] ), .B1(n29646), .B2(
        \xmem_data[81][6] ), .ZN(n7178) );
  AOI22_X1 U10851 ( .A1(n30664), .A2(\xmem_data[82][6] ), .B1(n30744), .B2(
        \xmem_data[83][6] ), .ZN(n7177) );
  AOI22_X1 U10852 ( .A1(n29436), .A2(\xmem_data[84][6] ), .B1(n30193), .B2(
        \xmem_data[85][6] ), .ZN(n7176) );
  AOI22_X1 U10853 ( .A1(n30747), .A2(\xmem_data[86][6] ), .B1(n20776), .B2(
        \xmem_data[87][6] ), .ZN(n7175) );
  NAND4_X1 U10854 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .ZN(n7179)
         );
  AOI22_X1 U10855 ( .A1(n3166), .A2(\xmem_data[24][6] ), .B1(n11426), .B2(
        \xmem_data[25][6] ), .ZN(n7183) );
  BUF_X1 U10856 ( .A(n15549), .Z(n29716) );
  AOI22_X1 U10857 ( .A1(n29716), .A2(\xmem_data[26][6] ), .B1(n29410), .B2(
        \xmem_data[27][6] ), .ZN(n7182) );
  AOI22_X1 U10858 ( .A1(n30766), .A2(\xmem_data[28][6] ), .B1(n29721), .B2(
        \xmem_data[29][6] ), .ZN(n7181) );
  AOI22_X1 U10859 ( .A1(n30646), .A2(\xmem_data[30][6] ), .B1(n30645), .B2(
        \xmem_data[31][6] ), .ZN(n7180) );
  NAND4_X1 U10860 ( .A1(n7183), .A2(n7182), .A3(n7181), .A4(n7180), .ZN(n7184)
         );
  NAND2_X1 U10861 ( .A1(n7184), .A2(n30741), .ZN(n7185) );
  NAND4_X1 U10862 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), .ZN(n7189)
         );
  OR4_X2 U10863 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n35114)
         );
  XNOR2_X1 U10864 ( .A(n35114), .B(\fmem_data[23][3] ), .ZN(n28266) );
  XOR2_X1 U10865 ( .A(\fmem_data[23][2] ), .B(\fmem_data[23][3] ), .Z(n7193)
         );
  OAI22_X1 U10866 ( .A1(n30464), .A2(n34412), .B1(n28266), .B2(n34410), .ZN(
        n34270) );
  BUF_X1 U10867 ( .A(n11439), .Z(n29395) );
  BUF_X1 U10868 ( .A(n8700), .Z(n29592) );
  AOI22_X1 U10869 ( .A1(n30250), .A2(\xmem_data[96][5] ), .B1(n29768), .B2(
        \xmem_data[97][5] ), .ZN(n7197) );
  NAND3_X1 U10870 ( .A1(n11343), .A2(n11342), .A3(n6173), .ZN(n7206) );
  NOR2_X1 U10871 ( .A1(n8000), .A2(n7206), .ZN(n29475) );
  BUF_X1 U10872 ( .A(n29187), .Z(n29396) );
  AOI22_X1 U10873 ( .A1(n29397), .A2(\xmem_data[98][5] ), .B1(n29605), .B2(
        \xmem_data[99][5] ), .ZN(n7196) );
  AOI22_X1 U10874 ( .A1(n3167), .A2(\xmem_data[100][5] ), .B1(n3188), .B2(
        \xmem_data[101][5] ), .ZN(n7195) );
  BUF_X1 U10875 ( .A(n14971), .Z(n29410) );
  AOI22_X1 U10876 ( .A1(n28689), .A2(\xmem_data[102][5] ), .B1(n29410), .B2(
        \xmem_data[103][5] ), .ZN(n7194) );
  NAND4_X1 U10877 ( .A1(n7197), .A2(n7196), .A3(n7195), .A4(n7194), .ZN(n7214)
         );
  AOI22_X1 U10878 ( .A1(n30063), .A2(\xmem_data[104][5] ), .B1(n30266), .B2(
        \xmem_data[105][5] ), .ZN(n7201) );
  NOR2_X2 U10879 ( .A1(n7010), .A2(n8005), .ZN(n7270) );
  BUF_X1 U10880 ( .A(n7270), .Z(n29380) );
  BUF_X1 U10881 ( .A(n14974), .Z(n29379) );
  AOI22_X1 U10882 ( .A1(n29380), .A2(\xmem_data[106][5] ), .B1(n29379), .B2(
        \xmem_data[107][5] ), .ZN(n7200) );
  BUF_X1 U10883 ( .A(n8073), .Z(n29382) );
  BUF_X1 U10884 ( .A(n8074), .Z(n29381) );
  AOI22_X1 U10885 ( .A1(n29382), .A2(\xmem_data[108][5] ), .B1(n29381), .B2(
        \xmem_data[109][5] ), .ZN(n7199) );
  NOR2_X1 U10886 ( .A1(n11360), .A2(n8005), .ZN(n8075) );
  BUF_X1 U10887 ( .A(n8075), .Z(n29384) );
  BUF_X1 U10888 ( .A(n13127), .Z(n29383) );
  AOI22_X1 U10889 ( .A1(n29384), .A2(\xmem_data[110][5] ), .B1(n29383), .B2(
        \xmem_data[111][5] ), .ZN(n7198) );
  NAND4_X1 U10890 ( .A1(n7201), .A2(n7200), .A3(n7199), .A4(n7198), .ZN(n7213)
         );
  NOR2_X1 U10891 ( .A1(n11361), .A2(n8010), .ZN(n7275) );
  AOI22_X1 U10892 ( .A1(n29419), .A2(\xmem_data[112][5] ), .B1(n29418), .B2(
        \xmem_data[113][5] ), .ZN(n7205) );
  NOR2_X1 U10893 ( .A1(n7206), .A2(n8010), .ZN(n7276) );
  BUF_X1 U10894 ( .A(n7276), .Z(n29420) );
  AOI22_X1 U10895 ( .A1(n29420), .A2(\xmem_data[114][5] ), .B1(n23732), .B2(
        \xmem_data[115][5] ), .ZN(n7204) );
  BUF_X2 U10896 ( .A(n11489), .Z(n29421) );
  BUF_X2 U10897 ( .A(n10861), .Z(n30290) );
  AOI22_X1 U10898 ( .A1(n30291), .A2(\xmem_data[116][5] ), .B1(n30290), .B2(
        \xmem_data[117][5] ), .ZN(n7203) );
  BUF_X1 U10899 ( .A(n11451), .Z(n29423) );
  BUF_X1 U10900 ( .A(n14988), .Z(n29422) );
  AOI22_X1 U10901 ( .A1(n29790), .A2(\xmem_data[118][5] ), .B1(n29422), .B2(
        \xmem_data[119][5] ), .ZN(n7202) );
  NAND4_X1 U10902 ( .A1(n7205), .A2(n7204), .A3(n7203), .A4(n7202), .ZN(n7212)
         );
  BUF_X1 U10903 ( .A(n11484), .Z(n29400) );
  AOI22_X1 U10904 ( .A1(n29400), .A2(\xmem_data[120][5] ), .B1(n29708), .B2(
        \xmem_data[121][5] ), .ZN(n7210) );
  NOR2_X1 U10905 ( .A1(n7206), .A2(n3447), .ZN(n7281) );
  BUF_X1 U10906 ( .A(n7281), .Z(n29402) );
  BUF_X1 U10907 ( .A(n14991), .Z(n29401) );
  AOI22_X1 U10908 ( .A1(n29402), .A2(\xmem_data[122][5] ), .B1(n3135), .B2(
        \xmem_data[123][5] ), .ZN(n7209) );
  BUF_X1 U10909 ( .A(n11436), .Z(n29390) );
  BUF_X1 U10910 ( .A(n11437), .Z(n29347) );
  AOI22_X1 U10911 ( .A1(n28180), .A2(\xmem_data[124][5] ), .B1(n29589), .B2(
        \xmem_data[125][5] ), .ZN(n7208) );
  NOR2_X1 U10912 ( .A1(n11360), .A2(n3445), .ZN(n7282) );
  BUF_X1 U10913 ( .A(n14997), .Z(n29403) );
  AOI22_X1 U10914 ( .A1(n29404), .A2(\xmem_data[126][5] ), .B1(n29403), .B2(
        \xmem_data[127][5] ), .ZN(n7207) );
  NAND4_X1 U10915 ( .A1(n7210), .A2(n7209), .A3(n7208), .A4(n7207), .ZN(n7211)
         );
  OR4_X1 U10916 ( .A1(n7214), .A2(n7213), .A3(n7212), .A4(n7211), .ZN(n7220)
         );
  NAND2_X1 U10917 ( .A1(n7423), .A2(n7216), .ZN(n7217) );
  AOI22_X1 U10918 ( .A1(n10973), .A2(n7423), .B1(n4499), .B2(n7217), .ZN(n7292) );
  INV_X1 U10919 ( .A(n7423), .ZN(n7218) );
  NOR2_X1 U10920 ( .A1(n11381), .A2(n7218), .ZN(n7219) );
  XOR2_X1 U10921 ( .A(n7219), .B(load_xaddr_val[6]), .Z(n7291) );
  AND2_X1 U10922 ( .A1(n7292), .A2(n7291), .ZN(n29428) );
  NAND2_X1 U10923 ( .A1(n7220), .A2(n29428), .ZN(n7297) );
  BUF_X1 U10924 ( .A(n11439), .Z(n29436) );
  AOI22_X1 U10925 ( .A1(n28685), .A2(\xmem_data[64][5] ), .B1(n28778), .B2(
        \xmem_data[65][5] ), .ZN(n7224) );
  BUF_X1 U10926 ( .A(n29187), .Z(n29437) );
  AOI22_X1 U10927 ( .A1(n29438), .A2(\xmem_data[66][5] ), .B1(n31354), .B2(
        \xmem_data[67][5] ), .ZN(n7223) );
  AOI22_X1 U10928 ( .A1(n3166), .A2(\xmem_data[68][5] ), .B1(n3183), .B2(
        \xmem_data[69][5] ), .ZN(n7222) );
  BUF_X1 U10929 ( .A(n14971), .Z(n29439) );
  AOI22_X1 U10930 ( .A1(n30062), .A2(\xmem_data[70][5] ), .B1(n29439), .B2(
        \xmem_data[71][5] ), .ZN(n7221) );
  AOI22_X1 U10931 ( .A1(n30766), .A2(\xmem_data[72][5] ), .B1(n29640), .B2(
        \xmem_data[73][5] ), .ZN(n7228) );
  BUF_X1 U10932 ( .A(n7270), .Z(n29461) );
  BUF_X1 U10933 ( .A(n14974), .Z(n29460) );
  AOI22_X1 U10934 ( .A1(n29461), .A2(\xmem_data[74][5] ), .B1(n3151), .B2(
        \xmem_data[75][5] ), .ZN(n7227) );
  BUF_X1 U10935 ( .A(n8073), .Z(n29463) );
  AOI22_X1 U10936 ( .A1(n29463), .A2(\xmem_data[76][5] ), .B1(n29462), .B2(
        \xmem_data[77][5] ), .ZN(n7226) );
  BUF_X1 U10937 ( .A(n8075), .Z(n29464) );
  AOI22_X1 U10938 ( .A1(n29464), .A2(\xmem_data[78][5] ), .B1(n28772), .B2(
        \xmem_data[79][5] ), .ZN(n7225) );
  NAND4_X1 U10939 ( .A1(n7228), .A2(n7227), .A3(n7226), .A4(n7225), .ZN(n7232)
         );
  BUF_X1 U10940 ( .A(n11436), .Z(n29446) );
  AOI22_X1 U10941 ( .A1(n28180), .A2(\xmem_data[92][5] ), .B1(n28738), .B2(
        \xmem_data[93][5] ), .ZN(n7230) );
  AOI22_X1 U10942 ( .A1(n3170), .A2(\xmem_data[89][5] ), .B1(n30777), .B2(
        \xmem_data[88][5] ), .ZN(n7229) );
  NAND2_X1 U10943 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  NOR2_X1 U10944 ( .A1(n7232), .A2(n7231), .ZN(n7242) );
  BUF_X2 U10945 ( .A(n10861), .Z(n29432) );
  AOI22_X1 U10946 ( .A1(n28734), .A2(\xmem_data[84][5] ), .B1(n30100), .B2(
        \xmem_data[85][5] ), .ZN(n7241) );
  BUF_X1 U10947 ( .A(n14988), .Z(n29431) );
  AOI22_X1 U10948 ( .A1(n30215), .A2(\xmem_data[86][5] ), .B1(n29431), .B2(
        \xmem_data[87][5] ), .ZN(n7233) );
  INV_X1 U10949 ( .A(n7233), .ZN(n7239) );
  BUF_X1 U10950 ( .A(n7276), .Z(n29449) );
  AOI22_X1 U10951 ( .A1(n29449), .A2(\xmem_data[82][5] ), .B1(n29661), .B2(
        \xmem_data[83][5] ), .ZN(n7237) );
  BUF_X1 U10952 ( .A(n7281), .Z(n29450) );
  BUF_X1 U10953 ( .A(n14991), .Z(n29350) );
  AOI22_X1 U10954 ( .A1(n29450), .A2(\xmem_data[90][5] ), .B1(n29350), .B2(
        \xmem_data[91][5] ), .ZN(n7236) );
  BUF_X1 U10955 ( .A(n7275), .Z(n29447) );
  AOI22_X1 U10956 ( .A1(n29447), .A2(\xmem_data[80][5] ), .B1(n27812), .B2(
        \xmem_data[81][5] ), .ZN(n7235) );
  BUF_X1 U10957 ( .A(n14997), .Z(n29451) );
  AOI22_X1 U10958 ( .A1(n29802), .A2(\xmem_data[94][5] ), .B1(n29451), .B2(
        \xmem_data[95][5] ), .ZN(n7234) );
  NAND4_X1 U10959 ( .A1(n7237), .A2(n7236), .A3(n7235), .A4(n7234), .ZN(n7238)
         );
  NOR2_X1 U10960 ( .A1(n7239), .A2(n7238), .ZN(n7240) );
  NAND4_X1 U10961 ( .A1(n3833), .A2(n7242), .A3(n7241), .A4(n7240), .ZN(n7243)
         );
  INV_X1 U10962 ( .A(n7291), .ZN(n7264) );
  NOR2_X1 U10963 ( .A1(n7292), .A2(n7264), .ZN(n29376) );
  NAND2_X1 U10964 ( .A1(n7243), .A2(n29376), .ZN(n7296) );
  BUF_X1 U10965 ( .A(n8700), .Z(n30634) );
  AOI22_X1 U10966 ( .A1(n30635), .A2(\xmem_data[32][5] ), .B1(n28684), .B2(
        \xmem_data[33][5] ), .ZN(n7247) );
  AOI22_X1 U10967 ( .A1(n29438), .A2(\xmem_data[34][5] ), .B1(n27818), .B2(
        \xmem_data[35][5] ), .ZN(n7246) );
  AOI22_X1 U10968 ( .A1(n3162), .A2(\xmem_data[36][5] ), .B1(n3186), .B2(
        \xmem_data[37][5] ), .ZN(n7245) );
  AOI22_X1 U10969 ( .A1(n29810), .A2(\xmem_data[38][5] ), .B1(n29439), .B2(
        \xmem_data[39][5] ), .ZN(n7244) );
  NAND4_X1 U10970 ( .A1(n7247), .A2(n7246), .A3(n7245), .A4(n7244), .ZN(n7263)
         );
  AOI22_X1 U10971 ( .A1(n30717), .A2(\xmem_data[40][5] ), .B1(n30765), .B2(
        \xmem_data[41][5] ), .ZN(n7251) );
  AOI22_X1 U10972 ( .A1(n29461), .A2(\xmem_data[42][5] ), .B1(n3151), .B2(
        \xmem_data[43][5] ), .ZN(n7250) );
  AOI22_X1 U10973 ( .A1(n29463), .A2(\xmem_data[44][5] ), .B1(n29462), .B2(
        \xmem_data[45][5] ), .ZN(n7249) );
  AOI22_X1 U10974 ( .A1(n29464), .A2(\xmem_data[46][5] ), .B1(n20567), .B2(
        \xmem_data[47][5] ), .ZN(n7248) );
  NAND4_X1 U10975 ( .A1(n7251), .A2(n7250), .A3(n7249), .A4(n7248), .ZN(n7262)
         );
  AOI22_X1 U10976 ( .A1(n29447), .A2(\xmem_data[48][5] ), .B1(n27743), .B2(
        \xmem_data[49][5] ), .ZN(n7255) );
  AOI22_X1 U10977 ( .A1(n29449), .A2(\xmem_data[50][5] ), .B1(n3333), .B2(
        \xmem_data[51][5] ), .ZN(n7254) );
  AOI22_X1 U10978 ( .A1(n28734), .A2(\xmem_data[52][5] ), .B1(n30654), .B2(
        \xmem_data[53][5] ), .ZN(n7253) );
  AOI22_X1 U10979 ( .A1(n3392), .A2(\xmem_data[54][5] ), .B1(n29431), .B2(
        \xmem_data[55][5] ), .ZN(n7252) );
  NAND4_X1 U10980 ( .A1(n7255), .A2(n7254), .A3(n7253), .A4(n7252), .ZN(n7261)
         );
  AOI22_X1 U10981 ( .A1(n30280), .A2(\xmem_data[56][5] ), .B1(n30293), .B2(
        \xmem_data[57][5] ), .ZN(n7259) );
  AOI22_X1 U10982 ( .A1(n29450), .A2(\xmem_data[58][5] ), .B1(n30295), .B2(
        \xmem_data[59][5] ), .ZN(n7258) );
  BUF_X1 U10983 ( .A(n11437), .Z(n29389) );
  AOI22_X1 U10984 ( .A1(n29602), .A2(\xmem_data[60][5] ), .B1(n27761), .B2(
        \xmem_data[61][5] ), .ZN(n7257) );
  AOI22_X1 U10985 ( .A1(n29802), .A2(\xmem_data[62][5] ), .B1(n29451), .B2(
        \xmem_data[63][5] ), .ZN(n7256) );
  NAND4_X1 U10986 ( .A1(n7259), .A2(n7258), .A3(n7257), .A4(n7256), .ZN(n7260)
         );
  AND2_X1 U10987 ( .A1(n7264), .A2(n7292), .ZN(n29471) );
  NAND2_X1 U10988 ( .A1(n7265), .A2(n29471), .ZN(n7295) );
  BUF_X1 U10989 ( .A(n11439), .Z(n29474) );
  AOI22_X1 U10990 ( .A1(n29395), .A2(\xmem_data[0][5] ), .B1(n26884), .B2(
        \xmem_data[1][5] ), .ZN(n7269) );
  AOI22_X1 U10991 ( .A1(n29397), .A2(\xmem_data[2][5] ), .B1(n30948), .B2(
        \xmem_data[3][5] ), .ZN(n7268) );
  AOI22_X1 U10992 ( .A1(n3167), .A2(\xmem_data[4][5] ), .B1(n3190), .B2(
        \xmem_data[5][5] ), .ZN(n7267) );
  AOI22_X1 U10993 ( .A1(n29810), .A2(\xmem_data[6][5] ), .B1(n28147), .B2(
        \xmem_data[7][5] ), .ZN(n7266) );
  NAND4_X1 U10994 ( .A1(n7269), .A2(n7268), .A3(n7267), .A4(n7266), .ZN(n7290)
         );
  AOI22_X1 U10995 ( .A1(n29547), .A2(\xmem_data[8][5] ), .B1(n30170), .B2(
        \xmem_data[9][5] ), .ZN(n7274) );
  AOI22_X1 U10996 ( .A1(n7270), .A2(\xmem_data[10][5] ), .B1(n29573), .B2(
        \xmem_data[11][5] ), .ZN(n7273) );
  AOI22_X1 U10997 ( .A1(n28725), .A2(\xmem_data[12][5] ), .B1(n28696), .B2(
        \xmem_data[13][5] ), .ZN(n7272) );
  BUF_X1 U10998 ( .A(n8075), .Z(n29489) );
  AOI22_X1 U10999 ( .A1(n29489), .A2(\xmem_data[14][5] ), .B1(n21060), .B2(
        \xmem_data[15][5] ), .ZN(n7271) );
  NAND4_X1 U11000 ( .A1(n7274), .A2(n7273), .A3(n7272), .A4(n7271), .ZN(n7289)
         );
  AOI22_X1 U11001 ( .A1(n7275), .A2(\xmem_data[16][5] ), .B1(n29497), .B2(
        \xmem_data[17][5] ), .ZN(n7280) );
  BUF_X1 U11002 ( .A(n7276), .Z(n29499) );
  AOI22_X1 U11003 ( .A1(n29499), .A2(\xmem_data[18][5] ), .B1(n3387), .B2(
        \xmem_data[19][5] ), .ZN(n7279) );
  AOI22_X1 U11004 ( .A1(n29421), .A2(\xmem_data[20][5] ), .B1(n28206), .B2(
        \xmem_data[21][5] ), .ZN(n7278) );
  BUF_X1 U11005 ( .A(n14988), .Z(n29494) );
  AOI22_X1 U11006 ( .A1(n29423), .A2(\xmem_data[22][5] ), .B1(n29494), .B2(
        \xmem_data[23][5] ), .ZN(n7277) );
  NAND4_X1 U11007 ( .A1(n7280), .A2(n7279), .A3(n7278), .A4(n7277), .ZN(n7288)
         );
  BUF_X1 U11008 ( .A(n11780), .Z(n29495) );
  AOI22_X1 U11009 ( .A1(n27771), .A2(\xmem_data[24][5] ), .B1(n28667), .B2(
        \xmem_data[25][5] ), .ZN(n7286) );
  BUF_X1 U11010 ( .A(n7281), .Z(n29501) );
  AOI22_X1 U11011 ( .A1(n29501), .A2(\xmem_data[26][5] ), .B1(n30698), .B2(
        \xmem_data[27][5] ), .ZN(n7285) );
  BUF_X1 U11012 ( .A(n11436), .Z(n29481) );
  AOI22_X1 U11013 ( .A1(n30191), .A2(\xmem_data[28][5] ), .B1(n28665), .B2(
        \xmem_data[29][5] ), .ZN(n7284) );
  AOI22_X1 U11014 ( .A1(n29500), .A2(\xmem_data[30][5] ), .B1(n28743), .B2(
        \xmem_data[31][5] ), .ZN(n7283) );
  NAND4_X1 U11015 ( .A1(n7286), .A2(n7285), .A3(n7284), .A4(n7283), .ZN(n7287)
         );
  NAND2_X1 U11016 ( .A1(n7293), .A2(n29511), .ZN(n7294) );
  XNOR2_X1 U11017 ( .A(n31402), .B(\fmem_data[3][5] ), .ZN(n33030) );
  AOI22_X1 U11018 ( .A1(n29626), .A2(\xmem_data[116][4] ), .B1(n29697), .B2(
        \xmem_data[117][4] ), .ZN(n7298) );
  INV_X1 U11019 ( .A(n7298), .ZN(n7301) );
  BUF_X1 U11020 ( .A(n11437), .Z(n29482) );
  AOI22_X1 U11021 ( .A1(n28739), .A2(\xmem_data[124][4] ), .B1(n27761), .B2(
        \xmem_data[125][4] ), .ZN(n7299) );
  INV_X1 U11022 ( .A(n7299), .ZN(n7300) );
  NOR2_X1 U11023 ( .A1(n7301), .A2(n7300), .ZN(n7315) );
  AOI22_X1 U11024 ( .A1(n28700), .A2(\xmem_data[118][4] ), .B1(n29422), .B2(
        \xmem_data[119][4] ), .ZN(n7314) );
  AOI22_X1 U11025 ( .A1(n29400), .A2(\xmem_data[120][4] ), .B1(n27833), .B2(
        \xmem_data[121][4] ), .ZN(n7302) );
  INV_X1 U11026 ( .A(n7302), .ZN(n7308) );
  AOI22_X1 U11027 ( .A1(n29420), .A2(\xmem_data[114][4] ), .B1(n16980), .B2(
        \xmem_data[115][4] ), .ZN(n7306) );
  AOI22_X1 U11028 ( .A1(n29402), .A2(\xmem_data[122][4] ), .B1(n29350), .B2(
        \xmem_data[123][4] ), .ZN(n7305) );
  AOI22_X1 U11029 ( .A1(n29419), .A2(\xmem_data[112][4] ), .B1(n29418), .B2(
        \xmem_data[113][4] ), .ZN(n7304) );
  AOI22_X1 U11030 ( .A1(n29404), .A2(\xmem_data[126][4] ), .B1(n29403), .B2(
        \xmem_data[127][4] ), .ZN(n7303) );
  NAND4_X1 U11031 ( .A1(n7306), .A2(n7305), .A3(n7304), .A4(n7303), .ZN(n7307)
         );
  NOR2_X1 U11032 ( .A1(n7308), .A2(n7307), .ZN(n7313) );
  AOI22_X1 U11033 ( .A1(n30717), .A2(\xmem_data[104][4] ), .B1(n30765), .B2(
        \xmem_data[105][4] ), .ZN(n7312) );
  AOI22_X1 U11034 ( .A1(n29380), .A2(\xmem_data[106][4] ), .B1(n29379), .B2(
        \xmem_data[107][4] ), .ZN(n7311) );
  AOI22_X1 U11035 ( .A1(n29382), .A2(\xmem_data[108][4] ), .B1(n29381), .B2(
        \xmem_data[109][4] ), .ZN(n7310) );
  AOI22_X1 U11036 ( .A1(n29384), .A2(\xmem_data[110][4] ), .B1(n29383), .B2(
        \xmem_data[111][4] ), .ZN(n7309) );
  NAND4_X1 U11037 ( .A1(n7315), .A2(n7314), .A3(n7313), .A4(n3768), .ZN(n7321)
         );
  AOI22_X1 U11038 ( .A1(n3174), .A2(\xmem_data[96][4] ), .B1(n27753), .B2(
        \xmem_data[97][4] ), .ZN(n7319) );
  AOI22_X1 U11039 ( .A1(n29397), .A2(\xmem_data[98][4] ), .B1(n30892), .B2(
        \xmem_data[99][4] ), .ZN(n7318) );
  AOI22_X1 U11040 ( .A1(n3164), .A2(\xmem_data[100][4] ), .B1(n3183), .B2(
        \xmem_data[101][4] ), .ZN(n7317) );
  BUF_X1 U11041 ( .A(n15549), .Z(n29610) );
  AOI22_X1 U11042 ( .A1(n29610), .A2(\xmem_data[102][4] ), .B1(n29410), .B2(
        \xmem_data[103][4] ), .ZN(n7316) );
  NAND4_X1 U11043 ( .A1(n7319), .A2(n7318), .A3(n7317), .A4(n7316), .ZN(n7320)
         );
  OAI21_X1 U11044 ( .B1(n7321), .B2(n7320), .A(n29428), .ZN(n7398) );
  AOI22_X1 U11045 ( .A1(n30302), .A2(\xmem_data[32][4] ), .B1(n29592), .B2(
        \xmem_data[33][4] ), .ZN(n7325) );
  AOI22_X1 U11046 ( .A1(n29438), .A2(\xmem_data[34][4] ), .B1(n29315), .B2(
        \xmem_data[35][4] ), .ZN(n7324) );
  AOI22_X1 U11047 ( .A1(n3165), .A2(\xmem_data[36][4] ), .B1(n3182), .B2(
        \xmem_data[37][4] ), .ZN(n7323) );
  AOI22_X1 U11048 ( .A1(n28755), .A2(\xmem_data[38][4] ), .B1(n29439), .B2(
        \xmem_data[39][4] ), .ZN(n7322) );
  AOI22_X1 U11049 ( .A1(n30063), .A2(\xmem_data[40][4] ), .B1(n29640), .B2(
        \xmem_data[41][4] ), .ZN(n7329) );
  AOI22_X1 U11050 ( .A1(n29461), .A2(\xmem_data[42][4] ), .B1(n3151), .B2(
        \xmem_data[43][4] ), .ZN(n7328) );
  AOI22_X1 U11051 ( .A1(n29463), .A2(\xmem_data[44][4] ), .B1(n29462), .B2(
        \xmem_data[45][4] ), .ZN(n7327) );
  AOI22_X1 U11052 ( .A1(n29464), .A2(\xmem_data[46][4] ), .B1(n30257), .B2(
        \xmem_data[47][4] ), .ZN(n7326) );
  NAND4_X1 U11053 ( .A1(n7329), .A2(n7328), .A3(n7327), .A4(n7326), .ZN(n7333)
         );
  AOI22_X1 U11054 ( .A1(n27740), .A2(\xmem_data[54][4] ), .B1(n29431), .B2(
        \xmem_data[55][4] ), .ZN(n7331) );
  AOI22_X1 U11055 ( .A1(n29433), .A2(\xmem_data[52][4] ), .B1(n29831), .B2(
        \xmem_data[53][4] ), .ZN(n7330) );
  NAND2_X1 U11056 ( .A1(n7331), .A2(n7330), .ZN(n7332) );
  NOR2_X1 U11057 ( .A1(n7333), .A2(n7332), .ZN(n7343) );
  AOI22_X1 U11058 ( .A1(n29630), .A2(\xmem_data[56][4] ), .B1(n29798), .B2(
        \xmem_data[57][4] ), .ZN(n7342) );
  AOI22_X1 U11059 ( .A1(n29801), .A2(\xmem_data[60][4] ), .B1(n28145), .B2(
        \xmem_data[61][4] ), .ZN(n7334) );
  INV_X1 U11060 ( .A(n7334), .ZN(n7340) );
  AOI22_X1 U11061 ( .A1(n29449), .A2(\xmem_data[50][4] ), .B1(n28039), .B2(
        \xmem_data[51][4] ), .ZN(n7338) );
  AOI22_X1 U11062 ( .A1(n29450), .A2(\xmem_data[58][4] ), .B1(n3135), .B2(
        \xmem_data[59][4] ), .ZN(n7337) );
  AOI22_X1 U11063 ( .A1(n29447), .A2(\xmem_data[48][4] ), .B1(n27743), .B2(
        \xmem_data[49][4] ), .ZN(n7336) );
  AOI22_X1 U11064 ( .A1(n29500), .A2(\xmem_data[62][4] ), .B1(n29451), .B2(
        \xmem_data[63][4] ), .ZN(n7335) );
  NAND4_X1 U11065 ( .A1(n7338), .A2(n7337), .A3(n7336), .A4(n7335), .ZN(n7339)
         );
  NOR2_X1 U11066 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  NAND4_X1 U11067 ( .A1(n7343), .A2(n3848), .A3(n7342), .A4(n7341), .ZN(n7344)
         );
  NAND2_X1 U11068 ( .A1(n7344), .A2(n29471), .ZN(n7397) );
  AOI22_X1 U11069 ( .A1(n29433), .A2(\xmem_data[20][4] ), .B1(n29672), .B2(
        \xmem_data[21][4] ), .ZN(n7348) );
  AOI22_X1 U11070 ( .A1(n29499), .A2(\xmem_data[18][4] ), .B1(n3414), .B2(
        \xmem_data[19][4] ), .ZN(n7347) );
  AOI22_X1 U11071 ( .A1(n29786), .A2(\xmem_data[16][4] ), .B1(n29497), .B2(
        \xmem_data[17][4] ), .ZN(n7346) );
  AOI22_X1 U11072 ( .A1(n28700), .A2(\xmem_data[22][4] ), .B1(n29494), .B2(
        \xmem_data[23][4] ), .ZN(n7345) );
  NAND4_X1 U11073 ( .A1(n7348), .A2(n7347), .A3(n7346), .A4(n7345), .ZN(n7349)
         );
  NAND2_X1 U11074 ( .A1(n7349), .A2(n29511), .ZN(n7374) );
  AOI22_X1 U11075 ( .A1(n29705), .A2(\xmem_data[28][4] ), .B1(n30730), .B2(
        \xmem_data[29][4] ), .ZN(n7353) );
  AOI22_X1 U11076 ( .A1(n29501), .A2(\xmem_data[26][4] ), .B1(n25451), .B2(
        \xmem_data[27][4] ), .ZN(n7352) );
  AOI22_X1 U11077 ( .A1(n30280), .A2(\xmem_data[24][4] ), .B1(n30293), .B2(
        \xmem_data[25][4] ), .ZN(n7351) );
  AOI22_X1 U11078 ( .A1(n29500), .A2(\xmem_data[30][4] ), .B1(n28233), .B2(
        \xmem_data[31][4] ), .ZN(n7350) );
  NAND4_X1 U11079 ( .A1(n7353), .A2(n7352), .A3(n7351), .A4(n7350), .ZN(n7359)
         );
  AOI22_X1 U11080 ( .A1(n29547), .A2(\xmem_data[8][4] ), .B1(n30685), .B2(
        \xmem_data[9][4] ), .ZN(n7357) );
  AOI22_X1 U11081 ( .A1(n7270), .A2(\xmem_data[10][4] ), .B1(n3151), .B2(
        \xmem_data[11][4] ), .ZN(n7356) );
  AOI22_X1 U11082 ( .A1(n29382), .A2(\xmem_data[12][4] ), .B1(n29462), .B2(
        \xmem_data[13][4] ), .ZN(n7355) );
  AOI22_X1 U11083 ( .A1(n29489), .A2(\xmem_data[14][4] ), .B1(n20770), .B2(
        \xmem_data[15][4] ), .ZN(n7354) );
  NAND4_X1 U11084 ( .A1(n7357), .A2(n7356), .A3(n7355), .A4(n7354), .ZN(n7358)
         );
  OAI21_X1 U11085 ( .B1(n7359), .B2(n7358), .A(n29511), .ZN(n7373) );
  BUF_X1 U11086 ( .A(n8700), .Z(n27753) );
  AOI22_X1 U11087 ( .A1(n28751), .A2(\xmem_data[0][4] ), .B1(n30634), .B2(
        \xmem_data[1][4] ), .ZN(n7363) );
  AOI22_X1 U11088 ( .A1(n29438), .A2(\xmem_data[2][4] ), .B1(n30948), .B2(
        \xmem_data[3][4] ), .ZN(n7362) );
  AOI22_X1 U11089 ( .A1(n3164), .A2(\xmem_data[4][4] ), .B1(n3188), .B2(
        \xmem_data[5][4] ), .ZN(n7361) );
  BUF_X1 U11090 ( .A(n15549), .Z(n30075) );
  AOI22_X1 U11091 ( .A1(n30075), .A2(\xmem_data[6][4] ), .B1(n24710), .B2(
        \xmem_data[7][4] ), .ZN(n7360) );
  NAND4_X1 U11092 ( .A1(n7363), .A2(n7362), .A3(n7361), .A4(n7360), .ZN(n7364)
         );
  NAND2_X1 U11093 ( .A1(n7364), .A2(n29511), .ZN(n7372) );
  AOI22_X1 U11094 ( .A1(n29447), .A2(\xmem_data[80][4] ), .B1(n27743), .B2(
        \xmem_data[81][4] ), .ZN(n7369) );
  AOI22_X1 U11095 ( .A1(n29449), .A2(\xmem_data[82][4] ), .B1(n3306), .B2(
        \xmem_data[83][4] ), .ZN(n7368) );
  AOI22_X1 U11096 ( .A1(n30708), .A2(\xmem_data[84][4] ), .B1(n30707), .B2(
        \xmem_data[85][4] ), .ZN(n7367) );
  AND2_X1 U11097 ( .A1(n29431), .A2(\xmem_data[87][4] ), .ZN(n7365) );
  AOI21_X1 U11098 ( .B1(n30215), .B2(\xmem_data[86][4] ), .A(n7365), .ZN(n7366) );
  NAND4_X1 U11099 ( .A1(n7369), .A2(n7368), .A3(n7367), .A4(n7366), .ZN(n7370)
         );
  NAND2_X1 U11100 ( .A1(n7370), .A2(n29376), .ZN(n7371) );
  AND4_X1 U11101 ( .A1(n7374), .A2(n7373), .A3(n7372), .A4(n7371), .ZN(n7396)
         );
  AOI22_X1 U11102 ( .A1(n29446), .A2(\xmem_data[92][4] ), .B1(n30730), .B2(
        \xmem_data[93][4] ), .ZN(n7377) );
  AOI22_X1 U11103 ( .A1(n29438), .A2(\xmem_data[66][4] ), .B1(n23795), .B2(
        \xmem_data[67][4] ), .ZN(n7376) );
  AOI22_X1 U11104 ( .A1(n3164), .A2(\xmem_data[68][4] ), .B1(n3185), .B2(
        \xmem_data[69][4] ), .ZN(n7375) );
  AOI22_X1 U11105 ( .A1(n29547), .A2(\xmem_data[72][4] ), .B1(n30685), .B2(
        \xmem_data[73][4] ), .ZN(n7381) );
  AOI22_X1 U11106 ( .A1(n29461), .A2(\xmem_data[74][4] ), .B1(n3151), .B2(
        \xmem_data[75][4] ), .ZN(n7380) );
  AOI22_X1 U11107 ( .A1(n29463), .A2(\xmem_data[76][4] ), .B1(n29462), .B2(
        \xmem_data[77][4] ), .ZN(n7379) );
  AOI22_X1 U11108 ( .A1(n29464), .A2(\xmem_data[78][4] ), .B1(n20708), .B2(
        \xmem_data[79][4] ), .ZN(n7378) );
  NAND4_X1 U11109 ( .A1(n7381), .A2(n7380), .A3(n7379), .A4(n7378), .ZN(n7382)
         );
  OR2_X1 U11110 ( .A1(n7383), .A2(n7382), .ZN(n7394) );
  AOI22_X1 U11111 ( .A1(n28219), .A2(\xmem_data[88][4] ), .B1(n28208), .B2(
        \xmem_data[89][4] ), .ZN(n7392) );
  AND2_X1 U11112 ( .A1(n29439), .A2(\xmem_data[71][4] ), .ZN(n7384) );
  AOI21_X1 U11113 ( .B1(n29610), .B2(\xmem_data[70][4] ), .A(n7384), .ZN(n7391) );
  AOI22_X1 U11114 ( .A1(n29769), .A2(\xmem_data[64][4] ), .B1(n26884), .B2(
        \xmem_data[65][4] ), .ZN(n7385) );
  INV_X1 U11115 ( .A(n7385), .ZN(n7389) );
  AOI22_X1 U11116 ( .A1(n29450), .A2(\xmem_data[90][4] ), .B1(n3375), .B2(
        \xmem_data[91][4] ), .ZN(n7387) );
  AOI22_X1 U11117 ( .A1(n29500), .A2(\xmem_data[94][4] ), .B1(n29451), .B2(
        \xmem_data[95][4] ), .ZN(n7386) );
  NAND2_X1 U11118 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  NOR2_X1 U11119 ( .A1(n7389), .A2(n7388), .ZN(n7390) );
  OAI21_X1 U11120 ( .B1(n7394), .B2(n7393), .A(n29376), .ZN(n7395) );
  NAND4_X1 U11121 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), .ZN(n32194) );
  XNOR2_X1 U11122 ( .A(n32194), .B(\fmem_data[3][5] ), .ZN(n27333) );
  XOR2_X1 U11123 ( .A(\fmem_data[3][4] ), .B(\fmem_data[3][5] ), .Z(n7399) );
  OAI22_X1 U11124 ( .A1(n33030), .A2(n34919), .B1(n27333), .B2(n34918), .ZN(
        n34269) );
  BUF_X1 U11125 ( .A(n11484), .Z(n27701) );
  AOI22_X1 U11126 ( .A1(n27701), .A2(\xmem_data[48][7] ), .B1(n30217), .B2(
        \xmem_data[49][7] ), .ZN(n7403) );
  NOR2_X1 U11127 ( .A1(n8011), .A2(n3445), .ZN(n26878) );
  BUF_X1 U11128 ( .A(n26878), .Z(n27702) );
  BUF_X1 U11129 ( .A(n14991), .Z(n27762) );
  AOI22_X1 U11130 ( .A1(n27702), .A2(\xmem_data[50][7] ), .B1(n3140), .B2(
        \xmem_data[51][7] ), .ZN(n7402) );
  BUF_X1 U11131 ( .A(n11436), .Z(n27703) );
  BUF_X2 U11132 ( .A(n11437), .Z(n27761) );
  AOI22_X1 U11133 ( .A1(n27703), .A2(\xmem_data[52][7] ), .B1(n28238), .B2(
        \xmem_data[53][7] ), .ZN(n7401) );
  NOR2_X1 U11134 ( .A1(n3377), .A2(n3446), .ZN(n26879) );
  BUF_X1 U11135 ( .A(n14997), .Z(n27763) );
  AOI22_X1 U11136 ( .A1(n29404), .A2(\xmem_data[54][7] ), .B1(n27763), .B2(
        \xmem_data[55][7] ), .ZN(n7400) );
  NAND4_X1 U11137 ( .A1(n7403), .A2(n7402), .A3(n7401), .A4(n7400), .ZN(n7420)
         );
  NOR2_X1 U11138 ( .A1(n11361), .A2(n8010), .ZN(n7451) );
  NOR2_X1 U11139 ( .A1(n3246), .A2(n8010), .ZN(n7452) );
  BUF_X1 U11140 ( .A(n7452), .Z(n27723) );
  AOI22_X1 U11141 ( .A1(n29786), .A2(\xmem_data[40][7] ), .B1(n27723), .B2(
        \xmem_data[41][7] ), .ZN(n7407) );
  NOR2_X1 U11142 ( .A1(n7206), .A2(n8010), .ZN(n11850) );
  BUF_X1 U11143 ( .A(n28973), .Z(n27724) );
  AOI22_X1 U11144 ( .A1(n27742), .A2(\xmem_data[42][7] ), .B1(n3149), .B2(
        \xmem_data[43][7] ), .ZN(n7406) );
  AOI22_X1 U11145 ( .A1(n27741), .A2(\xmem_data[44][7] ), .B1(n29672), .B2(
        \xmem_data[45][7] ), .ZN(n7405) );
  BUF_X1 U11146 ( .A(n14988), .Z(n27708) );
  AOI22_X1 U11147 ( .A1(n30279), .A2(\xmem_data[46][7] ), .B1(n27708), .B2(
        \xmem_data[47][7] ), .ZN(n7404) );
  NAND4_X1 U11148 ( .A1(n7407), .A2(n7406), .A3(n7405), .A4(n7404), .ZN(n7419)
         );
  BUF_X1 U11149 ( .A(n8700), .Z(n30249) );
  AOI22_X1 U11150 ( .A1(n27754), .A2(\xmem_data[56][7] ), .B1(n30301), .B2(
        \xmem_data[57][7] ), .ZN(n7412) );
  NOR2_X1 U11151 ( .A1(n7645), .A2(n3261), .ZN(n11846) );
  BUF_X1 U11152 ( .A(n11846), .Z(n27729) );
  BUF_X1 U11153 ( .A(n29187), .Z(n27818) );
  AOI22_X1 U11154 ( .A1(n27729), .A2(\xmem_data[58][7] ), .B1(n27755), .B2(
        \xmem_data[59][7] ), .ZN(n7411) );
  AOI22_X1 U11155 ( .A1(n3163), .A2(\xmem_data[60][7] ), .B1(n3190), .B2(
        \xmem_data[61][7] ), .ZN(n7410) );
  AOI22_X1 U11156 ( .A1(n23901), .A2(\xmem_data[62][7] ), .B1(n29439), .B2(
        \xmem_data[63][7] ), .ZN(n7409) );
  NAND4_X1 U11157 ( .A1(n7412), .A2(n7411), .A3(n7410), .A4(n7409), .ZN(n7418)
         );
  AOI22_X1 U11158 ( .A1(n29488), .A2(\xmem_data[32][7] ), .B1(n29721), .B2(
        \xmem_data[33][7] ), .ZN(n7416) );
  BUF_X1 U11159 ( .A(n7446), .Z(n27714) );
  AOI22_X1 U11160 ( .A1(n27714), .A2(\xmem_data[34][7] ), .B1(n3337), .B2(
        \xmem_data[35][7] ), .ZN(n7415) );
  BUF_X1 U11161 ( .A(n8073), .Z(n27716) );
  BUF_X1 U11162 ( .A(n8074), .Z(n27715) );
  AOI22_X1 U11163 ( .A1(n27716), .A2(\xmem_data[36][7] ), .B1(n27715), .B2(
        \xmem_data[37][7] ), .ZN(n7414) );
  BUF_X1 U11164 ( .A(n8075), .Z(n27718) );
  BUF_X1 U11165 ( .A(n13420), .Z(n27717) );
  AOI22_X1 U11166 ( .A1(n27718), .A2(\xmem_data[38][7] ), .B1(n27717), .B2(
        \xmem_data[39][7] ), .ZN(n7413) );
  NAND4_X1 U11167 ( .A1(n7416), .A2(n7415), .A3(n7414), .A4(n7413), .ZN(n7417)
         );
  INV_X1 U11168 ( .A(n7421), .ZN(n7422) );
  AOI22_X1 U11169 ( .A1(n7422), .A2(n39040), .B1(n14909), .B2(n7421), .ZN(
        n7469) );
  INV_X1 U11170 ( .A(n7469), .ZN(n7470) );
  INV_X1 U11171 ( .A(n10288), .ZN(n37190) );
  NAND2_X1 U11172 ( .A1(load_xaddr_val[5]), .A2(n37190), .ZN(n10287) );
  OAI22_X1 U11173 ( .A1(n7423), .A2(n10287), .B1(load_xaddr_val[5]), .B2(n7422), .ZN(n7471) );
  AOI22_X1 U11174 ( .A1(n30198), .A2(\xmem_data[0][7] ), .B1(n29640), .B2(
        \xmem_data[1][7] ), .ZN(n7427) );
  AOI22_X1 U11175 ( .A1(n27804), .A2(\xmem_data[2][7] ), .B1(n28955), .B2(
        \xmem_data[3][7] ), .ZN(n7426) );
  AOI22_X1 U11176 ( .A1(n28725), .A2(\xmem_data[4][7] ), .B1(n28696), .B2(
        \xmem_data[5][7] ), .ZN(n7425) );
  AOI22_X1 U11177 ( .A1(n29384), .A2(\xmem_data[6][7] ), .B1(n20708), .B2(
        \xmem_data[7][7] ), .ZN(n7424) );
  NAND4_X1 U11178 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n7443)
         );
  AOI22_X1 U11179 ( .A1(n29419), .A2(\xmem_data[8][7] ), .B1(n27743), .B2(
        \xmem_data[9][7] ), .ZN(n7431) );
  AOI22_X1 U11180 ( .A1(n27742), .A2(\xmem_data[10][7] ), .B1(n3153), .B2(
        \xmem_data[11][7] ), .ZN(n7430) );
  BUF_X1 U11181 ( .A(n11489), .Z(n27741) );
  AOI22_X1 U11182 ( .A1(n28734), .A2(\xmem_data[12][7] ), .B1(n28206), .B2(
        \xmem_data[13][7] ), .ZN(n7429) );
  BUF_X1 U11183 ( .A(n11451), .Z(n27740) );
  AOI22_X1 U11184 ( .A1(n28207), .A2(\xmem_data[14][7] ), .B1(n29832), .B2(
        \xmem_data[15][7] ), .ZN(n7428) );
  NAND4_X1 U11185 ( .A1(n7431), .A2(n7430), .A3(n7429), .A4(n7428), .ZN(n7442)
         );
  AOI22_X1 U11186 ( .A1(n28180), .A2(\xmem_data[20][7] ), .B1(n29347), .B2(
        \xmem_data[21][7] ), .ZN(n7435) );
  BUF_X1 U11187 ( .A(n14991), .Z(n27817) );
  AOI22_X1 U11188 ( .A1(n3223), .A2(\xmem_data[18][7] ), .B1(n3147), .B2(
        \xmem_data[19][7] ), .ZN(n7434) );
  BUF_X1 U11189 ( .A(n11484), .Z(n27771) );
  BUF_X2 U11190 ( .A(n11780), .Z(n27833) );
  AOI22_X1 U11191 ( .A1(n27771), .A2(\xmem_data[16][7] ), .B1(n29495), .B2(
        \xmem_data[17][7] ), .ZN(n7433) );
  AOI22_X1 U11192 ( .A1(n26879), .A2(\xmem_data[22][7] ), .B1(n29179), .B2(
        \xmem_data[23][7] ), .ZN(n7432) );
  NAND4_X1 U11193 ( .A1(n7435), .A2(n7434), .A3(n7433), .A4(n7432), .ZN(n7441)
         );
  AOI22_X1 U11194 ( .A1(n30302), .A2(\xmem_data[24][7] ), .B1(n28684), .B2(
        \xmem_data[25][7] ), .ZN(n7439) );
  BUF_X1 U11195 ( .A(n11846), .Z(n27756) );
  AOI22_X1 U11196 ( .A1(n27756), .A2(\xmem_data[26][7] ), .B1(n28516), .B2(
        \xmem_data[27][7] ), .ZN(n7438) );
  AOI22_X1 U11197 ( .A1(n3163), .A2(\xmem_data[28][7] ), .B1(n3189), .B2(
        \xmem_data[29][7] ), .ZN(n7437) );
  AOI22_X1 U11198 ( .A1(n30715), .A2(\xmem_data[30][7] ), .B1(n28232), .B2(
        \xmem_data[31][7] ), .ZN(n7436) );
  NAND4_X1 U11199 ( .A1(n7439), .A2(n7438), .A3(n7437), .A4(n7436), .ZN(n7440)
         );
  AOI22_X1 U11200 ( .A1(n30717), .A2(\xmem_data[96][7] ), .B1(n29640), .B2(
        \xmem_data[97][7] ), .ZN(n7450) );
  AOI22_X1 U11201 ( .A1(n27804), .A2(\xmem_data[98][7] ), .B1(n28202), .B2(
        \xmem_data[99][7] ), .ZN(n7449) );
  AOI22_X1 U11202 ( .A1(n27716), .A2(\xmem_data[100][7] ), .B1(n27805), .B2(
        \xmem_data[101][7] ), .ZN(n7448) );
  BUF_X1 U11203 ( .A(n8075), .Z(n27806) );
  AOI22_X1 U11204 ( .A1(n27806), .A2(\xmem_data[102][7] ), .B1(n20952), .B2(
        \xmem_data[103][7] ), .ZN(n7447) );
  NAND4_X1 U11205 ( .A1(n7450), .A2(n7449), .A3(n7448), .A4(n7447), .ZN(n7468)
         );
  AOI22_X1 U11206 ( .A1(n7451), .A2(\xmem_data[104][7] ), .B1(n27812), .B2(
        \xmem_data[105][7] ), .ZN(n7456) );
  BUF_X1 U11207 ( .A(n28973), .Z(n27813) );
  AOI22_X1 U11208 ( .A1(n27814), .A2(\xmem_data[106][7] ), .B1(n27813), .B2(
        \xmem_data[107][7] ), .ZN(n7455) );
  AOI22_X1 U11209 ( .A1(n29788), .A2(\xmem_data[108][7] ), .B1(n30707), .B2(
        \xmem_data[109][7] ), .ZN(n7454) );
  BUF_X1 U11210 ( .A(n14988), .Z(n27831) );
  AOI22_X1 U11211 ( .A1(n29423), .A2(\xmem_data[110][7] ), .B1(n27831), .B2(
        \xmem_data[111][7] ), .ZN(n7453) );
  NAND4_X1 U11212 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7467)
         );
  BUF_X1 U11213 ( .A(n11484), .Z(n27834) );
  AOI22_X1 U11214 ( .A1(n27834), .A2(\xmem_data[112][7] ), .B1(n29495), .B2(
        \xmem_data[113][7] ), .ZN(n7460) );
  AOI22_X1 U11215 ( .A1(n3223), .A2(\xmem_data[114][7] ), .B1(n3146), .B2(
        \xmem_data[115][7] ), .ZN(n7459) );
  AOI22_X1 U11216 ( .A1(n27703), .A2(\xmem_data[116][7] ), .B1(n29646), .B2(
        \xmem_data[117][7] ), .ZN(n7458) );
  AOI22_X1 U11217 ( .A1(n29500), .A2(\xmem_data[118][7] ), .B1(n30943), .B2(
        \xmem_data[119][7] ), .ZN(n7457) );
  NAND4_X1 U11218 ( .A1(n7460), .A2(n7459), .A3(n7458), .A4(n7457), .ZN(n7466)
         );
  BUF_X1 U11219 ( .A(n11439), .Z(n27811) );
  AOI22_X1 U11220 ( .A1(n30745), .A2(\xmem_data[120][7] ), .B1(n30249), .B2(
        \xmem_data[121][7] ), .ZN(n7464) );
  BUF_X1 U11221 ( .A(n11846), .Z(n27819) );
  BUF_X1 U11222 ( .A(n3464), .Z(n27755) );
  AOI22_X1 U11223 ( .A1(n27819), .A2(\xmem_data[122][7] ), .B1(n20718), .B2(
        \xmem_data[123][7] ), .ZN(n7463) );
  AOI22_X1 U11224 ( .A1(n3166), .A2(\xmem_data[124][7] ), .B1(n3187), .B2(
        \xmem_data[125][7] ), .ZN(n7462) );
  BUF_X1 U11225 ( .A(n14971), .Z(n27825) );
  AOI22_X1 U11226 ( .A1(n30310), .A2(\xmem_data[126][7] ), .B1(n27825), .B2(
        \xmem_data[127][7] ), .ZN(n7461) );
  NAND4_X1 U11227 ( .A1(n7464), .A2(n7463), .A3(n7462), .A4(n7461), .ZN(n7465)
         );
  OR4_X1 U11228 ( .A1(n7468), .A2(n7467), .A3(n7466), .A4(n7465), .ZN(n7494)
         );
  AND2_X1 U11229 ( .A1(n7471), .A2(n7469), .ZN(n27801) );
  AOI22_X1 U11230 ( .A1(n29786), .A2(\xmem_data[72][7] ), .B1(n27723), .B2(
        \xmem_data[73][7] ), .ZN(n7475) );
  AOI22_X1 U11231 ( .A1(n27742), .A2(\xmem_data[74][7] ), .B1(n3149), .B2(
        \xmem_data[75][7] ), .ZN(n7474) );
  AOI22_X1 U11232 ( .A1(n29788), .A2(\xmem_data[76][7] ), .B1(n26510), .B2(
        \xmem_data[77][7] ), .ZN(n7473) );
  AOI22_X1 U11233 ( .A1(n3392), .A2(\xmem_data[78][7] ), .B1(n27708), .B2(
        \xmem_data[79][7] ), .ZN(n7472) );
  NAND4_X1 U11234 ( .A1(n7475), .A2(n7474), .A3(n7473), .A4(n7472), .ZN(n7492)
         );
  AOI22_X1 U11235 ( .A1(n27701), .A2(\xmem_data[80][7] ), .B1(n30776), .B2(
        \xmem_data[81][7] ), .ZN(n7479) );
  AOI22_X1 U11236 ( .A1(n27702), .A2(\xmem_data[82][7] ), .B1(n3147), .B2(
        \xmem_data[83][7] ), .ZN(n7478) );
  AOI22_X1 U11237 ( .A1(n29390), .A2(\xmem_data[84][7] ), .B1(n29646), .B2(
        \xmem_data[85][7] ), .ZN(n7477) );
  AOI22_X1 U11238 ( .A1(n26879), .A2(\xmem_data[86][7] ), .B1(n28671), .B2(
        \xmem_data[87][7] ), .ZN(n7476) );
  NAND4_X1 U11239 ( .A1(n7479), .A2(n7478), .A3(n7477), .A4(n7476), .ZN(n7491)
         );
  AOI22_X1 U11240 ( .A1(n29769), .A2(\xmem_data[88][7] ), .B1(n29739), .B2(
        \xmem_data[89][7] ), .ZN(n7484) );
  AOI22_X1 U11241 ( .A1(n27729), .A2(\xmem_data[90][7] ), .B1(n30666), .B2(
        \xmem_data[91][7] ), .ZN(n7483) );
  AOI22_X1 U11242 ( .A1(n3164), .A2(\xmem_data[92][7] ), .B1(n3190), .B2(
        \xmem_data[93][7] ), .ZN(n7482) );
  AND2_X1 U11243 ( .A1(n30309), .A2(\xmem_data[95][7] ), .ZN(n7480) );
  AOI21_X1 U11244 ( .B1(n29610), .B2(\xmem_data[94][7] ), .A(n7480), .ZN(n7481) );
  NAND4_X1 U11245 ( .A1(n7484), .A2(n7483), .A3(n7482), .A4(n7481), .ZN(n7490)
         );
  AOI22_X1 U11246 ( .A1(n30076), .A2(\xmem_data[64][7] ), .B1(n29721), .B2(
        \xmem_data[65][7] ), .ZN(n7488) );
  AOI22_X1 U11247 ( .A1(n27714), .A2(\xmem_data[66][7] ), .B1(n3271), .B2(
        \xmem_data[67][7] ), .ZN(n7487) );
  AOI22_X1 U11248 ( .A1(n27716), .A2(\xmem_data[68][7] ), .B1(n27715), .B2(
        \xmem_data[69][7] ), .ZN(n7486) );
  AOI22_X1 U11249 ( .A1(n27718), .A2(\xmem_data[70][7] ), .B1(n27717), .B2(
        \xmem_data[71][7] ), .ZN(n7485) );
  NAND4_X1 U11250 ( .A1(n7488), .A2(n7487), .A3(n7486), .A4(n7485), .ZN(n7489)
         );
  AOI22_X1 U11251 ( .A1(n7494), .A2(n27801), .B1(n27839), .B2(n7493), .ZN(
        n7495) );
  XNOR2_X1 U11252 ( .A(n35242), .B(\fmem_data[27][3] ), .ZN(n30438) );
  AOI22_X1 U11253 ( .A1(n29419), .A2(\xmem_data[72][6] ), .B1(n27723), .B2(
        \xmem_data[73][6] ), .ZN(n7500) );
  AOI22_X1 U11254 ( .A1(n11850), .A2(\xmem_data[74][6] ), .B1(n3149), .B2(
        \xmem_data[75][6] ), .ZN(n7499) );
  AOI22_X1 U11255 ( .A1(n29626), .A2(\xmem_data[76][6] ), .B1(n30290), .B2(
        \xmem_data[77][6] ), .ZN(n7498) );
  AOI22_X1 U11256 ( .A1(n28138), .A2(\xmem_data[78][6] ), .B1(n27708), .B2(
        \xmem_data[79][6] ), .ZN(n7497) );
  NAND4_X1 U11257 ( .A1(n7500), .A2(n7499), .A3(n7498), .A4(n7497), .ZN(n7518)
         );
  BUF_X1 U11258 ( .A(n8700), .Z(n29648) );
  AOI22_X1 U11259 ( .A1(n29604), .A2(\xmem_data[88][6] ), .B1(n30084), .B2(
        \xmem_data[89][6] ), .ZN(n7505) );
  AOI22_X1 U11260 ( .A1(n27729), .A2(\xmem_data[90][6] ), .B1(n30892), .B2(
        \xmem_data[91][6] ), .ZN(n7504) );
  AOI22_X1 U11261 ( .A1(n3167), .A2(\xmem_data[92][6] ), .B1(n3185), .B2(
        \xmem_data[93][6] ), .ZN(n7503) );
  AND2_X1 U11262 ( .A1(n27825), .A2(\xmem_data[95][6] ), .ZN(n7501) );
  AOI21_X1 U11263 ( .B1(n30075), .B2(\xmem_data[94][6] ), .A(n7501), .ZN(n7502) );
  NAND4_X1 U11264 ( .A1(n7505), .A2(n7504), .A3(n7503), .A4(n7502), .ZN(n7516)
         );
  AOI22_X1 U11265 ( .A1(n27701), .A2(\xmem_data[80][6] ), .B1(n30696), .B2(
        \xmem_data[81][6] ), .ZN(n7509) );
  AOI22_X1 U11266 ( .A1(n27702), .A2(\xmem_data[82][6] ), .B1(n3147), .B2(
        \xmem_data[83][6] ), .ZN(n7508) );
  AOI22_X1 U11267 ( .A1(n3249), .A2(\xmem_data[84][6] ), .B1(n28238), .B2(
        \xmem_data[85][6] ), .ZN(n7507) );
  AOI22_X1 U11268 ( .A1(n26879), .A2(\xmem_data[86][6] ), .B1(n17013), .B2(
        \xmem_data[87][6] ), .ZN(n7506) );
  NAND4_X1 U11269 ( .A1(n7509), .A2(n7508), .A3(n7507), .A4(n7506), .ZN(n7515)
         );
  BUF_X1 U11270 ( .A(n10802), .Z(n28173) );
  BUF_X2 U11271 ( .A(n18518), .Z(n30685) );
  AOI22_X1 U11272 ( .A1(n29815), .A2(\xmem_data[64][6] ), .B1(n30266), .B2(
        \xmem_data[65][6] ), .ZN(n7513) );
  BUF_X1 U11273 ( .A(\xmem_data[66][6] ), .Z(n20682) );
  AOI22_X1 U11274 ( .A1(n27714), .A2(n20682), .B1(n3269), .B2(
        \xmem_data[67][6] ), .ZN(n7512) );
  AOI22_X1 U11275 ( .A1(n27716), .A2(\xmem_data[68][6] ), .B1(n27715), .B2(
        \xmem_data[69][6] ), .ZN(n7511) );
  AOI22_X1 U11276 ( .A1(n27718), .A2(\xmem_data[70][6] ), .B1(n27717), .B2(
        \xmem_data[71][6] ), .ZN(n7510) );
  NAND4_X1 U11277 ( .A1(n7513), .A2(n7512), .A3(n7511), .A4(n7510), .ZN(n7514)
         );
  OAI21_X1 U11278 ( .B1(n7518), .B2(n7517), .A(n27839), .ZN(n7593) );
  AOI22_X1 U11279 ( .A1(n30250), .A2(\xmem_data[56][6] ), .B1(n30090), .B2(
        \xmem_data[57][6] ), .ZN(n7522) );
  AOI22_X1 U11280 ( .A1(n27729), .A2(\xmem_data[58][6] ), .B1(n3465), .B2(
        \xmem_data[59][6] ), .ZN(n7521) );
  AOI22_X1 U11281 ( .A1(n3165), .A2(\xmem_data[60][6] ), .B1(n3184), .B2(
        \xmem_data[61][6] ), .ZN(n7520) );
  AOI22_X1 U11282 ( .A1(n29610), .A2(\xmem_data[62][6] ), .B1(n29239), .B2(
        \xmem_data[63][6] ), .ZN(n7519) );
  NAND4_X1 U11283 ( .A1(n7522), .A2(n7521), .A3(n7520), .A4(n7519), .ZN(n7528)
         );
  AOI22_X1 U11284 ( .A1(n27701), .A2(\xmem_data[48][6] ), .B1(n29761), .B2(
        \xmem_data[49][6] ), .ZN(n7526) );
  AOI22_X1 U11285 ( .A1(n27702), .A2(\xmem_data[50][6] ), .B1(n3147), .B2(
        \xmem_data[51][6] ), .ZN(n7525) );
  AOI22_X1 U11286 ( .A1(n29446), .A2(\xmem_data[52][6] ), .B1(n29646), .B2(
        \xmem_data[53][6] ), .ZN(n7524) );
  AOI22_X1 U11287 ( .A1(n29500), .A2(\xmem_data[54][6] ), .B1(n22738), .B2(
        \xmem_data[55][6] ), .ZN(n7523) );
  NAND4_X1 U11288 ( .A1(n7526), .A2(n7525), .A3(n7524), .A4(n7523), .ZN(n7527)
         );
  OR2_X1 U11289 ( .A1(n7528), .A2(n7527), .ZN(n7541) );
  BUF_X1 U11290 ( .A(n10802), .Z(n30076) );
  AOI22_X1 U11291 ( .A1(n29815), .A2(\xmem_data[32][6] ), .B1(n30765), .B2(
        \xmem_data[33][6] ), .ZN(n7532) );
  AOI22_X1 U11292 ( .A1(n27714), .A2(\xmem_data[34][6] ), .B1(n3269), .B2(
        \xmem_data[35][6] ), .ZN(n7531) );
  AOI22_X1 U11293 ( .A1(n27716), .A2(\xmem_data[36][6] ), .B1(n27715), .B2(
        \xmem_data[37][6] ), .ZN(n7530) );
  AOI22_X1 U11294 ( .A1(n27718), .A2(\xmem_data[38][6] ), .B1(n27717), .B2(
        \xmem_data[39][6] ), .ZN(n7529) );
  AOI22_X1 U11295 ( .A1(n29423), .A2(\xmem_data[46][6] ), .B1(n27708), .B2(
        \xmem_data[47][6] ), .ZN(n7533) );
  INV_X1 U11296 ( .A(n7533), .ZN(n7538) );
  BUF_X1 U11297 ( .A(n7903), .Z(n26510) );
  AOI22_X1 U11298 ( .A1(n27710), .A2(\xmem_data[44][6] ), .B1(n29672), .B2(
        \xmem_data[45][6] ), .ZN(n7536) );
  AOI22_X1 U11299 ( .A1(n27742), .A2(\xmem_data[42][6] ), .B1(n3149), .B2(
        \xmem_data[43][6] ), .ZN(n7535) );
  AOI22_X1 U11300 ( .A1(n29419), .A2(\xmem_data[40][6] ), .B1(n27723), .B2(
        \xmem_data[41][6] ), .ZN(n7534) );
  NOR2_X1 U11301 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  NAND2_X1 U11302 ( .A1(n3771), .A2(n7539), .ZN(n7540) );
  OAI21_X1 U11303 ( .B1(n7541), .B2(n7540), .A(n27737), .ZN(n7592) );
  AOI22_X1 U11304 ( .A1(n29395), .A2(\xmem_data[120][6] ), .B1(n30193), .B2(
        \xmem_data[121][6] ), .ZN(n7542) );
  INV_X1 U11305 ( .A(n7542), .ZN(n7547) );
  AOI22_X1 U11306 ( .A1(n27819), .A2(\xmem_data[122][6] ), .B1(n30666), .B2(
        \xmem_data[123][6] ), .ZN(n7545) );
  AOI22_X1 U11307 ( .A1(n27814), .A2(\xmem_data[106][6] ), .B1(n27813), .B2(
        \xmem_data[107][6] ), .ZN(n7544) );
  AOI22_X1 U11308 ( .A1(n7451), .A2(\xmem_data[104][6] ), .B1(n27812), .B2(
        \xmem_data[105][6] ), .ZN(n7543) );
  NAND3_X1 U11309 ( .A1(n7545), .A2(n7544), .A3(n7543), .ZN(n7546) );
  NOR2_X1 U11310 ( .A1(n7547), .A2(n7546), .ZN(n7550) );
  AOI22_X1 U11311 ( .A1(n28734), .A2(\xmem_data[108][6] ), .B1(n30290), .B2(
        \xmem_data[109][6] ), .ZN(n7549) );
  AOI22_X1 U11312 ( .A1(n3165), .A2(\xmem_data[124][6] ), .B1(n3187), .B2(
        \xmem_data[125][6] ), .ZN(n7548) );
  NAND3_X1 U11313 ( .A1(n7550), .A2(n7549), .A3(n7548), .ZN(n7556) );
  AOI22_X1 U11314 ( .A1(n27834), .A2(\xmem_data[112][6] ), .B1(n29495), .B2(
        \xmem_data[113][6] ), .ZN(n7554) );
  AOI22_X1 U11315 ( .A1(n3223), .A2(\xmem_data[114][6] ), .B1(n3140), .B2(
        \xmem_data[115][6] ), .ZN(n7553) );
  AOI22_X1 U11316 ( .A1(n29390), .A2(\xmem_data[116][6] ), .B1(n29646), .B2(
        \xmem_data[117][6] ), .ZN(n7552) );
  AOI22_X1 U11317 ( .A1(n29500), .A2(\xmem_data[118][6] ), .B1(n27763), .B2(
        \xmem_data[119][6] ), .ZN(n7551) );
  NAND4_X1 U11318 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n7555)
         );
  AOI22_X1 U11319 ( .A1(n27713), .A2(\xmem_data[96][6] ), .B1(n29721), .B2(
        \xmem_data[97][6] ), .ZN(n7560) );
  AOI22_X1 U11320 ( .A1(n27804), .A2(\xmem_data[98][6] ), .B1(n17004), .B2(
        \xmem_data[99][6] ), .ZN(n7559) );
  AOI22_X1 U11321 ( .A1(n29819), .A2(\xmem_data[100][6] ), .B1(n27805), .B2(
        \xmem_data[101][6] ), .ZN(n7558) );
  AOI22_X1 U11322 ( .A1(n27806), .A2(\xmem_data[102][6] ), .B1(n25584), .B2(
        \xmem_data[103][6] ), .ZN(n7557) );
  AOI22_X1 U11323 ( .A1(n28207), .A2(\xmem_data[110][6] ), .B1(n27831), .B2(
        \xmem_data[111][6] ), .ZN(n7562) );
  AOI22_X1 U11324 ( .A1(n30062), .A2(\xmem_data[126][6] ), .B1(n27825), .B2(
        \xmem_data[127][6] ), .ZN(n7561) );
  NAND3_X1 U11325 ( .A1(n3526), .A2(n7562), .A3(n7561), .ZN(n7563) );
  AOI22_X1 U11326 ( .A1(n30708), .A2(\xmem_data[12][6] ), .B1(n30100), .B2(
        \xmem_data[13][6] ), .ZN(n7565) );
  INV_X1 U11327 ( .A(n7565), .ZN(n7575) );
  AOI22_X1 U11328 ( .A1(n3223), .A2(\xmem_data[18][6] ), .B1(n3146), .B2(
        \xmem_data[19][6] ), .ZN(n7568) );
  AOI22_X1 U11329 ( .A1(n29419), .A2(\xmem_data[8][6] ), .B1(n27743), .B2(
        \xmem_data[9][6] ), .ZN(n7567) );
  AOI22_X1 U11330 ( .A1(n26879), .A2(\xmem_data[22][6] ), .B1(n31327), .B2(
        \xmem_data[23][6] ), .ZN(n7566) );
  NAND3_X1 U11331 ( .A1(n7568), .A2(n7567), .A3(n7566), .ZN(n7574) );
  AOI22_X1 U11332 ( .A1(n27756), .A2(\xmem_data[26][6] ), .B1(n30303), .B2(
        \xmem_data[27][6] ), .ZN(n7570) );
  AOI22_X1 U11333 ( .A1(n27742), .A2(\xmem_data[10][6] ), .B1(n3149), .B2(
        \xmem_data[11][6] ), .ZN(n7569) );
  NAND2_X1 U11334 ( .A1(n7570), .A2(n7569), .ZN(n7573) );
  AOI22_X1 U11335 ( .A1(n28685), .A2(\xmem_data[24][6] ), .B1(n30237), .B2(
        \xmem_data[25][6] ), .ZN(n7571) );
  INV_X1 U11336 ( .A(n7571), .ZN(n7572) );
  NOR4_X1 U11337 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n7588)
         );
  AOI22_X1 U11338 ( .A1(n30063), .A2(\xmem_data[0][6] ), .B1(n30170), .B2(
        \xmem_data[1][6] ), .ZN(n7579) );
  AOI22_X1 U11339 ( .A1(n7446), .A2(\xmem_data[2][6] ), .B1(n3308), .B2(
        \xmem_data[3][6] ), .ZN(n7578) );
  AOI22_X1 U11340 ( .A1(n29463), .A2(\xmem_data[4][6] ), .B1(n27715), .B2(
        \xmem_data[5][6] ), .ZN(n7577) );
  AOI22_X1 U11341 ( .A1(n28727), .A2(\xmem_data[6][6] ), .B1(n25407), .B2(
        \xmem_data[7][6] ), .ZN(n7576) );
  BUF_X1 U11342 ( .A(n15549), .Z(n30070) );
  AOI22_X1 U11343 ( .A1(n30070), .A2(\xmem_data[30][6] ), .B1(n28754), .B2(
        \xmem_data[31][6] ), .ZN(n7581) );
  AOI22_X1 U11344 ( .A1(n3168), .A2(\xmem_data[28][6] ), .B1(n3182), .B2(
        \xmem_data[29][6] ), .ZN(n7580) );
  AOI22_X1 U11345 ( .A1(n29628), .A2(\xmem_data[14][6] ), .B1(n30292), .B2(
        \xmem_data[15][6] ), .ZN(n7582) );
  INV_X1 U11346 ( .A(n7582), .ZN(n7586) );
  AOI22_X1 U11347 ( .A1(n27771), .A2(\xmem_data[16][6] ), .B1(n29629), .B2(
        \xmem_data[17][6] ), .ZN(n7584) );
  AOI22_X1 U11348 ( .A1(n29705), .A2(\xmem_data[20][6] ), .B1(n27761), .B2(
        \xmem_data[21][6] ), .ZN(n7583) );
  NAND2_X1 U11349 ( .A1(n7584), .A2(n7583), .ZN(n7585) );
  NOR2_X1 U11350 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  NAND4_X1 U11351 ( .A1(n7588), .A2(n3534), .A3(n3929), .A4(n7587), .ZN(n7589)
         );
  NAND2_X1 U11352 ( .A1(n7589), .A2(n27778), .ZN(n7590) );
  XNOR2_X1 U11353 ( .A(n35145), .B(\fmem_data[27][3] ), .ZN(n22453) );
  XOR2_X1 U11354 ( .A(\fmem_data[27][2] ), .B(\fmem_data[27][3] ), .Z(n7594)
         );
  OAI22_X1 U11355 ( .A1(n30438), .A2(n34463), .B1(n22453), .B2(n34462), .ZN(
        n34268) );
  NOR2_X1 U11356 ( .A1(n11361), .A2(n8010), .ZN(n8088) );
  NOR2_X1 U11357 ( .A1(n8010), .A2(n3246), .ZN(n7691) );
  AOI22_X1 U11358 ( .A1(n29786), .A2(\xmem_data[32][6] ), .B1(n29785), .B2(
        \xmem_data[33][6] ), .ZN(n7598) );
  NAND3_X1 U11359 ( .A1(n11343), .A2(n11342), .A3(n6173), .ZN(n7645) );
  NOR2_X1 U11360 ( .A1(n8010), .A2(n7645), .ZN(n7692) );
  BUF_X1 U11361 ( .A(n7692), .Z(n29787) );
  AOI22_X1 U11362 ( .A1(n29787), .A2(\xmem_data[34][6] ), .B1(n25725), .B2(
        \xmem_data[35][6] ), .ZN(n7597) );
  AOI22_X1 U11363 ( .A1(n28734), .A2(\xmem_data[36][6] ), .B1(n27832), .B2(
        \xmem_data[37][6] ), .ZN(n7596) );
  BUF_X2 U11364 ( .A(n11451), .Z(n29790) );
  BUF_X1 U11365 ( .A(n14988), .Z(n29789) );
  AOI22_X1 U11366 ( .A1(n29423), .A2(\xmem_data[38][6] ), .B1(n29789), .B2(
        \xmem_data[39][6] ), .ZN(n7595) );
  NAND4_X1 U11367 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n7607)
         );
  NOR2_X1 U11368 ( .A1(n7601), .A2(n39041), .ZN(n7600) );
  OAI22_X1 U11369 ( .A1(n7601), .A2(n20978), .B1(n7600), .B2(n39040), .ZN(
        n7612) );
  INV_X1 U11370 ( .A(n7612), .ZN(n7618) );
  AOI21_X1 U11371 ( .B1(n7601), .B2(n39041), .A(n7600), .ZN(n7619) );
  AND2_X1 U11372 ( .A1(n7618), .A2(n7619), .ZN(n29795) );
  AOI22_X1 U11373 ( .A1(n29722), .A2(\xmem_data[24][6] ), .B1(n29640), .B2(
        \xmem_data[25][6] ), .ZN(n7605) );
  AOI22_X1 U11374 ( .A1(n3226), .A2(\xmem_data[26][6] ), .B1(n28701), .B2(
        \xmem_data[27][6] ), .ZN(n7604) );
  BUF_X1 U11375 ( .A(n8073), .Z(n29724) );
  BUF_X1 U11376 ( .A(n8074), .Z(n29723) );
  AOI22_X1 U11377 ( .A1(n29724), .A2(\xmem_data[28][6] ), .B1(n29723), .B2(
        \xmem_data[29][6] ), .ZN(n7603) );
  BUF_X1 U11378 ( .A(n8075), .Z(n29726) );
  BUF_X1 U11379 ( .A(n13127), .Z(n29725) );
  AOI22_X1 U11380 ( .A1(n29726), .A2(\xmem_data[30][6] ), .B1(n29725), .B2(
        \xmem_data[31][6] ), .ZN(n7602) );
  NAND4_X1 U11381 ( .A1(n7605), .A2(n7604), .A3(n7603), .A4(n7602), .ZN(n7606)
         );
  AOI22_X1 U11382 ( .A1(n7607), .A2(n29795), .B1(n7606), .B2(n29733), .ZN(
        n7629) );
  BUF_X2 U11383 ( .A(n8088), .Z(n29829) );
  AOI22_X1 U11384 ( .A1(n28765), .A2(\xmem_data[96][6] ), .B1(n29785), .B2(
        \xmem_data[97][6] ), .ZN(n7611) );
  BUF_X1 U11385 ( .A(n7692), .Z(n29830) );
  AOI22_X1 U11386 ( .A1(n29830), .A2(\xmem_data[98][6] ), .B1(n30864), .B2(
        \xmem_data[99][6] ), .ZN(n7610) );
  AOI22_X1 U11387 ( .A1(n29421), .A2(\xmem_data[100][6] ), .B1(n30106), .B2(
        \xmem_data[101][6] ), .ZN(n7609) );
  BUF_X1 U11388 ( .A(n14988), .Z(n29832) );
  AOI22_X1 U11389 ( .A1(n28138), .A2(\xmem_data[102][6] ), .B1(n29832), .B2(
        \xmem_data[103][6] ), .ZN(n7608) );
  NAND4_X1 U11390 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n7613)
         );
  AND2_X1 U11391 ( .A1(n7619), .A2(n7612), .ZN(n29837) );
  NAND2_X1 U11392 ( .A1(n7613), .A2(n29837), .ZN(n7628) );
  AOI22_X1 U11393 ( .A1(n29829), .A2(\xmem_data[64][6] ), .B1(n29785), .B2(
        \xmem_data[65][6] ), .ZN(n7617) );
  AOI22_X1 U11394 ( .A1(n29787), .A2(\xmem_data[66][6] ), .B1(n23732), .B2(
        \xmem_data[67][6] ), .ZN(n7616) );
  AOI22_X1 U11395 ( .A1(n29433), .A2(\xmem_data[68][6] ), .B1(n29432), .B2(
        \xmem_data[69][6] ), .ZN(n7615) );
  AOI22_X1 U11396 ( .A1(n28700), .A2(\xmem_data[70][6] ), .B1(n29789), .B2(
        \xmem_data[71][6] ), .ZN(n7614) );
  NAND4_X1 U11397 ( .A1(n7617), .A2(n7616), .A3(n7615), .A4(n7614), .ZN(n7620)
         );
  NAND2_X1 U11398 ( .A1(n7620), .A2(n29758), .ZN(n7627) );
  BUF_X1 U11399 ( .A(n11780), .Z(n29761) );
  AOI22_X1 U11400 ( .A1(n29799), .A2(\xmem_data[40][6] ), .B1(n30776), .B2(
        \xmem_data[41][6] ), .ZN(n7624) );
  NOR2_X1 U11401 ( .A1(n7010), .A2(n3445), .ZN(n7658) );
  AOI22_X1 U11402 ( .A1(n29707), .A2(\xmem_data[42][6] ), .B1(n3375), .B2(
        \xmem_data[43][6] ), .ZN(n7623) );
  AOI22_X1 U11403 ( .A1(n28146), .A2(\xmem_data[44][6] ), .B1(n29347), .B2(
        \xmem_data[45][6] ), .ZN(n7622) );
  NOR2_X1 U11404 ( .A1(n11360), .A2(n3445), .ZN(n7659) );
  BUF_X1 U11405 ( .A(n7659), .Z(n29763) );
  AOI22_X1 U11406 ( .A1(n29763), .A2(\xmem_data[46][6] ), .B1(n20587), .B2(
        \xmem_data[47][6] ), .ZN(n7621) );
  NAND4_X1 U11407 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n7625)
         );
  NAND2_X1 U11408 ( .A1(n7625), .A2(n29795), .ZN(n7626) );
  NAND4_X1 U11409 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n7704)
         );
  AOI22_X1 U11410 ( .A1(n30076), .A2(\xmem_data[88][6] ), .B1(n30765), .B2(
        \xmem_data[89][6] ), .ZN(n7633) );
  AOI22_X1 U11411 ( .A1(n3226), .A2(\xmem_data[90][6] ), .B1(n28701), .B2(
        \xmem_data[91][6] ), .ZN(n7632) );
  BUF_X1 U11412 ( .A(n8073), .Z(n29777) );
  BUF_X1 U11413 ( .A(n8074), .Z(n29776) );
  AOI22_X1 U11414 ( .A1(n29777), .A2(\xmem_data[92][6] ), .B1(n29776), .B2(
        \xmem_data[93][6] ), .ZN(n7631) );
  AOI22_X1 U11415 ( .A1(n28727), .A2(\xmem_data[94][6] ), .B1(n29327), .B2(
        \xmem_data[95][6] ), .ZN(n7630) );
  NAND4_X1 U11416 ( .A1(n7633), .A2(n7632), .A3(n7631), .A4(n7630), .ZN(n7639)
         );
  BUF_X1 U11417 ( .A(n10802), .Z(n27713) );
  AOI22_X1 U11418 ( .A1(n30717), .A2(\xmem_data[56][6] ), .B1(n30716), .B2(
        \xmem_data[57][6] ), .ZN(n7637) );
  BUF_X1 U11419 ( .A(n14974), .Z(n29816) );
  AOI22_X1 U11420 ( .A1(n3226), .A2(\xmem_data[58][6] ), .B1(n29816), .B2(
        \xmem_data[59][6] ), .ZN(n7636) );
  BUF_X1 U11421 ( .A(n8073), .Z(n29819) );
  BUF_X1 U11422 ( .A(n8074), .Z(n29818) );
  AOI22_X1 U11423 ( .A1(n29819), .A2(\xmem_data[60][6] ), .B1(n29818), .B2(
        \xmem_data[61][6] ), .ZN(n7635) );
  BUF_X1 U11424 ( .A(n8075), .Z(n29821) );
  BUF_X1 U11425 ( .A(n13420), .Z(n29820) );
  AOI22_X1 U11426 ( .A1(n29821), .A2(\xmem_data[62][6] ), .B1(n29820), .B2(
        \xmem_data[63][6] ), .ZN(n7634) );
  NAND4_X1 U11427 ( .A1(n7637), .A2(n7636), .A3(n7635), .A4(n7634), .ZN(n7638)
         );
  AOI22_X1 U11428 ( .A1(n29758), .A2(n7639), .B1(n7638), .B2(n29795), .ZN(
        n7668) );
  BUF_X1 U11429 ( .A(n10802), .Z(n29815) );
  AOI22_X1 U11430 ( .A1(n29363), .A2(\xmem_data[120][6] ), .B1(n30765), .B2(
        \xmem_data[121][6] ), .ZN(n7644) );
  BUF_X1 U11431 ( .A(n7640), .Z(n29817) );
  AOI22_X1 U11432 ( .A1(n29817), .A2(\xmem_data[122][6] ), .B1(n3151), .B2(
        \xmem_data[123][6] ), .ZN(n7643) );
  AOI22_X1 U11433 ( .A1(n29724), .A2(\xmem_data[124][6] ), .B1(n29723), .B2(
        \xmem_data[125][6] ), .ZN(n7642) );
  AOI22_X1 U11434 ( .A1(n29726), .A2(\xmem_data[126][6] ), .B1(n29725), .B2(
        \xmem_data[127][6] ), .ZN(n7641) );
  NAND4_X1 U11435 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7652)
         );
  BUF_X1 U11436 ( .A(n11439), .Z(n29714) );
  AOI22_X1 U11437 ( .A1(n27754), .A2(\xmem_data[16][6] ), .B1(n30634), .B2(
        \xmem_data[17][6] ), .ZN(n7650) );
  NOR2_X1 U11438 ( .A1(n7010), .A2(n8000), .ZN(n15525) );
  BUF_X1 U11439 ( .A(n15525), .Z(n29771) );
  AOI22_X1 U11440 ( .A1(n29771), .A2(\xmem_data[18][6] ), .B1(n28154), .B2(
        \xmem_data[19][6] ), .ZN(n7649) );
  AOI22_X1 U11441 ( .A1(n3165), .A2(\xmem_data[20][6] ), .B1(n3189), .B2(
        \xmem_data[21][6] ), .ZN(n7648) );
  AND2_X1 U11442 ( .A1(n28781), .A2(\xmem_data[23][6] ), .ZN(n7646) );
  AOI21_X1 U11443 ( .B1(n29716), .B2(\xmem_data[22][6] ), .A(n7646), .ZN(n7647) );
  NAND4_X1 U11444 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .ZN(n7651)
         );
  AOI22_X1 U11445 ( .A1(n29837), .A2(n7652), .B1(n7651), .B2(n29733), .ZN(
        n7667) );
  BUF_X1 U11446 ( .A(n11484), .Z(n29799) );
  AOI22_X1 U11447 ( .A1(n29799), .A2(\xmem_data[104][6] ), .B1(n30293), .B2(
        \xmem_data[105][6] ), .ZN(n7656) );
  BUF_X1 U11448 ( .A(n7658), .Z(n29800) );
  BUF_X1 U11449 ( .A(n14991), .Z(n29706) );
  AOI22_X1 U11450 ( .A1(n29800), .A2(\xmem_data[106][6] ), .B1(n29706), .B2(
        \xmem_data[107][6] ), .ZN(n7655) );
  BUF_X1 U11451 ( .A(n11436), .Z(n29801) );
  BUF_X1 U11452 ( .A(n11437), .Z(n29704) );
  AOI22_X1 U11453 ( .A1(n29801), .A2(\xmem_data[108][6] ), .B1(n29646), .B2(
        \xmem_data[109][6] ), .ZN(n7654) );
  BUF_X1 U11454 ( .A(n7659), .Z(n29802) );
  AOI22_X1 U11455 ( .A1(n29802), .A2(\xmem_data[110][6] ), .B1(n31353), .B2(
        \xmem_data[111][6] ), .ZN(n7653) );
  NAND4_X1 U11456 ( .A1(n7656), .A2(n7655), .A3(n7654), .A4(n7653), .ZN(n7657)
         );
  NAND2_X1 U11457 ( .A1(n7657), .A2(n29837), .ZN(n7666) );
  BUF_X1 U11458 ( .A(n11780), .Z(n29708) );
  AOI22_X1 U11459 ( .A1(n29630), .A2(\xmem_data[8][6] ), .B1(n30696), .B2(
        \xmem_data[9][6] ), .ZN(n7663) );
  AOI22_X1 U11460 ( .A1(n29707), .A2(\xmem_data[10][6] ), .B1(n29706), .B2(
        \xmem_data[11][6] ), .ZN(n7662) );
  BUF_X1 U11461 ( .A(n11436), .Z(n29705) );
  AOI22_X1 U11462 ( .A1(n29705), .A2(\xmem_data[12][6] ), .B1(n28665), .B2(
        \xmem_data[13][6] ), .ZN(n7661) );
  AOI22_X1 U11463 ( .A1(n29709), .A2(\xmem_data[14][6] ), .B1(n30508), .B2(
        \xmem_data[15][6] ), .ZN(n7660) );
  NAND4_X1 U11464 ( .A1(n7663), .A2(n7662), .A3(n7661), .A4(n7660), .ZN(n7664)
         );
  NAND2_X1 U11465 ( .A1(n7664), .A2(n29733), .ZN(n7665) );
  NAND4_X1 U11466 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7665), .ZN(n7703)
         );
  BUF_X1 U11467 ( .A(n11439), .Z(n29769) );
  AOI22_X1 U11468 ( .A1(n27754), .A2(\xmem_data[80][6] ), .B1(n30249), .B2(
        \xmem_data[81][6] ), .ZN(n7673) );
  BUF_X1 U11469 ( .A(n15525), .Z(n29808) );
  BUF_X1 U11470 ( .A(n3464), .Z(n29770) );
  AOI22_X1 U11471 ( .A1(n29808), .A2(\xmem_data[82][6] ), .B1(n31354), .B2(
        \xmem_data[83][6] ), .ZN(n7672) );
  AOI22_X1 U11472 ( .A1(n3168), .A2(\xmem_data[84][6] ), .B1(n3183), .B2(
        \xmem_data[85][6] ), .ZN(n7671) );
  AND2_X1 U11473 ( .A1(n28232), .A2(\xmem_data[87][6] ), .ZN(n7669) );
  AOI21_X1 U11474 ( .B1(n28755), .B2(\xmem_data[86][6] ), .A(n7669), .ZN(n7670) );
  NAND4_X1 U11475 ( .A1(n7673), .A2(n7672), .A3(n7671), .A4(n7670), .ZN(n7679)
         );
  AOI22_X1 U11476 ( .A1(n29604), .A2(\xmem_data[48][6] ), .B1(n29739), .B2(
        \xmem_data[49][6] ), .ZN(n7677) );
  AOI22_X1 U11477 ( .A1(n29771), .A2(\xmem_data[50][6] ), .B1(n29315), .B2(
        \xmem_data[51][6] ), .ZN(n7676) );
  AOI22_X1 U11478 ( .A1(n3163), .A2(\xmem_data[52][6] ), .B1(n3187), .B2(
        \xmem_data[53][6] ), .ZN(n7675) );
  BUF_X1 U11479 ( .A(n15549), .Z(n30310) );
  AOI22_X1 U11480 ( .A1(n30310), .A2(\xmem_data[54][6] ), .B1(n21008), .B2(
        \xmem_data[55][6] ), .ZN(n7674) );
  NAND4_X1 U11481 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n7678)
         );
  AOI22_X1 U11482 ( .A1(n29758), .A2(n7679), .B1(n7678), .B2(n29795), .ZN(
        n7701) );
  AOI22_X1 U11483 ( .A1(n30697), .A2(\xmem_data[72][6] ), .B1(n27833), .B2(
        \xmem_data[73][6] ), .ZN(n7683) );
  BUF_X1 U11484 ( .A(n14991), .Z(n29762) );
  AOI22_X1 U11485 ( .A1(n29707), .A2(\xmem_data[74][6] ), .B1(n29762), .B2(
        \xmem_data[75][6] ), .ZN(n7682) );
  AOI22_X1 U11486 ( .A1(n27703), .A2(\xmem_data[76][6] ), .B1(n29704), .B2(
        \xmem_data[77][6] ), .ZN(n7681) );
  AOI22_X1 U11487 ( .A1(n29763), .A2(\xmem_data[78][6] ), .B1(n30886), .B2(
        \xmem_data[79][6] ), .ZN(n7680) );
  NAND4_X1 U11488 ( .A1(n7683), .A2(n7682), .A3(n7681), .A4(n7680), .ZN(n7684)
         );
  NAND2_X1 U11489 ( .A1(n7684), .A2(n29758), .ZN(n7700) );
  AOI22_X1 U11490 ( .A1(n3166), .A2(\xmem_data[116][6] ), .B1(n3183), .B2(
        \xmem_data[117][6] ), .ZN(n7689) );
  BUF_X1 U11491 ( .A(n3464), .Z(n29807) );
  AOI22_X1 U11492 ( .A1(n29808), .A2(\xmem_data[114][6] ), .B1(n29807), .B2(
        \xmem_data[115][6] ), .ZN(n7688) );
  AOI22_X1 U11493 ( .A1(n29604), .A2(\xmem_data[112][6] ), .B1(n27753), .B2(
        \xmem_data[113][6] ), .ZN(n7687) );
  AND2_X1 U11494 ( .A1(n29439), .A2(\xmem_data[119][6] ), .ZN(n7685) );
  AOI21_X1 U11495 ( .B1(n30715), .B2(\xmem_data[118][6] ), .A(n7685), .ZN(
        n7686) );
  NAND4_X1 U11496 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .ZN(n7690)
         );
  NAND2_X1 U11497 ( .A1(n7690), .A2(n29837), .ZN(n7699) );
  BUF_X1 U11498 ( .A(n7691), .Z(n29695) );
  AOI22_X1 U11499 ( .A1(n29829), .A2(\xmem_data[0][6] ), .B1(n29695), .B2(
        \xmem_data[1][6] ), .ZN(n7696) );
  BUF_X1 U11500 ( .A(n7692), .Z(n29696) );
  AOI22_X1 U11501 ( .A1(n29696), .A2(\xmem_data[2][6] ), .B1(n3149), .B2(
        \xmem_data[3][6] ), .ZN(n7695) );
  AOI22_X1 U11502 ( .A1(n29626), .A2(\xmem_data[4][6] ), .B1(n30222), .B2(
        \xmem_data[5][6] ), .ZN(n7694) );
  BUF_X1 U11503 ( .A(n11451), .Z(n29699) );
  BUF_X1 U11504 ( .A(n14988), .Z(n29698) );
  AOI22_X1 U11505 ( .A1(n30279), .A2(\xmem_data[6][6] ), .B1(n29698), .B2(
        \xmem_data[7][6] ), .ZN(n7693) );
  NAND4_X1 U11506 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7693), .ZN(n7697)
         );
  NAND2_X1 U11507 ( .A1(n7697), .A2(n29733), .ZN(n7698) );
  NAND4_X1 U11508 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n7702)
         );
  XNOR2_X1 U11509 ( .A(n31817), .B(\fmem_data[19][3] ), .ZN(n30984) );
  XOR2_X1 U11510 ( .A(\fmem_data[19][2] ), .B(\fmem_data[19][3] ), .Z(n7705)
         );
  AOI22_X1 U11511 ( .A1(n29400), .A2(\xmem_data[40][7] ), .B1(n28208), .B2(
        \xmem_data[41][7] ), .ZN(n7709) );
  AOI22_X1 U11512 ( .A1(n29707), .A2(\xmem_data[42][7] ), .B1(n3375), .B2(
        \xmem_data[43][7] ), .ZN(n7708) );
  AOI22_X1 U11513 ( .A1(n29801), .A2(\xmem_data[44][7] ), .B1(n3369), .B2(
        \xmem_data[45][7] ), .ZN(n7707) );
  AOI22_X1 U11514 ( .A1(n29763), .A2(\xmem_data[46][7] ), .B1(n27514), .B2(
        \xmem_data[47][7] ), .ZN(n7706) );
  AOI22_X1 U11515 ( .A1(n29815), .A2(\xmem_data[56][7] ), .B1(n30685), .B2(
        \xmem_data[57][7] ), .ZN(n7713) );
  AOI22_X1 U11516 ( .A1(n3226), .A2(\xmem_data[58][7] ), .B1(n29816), .B2(
        \xmem_data[59][7] ), .ZN(n7712) );
  AOI22_X1 U11517 ( .A1(n29819), .A2(\xmem_data[60][7] ), .B1(n29818), .B2(
        \xmem_data[61][7] ), .ZN(n7711) );
  AOI22_X1 U11518 ( .A1(n29821), .A2(\xmem_data[62][7] ), .B1(n29820), .B2(
        \xmem_data[63][7] ), .ZN(n7710) );
  NAND4_X1 U11519 ( .A1(n7713), .A2(n7712), .A3(n7711), .A4(n7710), .ZN(n7719)
         );
  AOI22_X1 U11520 ( .A1(n28689), .A2(\xmem_data[54][7] ), .B1(n29639), .B2(
        \xmem_data[55][7] ), .ZN(n7717) );
  AOI22_X1 U11521 ( .A1(n28779), .A2(\xmem_data[48][7] ), .B1(n27753), .B2(
        \xmem_data[49][7] ), .ZN(n7716) );
  AOI22_X1 U11522 ( .A1(n3163), .A2(\xmem_data[52][7] ), .B1(n3186), .B2(
        \xmem_data[53][7] ), .ZN(n7715) );
  AOI22_X1 U11523 ( .A1(n29771), .A2(\xmem_data[50][7] ), .B1(n24213), .B2(
        \xmem_data[51][7] ), .ZN(n7714) );
  NAND4_X1 U11524 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), .ZN(n7718)
         );
  NOR2_X1 U11525 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  NAND2_X1 U11526 ( .A1(n7721), .A2(n7720), .ZN(n7727) );
  AOI22_X1 U11527 ( .A1(n28765), .A2(\xmem_data[32][7] ), .B1(n29785), .B2(
        \xmem_data[33][7] ), .ZN(n7725) );
  AOI22_X1 U11528 ( .A1(n29787), .A2(\xmem_data[34][7] ), .B1(n3348), .B2(
        \xmem_data[35][7] ), .ZN(n7724) );
  BUF_X2 U11529 ( .A(n7903), .Z(n28766) );
  AOI22_X1 U11530 ( .A1(n29626), .A2(\xmem_data[36][7] ), .B1(n28766), .B2(
        \xmem_data[37][7] ), .ZN(n7723) );
  AOI22_X1 U11531 ( .A1(n29628), .A2(\xmem_data[38][7] ), .B1(n29789), .B2(
        \xmem_data[39][7] ), .ZN(n7722) );
  NAND4_X1 U11532 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n7726)
         );
  OAI21_X1 U11533 ( .B1(n7727), .B2(n7726), .A(n29795), .ZN(n7796) );
  AOI22_X1 U11534 ( .A1(n29799), .A2(\xmem_data[104][7] ), .B1(n30776), .B2(
        \xmem_data[105][7] ), .ZN(n7731) );
  AOI22_X1 U11535 ( .A1(n29800), .A2(\xmem_data[106][7] ), .B1(n29706), .B2(
        \xmem_data[107][7] ), .ZN(n7730) );
  AOI22_X1 U11536 ( .A1(n28739), .A2(\xmem_data[108][7] ), .B1(n29482), .B2(
        \xmem_data[109][7] ), .ZN(n7729) );
  AOI22_X1 U11537 ( .A1(n29802), .A2(\xmem_data[110][7] ), .B1(n28743), .B2(
        \xmem_data[111][7] ), .ZN(n7728) );
  AOI22_X1 U11538 ( .A1(n27713), .A2(\xmem_data[120][7] ), .B1(n30266), .B2(
        \xmem_data[121][7] ), .ZN(n7735) );
  AOI22_X1 U11539 ( .A1(n29817), .A2(\xmem_data[122][7] ), .B1(n30311), .B2(
        \xmem_data[123][7] ), .ZN(n7734) );
  AOI22_X1 U11540 ( .A1(n29724), .A2(\xmem_data[124][7] ), .B1(n29723), .B2(
        \xmem_data[125][7] ), .ZN(n7733) );
  AOI22_X1 U11541 ( .A1(n29726), .A2(\xmem_data[126][7] ), .B1(n29725), .B2(
        \xmem_data[127][7] ), .ZN(n7732) );
  NAND4_X1 U11542 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7732), .ZN(n7741)
         );
  AOI22_X1 U11543 ( .A1(n27031), .A2(\xmem_data[118][7] ), .B1(n30950), .B2(
        \xmem_data[119][7] ), .ZN(n7739) );
  AOI22_X1 U11544 ( .A1(n3167), .A2(\xmem_data[116][7] ), .B1(n3182), .B2(
        \xmem_data[117][7] ), .ZN(n7738) );
  AOI22_X1 U11545 ( .A1(n30745), .A2(\xmem_data[112][7] ), .B1(n29648), .B2(
        \xmem_data[113][7] ), .ZN(n7737) );
  AOI22_X1 U11546 ( .A1(n29808), .A2(\xmem_data[114][7] ), .B1(n29807), .B2(
        \xmem_data[115][7] ), .ZN(n7736) );
  NAND4_X1 U11547 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n7740)
         );
  NOR2_X1 U11548 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  NAND2_X1 U11549 ( .A1(n3798), .A2(n7742), .ZN(n7748) );
  AOI22_X1 U11550 ( .A1(n29786), .A2(\xmem_data[96][7] ), .B1(n29695), .B2(
        \xmem_data[97][7] ), .ZN(n7746) );
  AOI22_X1 U11551 ( .A1(n29830), .A2(\xmem_data[98][7] ), .B1(n28164), .B2(
        \xmem_data[99][7] ), .ZN(n7745) );
  BUF_X2 U11552 ( .A(n11489), .Z(n29626) );
  AOI22_X1 U11553 ( .A1(n28136), .A2(\xmem_data[100][7] ), .B1(n30222), .B2(
        \xmem_data[101][7] ), .ZN(n7744) );
  AOI22_X1 U11554 ( .A1(n29423), .A2(\xmem_data[102][7] ), .B1(n29832), .B2(
        \xmem_data[103][7] ), .ZN(n7743) );
  NAND4_X1 U11555 ( .A1(n7746), .A2(n7745), .A3(n7744), .A4(n7743), .ZN(n7747)
         );
  OAI21_X1 U11556 ( .B1(n7748), .B2(n7747), .A(n29837), .ZN(n7795) );
  AOI22_X1 U11557 ( .A1(n30062), .A2(\xmem_data[86][7] ), .B1(n24115), .B2(
        \xmem_data[87][7] ), .ZN(n7752) );
  BUF_X1 U11558 ( .A(n8700), .Z(n29739) );
  AOI22_X1 U11559 ( .A1(n29604), .A2(\xmem_data[80][7] ), .B1(n29648), .B2(
        \xmem_data[81][7] ), .ZN(n7751) );
  AOI22_X1 U11560 ( .A1(n3161), .A2(\xmem_data[84][7] ), .B1(n3189), .B2(
        \xmem_data[85][7] ), .ZN(n7750) );
  AOI22_X1 U11561 ( .A1(n29771), .A2(\xmem_data[82][7] ), .B1(n27517), .B2(
        \xmem_data[83][7] ), .ZN(n7749) );
  NAND4_X1 U11562 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7758)
         );
  AOI22_X1 U11563 ( .A1(n30076), .A2(\xmem_data[88][7] ), .B1(n29640), .B2(
        \xmem_data[89][7] ), .ZN(n7756) );
  AOI22_X1 U11564 ( .A1(n3226), .A2(\xmem_data[90][7] ), .B1(n29816), .B2(
        \xmem_data[91][7] ), .ZN(n7755) );
  AOI22_X1 U11565 ( .A1(n29819), .A2(\xmem_data[92][7] ), .B1(n29818), .B2(
        \xmem_data[93][7] ), .ZN(n7754) );
  AOI22_X1 U11566 ( .A1(n29821), .A2(\xmem_data[94][7] ), .B1(n29820), .B2(
        \xmem_data[95][7] ), .ZN(n7753) );
  NAND4_X1 U11567 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n7757)
         );
  NOR2_X1 U11568 ( .A1(n7758), .A2(n7757), .ZN(n7764) );
  AOI22_X1 U11569 ( .A1(n27701), .A2(\xmem_data[72][7] ), .B1(n29495), .B2(
        \xmem_data[73][7] ), .ZN(n7762) );
  AOI22_X1 U11570 ( .A1(n29707), .A2(\xmem_data[74][7] ), .B1(n3375), .B2(
        \xmem_data[75][7] ), .ZN(n7761) );
  AOI22_X1 U11571 ( .A1(n28146), .A2(\xmem_data[76][7] ), .B1(n29589), .B2(
        \xmem_data[77][7] ), .ZN(n7760) );
  AOI22_X1 U11572 ( .A1(n29763), .A2(\xmem_data[78][7] ), .B1(n27944), .B2(
        \xmem_data[79][7] ), .ZN(n7759) );
  AND4_X1 U11573 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n7763)
         );
  NAND2_X1 U11574 ( .A1(n7764), .A2(n7763), .ZN(n7770) );
  AOI22_X1 U11575 ( .A1(n29786), .A2(\xmem_data[64][7] ), .B1(n29785), .B2(
        \xmem_data[65][7] ), .ZN(n7768) );
  AOI22_X1 U11576 ( .A1(n29787), .A2(\xmem_data[66][7] ), .B1(n3413), .B2(
        \xmem_data[67][7] ), .ZN(n7767) );
  AOI22_X1 U11577 ( .A1(n29421), .A2(\xmem_data[68][7] ), .B1(n29831), .B2(
        \xmem_data[69][7] ), .ZN(n7766) );
  AOI22_X1 U11578 ( .A1(n30279), .A2(\xmem_data[70][7] ), .B1(n29789), .B2(
        \xmem_data[71][7] ), .ZN(n7765) );
  NAND4_X1 U11579 ( .A1(n7768), .A2(n7767), .A3(n7766), .A4(n7765), .ZN(n7769)
         );
  OAI21_X1 U11580 ( .B1(n7770), .B2(n7769), .A(n29758), .ZN(n7794) );
  AOI22_X1 U11581 ( .A1(n28717), .A2(\xmem_data[0][7] ), .B1(n29695), .B2(
        \xmem_data[1][7] ), .ZN(n7774) );
  AOI22_X1 U11582 ( .A1(n29696), .A2(\xmem_data[2][7] ), .B1(n3433), .B2(
        \xmem_data[3][7] ), .ZN(n7773) );
  AOI22_X1 U11583 ( .A1(n27710), .A2(\xmem_data[4][7] ), .B1(n26510), .B2(
        \xmem_data[5][7] ), .ZN(n7772) );
  AOI22_X1 U11584 ( .A1(n28207), .A2(\xmem_data[6][7] ), .B1(n29698), .B2(
        \xmem_data[7][7] ), .ZN(n7771) );
  NAND4_X1 U11585 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .ZN(n7780)
         );
  AOI22_X1 U11586 ( .A1(n30777), .A2(\xmem_data[8][7] ), .B1(n29629), .B2(
        \xmem_data[9][7] ), .ZN(n7778) );
  AOI22_X1 U11587 ( .A1(n29707), .A2(\xmem_data[10][7] ), .B1(n29762), .B2(
        \xmem_data[11][7] ), .ZN(n7777) );
  AOI22_X1 U11588 ( .A1(n29602), .A2(\xmem_data[12][7] ), .B1(n30662), .B2(
        \xmem_data[13][7] ), .ZN(n7776) );
  AOI22_X1 U11589 ( .A1(n29709), .A2(\xmem_data[14][7] ), .B1(n23762), .B2(
        \xmem_data[15][7] ), .ZN(n7775) );
  NAND4_X1 U11590 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .ZN(n7779)
         );
  OR2_X1 U11591 ( .A1(n7780), .A2(n7779), .ZN(n7792) );
  AOI22_X1 U11592 ( .A1(n29610), .A2(\xmem_data[22][7] ), .B1(n29639), .B2(
        \xmem_data[23][7] ), .ZN(n7784) );
  AOI22_X1 U11593 ( .A1(n27811), .A2(\xmem_data[16][7] ), .B1(n27728), .B2(
        \xmem_data[17][7] ), .ZN(n7783) );
  AOI22_X1 U11594 ( .A1(n3164), .A2(\xmem_data[20][7] ), .B1(n3185), .B2(
        \xmem_data[21][7] ), .ZN(n7782) );
  AOI22_X1 U11595 ( .A1(n29808), .A2(\xmem_data[18][7] ), .B1(n30543), .B2(
        \xmem_data[19][7] ), .ZN(n7781) );
  NAND4_X1 U11596 ( .A1(n7784), .A2(n7783), .A3(n7782), .A4(n7781), .ZN(n7790)
         );
  AOI22_X1 U11597 ( .A1(n29363), .A2(\xmem_data[24][7] ), .B1(n30644), .B2(
        \xmem_data[25][7] ), .ZN(n7788) );
  AOI22_X1 U11598 ( .A1(n3226), .A2(\xmem_data[26][7] ), .B1(n29379), .B2(
        \xmem_data[27][7] ), .ZN(n7787) );
  AOI22_X1 U11599 ( .A1(n29777), .A2(\xmem_data[28][7] ), .B1(n29776), .B2(
        \xmem_data[29][7] ), .ZN(n7786) );
  AOI22_X1 U11600 ( .A1(n28681), .A2(\xmem_data[30][7] ), .B1(n20708), .B2(
        \xmem_data[31][7] ), .ZN(n7785) );
  NAND4_X1 U11601 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n7789)
         );
  OR2_X1 U11602 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  OAI21_X1 U11603 ( .B1(n7792), .B2(n7791), .A(n29733), .ZN(n7793) );
  XNOR2_X1 U11604 ( .A(n35270), .B(\fmem_data[19][3] ), .ZN(n30350) );
  OAI22_X1 U11605 ( .A1(n30984), .A2(n34474), .B1(n34472), .B2(n30350), .ZN(
        n34260) );
  AOI22_X1 U11606 ( .A1(n30635), .A2(\xmem_data[96][3] ), .B1(n30301), .B2(
        \xmem_data[97][3] ), .ZN(n7800) );
  AOI22_X1 U11607 ( .A1(n29397), .A2(\xmem_data[98][3] ), .B1(n30746), .B2(
        \xmem_data[99][3] ), .ZN(n7799) );
  AOI22_X1 U11608 ( .A1(n3164), .A2(\xmem_data[100][3] ), .B1(n3187), .B2(
        \xmem_data[101][3] ), .ZN(n7798) );
  AOI22_X1 U11609 ( .A1(n23901), .A2(\xmem_data[102][3] ), .B1(n29410), .B2(
        \xmem_data[103][3] ), .ZN(n7797) );
  NAND4_X1 U11610 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n7816)
         );
  AOI22_X1 U11611 ( .A1(n30766), .A2(\xmem_data[104][3] ), .B1(n29721), .B2(
        \xmem_data[105][3] ), .ZN(n7804) );
  AOI22_X1 U11612 ( .A1(n29380), .A2(\xmem_data[106][3] ), .B1(n29379), .B2(
        \xmem_data[107][3] ), .ZN(n7803) );
  AOI22_X1 U11613 ( .A1(n29382), .A2(\xmem_data[108][3] ), .B1(n29381), .B2(
        \xmem_data[109][3] ), .ZN(n7802) );
  AOI22_X1 U11614 ( .A1(n29384), .A2(\xmem_data[110][3] ), .B1(n29383), .B2(
        \xmem_data[111][3] ), .ZN(n7801) );
  NAND4_X1 U11615 ( .A1(n7804), .A2(n7803), .A3(n7802), .A4(n7801), .ZN(n7815)
         );
  AOI22_X1 U11616 ( .A1(n29419), .A2(\xmem_data[112][3] ), .B1(n29418), .B2(
        \xmem_data[113][3] ), .ZN(n7808) );
  AOI22_X1 U11617 ( .A1(n29420), .A2(\xmem_data[114][3] ), .B1(n29661), .B2(
        \xmem_data[115][3] ), .ZN(n7807) );
  AOI22_X1 U11618 ( .A1(n28734), .A2(\xmem_data[116][3] ), .B1(n26510), .B2(
        \xmem_data[117][3] ), .ZN(n7806) );
  AOI22_X1 U11619 ( .A1(n27740), .A2(\xmem_data[118][3] ), .B1(n29422), .B2(
        \xmem_data[119][3] ), .ZN(n7805) );
  NAND4_X1 U11620 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n7814)
         );
  AOI22_X1 U11621 ( .A1(n29400), .A2(\xmem_data[120][3] ), .B1(n3198), .B2(
        \xmem_data[121][3] ), .ZN(n7812) );
  AOI22_X1 U11622 ( .A1(n29402), .A2(\xmem_data[122][3] ), .B1(n3134), .B2(
        \xmem_data[123][3] ), .ZN(n7811) );
  AOI22_X1 U11623 ( .A1(n29590), .A2(\xmem_data[124][3] ), .B1(n28145), .B2(
        \xmem_data[125][3] ), .ZN(n7810) );
  AOI22_X1 U11624 ( .A1(n29404), .A2(\xmem_data[126][3] ), .B1(n29403), .B2(
        \xmem_data[127][3] ), .ZN(n7809) );
  NAND4_X1 U11625 ( .A1(n7812), .A2(n7811), .A3(n7810), .A4(n7809), .ZN(n7813)
         );
  OR4_X2 U11626 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n7838)
         );
  AOI22_X1 U11627 ( .A1(n29419), .A2(\xmem_data[80][3] ), .B1(n29418), .B2(
        \xmem_data[81][3] ), .ZN(n7820) );
  AOI22_X1 U11628 ( .A1(n29420), .A2(\xmem_data[82][3] ), .B1(n3351), .B2(
        \xmem_data[83][3] ), .ZN(n7819) );
  AOI22_X1 U11629 ( .A1(n29626), .A2(\xmem_data[84][3] ), .B1(n30695), .B2(
        \xmem_data[85][3] ), .ZN(n7818) );
  AOI22_X1 U11630 ( .A1(n29628), .A2(\xmem_data[86][3] ), .B1(n29422), .B2(
        \xmem_data[87][3] ), .ZN(n7817) );
  NAND4_X1 U11631 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n7836)
         );
  AOI22_X1 U11632 ( .A1(n30635), .A2(\xmem_data[64][3] ), .B1(n30634), .B2(
        \xmem_data[65][3] ), .ZN(n7824) );
  AOI22_X1 U11633 ( .A1(n29397), .A2(\xmem_data[66][3] ), .B1(n29437), .B2(
        \xmem_data[67][3] ), .ZN(n7823) );
  AOI22_X1 U11634 ( .A1(n3168), .A2(\xmem_data[68][3] ), .B1(n3187), .B2(
        \xmem_data[69][3] ), .ZN(n7822) );
  AOI22_X1 U11635 ( .A1(n26812), .A2(\xmem_data[70][3] ), .B1(n29410), .B2(
        \xmem_data[71][3] ), .ZN(n7821) );
  NAND4_X1 U11636 ( .A1(n7824), .A2(n7823), .A3(n7822), .A4(n7821), .ZN(n7835)
         );
  AOI22_X1 U11637 ( .A1(n28146), .A2(\xmem_data[92][3] ), .B1(n27761), .B2(
        \xmem_data[93][3] ), .ZN(n7828) );
  AOI22_X1 U11638 ( .A1(n29402), .A2(\xmem_data[90][3] ), .B1(n3135), .B2(
        \xmem_data[91][3] ), .ZN(n7827) );
  AOI22_X1 U11639 ( .A1(n29400), .A2(\xmem_data[88][3] ), .B1(n28786), .B2(
        \xmem_data[89][3] ), .ZN(n7826) );
  AOI22_X1 U11640 ( .A1(n29404), .A2(\xmem_data[94][3] ), .B1(n29403), .B2(
        \xmem_data[95][3] ), .ZN(n7825) );
  NAND4_X1 U11641 ( .A1(n7826), .A2(n7827), .A3(n7828), .A4(n7825), .ZN(n7834)
         );
  AOI22_X1 U11642 ( .A1(n29722), .A2(\xmem_data[72][3] ), .B1(n30716), .B2(
        \xmem_data[73][3] ), .ZN(n7832) );
  AOI22_X1 U11643 ( .A1(n29380), .A2(\xmem_data[74][3] ), .B1(n29379), .B2(
        \xmem_data[75][3] ), .ZN(n7831) );
  AOI22_X1 U11644 ( .A1(n29382), .A2(\xmem_data[76][3] ), .B1(n29381), .B2(
        \xmem_data[77][3] ), .ZN(n7830) );
  AOI22_X1 U11645 ( .A1(n29384), .A2(\xmem_data[78][3] ), .B1(n29383), .B2(
        \xmem_data[79][3] ), .ZN(n7829) );
  NAND4_X1 U11646 ( .A1(n7832), .A2(n7831), .A3(n7830), .A4(n7829), .ZN(n7833)
         );
  AOI22_X1 U11647 ( .A1(n29423), .A2(\xmem_data[54][3] ), .B1(n29431), .B2(
        \xmem_data[55][3] ), .ZN(n7844) );
  AOI22_X1 U11648 ( .A1(n29449), .A2(\xmem_data[50][3] ), .B1(n28245), .B2(
        \xmem_data[51][3] ), .ZN(n7841) );
  AOI22_X1 U11649 ( .A1(n29447), .A2(\xmem_data[48][3] ), .B1(n27812), .B2(
        \xmem_data[49][3] ), .ZN(n7840) );
  NAND2_X1 U11650 ( .A1(n29753), .A2(\xmem_data[53][3] ), .ZN(n7839) );
  AOI21_X1 U11651 ( .B1(n27710), .B2(\xmem_data[52][3] ), .A(n7842), .ZN(n7843) );
  AOI22_X1 U11652 ( .A1(n28173), .A2(\xmem_data[40][3] ), .B1(n30266), .B2(
        \xmem_data[41][3] ), .ZN(n7848) );
  AOI22_X1 U11653 ( .A1(n29461), .A2(\xmem_data[42][3] ), .B1(n3151), .B2(
        \xmem_data[43][3] ), .ZN(n7847) );
  AOI22_X1 U11654 ( .A1(n29463), .A2(\xmem_data[44][3] ), .B1(n29462), .B2(
        \xmem_data[45][3] ), .ZN(n7846) );
  AOI22_X1 U11655 ( .A1(n29464), .A2(\xmem_data[46][3] ), .B1(n30901), .B2(
        \xmem_data[47][3] ), .ZN(n7845) );
  NAND4_X1 U11656 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n7855)
         );
  AOI22_X1 U11657 ( .A1(n29566), .A2(\xmem_data[56][3] ), .B1(n29708), .B2(
        \xmem_data[57][3] ), .ZN(n7849) );
  INV_X1 U11658 ( .A(n7849), .ZN(n7854) );
  AOI22_X1 U11659 ( .A1(n28146), .A2(\xmem_data[60][3] ), .B1(n29482), .B2(
        \xmem_data[61][3] ), .ZN(n7852) );
  AOI22_X1 U11660 ( .A1(n29500), .A2(\xmem_data[62][3] ), .B1(n29451), .B2(
        \xmem_data[63][3] ), .ZN(n7851) );
  AOI22_X1 U11661 ( .A1(n29450), .A2(\xmem_data[58][3] ), .B1(n3345), .B2(
        \xmem_data[59][3] ), .ZN(n7850) );
  NAND3_X1 U11662 ( .A1(n7852), .A2(n7851), .A3(n7850), .ZN(n7853) );
  NOR3_X1 U11663 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(n7860) );
  AOI22_X1 U11664 ( .A1(n27811), .A2(\xmem_data[32][3] ), .B1(n26884), .B2(
        \xmem_data[33][3] ), .ZN(n7859) );
  AOI22_X1 U11665 ( .A1(n29438), .A2(\xmem_data[34][3] ), .B1(n17018), .B2(
        \xmem_data[35][3] ), .ZN(n7858) );
  AOI22_X1 U11666 ( .A1(n3166), .A2(\xmem_data[36][3] ), .B1(n3189), .B2(
        \xmem_data[37][3] ), .ZN(n7857) );
  AOI22_X1 U11667 ( .A1(n28755), .A2(\xmem_data[38][3] ), .B1(n29439), .B2(
        \xmem_data[39][3] ), .ZN(n7856) );
  NAND3_X1 U11668 ( .A1(n3934), .A2(n7860), .A3(n3524), .ZN(n7882) );
  AOI22_X1 U11669 ( .A1(n28751), .A2(\xmem_data[0][3] ), .B1(n27728), .B2(
        \xmem_data[1][3] ), .ZN(n7864) );
  AOI22_X1 U11670 ( .A1(n29475), .A2(\xmem_data[2][3] ), .B1(n3120), .B2(
        \xmem_data[3][3] ), .ZN(n7863) );
  AOI22_X1 U11671 ( .A1(n3167), .A2(\xmem_data[4][3] ), .B1(n3189), .B2(
        \xmem_data[5][3] ), .ZN(n7862) );
  AOI22_X1 U11672 ( .A1(n26812), .A2(\xmem_data[6][3] ), .B1(n28232), .B2(
        \xmem_data[7][3] ), .ZN(n7861) );
  AND4_X1 U11673 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7880)
         );
  AOI22_X1 U11674 ( .A1(n29363), .A2(\xmem_data[8][3] ), .B1(n30765), .B2(
        \xmem_data[9][3] ), .ZN(n7868) );
  AOI22_X1 U11675 ( .A1(n7270), .A2(\xmem_data[10][3] ), .B1(n30311), .B2(
        \xmem_data[11][3] ), .ZN(n7867) );
  AOI22_X1 U11676 ( .A1(n28725), .A2(\xmem_data[12][3] ), .B1(n27805), .B2(
        \xmem_data[13][3] ), .ZN(n7866) );
  AOI22_X1 U11677 ( .A1(n29489), .A2(\xmem_data[14][3] ), .B1(n31345), .B2(
        \xmem_data[15][3] ), .ZN(n7865) );
  AND4_X1 U11678 ( .A1(n7868), .A2(n7867), .A3(n7866), .A4(n7865), .ZN(n7879)
         );
  AOI22_X1 U11679 ( .A1(n29829), .A2(\xmem_data[16][3] ), .B1(n29497), .B2(
        \xmem_data[17][3] ), .ZN(n7872) );
  AOI22_X1 U11680 ( .A1(n29499), .A2(\xmem_data[18][3] ), .B1(n28164), .B2(
        \xmem_data[19][3] ), .ZN(n7871) );
  AOI22_X1 U11681 ( .A1(n29788), .A2(\xmem_data[20][3] ), .B1(n30707), .B2(
        \xmem_data[21][3] ), .ZN(n7870) );
  AOI22_X1 U11682 ( .A1(n28138), .A2(\xmem_data[22][3] ), .B1(n29494), .B2(
        \xmem_data[23][3] ), .ZN(n7869) );
  AND4_X1 U11683 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n7878)
         );
  AOI22_X1 U11684 ( .A1(n30294), .A2(\xmem_data[24][3] ), .B1(n28208), .B2(
        \xmem_data[25][3] ), .ZN(n7876) );
  AOI22_X1 U11685 ( .A1(n29501), .A2(\xmem_data[26][3] ), .B1(n3134), .B2(
        \xmem_data[27][3] ), .ZN(n7875) );
  AOI22_X1 U11686 ( .A1(n30633), .A2(\xmem_data[28][3] ), .B1(n29704), .B2(
        \xmem_data[29][3] ), .ZN(n7874) );
  AOI22_X1 U11687 ( .A1(n29500), .A2(\xmem_data[30][3] ), .B1(n30083), .B2(
        \xmem_data[31][3] ), .ZN(n7873) );
  AND4_X1 U11688 ( .A1(n7876), .A2(n7875), .A3(n7874), .A4(n7873), .ZN(n7877)
         );
  NAND4_X1 U11689 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n7881)
         );
  XNOR2_X1 U11690 ( .A(n3450), .B(\fmem_data[3][7] ), .ZN(n31983) );
  AOI22_X1 U11691 ( .A1(n29400), .A2(\xmem_data[88][2] ), .B1(n29556), .B2(
        \xmem_data[89][2] ), .ZN(n7883) );
  INV_X1 U11692 ( .A(n7883), .ZN(n7893) );
  AOI22_X1 U11693 ( .A1(n30248), .A2(\xmem_data[92][2] ), .B1(n28665), .B2(
        \xmem_data[93][2] ), .ZN(n7891) );
  AOI22_X1 U11694 ( .A1(n29419), .A2(\xmem_data[80][2] ), .B1(n29418), .B2(
        \xmem_data[81][2] ), .ZN(n7884) );
  INV_X1 U11695 ( .A(n7884), .ZN(n7889) );
  AOI22_X1 U11696 ( .A1(n29420), .A2(\xmem_data[82][2] ), .B1(n24693), .B2(
        \xmem_data[83][2] ), .ZN(n7887) );
  AOI22_X1 U11697 ( .A1(n29404), .A2(\xmem_data[94][2] ), .B1(n29403), .B2(
        \xmem_data[95][2] ), .ZN(n7886) );
  AOI22_X1 U11698 ( .A1(n29402), .A2(\xmem_data[90][2] ), .B1(n3134), .B2(
        \xmem_data[91][2] ), .ZN(n7885) );
  NOR2_X1 U11699 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U11700 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NOR2_X1 U11701 ( .A1(n7893), .A2(n7892), .ZN(n7910) );
  AOI22_X1 U11702 ( .A1(n27754), .A2(\xmem_data[64][2] ), .B1(n30301), .B2(
        \xmem_data[65][2] ), .ZN(n7898) );
  AOI22_X1 U11703 ( .A1(n29397), .A2(\xmem_data[66][2] ), .B1(n30543), .B2(
        \xmem_data[67][2] ), .ZN(n7897) );
  AOI22_X1 U11704 ( .A1(n3161), .A2(\xmem_data[68][2] ), .B1(n3190), .B2(
        \xmem_data[69][2] ), .ZN(n7896) );
  AND2_X1 U11705 ( .A1(n29410), .A2(\xmem_data[71][2] ), .ZN(n7894) );
  AOI21_X1 U11706 ( .B1(n30070), .B2(\xmem_data[70][2] ), .A(n7894), .ZN(n7895) );
  BUF_X1 U11707 ( .A(n10802), .Z(n29488) );
  AOI22_X1 U11708 ( .A1(n28680), .A2(\xmem_data[72][2] ), .B1(n29640), .B2(
        \xmem_data[73][2] ), .ZN(n7902) );
  AOI22_X1 U11709 ( .A1(n29380), .A2(\xmem_data[74][2] ), .B1(n29379), .B2(
        \xmem_data[75][2] ), .ZN(n7901) );
  AOI22_X1 U11710 ( .A1(n29382), .A2(\xmem_data[76][2] ), .B1(n29381), .B2(
        \xmem_data[77][2] ), .ZN(n7900) );
  AOI22_X1 U11711 ( .A1(n29384), .A2(\xmem_data[78][2] ), .B1(n29383), .B2(
        \xmem_data[79][2] ), .ZN(n7899) );
  AND2_X1 U11712 ( .A1(n28700), .A2(\xmem_data[86][2] ), .ZN(n7908) );
  NAND2_X1 U11713 ( .A1(n29831), .A2(\xmem_data[85][2] ), .ZN(n7905) );
  NAND2_X1 U11714 ( .A1(n29422), .A2(\xmem_data[87][2] ), .ZN(n7904) );
  NAND2_X1 U11715 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  NOR3_X1 U11716 ( .A1(n7908), .A2(n7907), .A3(n7906), .ZN(n7909) );
  NAND4_X1 U11717 ( .A1(n7910), .A2(n3812), .A3(n3518), .A4(n7909), .ZN(n7911)
         );
  NAND2_X1 U11718 ( .A1(n7911), .A2(n29376), .ZN(n7990) );
  NAND2_X1 U11719 ( .A1(n29629), .A2(\xmem_data[57][2] ), .ZN(n7913) );
  NAND2_X1 U11720 ( .A1(n28740), .A2(\xmem_data[56][2] ), .ZN(n7912) );
  NAND2_X1 U11721 ( .A1(n7913), .A2(n7912), .ZN(n7923) );
  AOI22_X1 U11722 ( .A1(n28146), .A2(\xmem_data[60][2] ), .B1(n30730), .B2(
        \xmem_data[61][2] ), .ZN(n7921) );
  AOI22_X1 U11723 ( .A1(n29447), .A2(\xmem_data[48][2] ), .B1(n27743), .B2(
        \xmem_data[49][2] ), .ZN(n7914) );
  INV_X1 U11724 ( .A(n7914), .ZN(n7919) );
  AOI22_X1 U11725 ( .A1(n29449), .A2(\xmem_data[50][2] ), .B1(n3351), .B2(
        \xmem_data[51][2] ), .ZN(n7917) );
  AOI22_X1 U11726 ( .A1(n7282), .A2(\xmem_data[62][2] ), .B1(n29451), .B2(
        \xmem_data[63][2] ), .ZN(n7916) );
  AOI22_X1 U11727 ( .A1(n29450), .A2(\xmem_data[58][2] ), .B1(n3134), .B2(
        \xmem_data[59][2] ), .ZN(n7915) );
  NOR2_X1 U11728 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U11729 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  NOR2_X1 U11730 ( .A1(n7923), .A2(n7922), .ZN(n7935) );
  AOI22_X1 U11731 ( .A1(n29363), .A2(\xmem_data[40][2] ), .B1(n30644), .B2(
        \xmem_data[41][2] ), .ZN(n7927) );
  AOI22_X1 U11732 ( .A1(n29461), .A2(\xmem_data[42][2] ), .B1(n3151), .B2(
        \xmem_data[43][2] ), .ZN(n7926) );
  AOI22_X1 U11733 ( .A1(n29463), .A2(\xmem_data[44][2] ), .B1(n29462), .B2(
        \xmem_data[45][2] ), .ZN(n7925) );
  AOI22_X1 U11734 ( .A1(n29464), .A2(\xmem_data[46][2] ), .B1(n30901), .B2(
        \xmem_data[47][2] ), .ZN(n7924) );
  AOI22_X1 U11735 ( .A1(n30745), .A2(\xmem_data[32][2] ), .B1(n29648), .B2(
        \xmem_data[33][2] ), .ZN(n7931) );
  AOI22_X1 U11736 ( .A1(n29438), .A2(\xmem_data[34][2] ), .B1(n28516), .B2(
        \xmem_data[35][2] ), .ZN(n7930) );
  AOI22_X1 U11737 ( .A1(n3163), .A2(\xmem_data[36][2] ), .B1(n3188), .B2(
        \xmem_data[37][2] ), .ZN(n7929) );
  BUF_X1 U11738 ( .A(n15549), .Z(n30684) );
  AOI22_X1 U11739 ( .A1(n30684), .A2(\xmem_data[38][2] ), .B1(n29439), .B2(
        \xmem_data[39][2] ), .ZN(n7928) );
  AOI22_X1 U11740 ( .A1(n29628), .A2(\xmem_data[54][2] ), .B1(n29431), .B2(
        \xmem_data[55][2] ), .ZN(n7933) );
  AOI22_X1 U11741 ( .A1(n29788), .A2(\xmem_data[52][2] ), .B1(n29831), .B2(
        \xmem_data[53][2] ), .ZN(n7932) );
  NAND4_X1 U11742 ( .A1(n7935), .A2(n3813), .A3(n3519), .A4(n7934), .ZN(n7936)
         );
  NAND2_X1 U11743 ( .A1(n7936), .A2(n29471), .ZN(n7989) );
  AOI22_X1 U11744 ( .A1(n27754), .A2(\xmem_data[96][2] ), .B1(n30634), .B2(
        \xmem_data[97][2] ), .ZN(n7940) );
  AOI22_X1 U11745 ( .A1(n29397), .A2(\xmem_data[98][2] ), .B1(n25461), .B2(
        \xmem_data[99][2] ), .ZN(n7939) );
  AOI22_X1 U11746 ( .A1(n3168), .A2(\xmem_data[100][2] ), .B1(n3182), .B2(
        \xmem_data[101][2] ), .ZN(n7938) );
  AOI22_X1 U11747 ( .A1(n23901), .A2(\xmem_data[102][2] ), .B1(n29410), .B2(
        \xmem_data[103][2] ), .ZN(n7937) );
  AOI22_X1 U11748 ( .A1(n29400), .A2(\xmem_data[120][2] ), .B1(n29761), .B2(
        \xmem_data[121][2] ), .ZN(n7941) );
  INV_X1 U11749 ( .A(n7941), .ZN(n7951) );
  AOI22_X1 U11750 ( .A1(n30633), .A2(\xmem_data[124][2] ), .B1(n3369), .B2(
        \xmem_data[125][2] ), .ZN(n7949) );
  AOI22_X1 U11751 ( .A1(n29419), .A2(\xmem_data[112][2] ), .B1(n29418), .B2(
        \xmem_data[113][2] ), .ZN(n7942) );
  INV_X1 U11752 ( .A(n7942), .ZN(n7947) );
  AOI22_X1 U11753 ( .A1(n29420), .A2(\xmem_data[114][2] ), .B1(n23732), .B2(
        \xmem_data[115][2] ), .ZN(n7945) );
  AOI22_X1 U11754 ( .A1(n29404), .A2(\xmem_data[126][2] ), .B1(n29403), .B2(
        \xmem_data[127][2] ), .ZN(n7944) );
  AOI22_X1 U11755 ( .A1(n29402), .A2(\xmem_data[122][2] ), .B1(n29350), .B2(
        \xmem_data[123][2] ), .ZN(n7943) );
  NAND3_X1 U11756 ( .A1(n7945), .A2(n7944), .A3(n7943), .ZN(n7946) );
  NOR2_X1 U11757 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  NAND2_X1 U11758 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  NOR2_X1 U11759 ( .A1(n7951), .A2(n7950), .ZN(n7962) );
  AOI22_X1 U11760 ( .A1(n30063), .A2(\xmem_data[104][2] ), .B1(n30685), .B2(
        \xmem_data[105][2] ), .ZN(n7955) );
  AOI22_X1 U11761 ( .A1(n29380), .A2(\xmem_data[106][2] ), .B1(n29379), .B2(
        \xmem_data[107][2] ), .ZN(n7954) );
  AOI22_X1 U11762 ( .A1(n29382), .A2(\xmem_data[108][2] ), .B1(n29381), .B2(
        \xmem_data[109][2] ), .ZN(n7953) );
  AOI22_X1 U11763 ( .A1(n29384), .A2(\xmem_data[110][2] ), .B1(n29383), .B2(
        \xmem_data[111][2] ), .ZN(n7952) );
  AND2_X1 U11764 ( .A1(n3392), .A2(\xmem_data[118][2] ), .ZN(n7960) );
  NAND2_X1 U11765 ( .A1(n28766), .A2(\xmem_data[117][2] ), .ZN(n7957) );
  NAND2_X1 U11766 ( .A1(n29422), .A2(\xmem_data[119][2] ), .ZN(n7956) );
  NAND2_X1 U11767 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NOR3_X1 U11768 ( .A1(n7960), .A2(n7959), .A3(n7958), .ZN(n7961) );
  NAND4_X1 U11769 ( .A1(n3842), .A2(n7962), .A3(n3520), .A4(n7961), .ZN(n7963)
         );
  NAND2_X1 U11770 ( .A1(n7963), .A2(n29428), .ZN(n7988) );
  AOI22_X1 U11771 ( .A1(n28717), .A2(\xmem_data[16][2] ), .B1(n29497), .B2(
        \xmem_data[17][2] ), .ZN(n7967) );
  AOI22_X1 U11772 ( .A1(n29499), .A2(\xmem_data[18][2] ), .B1(n3153), .B2(
        \xmem_data[19][2] ), .ZN(n7966) );
  AOI22_X1 U11773 ( .A1(n27741), .A2(\xmem_data[20][2] ), .B1(n30182), .B2(
        \xmem_data[21][2] ), .ZN(n7965) );
  AOI22_X1 U11774 ( .A1(n28700), .A2(\xmem_data[22][2] ), .B1(n29494), .B2(
        \xmem_data[23][2] ), .ZN(n7964) );
  AOI22_X1 U11775 ( .A1(n30633), .A2(\xmem_data[28][2] ), .B1(n28665), .B2(
        \xmem_data[29][2] ), .ZN(n7985) );
  AOI22_X1 U11776 ( .A1(n27771), .A2(\xmem_data[24][2] ), .B1(n28667), .B2(
        \xmem_data[25][2] ), .ZN(n7968) );
  INV_X1 U11777 ( .A(n7968), .ZN(n7972) );
  AOI22_X1 U11778 ( .A1(n29501), .A2(\xmem_data[26][2] ), .B1(n29350), .B2(
        \xmem_data[27][2] ), .ZN(n7970) );
  AOI22_X1 U11779 ( .A1(n29500), .A2(\xmem_data[30][2] ), .B1(n28152), .B2(
        \xmem_data[31][2] ), .ZN(n7969) );
  NAND2_X1 U11780 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  NOR2_X1 U11781 ( .A1(n7972), .A2(n7971), .ZN(n7984) );
  AOI22_X1 U11782 ( .A1(n30302), .A2(\xmem_data[0][2] ), .B1(n30634), .B2(
        \xmem_data[1][2] ), .ZN(n7976) );
  AOI22_X1 U11783 ( .A1(n29438), .A2(\xmem_data[2][2] ), .B1(n3465), .B2(
        \xmem_data[3][2] ), .ZN(n7975) );
  AOI22_X1 U11784 ( .A1(n3168), .A2(\xmem_data[4][2] ), .B1(n3184), .B2(
        \xmem_data[5][2] ), .ZN(n7974) );
  AOI22_X1 U11785 ( .A1(n27031), .A2(\xmem_data[6][2] ), .B1(n29639), .B2(
        \xmem_data[7][2] ), .ZN(n7973) );
  NAND4_X1 U11786 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n7982)
         );
  AOI22_X1 U11787 ( .A1(n30766), .A2(\xmem_data[8][2] ), .B1(n29640), .B2(
        \xmem_data[9][2] ), .ZN(n7980) );
  AOI22_X1 U11788 ( .A1(n7270), .A2(\xmem_data[10][2] ), .B1(n29379), .B2(
        \xmem_data[11][2] ), .ZN(n7979) );
  AOI22_X1 U11789 ( .A1(n28725), .A2(\xmem_data[12][2] ), .B1(n29723), .B2(
        \xmem_data[13][2] ), .ZN(n7978) );
  AOI22_X1 U11790 ( .A1(n29489), .A2(\xmem_data[14][2] ), .B1(n28772), .B2(
        \xmem_data[15][2] ), .ZN(n7977) );
  NAND4_X1 U11791 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n7981)
         );
  NOR2_X1 U11792 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  NAND4_X1 U11793 ( .A1(n3860), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n7986)
         );
  NAND2_X1 U11794 ( .A1(n7986), .A2(n29511), .ZN(n7987) );
  XNOR2_X1 U11795 ( .A(n33720), .B(\fmem_data[3][7] ), .ZN(n30407) );
  XOR2_X1 U11796 ( .A(\fmem_data[3][6] ), .B(\fmem_data[3][7] ), .Z(n7991) );
  OAI22_X1 U11797 ( .A1(n31983), .A2(n35638), .B1(n30407), .B2(n35637), .ZN(
        n34259) );
  BUF_X1 U11798 ( .A(n11436), .Z(n28739) );
  BUF_X1 U11799 ( .A(n11437), .Z(n28738) );
  AOI22_X1 U11800 ( .A1(n30248), .A2(\xmem_data[100][5] ), .B1(n28145), .B2(
        \xmem_data[101][5] ), .ZN(n7999) );
  BUF_X1 U11801 ( .A(n11484), .Z(n28740) );
  AOI22_X1 U11802 ( .A1(n28740), .A2(\xmem_data[96][5] ), .B1(n27833), .B2(
        \xmem_data[97][5] ), .ZN(n7998) );
  NAND3_X1 U11803 ( .A1(n11343), .A2(n11342), .A3(n6173), .ZN(n8011) );
  NOR2_X1 U11804 ( .A1(n3447), .A2(n8011), .ZN(n8080) );
  BUF_X1 U11805 ( .A(n14991), .Z(n28741) );
  AOI22_X1 U11806 ( .A1(n3244), .A2(\xmem_data[98][5] ), .B1(n3126), .B2(
        \xmem_data[99][5] ), .ZN(n7992) );
  NOR2_X1 U11807 ( .A1(n3445), .A2(n11360), .ZN(n8081) );
  BUF_X2 U11808 ( .A(n8081), .Z(n28744) );
  BUF_X1 U11809 ( .A(n14997), .Z(n28743) );
  AOI22_X1 U11810 ( .A1(n28744), .A2(\xmem_data[102][5] ), .B1(n28743), .B2(
        \xmem_data[103][5] ), .ZN(n7994) );
  NAND3_X1 U11811 ( .A1(n7999), .A2(n7998), .A3(n7997), .ZN(n8019) );
  BUF_X1 U11812 ( .A(n11439), .Z(n28751) );
  AOI22_X1 U11813 ( .A1(n30302), .A2(\xmem_data[104][5] ), .B1(n29592), .B2(
        \xmem_data[105][5] ), .ZN(n8004) );
  NOR2_X1 U11814 ( .A1(n8000), .A2(n8011), .ZN(n28780) );
  BUF_X1 U11815 ( .A(n28780), .Z(n28753) );
  BUF_X1 U11816 ( .A(n29187), .Z(n28752) );
  AOI22_X1 U11817 ( .A1(n28753), .A2(\xmem_data[106][5] ), .B1(n28154), .B2(
        \xmem_data[107][5] ), .ZN(n8003) );
  AOI22_X1 U11818 ( .A1(n3163), .A2(\xmem_data[108][5] ), .B1(n3187), .B2(
        \xmem_data[109][5] ), .ZN(n8002) );
  BUF_X1 U11819 ( .A(n14971), .Z(n28781) );
  AOI22_X1 U11820 ( .A1(n29716), .A2(\xmem_data[110][5] ), .B1(n28781), .B2(
        \xmem_data[111][5] ), .ZN(n8001) );
  NAND4_X1 U11821 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n8018)
         );
  AOI22_X1 U11822 ( .A1(n28173), .A2(\xmem_data[112][5] ), .B1(n30170), .B2(
        \xmem_data[113][5] ), .ZN(n8009) );
  NOR2_X1 U11823 ( .A1(n8011), .A2(n8005), .ZN(n8072) );
  BUF_X1 U11824 ( .A(n8072), .Z(n28720) );
  AOI22_X1 U11825 ( .A1(n28720), .A2(\xmem_data[114][5] ), .B1(n3330), .B2(
        \xmem_data[115][5] ), .ZN(n8008) );
  BUF_X1 U11826 ( .A(n8074), .Z(n28724) );
  AOI22_X1 U11827 ( .A1(n28725), .A2(\xmem_data[116][5] ), .B1(n28724), .B2(
        \xmem_data[117][5] ), .ZN(n8007) );
  BUF_X1 U11828 ( .A(n8075), .Z(n28727) );
  AOI22_X1 U11829 ( .A1(n28727), .A2(\xmem_data[118][5] ), .B1(n30901), .B2(
        \xmem_data[119][5] ), .ZN(n8006) );
  NAND4_X1 U11830 ( .A1(n8009), .A2(n8008), .A3(n8007), .A4(n8006), .ZN(n8017)
         );
  BUF_X1 U11831 ( .A(n8088), .Z(n28717) );
  NOR2_X1 U11832 ( .A1(n3246), .A2(n8010), .ZN(n8089) );
  AOI22_X1 U11833 ( .A1(n29786), .A2(\xmem_data[120][5] ), .B1(n3124), .B2(
        \xmem_data[121][5] ), .ZN(n8015) );
  NOR2_X1 U11834 ( .A1(n8011), .A2(n8010), .ZN(n8090) );
  BUF_X1 U11835 ( .A(n8090), .Z(n28719) );
  BUF_X1 U11836 ( .A(n28973), .Z(n28718) );
  AOI22_X1 U11837 ( .A1(n28719), .A2(\xmem_data[122][5] ), .B1(n28718), .B2(
        \xmem_data[123][5] ), .ZN(n8014) );
  BUF_X2 U11838 ( .A(n11489), .Z(n28734) );
  AOI22_X1 U11839 ( .A1(n30223), .A2(\xmem_data[124][5] ), .B1(n30290), .B2(
        \xmem_data[125][5] ), .ZN(n8013) );
  BUF_X1 U11840 ( .A(n14988), .Z(n28733) );
  AOI22_X1 U11841 ( .A1(n29628), .A2(\xmem_data[126][5] ), .B1(n28733), .B2(
        \xmem_data[127][5] ), .ZN(n8012) );
  NAND4_X1 U11842 ( .A1(n8015), .A2(n8014), .A3(n8013), .A4(n8012), .ZN(n8016)
         );
  NOR2_X1 U11843 ( .A1(n39041), .A2(n3444), .ZN(n8021) );
  AOI21_X1 U11844 ( .B1(n4499), .B2(n3444), .A(n8021), .ZN(n8067) );
  XOR2_X1 U11845 ( .A(n8021), .B(load_xaddr_val[6]), .Z(n8066) );
  AND2_X1 U11846 ( .A1(n8067), .A2(n8066), .ZN(n28762) );
  INV_X1 U11847 ( .A(n8066), .ZN(n8045) );
  BUF_X1 U11848 ( .A(n11780), .Z(n28667) );
  AOI22_X1 U11849 ( .A1(n28740), .A2(\xmem_data[64][5] ), .B1(n28667), .B2(
        \xmem_data[65][5] ), .ZN(n8025) );
  BUF_X1 U11850 ( .A(n8080), .Z(n28670) );
  AOI22_X1 U11851 ( .A1(n28670), .A2(\xmem_data[66][5] ), .B1(n3140), .B2(
        \xmem_data[67][5] ), .ZN(n8024) );
  BUF_X2 U11852 ( .A(n11437), .Z(n28665) );
  AOI22_X1 U11853 ( .A1(n29801), .A2(\xmem_data[68][5] ), .B1(n28238), .B2(
        \xmem_data[69][5] ), .ZN(n8023) );
  BUF_X1 U11854 ( .A(n14997), .Z(n28671) );
  AOI22_X1 U11855 ( .A1(n28744), .A2(\xmem_data[70][5] ), .B1(n28671), .B2(
        \xmem_data[71][5] ), .ZN(n8022) );
  NAND4_X1 U11856 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), .ZN(n8042)
         );
  BUF_X1 U11857 ( .A(n11439), .Z(n28685) );
  AOI22_X1 U11858 ( .A1(n28751), .A2(\xmem_data[72][5] ), .B1(n30237), .B2(
        \xmem_data[73][5] ), .ZN(n8030) );
  BUF_X1 U11859 ( .A(n28780), .Z(n28686) );
  AOI22_X1 U11860 ( .A1(n28686), .A2(\xmem_data[74][5] ), .B1(n24213), .B2(
        \xmem_data[75][5] ), .ZN(n8029) );
  AOI22_X1 U11861 ( .A1(n3165), .A2(\xmem_data[76][5] ), .B1(n3189), .B2(
        \xmem_data[77][5] ), .ZN(n8028) );
  BUF_X1 U11862 ( .A(n14971), .Z(n28687) );
  AND2_X1 U11863 ( .A1(n28687), .A2(\xmem_data[79][5] ), .ZN(n8026) );
  AOI21_X1 U11864 ( .B1(n29610), .B2(\xmem_data[78][5] ), .A(n8026), .ZN(n8027) );
  NAND4_X1 U11865 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n8041)
         );
  AOI22_X1 U11866 ( .A1(n29786), .A2(\xmem_data[88][5] ), .B1(n29418), .B2(
        \xmem_data[89][5] ), .ZN(n8034) );
  BUF_X1 U11867 ( .A(n28973), .Z(n28677) );
  AOI22_X1 U11868 ( .A1(n3227), .A2(\xmem_data[90][5] ), .B1(n28677), .B2(
        \xmem_data[91][5] ), .ZN(n8033) );
  AOI22_X1 U11869 ( .A1(n29421), .A2(\xmem_data[92][5] ), .B1(n30654), .B2(
        \xmem_data[93][5] ), .ZN(n8032) );
  BUF_X2 U11870 ( .A(n11451), .Z(n28700) );
  AOI22_X1 U11871 ( .A1(n30215), .A2(\xmem_data[94][5] ), .B1(n29832), .B2(
        \xmem_data[95][5] ), .ZN(n8031) );
  NAND4_X1 U11872 ( .A1(n8032), .A2(n8033), .A3(n8034), .A4(n8031), .ZN(n8040)
         );
  AOI22_X1 U11873 ( .A1(n30766), .A2(\xmem_data[80][5] ), .B1(n29487), .B2(
        \xmem_data[81][5] ), .ZN(n8038) );
  BUF_X1 U11874 ( .A(n14974), .Z(n28701) );
  AOI22_X1 U11875 ( .A1(n28702), .A2(\xmem_data[82][5] ), .B1(n28701), .B2(
        \xmem_data[83][5] ), .ZN(n8037) );
  BUF_X1 U11876 ( .A(n8074), .Z(n28696) );
  AOI22_X1 U11877 ( .A1(n28725), .A2(\xmem_data[84][5] ), .B1(n28696), .B2(
        \xmem_data[85][5] ), .ZN(n8036) );
  AOI22_X1 U11878 ( .A1(n28681), .A2(\xmem_data[86][5] ), .B1(n28192), .B2(
        \xmem_data[87][5] ), .ZN(n8035) );
  NAND4_X1 U11879 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8039)
         );
  AND2_X1 U11880 ( .A1(n8045), .A2(n8067), .ZN(n28713) );
  AOI22_X1 U11881 ( .A1(n27834), .A2(\xmem_data[32][5] ), .B1(n30293), .B2(
        \xmem_data[33][5] ), .ZN(n8049) );
  AOI22_X1 U11882 ( .A1(n28670), .A2(\xmem_data[34][5] ), .B1(n28308), .B2(
        \xmem_data[35][5] ), .ZN(n8048) );
  AOI22_X1 U11883 ( .A1(n3249), .A2(\xmem_data[36][5] ), .B1(n29646), .B2(
        \xmem_data[37][5] ), .ZN(n8047) );
  AOI22_X1 U11884 ( .A1(n28744), .A2(\xmem_data[38][5] ), .B1(n28671), .B2(
        \xmem_data[39][5] ), .ZN(n8046) );
  NAND4_X1 U11885 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n8065)
         );
  AOI22_X1 U11886 ( .A1(n29395), .A2(\xmem_data[40][5] ), .B1(n30084), .B2(
        \xmem_data[41][5] ), .ZN(n8053) );
  AOI22_X1 U11887 ( .A1(n28686), .A2(\xmem_data[42][5] ), .B1(n20718), .B2(
        \xmem_data[43][5] ), .ZN(n8052) );
  AOI22_X1 U11888 ( .A1(n3161), .A2(\xmem_data[44][5] ), .B1(n11426), .B2(
        \xmem_data[45][5] ), .ZN(n8051) );
  AOI22_X1 U11889 ( .A1(n30684), .A2(\xmem_data[46][5] ), .B1(n28687), .B2(
        \xmem_data[47][5] ), .ZN(n8050) );
  NAND4_X1 U11890 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n8064)
         );
  AOI22_X1 U11891 ( .A1(n30766), .A2(\xmem_data[48][5] ), .B1(n30170), .B2(
        \xmem_data[49][5] ), .ZN(n8057) );
  AOI22_X1 U11892 ( .A1(n28702), .A2(\xmem_data[50][5] ), .B1(n28701), .B2(
        \xmem_data[51][5] ), .ZN(n8056) );
  AOI22_X1 U11893 ( .A1(n28725), .A2(\xmem_data[52][5] ), .B1(n28696), .B2(
        \xmem_data[53][5] ), .ZN(n8055) );
  AOI22_X1 U11894 ( .A1(n28681), .A2(\xmem_data[54][5] ), .B1(n17051), .B2(
        \xmem_data[55][5] ), .ZN(n8054) );
  NAND4_X1 U11895 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n8063)
         );
  AOI22_X1 U11896 ( .A1(n28765), .A2(\xmem_data[56][5] ), .B1(n27723), .B2(
        \xmem_data[57][5] ), .ZN(n8061) );
  AOI22_X1 U11897 ( .A1(n3227), .A2(\xmem_data[58][5] ), .B1(n28677), .B2(
        \xmem_data[59][5] ), .ZN(n8060) );
  AOI22_X1 U11898 ( .A1(n29626), .A2(\xmem_data[60][5] ), .B1(n26616), .B2(
        \xmem_data[61][5] ), .ZN(n8059) );
  AOI22_X1 U11899 ( .A1(n29790), .A2(\xmem_data[62][5] ), .B1(n28218), .B2(
        \xmem_data[63][5] ), .ZN(n8058) );
  NAND4_X1 U11900 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n8062)
         );
  BUF_X1 U11901 ( .A(n11439), .Z(n28779) );
  AOI22_X1 U11902 ( .A1(n3173), .A2(\xmem_data[8][5] ), .B1(n29648), .B2(
        \xmem_data[9][5] ), .ZN(n8071) );
  AOI22_X1 U11903 ( .A1(n28780), .A2(\xmem_data[10][5] ), .B1(n30746), .B2(
        \xmem_data[11][5] ), .ZN(n8070) );
  AOI22_X1 U11904 ( .A1(n3162), .A2(\xmem_data[12][5] ), .B1(n3187), .B2(
        \xmem_data[13][5] ), .ZN(n8069) );
  BUF_X1 U11905 ( .A(n15549), .Z(n28755) );
  BUF_X1 U11906 ( .A(n14971), .Z(n28754) );
  AOI22_X1 U11907 ( .A1(n28755), .A2(\xmem_data[14][5] ), .B1(n28754), .B2(
        \xmem_data[15][5] ), .ZN(n8068) );
  AOI22_X1 U11908 ( .A1(n29722), .A2(\xmem_data[16][5] ), .B1(n29721), .B2(
        \xmem_data[17][5] ), .ZN(n8079) );
  AOI22_X1 U11909 ( .A1(n28702), .A2(\xmem_data[18][5] ), .B1(n29816), .B2(
        \xmem_data[19][5] ), .ZN(n8078) );
  AOI22_X1 U11910 ( .A1(n28725), .A2(\xmem_data[20][5] ), .B1(n29381), .B2(
        \xmem_data[21][5] ), .ZN(n8077) );
  BUF_X1 U11911 ( .A(n13420), .Z(n28772) );
  AOI22_X1 U11912 ( .A1(n29489), .A2(\xmem_data[22][5] ), .B1(n28772), .B2(
        \xmem_data[23][5] ), .ZN(n8076) );
  BUF_X1 U11913 ( .A(n11484), .Z(n28787) );
  BUF_X1 U11914 ( .A(n11780), .Z(n28786) );
  AOI22_X1 U11915 ( .A1(n28787), .A2(\xmem_data[0][5] ), .B1(n29495), .B2(
        \xmem_data[1][5] ), .ZN(n8085) );
  AOI22_X1 U11916 ( .A1(n3244), .A2(\xmem_data[2][5] ), .B1(n29706), .B2(
        \xmem_data[3][5] ), .ZN(n8084) );
  AOI22_X1 U11917 ( .A1(n29390), .A2(\xmem_data[4][5] ), .B1(n27761), .B2(
        \xmem_data[5][5] ), .ZN(n8083) );
  BUF_X1 U11918 ( .A(n8081), .Z(n28788) );
  AOI22_X1 U11919 ( .A1(n28788), .A2(\xmem_data[6][5] ), .B1(n30083), .B2(
        \xmem_data[7][5] ), .ZN(n8082) );
  AOI22_X1 U11920 ( .A1(n27710), .A2(\xmem_data[28][5] ), .B1(n28766), .B2(
        \xmem_data[29][5] ), .ZN(n8086) );
  INV_X1 U11921 ( .A(n8086), .ZN(n8095) );
  AOI22_X1 U11922 ( .A1(n29699), .A2(\xmem_data[30][5] ), .B1(n29832), .B2(
        \xmem_data[31][5] ), .ZN(n8087) );
  INV_X1 U11923 ( .A(n8087), .ZN(n8094) );
  AOI22_X1 U11924 ( .A1(n28765), .A2(\xmem_data[24][5] ), .B1(n27723), .B2(
        \xmem_data[25][5] ), .ZN(n8092) );
  AOI22_X1 U11925 ( .A1(n3227), .A2(\xmem_data[26][5] ), .B1(n24630), .B2(
        \xmem_data[27][5] ), .ZN(n8091) );
  NAND2_X1 U11926 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  NOR3_X1 U11927 ( .A1(n8095), .A2(n8094), .A3(n8093), .ZN(n8096) );
  NAND4_X1 U11928 ( .A1(n3840), .A2(n3541), .A3(n3476), .A4(n8096), .ZN(n8097)
         );
  AOI22_X1 U11929 ( .A1(n28713), .A2(n8098), .B1(n28794), .B2(n8097), .ZN(
        n8099) );
  AOI22_X1 U11930 ( .A1(n29786), .A2(\xmem_data[120][4] ), .B1(n3124), .B2(
        \xmem_data[121][4] ), .ZN(n8104) );
  AOI22_X1 U11931 ( .A1(n28719), .A2(\xmem_data[122][4] ), .B1(n28718), .B2(
        \xmem_data[123][4] ), .ZN(n8103) );
  AOI22_X1 U11932 ( .A1(n27710), .A2(\xmem_data[124][4] ), .B1(n30707), .B2(
        \xmem_data[125][4] ), .ZN(n8102) );
  AOI22_X1 U11933 ( .A1(n29628), .A2(\xmem_data[126][4] ), .B1(n28733), .B2(
        \xmem_data[127][4] ), .ZN(n8101) );
  NAND4_X1 U11934 ( .A1(n8104), .A2(n8103), .A3(n8102), .A4(n8101), .ZN(n8121)
         );
  AOI22_X1 U11935 ( .A1(n28740), .A2(\xmem_data[96][4] ), .B1(n28208), .B2(
        \xmem_data[97][4] ), .ZN(n8108) );
  AOI22_X1 U11936 ( .A1(n3244), .A2(\xmem_data[98][4] ), .B1(n3126), .B2(
        \xmem_data[99][4] ), .ZN(n8107) );
  AOI22_X1 U11937 ( .A1(n30633), .A2(\xmem_data[100][4] ), .B1(n28145), .B2(
        \xmem_data[101][4] ), .ZN(n8106) );
  AOI22_X1 U11938 ( .A1(n28744), .A2(\xmem_data[102][4] ), .B1(n28743), .B2(
        \xmem_data[103][4] ), .ZN(n8105) );
  NAND4_X1 U11939 ( .A1(n8108), .A2(n8107), .A3(n8106), .A4(n8105), .ZN(n8120)
         );
  AOI22_X1 U11940 ( .A1(n29363), .A2(\xmem_data[112][4] ), .B1(n30266), .B2(
        \xmem_data[113][4] ), .ZN(n8112) );
  AOI22_X1 U11941 ( .A1(n28720), .A2(\xmem_data[114][4] ), .B1(n28701), .B2(
        \xmem_data[115][4] ), .ZN(n8111) );
  AOI22_X1 U11942 ( .A1(n28725), .A2(\xmem_data[116][4] ), .B1(n28724), .B2(
        \xmem_data[117][4] ), .ZN(n8110) );
  AOI22_X1 U11943 ( .A1(n28727), .A2(\xmem_data[118][4] ), .B1(n29298), .B2(
        \xmem_data[119][4] ), .ZN(n8109) );
  NAND4_X1 U11944 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8119)
         );
  AOI22_X1 U11945 ( .A1(n27754), .A2(\xmem_data[104][4] ), .B1(n29739), .B2(
        \xmem_data[105][4] ), .ZN(n8117) );
  AOI22_X1 U11946 ( .A1(n28753), .A2(\xmem_data[106][4] ), .B1(n29437), .B2(
        \xmem_data[107][4] ), .ZN(n8116) );
  AOI22_X1 U11947 ( .A1(n3164), .A2(\xmem_data[108][4] ), .B1(n3188), .B2(
        \xmem_data[109][4] ), .ZN(n8115) );
  AND2_X1 U11948 ( .A1(n28781), .A2(\xmem_data[111][4] ), .ZN(n8113) );
  AOI21_X1 U11949 ( .B1(n29810), .B2(\xmem_data[110][4] ), .A(n8113), .ZN(
        n8114) );
  NAND4_X1 U11950 ( .A1(n8117), .A2(n8116), .A3(n8115), .A4(n8114), .ZN(n8118)
         );
  NAND2_X1 U11951 ( .A1(n8122), .A2(n28762), .ZN(n8196) );
  AOI22_X1 U11952 ( .A1(n30294), .A2(\xmem_data[32][4] ), .B1(n29761), .B2(
        \xmem_data[33][4] ), .ZN(n8126) );
  AOI22_X1 U11953 ( .A1(n28670), .A2(\xmem_data[34][4] ), .B1(n29350), .B2(
        \xmem_data[35][4] ), .ZN(n8125) );
  AOI22_X1 U11954 ( .A1(n28180), .A2(\xmem_data[36][4] ), .B1(n28238), .B2(
        \xmem_data[37][4] ), .ZN(n8124) );
  AOI22_X1 U11955 ( .A1(n28788), .A2(\xmem_data[38][4] ), .B1(n28671), .B2(
        \xmem_data[39][4] ), .ZN(n8123) );
  NAND4_X1 U11956 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n8143)
         );
  AOI22_X1 U11957 ( .A1(n3174), .A2(\xmem_data[40][4] ), .B1(n30301), .B2(
        \xmem_data[41][4] ), .ZN(n8130) );
  AOI22_X1 U11958 ( .A1(n28686), .A2(\xmem_data[42][4] ), .B1(n29237), .B2(
        \xmem_data[43][4] ), .ZN(n8129) );
  AOI22_X1 U11959 ( .A1(n3168), .A2(\xmem_data[44][4] ), .B1(n3184), .B2(
        \xmem_data[45][4] ), .ZN(n8128) );
  AOI22_X1 U11960 ( .A1(n23901), .A2(\xmem_data[46][4] ), .B1(n28754), .B2(
        \xmem_data[47][4] ), .ZN(n8127) );
  NAND4_X1 U11961 ( .A1(n8130), .A2(n8129), .A3(n8128), .A4(n8127), .ZN(n8142)
         );
  AOI22_X1 U11962 ( .A1(n29722), .A2(\xmem_data[48][4] ), .B1(n30685), .B2(
        \xmem_data[49][4] ), .ZN(n8134) );
  AOI22_X1 U11963 ( .A1(n28702), .A2(\xmem_data[50][4] ), .B1(n28701), .B2(
        \xmem_data[51][4] ), .ZN(n8133) );
  AOI22_X1 U11964 ( .A1(n29724), .A2(\xmem_data[52][4] ), .B1(n28696), .B2(
        \xmem_data[53][4] ), .ZN(n8132) );
  AOI22_X1 U11965 ( .A1(n28681), .A2(\xmem_data[54][4] ), .B1(n25684), .B2(
        \xmem_data[55][4] ), .ZN(n8131) );
  NAND4_X1 U11966 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n8141)
         );
  AOI22_X1 U11967 ( .A1(n29786), .A2(\xmem_data[56][4] ), .B1(n29418), .B2(
        \xmem_data[57][4] ), .ZN(n8139) );
  AOI22_X1 U11968 ( .A1(n3227), .A2(\xmem_data[58][4] ), .B1(n28677), .B2(
        \xmem_data[59][4] ), .ZN(n8138) );
  AOI22_X1 U11969 ( .A1(n29626), .A2(\xmem_data[60][4] ), .B1(n29672), .B2(
        \xmem_data[61][4] ), .ZN(n8137) );
  AND2_X1 U11970 ( .A1(n30292), .A2(\xmem_data[63][4] ), .ZN(n8135) );
  AOI21_X1 U11971 ( .B1(n29423), .B2(\xmem_data[62][4] ), .A(n8135), .ZN(n8136) );
  NAND4_X1 U11972 ( .A1(n8137), .A2(n8138), .A3(n8139), .A4(n8136), .ZN(n8140)
         );
  NAND2_X1 U11973 ( .A1(n8144), .A2(n28713), .ZN(n8195) );
  NAND2_X1 U11974 ( .A1(n27833), .A2(\xmem_data[65][4] ), .ZN(n8146) );
  NAND2_X1 U11975 ( .A1(n28740), .A2(\xmem_data[64][4] ), .ZN(n8145) );
  NAND2_X1 U11976 ( .A1(n8146), .A2(n8145), .ZN(n8152) );
  AOI22_X1 U11977 ( .A1(n30633), .A2(\xmem_data[68][4] ), .B1(n29704), .B2(
        \xmem_data[69][4] ), .ZN(n8147) );
  INV_X1 U11978 ( .A(n8147), .ZN(n8151) );
  AOI22_X1 U11979 ( .A1(n28670), .A2(\xmem_data[66][4] ), .B1(n14991), .B2(
        \xmem_data[67][4] ), .ZN(n8149) );
  AOI22_X1 U11980 ( .A1(n28744), .A2(\xmem_data[70][4] ), .B1(n28671), .B2(
        \xmem_data[71][4] ), .ZN(n8148) );
  NAND2_X1 U11981 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  NOR3_X1 U11982 ( .A1(n8152), .A2(n8151), .A3(n8150), .ZN(n8170) );
  NAND2_X1 U11983 ( .A1(n29433), .A2(\xmem_data[92][4] ), .ZN(n8154) );
  NAND2_X1 U11984 ( .A1(n30100), .A2(\xmem_data[93][4] ), .ZN(n8153) );
  NAND2_X1 U11985 ( .A1(n8154), .A2(n8153), .ZN(n8159) );
  AOI22_X1 U11986 ( .A1(n29628), .A2(\xmem_data[94][4] ), .B1(n29565), .B2(
        \xmem_data[95][4] ), .ZN(n8157) );
  AOI22_X1 U11987 ( .A1(n3227), .A2(\xmem_data[90][4] ), .B1(n28677), .B2(
        \xmem_data[91][4] ), .ZN(n8156) );
  AOI22_X1 U11988 ( .A1(n29829), .A2(\xmem_data[88][4] ), .B1(n27743), .B2(
        \xmem_data[89][4] ), .ZN(n8155) );
  NAND3_X1 U11989 ( .A1(n8157), .A2(n8156), .A3(n8155), .ZN(n8158) );
  NOR2_X1 U11990 ( .A1(n8159), .A2(n8158), .ZN(n8169) );
  AOI22_X1 U11991 ( .A1(n27754), .A2(\xmem_data[72][4] ), .B1(n30193), .B2(
        \xmem_data[73][4] ), .ZN(n8164) );
  AOI22_X1 U11992 ( .A1(n28686), .A2(\xmem_data[74][4] ), .B1(n27818), .B2(
        \xmem_data[75][4] ), .ZN(n8163) );
  AOI22_X1 U11993 ( .A1(n3161), .A2(\xmem_data[76][4] ), .B1(n3184), .B2(
        \xmem_data[77][4] ), .ZN(n8162) );
  AND2_X1 U11994 ( .A1(n28781), .A2(\xmem_data[79][4] ), .ZN(n8160) );
  AOI21_X1 U11995 ( .B1(n29716), .B2(\xmem_data[78][4] ), .A(n8160), .ZN(n8161) );
  AOI22_X1 U11996 ( .A1(n27713), .A2(\xmem_data[80][4] ), .B1(n29640), .B2(
        \xmem_data[81][4] ), .ZN(n8168) );
  AOI22_X1 U11997 ( .A1(n28702), .A2(\xmem_data[82][4] ), .B1(n28701), .B2(
        \xmem_data[83][4] ), .ZN(n8167) );
  AOI22_X1 U11998 ( .A1(n28725), .A2(\xmem_data[84][4] ), .B1(n28696), .B2(
        \xmem_data[85][4] ), .ZN(n8166) );
  AOI22_X1 U11999 ( .A1(n28681), .A2(\xmem_data[86][4] ), .B1(n29298), .B2(
        \xmem_data[87][4] ), .ZN(n8165) );
  NAND4_X1 U12000 ( .A1(n8170), .A2(n8169), .A3(n3794), .A4(n3507), .ZN(n8171)
         );
  NAND2_X1 U12001 ( .A1(n8171), .A2(n28662), .ZN(n8194) );
  AOI22_X1 U12002 ( .A1(n29829), .A2(\xmem_data[24][4] ), .B1(n27743), .B2(
        \xmem_data[25][4] ), .ZN(n8175) );
  AOI22_X1 U12003 ( .A1(n3227), .A2(\xmem_data[26][4] ), .B1(n3149), .B2(
        \xmem_data[27][4] ), .ZN(n8174) );
  AOI22_X1 U12004 ( .A1(n29628), .A2(\xmem_data[30][4] ), .B1(n30278), .B2(
        \xmem_data[31][4] ), .ZN(n8172) );
  NAND4_X1 U12005 ( .A1(n8175), .A2(n8174), .A3(n8173), .A4(n8172), .ZN(n8191)
         );
  AOI22_X1 U12006 ( .A1(n29436), .A2(\xmem_data[8][4] ), .B1(n29768), .B2(
        \xmem_data[9][4] ), .ZN(n8179) );
  AOI22_X1 U12007 ( .A1(n28780), .A2(\xmem_data[10][4] ), .B1(n27945), .B2(
        \xmem_data[11][4] ), .ZN(n8178) );
  AOI22_X1 U12008 ( .A1(n3164), .A2(\xmem_data[12][4] ), .B1(n3184), .B2(
        \xmem_data[13][4] ), .ZN(n8177) );
  AOI22_X1 U12009 ( .A1(n26812), .A2(\xmem_data[14][4] ), .B1(n28754), .B2(
        \xmem_data[15][4] ), .ZN(n8176) );
  NAND4_X1 U12010 ( .A1(n8179), .A2(n8178), .A3(n8177), .A4(n8176), .ZN(n8190)
         );
  AOI22_X1 U12011 ( .A1(n29722), .A2(\xmem_data[16][4] ), .B1(n30716), .B2(
        \xmem_data[17][4] ), .ZN(n8183) );
  AOI22_X1 U12012 ( .A1(n28702), .A2(\xmem_data[18][4] ), .B1(n29379), .B2(
        \xmem_data[19][4] ), .ZN(n8182) );
  AOI22_X1 U12013 ( .A1(n29724), .A2(\xmem_data[20][4] ), .B1(n27805), .B2(
        \xmem_data[21][4] ), .ZN(n8181) );
  AOI22_X1 U12014 ( .A1(n29489), .A2(\xmem_data[22][4] ), .B1(n28772), .B2(
        \xmem_data[23][4] ), .ZN(n8180) );
  NAND4_X1 U12015 ( .A1(n8183), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(n8189)
         );
  AOI22_X1 U12016 ( .A1(n28787), .A2(\xmem_data[0][4] ), .B1(n28208), .B2(
        \xmem_data[1][4] ), .ZN(n8187) );
  AOI22_X1 U12017 ( .A1(n3244), .A2(\xmem_data[2][4] ), .B1(n3146), .B2(
        \xmem_data[3][4] ), .ZN(n8186) );
  AOI22_X1 U12018 ( .A1(n29590), .A2(\xmem_data[4][4] ), .B1(n28738), .B2(
        \xmem_data[5][4] ), .ZN(n8185) );
  AOI22_X1 U12019 ( .A1(n28788), .A2(\xmem_data[6][4] ), .B1(n30083), .B2(
        \xmem_data[7][4] ), .ZN(n8184) );
  NAND4_X1 U12020 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n8188)
         );
  NAND2_X1 U12021 ( .A1(n8192), .A2(n28794), .ZN(n8193) );
  XNOR2_X1 U12022 ( .A(n3316), .B(\fmem_data[11][5] ), .ZN(n32024) );
  XOR2_X1 U12023 ( .A(\fmem_data[11][4] ), .B(\fmem_data[11][5] ), .Z(n8197)
         );
  AOI22_X1 U12024 ( .A1(n3163), .A2(\xmem_data[96][7] ), .B1(n3184), .B2(
        \xmem_data[97][7] ), .ZN(n8203) );
  BUF_X1 U12025 ( .A(n14971), .Z(n28232) );
  AOI22_X1 U12026 ( .A1(n30715), .A2(\xmem_data[98][7] ), .B1(n28232), .B2(
        \xmem_data[99][7] ), .ZN(n8202) );
  BUF_X1 U12027 ( .A(n10802), .Z(n28680) );
  AOI22_X1 U12028 ( .A1(n29488), .A2(\xmem_data[100][7] ), .B1(n30170), .B2(
        \xmem_data[101][7] ), .ZN(n8201) );
  NAND2_X1 U12029 ( .A1(n8204), .A2(n11350), .ZN(n8199) );
  AND2_X1 U12030 ( .A1(n11343), .A2(n6173), .ZN(n8198) );
  NAND2_X1 U12031 ( .A1(n11342), .A2(n8198), .ZN(n8218) );
  NOR2_X1 U12032 ( .A1(n8199), .A2(n8218), .ZN(n8253) );
  BUF_X1 U12033 ( .A(n14974), .Z(n28226) );
  AOI22_X1 U12034 ( .A1(n3233), .A2(\xmem_data[102][7] ), .B1(n28226), .B2(
        \xmem_data[103][7] ), .ZN(n8200) );
  NAND4_X1 U12035 ( .A1(n8203), .A2(n8202), .A3(n8201), .A4(n8200), .ZN(n8226)
         );
  NAND2_X1 U12036 ( .A1(n8204), .A2(n11357), .ZN(n8205) );
  NOR2_X1 U12037 ( .A1(n11358), .A2(n8205), .ZN(n8264) );
  BUF_X1 U12038 ( .A(n8264), .Z(n28240) );
  NOR2_X1 U12039 ( .A1(n11359), .A2(n8205), .ZN(n8368) );
  BUF_X2 U12040 ( .A(n8368), .Z(n28159) );
  AOI22_X1 U12041 ( .A1(n28240), .A2(\xmem_data[104][7] ), .B1(n28159), .B2(
        \xmem_data[105][7] ), .ZN(n8209) );
  NOR2_X1 U12042 ( .A1(n3378), .A2(n8205), .ZN(n8265) );
  BUF_X1 U12043 ( .A(n8265), .Z(n28242) );
  BUF_X1 U12044 ( .A(n13420), .Z(n28241) );
  AOI22_X1 U12045 ( .A1(n28242), .A2(\xmem_data[106][7] ), .B1(n28241), .B2(
        \xmem_data[107][7] ), .ZN(n8208) );
  NOR2_X1 U12046 ( .A1(n11361), .A2(n8205), .ZN(n8266) );
  NOR2_X1 U12047 ( .A1(n8205), .A2(n3246), .ZN(n8267) );
  AOI22_X1 U12048 ( .A1(n28244), .A2(\xmem_data[108][7] ), .B1(n28243), .B2(
        \xmem_data[109][7] ), .ZN(n8207) );
  NOR2_X1 U12049 ( .A1(n8218), .A2(n8205), .ZN(n28111) );
  BUF_X1 U12050 ( .A(n28111), .Z(n28246) );
  BUF_X1 U12051 ( .A(n28973), .Z(n28245) );
  AOI22_X1 U12052 ( .A1(n28246), .A2(\xmem_data[110][7] ), .B1(n28245), .B2(
        \xmem_data[111][7] ), .ZN(n8206) );
  NAND4_X1 U12053 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8225)
         );
  AOI22_X1 U12054 ( .A1(n28136), .A2(\xmem_data[112][7] ), .B1(n30106), .B2(
        \xmem_data[113][7] ), .ZN(n8215) );
  BUF_X1 U12055 ( .A(n14988), .Z(n28218) );
  AOI22_X1 U12056 ( .A1(n28138), .A2(\xmem_data[114][7] ), .B1(n28218), .B2(
        \xmem_data[115][7] ), .ZN(n8214) );
  BUF_X1 U12057 ( .A(n11484), .Z(n28219) );
  AOI22_X1 U12058 ( .A1(n28219), .A2(\xmem_data[116][7] ), .B1(n28786), .B2(
        \xmem_data[117][7] ), .ZN(n8213) );
  NAND2_X1 U12059 ( .A1(n8210), .A2(n11350), .ZN(n8211) );
  NOR2_X1 U12060 ( .A1(n8218), .A2(n8211), .ZN(n8272) );
  BUF_X1 U12061 ( .A(n8272), .Z(n28220) );
  AOI22_X1 U12062 ( .A1(n28220), .A2(\xmem_data[118][7] ), .B1(n3126), .B2(
        \xmem_data[119][7] ), .ZN(n8212) );
  NAND4_X1 U12063 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n8212), .ZN(n8224)
         );
  BUF_X1 U12064 ( .A(n11437), .Z(n28238) );
  AOI22_X1 U12065 ( .A1(n29390), .A2(\xmem_data[120][7] ), .B1(n28665), .B2(
        \xmem_data[121][7] ), .ZN(n8222) );
  NAND2_X1 U12066 ( .A1(n8216), .A2(n11357), .ZN(n8217) );
  NOR2_X1 U12067 ( .A1(n3378), .A2(n8217), .ZN(n8258) );
  BUF_X1 U12068 ( .A(n14997), .Z(n28233) );
  AOI22_X1 U12069 ( .A1(n3241), .A2(\xmem_data[122][7] ), .B1(n28233), .B2(
        \xmem_data[123][7] ), .ZN(n8221) );
  BUF_X1 U12070 ( .A(n8700), .Z(n30090) );
  AOI22_X1 U12071 ( .A1(n30665), .A2(\xmem_data[124][7] ), .B1(n30084), .B2(
        \xmem_data[125][7] ), .ZN(n8220) );
  NOR2_X1 U12072 ( .A1(n8218), .A2(n8217), .ZN(n8259) );
  BUF_X1 U12073 ( .A(n3464), .Z(n28231) );
  AOI22_X1 U12074 ( .A1(n3240), .A2(\xmem_data[126][7] ), .B1(n28231), .B2(
        \xmem_data[127][7] ), .ZN(n8219) );
  NAND4_X1 U12075 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n8223)
         );
  INV_X1 U12076 ( .A(n3464), .ZN(n8228) );
  NOR3_X1 U12077 ( .A1(n37191), .A2(n8409), .A3(n8227), .ZN(n9418) );
  AOI22_X1 U12078 ( .A1(load_xaddr_val[5]), .A2(n8228), .B1(n9418), .B2(n3248), 
        .ZN(n8303) );
  INV_X1 U12079 ( .A(n14909), .ZN(n8230) );
  NAND2_X1 U12080 ( .A1(n3464), .A2(n39040), .ZN(n8229) );
  OAI21_X1 U12081 ( .B1(n21005), .B2(n8230), .A(n8229), .ZN(n8302) );
  INV_X1 U12082 ( .A(n8302), .ZN(n8283) );
  AND2_X1 U12083 ( .A1(n8303), .A2(n8283), .ZN(n28133) );
  NAND2_X1 U12084 ( .A1(n8231), .A2(n28133), .ZN(n8308) );
  AOI22_X1 U12085 ( .A1(n3164), .A2(\xmem_data[32][7] ), .B1(n3189), .B2(
        \xmem_data[33][7] ), .ZN(n8235) );
  BUF_X1 U12086 ( .A(n14971), .Z(n28147) );
  AOI22_X1 U12087 ( .A1(n30684), .A2(\xmem_data[34][7] ), .B1(n28147), .B2(
        \xmem_data[35][7] ), .ZN(n8234) );
  AOI22_X1 U12088 ( .A1(n29488), .A2(\xmem_data[36][7] ), .B1(n30266), .B2(
        \xmem_data[37][7] ), .ZN(n8233) );
  BUF_X1 U12089 ( .A(n8253), .Z(n28151) );
  AOI22_X1 U12090 ( .A1(n28151), .A2(\xmem_data[38][7] ), .B1(n29573), .B2(
        \xmem_data[39][7] ), .ZN(n8232) );
  NAND4_X1 U12091 ( .A1(n8235), .A2(n8234), .A3(n8233), .A4(n8232), .ZN(n8251)
         );
  BUF_X1 U12092 ( .A(n8264), .Z(n28160) );
  AOI22_X1 U12093 ( .A1(n28160), .A2(\xmem_data[40][7] ), .B1(n28159), .B2(
        \xmem_data[41][7] ), .ZN(n8239) );
  BUF_X1 U12094 ( .A(n8265), .Z(n28161) );
  AOI22_X1 U12095 ( .A1(n28161), .A2(\xmem_data[42][7] ), .B1(n28192), .B2(
        \xmem_data[43][7] ), .ZN(n8238) );
  AOI22_X1 U12096 ( .A1(n28163), .A2(\xmem_data[44][7] ), .B1(n28162), .B2(
        \xmem_data[45][7] ), .ZN(n8237) );
  BUF_X1 U12097 ( .A(n28973), .Z(n28164) );
  AOI22_X1 U12098 ( .A1(n28165), .A2(\xmem_data[46][7] ), .B1(n28164), .B2(
        \xmem_data[47][7] ), .ZN(n8236) );
  NAND4_X1 U12099 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n8250)
         );
  BUF_X2 U12100 ( .A(n11451), .Z(n28138) );
  BUF_X1 U12101 ( .A(n14988), .Z(n28137) );
  AOI22_X1 U12102 ( .A1(n28700), .A2(\xmem_data[50][7] ), .B1(n28137), .B2(
        \xmem_data[51][7] ), .ZN(n8243) );
  AOI22_X1 U12103 ( .A1(n30708), .A2(\xmem_data[48][7] ), .B1(n28766), .B2(
        \xmem_data[49][7] ), .ZN(n8242) );
  BUF_X1 U12104 ( .A(n11484), .Z(n28139) );
  AOI22_X1 U12105 ( .A1(n28139), .A2(\xmem_data[52][7] ), .B1(n30776), .B2(
        \xmem_data[53][7] ), .ZN(n8241) );
  BUF_X1 U12106 ( .A(n8272), .Z(n28140) );
  AOI22_X1 U12107 ( .A1(n28140), .A2(\xmem_data[54][7] ), .B1(n27905), .B2(
        \xmem_data[55][7] ), .ZN(n8240) );
  NAND4_X1 U12108 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n8249)
         );
  BUF_X1 U12109 ( .A(n11436), .Z(n28146) );
  AOI22_X1 U12110 ( .A1(n29602), .A2(\xmem_data[56][7] ), .B1(n3369), .B2(
        \xmem_data[57][7] ), .ZN(n8247) );
  BUF_X1 U12111 ( .A(n8258), .Z(n28153) );
  BUF_X1 U12112 ( .A(n14997), .Z(n28152) );
  AOI22_X1 U12113 ( .A1(n28153), .A2(\xmem_data[58][7] ), .B1(n28152), .B2(
        \xmem_data[59][7] ), .ZN(n8246) );
  BUF_X1 U12114 ( .A(n8700), .Z(n30084) );
  AOI22_X1 U12115 ( .A1(n29604), .A2(\xmem_data[60][7] ), .B1(n26884), .B2(
        \xmem_data[61][7] ), .ZN(n8245) );
  BUF_X1 U12116 ( .A(n8259), .Z(n28155) );
  BUF_X1 U12117 ( .A(n3464), .Z(n28154) );
  AOI22_X1 U12118 ( .A1(n28155), .A2(\xmem_data[62][7] ), .B1(n28154), .B2(
        \xmem_data[63][7] ), .ZN(n8244) );
  NAND4_X1 U12119 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(n8248)
         );
  OR4_X1 U12120 ( .A1(n8251), .A2(n8249), .A3(n8250), .A4(n8248), .ZN(n8252)
         );
  NAND2_X1 U12121 ( .A1(n8252), .A2(n28177), .ZN(n8307) );
  AOI22_X1 U12122 ( .A1(n3160), .A2(\xmem_data[0][7] ), .B1(n3185), .B2(
        \xmem_data[1][7] ), .ZN(n8257) );
  AOI22_X1 U12123 ( .A1(n30684), .A2(\xmem_data[2][7] ), .B1(n24115), .B2(
        \xmem_data[3][7] ), .ZN(n8256) );
  AOI22_X1 U12124 ( .A1(n30717), .A2(\xmem_data[4][7] ), .B1(n30266), .B2(
        \xmem_data[5][7] ), .ZN(n8255) );
  BUF_X1 U12125 ( .A(n14974), .Z(n28202) );
  AOI22_X1 U12126 ( .A1(n3233), .A2(\xmem_data[6][7] ), .B1(n28202), .B2(
        \xmem_data[7][7] ), .ZN(n8254) );
  BUF_X1 U12127 ( .A(n11436), .Z(n28180) );
  AOI22_X1 U12128 ( .A1(n28739), .A2(\xmem_data[24][7] ), .B1(n28738), .B2(
        \xmem_data[25][7] ), .ZN(n8263) );
  AOI22_X1 U12129 ( .A1(n3241), .A2(\xmem_data[26][7] ), .B1(n30083), .B2(
        \xmem_data[27][7] ), .ZN(n8262) );
  AOI22_X1 U12130 ( .A1(n27811), .A2(\xmem_data[28][7] ), .B1(n27728), .B2(
        \xmem_data[29][7] ), .ZN(n8261) );
  AOI22_X1 U12131 ( .A1(n3240), .A2(\xmem_data[30][7] ), .B1(n21005), .B2(
        \xmem_data[31][7] ), .ZN(n8260) );
  NAND4_X1 U12132 ( .A1(n8263), .A2(n8262), .A3(n8261), .A4(n8260), .ZN(n8279)
         );
  BUF_X1 U12133 ( .A(n11484), .Z(n28209) );
  BUF_X1 U12134 ( .A(n11780), .Z(n28208) );
  AOI22_X1 U12135 ( .A1(n28209), .A2(\xmem_data[20][7] ), .B1(n3198), .B2(
        \xmem_data[21][7] ), .ZN(n8277) );
  BUF_X1 U12136 ( .A(n8264), .Z(n28191) );
  BUF_X1 U12137 ( .A(n8368), .Z(n28190) );
  AOI22_X1 U12138 ( .A1(n28191), .A2(\xmem_data[8][7] ), .B1(n28190), .B2(
        \xmem_data[9][7] ), .ZN(n8271) );
  BUF_X1 U12139 ( .A(n8265), .Z(n28193) );
  BUF_X1 U12140 ( .A(n13127), .Z(n28192) );
  AOI22_X1 U12141 ( .A1(n28193), .A2(\xmem_data[10][7] ), .B1(n28192), .B2(
        \xmem_data[11][7] ), .ZN(n8270) );
  BUF_X1 U12142 ( .A(n8266), .Z(n28195) );
  AOI22_X1 U12143 ( .A1(n28195), .A2(\xmem_data[12][7] ), .B1(n28194), .B2(
        \xmem_data[13][7] ), .ZN(n8269) );
  AOI22_X1 U12144 ( .A1(n28196), .A2(\xmem_data[14][7] ), .B1(n28677), .B2(
        \xmem_data[15][7] ), .ZN(n8268) );
  NAND4_X1 U12145 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(n8275)
         );
  BUF_X1 U12146 ( .A(n8272), .Z(n28210) );
  AOI22_X1 U12147 ( .A1(n28210), .A2(\xmem_data[22][7] ), .B1(n30698), .B2(
        \xmem_data[23][7] ), .ZN(n8273) );
  INV_X1 U12148 ( .A(n8273), .ZN(n8274) );
  NOR2_X1 U12149 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  NAND2_X1 U12150 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  NOR2_X1 U12151 ( .A1(n8279), .A2(n8278), .ZN(n8282) );
  BUF_X1 U12152 ( .A(n11451), .Z(n28207) );
  AOI22_X1 U12153 ( .A1(n29790), .A2(\xmem_data[18][7] ), .B1(n29565), .B2(
        \xmem_data[19][7] ), .ZN(n8281) );
  AOI22_X1 U12154 ( .A1(n29433), .A2(\xmem_data[16][7] ), .B1(n30290), .B2(
        \xmem_data[17][7] ), .ZN(n8280) );
  NAND4_X1 U12155 ( .A1(n3826), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n8284)
         );
  NOR2_X1 U12156 ( .A1(n8303), .A2(n8283), .ZN(n28215) );
  NAND2_X1 U12157 ( .A1(n8284), .A2(n28215), .ZN(n8306) );
  AOI22_X1 U12158 ( .A1(n3164), .A2(\xmem_data[64][7] ), .B1(n3181), .B2(
        \xmem_data[65][7] ), .ZN(n8288) );
  AOI22_X1 U12159 ( .A1(n30070), .A2(\xmem_data[66][7] ), .B1(n28147), .B2(
        \xmem_data[67][7] ), .ZN(n8287) );
  AOI22_X1 U12160 ( .A1(n29363), .A2(\xmem_data[68][7] ), .B1(n30716), .B2(
        \xmem_data[69][7] ), .ZN(n8286) );
  AOI22_X1 U12161 ( .A1(n28151), .A2(\xmem_data[70][7] ), .B1(n30645), .B2(
        \xmem_data[71][7] ), .ZN(n8285) );
  AOI22_X1 U12162 ( .A1(n28160), .A2(\xmem_data[72][7] ), .B1(n28159), .B2(
        \xmem_data[73][7] ), .ZN(n8292) );
  AOI22_X1 U12163 ( .A1(n28161), .A2(\xmem_data[74][7] ), .B1(n14982), .B2(
        \xmem_data[75][7] ), .ZN(n8291) );
  AOI22_X1 U12164 ( .A1(n28163), .A2(\xmem_data[76][7] ), .B1(n28162), .B2(
        \xmem_data[77][7] ), .ZN(n8290) );
  AOI22_X1 U12165 ( .A1(n28165), .A2(\xmem_data[78][7] ), .B1(n28164), .B2(
        \xmem_data[79][7] ), .ZN(n8289) );
  AOI22_X1 U12166 ( .A1(n28138), .A2(\xmem_data[82][7] ), .B1(n28137), .B2(
        \xmem_data[83][7] ), .ZN(n8297) );
  AOI22_X1 U12167 ( .A1(n28139), .A2(\xmem_data[84][7] ), .B1(n28786), .B2(
        \xmem_data[85][7] ), .ZN(n8296) );
  AOI22_X1 U12168 ( .A1(n30291), .A2(\xmem_data[80][7] ), .B1(n28206), .B2(
        \xmem_data[81][7] ), .ZN(n8295) );
  AOI22_X1 U12169 ( .A1(n28140), .A2(\xmem_data[86][7] ), .B1(n30295), .B2(
        \xmem_data[87][7] ), .ZN(n8294) );
  AOI22_X1 U12170 ( .A1(n30633), .A2(\xmem_data[88][7] ), .B1(n29482), .B2(
        \xmem_data[89][7] ), .ZN(n8301) );
  AOI22_X1 U12171 ( .A1(n28153), .A2(\xmem_data[90][7] ), .B1(n28152), .B2(
        \xmem_data[91][7] ), .ZN(n8300) );
  AOI22_X1 U12172 ( .A1(n30302), .A2(\xmem_data[92][7] ), .B1(n30084), .B2(
        \xmem_data[93][7] ), .ZN(n8299) );
  AOI22_X1 U12173 ( .A1(n28155), .A2(\xmem_data[94][7] ), .B1(n28154), .B2(
        \xmem_data[95][7] ), .ZN(n8298) );
  NOR2_X1 U12174 ( .A1(n8303), .A2(n8302), .ZN(n28258) );
  NAND2_X1 U12175 ( .A1(n8304), .A2(n28258), .ZN(n8305) );
  NAND4_X2 U12176 ( .A1(n8308), .A2(n8305), .A3(n8307), .A4(n8306), .ZN(n35256) );
  XNOR2_X1 U12177 ( .A(n35256), .B(\fmem_data[31][3] ), .ZN(n30364) );
  AOI22_X1 U12178 ( .A1(n3163), .A2(\xmem_data[32][6] ), .B1(n3186), .B2(
        \xmem_data[33][6] ), .ZN(n8312) );
  AOI22_X1 U12179 ( .A1(n30075), .A2(\xmem_data[34][6] ), .B1(n28147), .B2(
        \xmem_data[35][6] ), .ZN(n8311) );
  AOI22_X1 U12180 ( .A1(n29488), .A2(\xmem_data[36][6] ), .B1(n29487), .B2(
        \xmem_data[37][6] ), .ZN(n8310) );
  AOI22_X1 U12181 ( .A1(n28151), .A2(\xmem_data[38][6] ), .B1(n29297), .B2(
        \xmem_data[39][6] ), .ZN(n8309) );
  AOI22_X1 U12182 ( .A1(n29390), .A2(\xmem_data[56][6] ), .B1(n30730), .B2(
        \xmem_data[57][6] ), .ZN(n8316) );
  AOI22_X1 U12183 ( .A1(n28153), .A2(\xmem_data[58][6] ), .B1(n28152), .B2(
        \xmem_data[59][6] ), .ZN(n8315) );
  AOI22_X1 U12184 ( .A1(n30250), .A2(\xmem_data[60][6] ), .B1(n30084), .B2(
        \xmem_data[61][6] ), .ZN(n8314) );
  AOI22_X1 U12185 ( .A1(n28155), .A2(\xmem_data[62][6] ), .B1(n28154), .B2(
        \xmem_data[63][6] ), .ZN(n8313) );
  NAND4_X1 U12186 ( .A1(n8316), .A2(n8315), .A3(n8314), .A4(n8313), .ZN(n8329)
         );
  AOI22_X1 U12187 ( .A1(n29790), .A2(\xmem_data[50][6] ), .B1(n28137), .B2(
        \xmem_data[51][6] ), .ZN(n8327) );
  AOI22_X1 U12188 ( .A1(n30708), .A2(\xmem_data[48][6] ), .B1(n29753), .B2(
        \xmem_data[49][6] ), .ZN(n8326) );
  AOI22_X1 U12189 ( .A1(n28139), .A2(\xmem_data[52][6] ), .B1(n29798), .B2(
        \xmem_data[53][6] ), .ZN(n8325) );
  AOI22_X1 U12190 ( .A1(n28161), .A2(\xmem_data[42][6] ), .B1(n30674), .B2(
        \xmem_data[43][6] ), .ZN(n8320) );
  AOI22_X1 U12191 ( .A1(n28160), .A2(\xmem_data[40][6] ), .B1(n28159), .B2(
        \xmem_data[41][6] ), .ZN(n8319) );
  AOI22_X1 U12192 ( .A1(n28163), .A2(\xmem_data[44][6] ), .B1(n28162), .B2(
        \xmem_data[45][6] ), .ZN(n8318) );
  AOI22_X1 U12193 ( .A1(n28165), .A2(\xmem_data[46][6] ), .B1(n28164), .B2(
        \xmem_data[47][6] ), .ZN(n8317) );
  NAND4_X1 U12194 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n8323)
         );
  AOI22_X1 U12195 ( .A1(n28140), .A2(\xmem_data[54][6] ), .B1(n23742), .B2(
        \xmem_data[55][6] ), .ZN(n8321) );
  INV_X1 U12196 ( .A(n8321), .ZN(n8322) );
  NOR2_X1 U12197 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND4_X1 U12198 ( .A1(n8327), .A2(n8326), .A3(n8325), .A4(n8324), .ZN(n8328)
         );
  NOR2_X1 U12199 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  NAND2_X1 U12200 ( .A1(n3772), .A2(n8330), .ZN(n8355) );
  AOI22_X1 U12201 ( .A1(n3166), .A2(\xmem_data[0][6] ), .B1(n3189), .B2(
        \xmem_data[1][6] ), .ZN(n8334) );
  AOI22_X1 U12202 ( .A1(n27031), .A2(\xmem_data[2][6] ), .B1(n29639), .B2(
        \xmem_data[3][6] ), .ZN(n8333) );
  AOI22_X1 U12203 ( .A1(n30766), .A2(\xmem_data[4][6] ), .B1(n29487), .B2(
        \xmem_data[5][6] ), .ZN(n8332) );
  AOI22_X1 U12204 ( .A1(n3233), .A2(\xmem_data[6][6] ), .B1(n28202), .B2(
        \xmem_data[7][6] ), .ZN(n8331) );
  AOI22_X1 U12205 ( .A1(n29433), .A2(\xmem_data[16][6] ), .B1(n29432), .B2(
        \xmem_data[17][6] ), .ZN(n8353) );
  AND2_X1 U12206 ( .A1(n28218), .A2(\xmem_data[19][6] ), .ZN(n8335) );
  AOI21_X1 U12207 ( .B1(n28138), .B2(\xmem_data[18][6] ), .A(n8335), .ZN(n8352) );
  AOI22_X1 U12208 ( .A1(n28739), .A2(\xmem_data[24][6] ), .B1(n28738), .B2(
        \xmem_data[25][6] ), .ZN(n8339) );
  AOI22_X1 U12209 ( .A1(n3241), .A2(\xmem_data[26][6] ), .B1(n30083), .B2(
        \xmem_data[27][6] ), .ZN(n8338) );
  AOI22_X1 U12210 ( .A1(n28779), .A2(\xmem_data[28][6] ), .B1(n30090), .B2(
        \xmem_data[29][6] ), .ZN(n8337) );
  AOI22_X1 U12211 ( .A1(n3240), .A2(\xmem_data[30][6] ), .B1(n3158), .B2(
        \xmem_data[31][6] ), .ZN(n8336) );
  NAND4_X1 U12212 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(n8350)
         );
  AOI22_X1 U12213 ( .A1(n28209), .A2(\xmem_data[20][6] ), .B1(n29798), .B2(
        \xmem_data[21][6] ), .ZN(n8348) );
  AOI22_X1 U12214 ( .A1(n28191), .A2(\xmem_data[8][6] ), .B1(n28190), .B2(
        \xmem_data[9][6] ), .ZN(n8343) );
  AOI22_X1 U12215 ( .A1(n28193), .A2(\xmem_data[10][6] ), .B1(n28192), .B2(
        \xmem_data[11][6] ), .ZN(n8342) );
  AOI22_X1 U12216 ( .A1(n28195), .A2(\xmem_data[12][6] ), .B1(n28194), .B2(
        \xmem_data[13][6] ), .ZN(n8341) );
  AOI22_X1 U12217 ( .A1(n28196), .A2(\xmem_data[14][6] ), .B1(n3142), .B2(
        \xmem_data[15][6] ), .ZN(n8340) );
  NAND4_X1 U12218 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n8346)
         );
  AOI22_X1 U12219 ( .A1(n28210), .A2(\xmem_data[22][6] ), .B1(n3147), .B2(
        \xmem_data[23][6] ), .ZN(n8344) );
  INV_X1 U12220 ( .A(n8344), .ZN(n8345) );
  NOR2_X1 U12221 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NAND2_X1 U12222 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NOR2_X1 U12223 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  AOI22_X1 U12224 ( .A1(n28177), .A2(n8355), .B1(n8354), .B2(n28215), .ZN(
        n8404) );
  AOI22_X1 U12225 ( .A1(n30248), .A2(\xmem_data[120][6] ), .B1(n30730), .B2(
        \xmem_data[121][6] ), .ZN(n8359) );
  AOI22_X1 U12226 ( .A1(n3241), .A2(\xmem_data[122][6] ), .B1(n28233), .B2(
        \xmem_data[123][6] ), .ZN(n8358) );
  AOI22_X1 U12227 ( .A1(n30745), .A2(\xmem_data[124][6] ), .B1(n28110), .B2(
        \xmem_data[125][6] ), .ZN(n8357) );
  AOI22_X1 U12228 ( .A1(n3240), .A2(\xmem_data[126][6] ), .B1(n28231), .B2(
        \xmem_data[127][6] ), .ZN(n8356) );
  AOI22_X1 U12229 ( .A1(n3167), .A2(\xmem_data[96][6] ), .B1(n3188), .B2(
        \xmem_data[97][6] ), .ZN(n8363) );
  BUF_X2 U12230 ( .A(n15549), .Z(n30062) );
  AOI22_X1 U12231 ( .A1(n30062), .A2(\xmem_data[98][6] ), .B1(n28232), .B2(
        \xmem_data[99][6] ), .ZN(n8362) );
  AOI22_X1 U12232 ( .A1(n30766), .A2(\xmem_data[100][6] ), .B1(n30266), .B2(
        \xmem_data[101][6] ), .ZN(n8361) );
  AOI22_X1 U12233 ( .A1(n3233), .A2(\xmem_data[102][6] ), .B1(n28226), .B2(
        \xmem_data[103][6] ), .ZN(n8360) );
  AOI22_X1 U12234 ( .A1(n29790), .A2(\xmem_data[114][6] ), .B1(n28218), .B2(
        \xmem_data[115][6] ), .ZN(n8365) );
  AOI22_X1 U12235 ( .A1(n29433), .A2(\xmem_data[112][6] ), .B1(n30695), .B2(
        \xmem_data[113][6] ), .ZN(n8364) );
  NAND2_X1 U12236 ( .A1(n28786), .A2(\xmem_data[117][6] ), .ZN(n8367) );
  NAND2_X1 U12237 ( .A1(n28219), .A2(\xmem_data[116][6] ), .ZN(n8366) );
  NAND2_X1 U12238 ( .A1(n8367), .A2(n8366), .ZN(n8376) );
  BUF_X1 U12239 ( .A(n8368), .Z(n28239) );
  AOI22_X1 U12240 ( .A1(n28240), .A2(\xmem_data[104][6] ), .B1(n28239), .B2(
        \xmem_data[105][6] ), .ZN(n8372) );
  AOI22_X1 U12241 ( .A1(n28242), .A2(\xmem_data[106][6] ), .B1(n28241), .B2(
        \xmem_data[107][6] ), .ZN(n8371) );
  AOI22_X1 U12242 ( .A1(n28244), .A2(\xmem_data[108][6] ), .B1(n28194), .B2(
        \xmem_data[109][6] ), .ZN(n8370) );
  AOI22_X1 U12243 ( .A1(n28246), .A2(\xmem_data[110][6] ), .B1(n28245), .B2(
        \xmem_data[111][6] ), .ZN(n8369) );
  NAND4_X1 U12244 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n8375)
         );
  AOI22_X1 U12245 ( .A1(n28220), .A2(\xmem_data[118][6] ), .B1(n24702), .B2(
        \xmem_data[119][6] ), .ZN(n8373) );
  INV_X1 U12246 ( .A(n8373), .ZN(n8374) );
  NOR3_X1 U12247 ( .A1(n8376), .A2(n8375), .A3(n8374), .ZN(n8377) );
  NAND4_X1 U12248 ( .A1(n8379), .A2(n3781), .A3(n8378), .A4(n8377), .ZN(n8380)
         );
  NAND2_X1 U12249 ( .A1(n8380), .A2(n28133), .ZN(n8403) );
  AOI22_X1 U12250 ( .A1(n29628), .A2(\xmem_data[82][6] ), .B1(n28137), .B2(
        \xmem_data[83][6] ), .ZN(n8384) );
  AOI22_X1 U12251 ( .A1(n28136), .A2(\xmem_data[80][6] ), .B1(n29697), .B2(
        \xmem_data[81][6] ), .ZN(n8383) );
  AOI22_X1 U12252 ( .A1(n28139), .A2(\xmem_data[84][6] ), .B1(n27833), .B2(
        \xmem_data[85][6] ), .ZN(n8382) );
  AOI22_X1 U12253 ( .A1(n28140), .A2(\xmem_data[86][6] ), .B1(n3137), .B2(
        \xmem_data[87][6] ), .ZN(n8381) );
  NAND4_X1 U12254 ( .A1(n8384), .A2(n8383), .A3(n8382), .A4(n8381), .ZN(n8400)
         );
  AOI22_X1 U12255 ( .A1(n29602), .A2(\xmem_data[88][6] ), .B1(n29389), .B2(
        \xmem_data[89][6] ), .ZN(n8388) );
  AOI22_X1 U12256 ( .A1(n28153), .A2(\xmem_data[90][6] ), .B1(n28152), .B2(
        \xmem_data[91][6] ), .ZN(n8387) );
  AOI22_X1 U12257 ( .A1(n29395), .A2(\xmem_data[92][6] ), .B1(n29739), .B2(
        \xmem_data[93][6] ), .ZN(n8386) );
  AOI22_X1 U12258 ( .A1(n28155), .A2(\xmem_data[94][6] ), .B1(n28154), .B2(
        \xmem_data[95][6] ), .ZN(n8385) );
  NAND4_X1 U12259 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n8399)
         );
  AOI22_X1 U12260 ( .A1(n30075), .A2(n20682), .B1(n28147), .B2(
        \xmem_data[67][6] ), .ZN(n8392) );
  AOI22_X1 U12261 ( .A1(n3166), .A2(\xmem_data[64][6] ), .B1(n3189), .B2(
        \xmem_data[65][6] ), .ZN(n8391) );
  AOI22_X1 U12262 ( .A1(n28173), .A2(\xmem_data[68][6] ), .B1(n29487), .B2(
        \xmem_data[69][6] ), .ZN(n8390) );
  AOI22_X1 U12263 ( .A1(n28151), .A2(\xmem_data[70][6] ), .B1(n23724), .B2(
        \xmem_data[71][6] ), .ZN(n8389) );
  NAND4_X1 U12264 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n8398)
         );
  AOI22_X1 U12265 ( .A1(n28160), .A2(\xmem_data[72][6] ), .B1(n28159), .B2(
        \xmem_data[73][6] ), .ZN(n8396) );
  AOI22_X1 U12266 ( .A1(n28161), .A2(\xmem_data[74][6] ), .B1(n30674), .B2(
        \xmem_data[75][6] ), .ZN(n8395) );
  AOI22_X1 U12267 ( .A1(n28163), .A2(\xmem_data[76][6] ), .B1(n28162), .B2(
        \xmem_data[77][6] ), .ZN(n8394) );
  AOI22_X1 U12268 ( .A1(n28165), .A2(\xmem_data[78][6] ), .B1(n28164), .B2(
        \xmem_data[79][6] ), .ZN(n8393) );
  NAND4_X1 U12269 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n8397)
         );
  XNOR2_X1 U12270 ( .A(n35110), .B(\fmem_data[31][3] ), .ZN(n29210) );
  XOR2_X1 U12271 ( .A(\fmem_data[31][2] ), .B(\fmem_data[31][3] ), .Z(n8405)
         );
  OAI22_X1 U12272 ( .A1(n30364), .A2(n34470), .B1(n29210), .B2(n34468), .ZN(
        n34273) );
  INV_X1 U12273 ( .A(\add_x_2/A[0] ), .ZN(n8410) );
  XOR2_X1 U12274 ( .A(n8407), .B(load_xaddr_val[6]), .Z(n8483) );
  INV_X1 U12275 ( .A(n8483), .ZN(n37315) );
  HA_X1 U12276 ( .A(n8408), .B(n37191), .CO(n8407), .S(n38992) );
  AND2_X1 U12277 ( .A1(n37315), .A2(n38992), .ZN(n29937) );
  NOR2_X1 U12278 ( .A1(n8422), .A2(n3248), .ZN(n8421) );
  INV_X1 U12279 ( .A(n8423), .ZN(n38990) );
  NAND2_X1 U12280 ( .A1(n8421), .A2(n38990), .ZN(n8440) );
  INV_X1 U12281 ( .A(n10589), .ZN(n8414) );
  NOR3_X1 U12282 ( .A1(n6486), .A2(n8416), .A3(n10589), .ZN(n8411) );
  NAND2_X1 U12283 ( .A1(n6172), .A2(n8411), .ZN(n8413) );
  NAND2_X1 U12284 ( .A1(n8417), .A2(n10589), .ZN(n8412) );
  NOR2_X1 U12285 ( .A1(n8417), .A2(n8416), .ZN(n8419) );
  XNOR2_X1 U12286 ( .A(n8419), .B(n8418), .ZN(n8429) );
  OR2_X2 U12287 ( .A1(n8448), .A2(n8420), .ZN(n8424) );
  NOR2_X1 U12288 ( .A1(n8440), .A2(n8424), .ZN(n8484) );
  BUF_X1 U12289 ( .A(n8484), .Z(n29849) );
  INV_X1 U12290 ( .A(n8422), .ZN(n37198) );
  NAND3_X1 U12291 ( .A1(n3248), .A2(n38990), .A3(n37198), .ZN(n8441) );
  NOR2_X1 U12292 ( .A1(n8424), .A2(n8441), .ZN(n8485) );
  BUF_X1 U12293 ( .A(n8485), .Z(n29848) );
  AOI22_X1 U12294 ( .A1(n29849), .A2(\xmem_data[32][5] ), .B1(n29848), .B2(
        \xmem_data[33][5] ), .ZN(n8428) );
  NAND3_X1 U12295 ( .A1(n8422), .A2(n38990), .A3(n6173), .ZN(n8442) );
  NOR2_X1 U12296 ( .A1(n8424), .A2(n8442), .ZN(n8486) );
  BUF_X1 U12297 ( .A(n8486), .Z(n29851) );
  NAND3_X1 U12298 ( .A1(n8422), .A2(n8410), .A3(n38990), .ZN(n8443) );
  NOR2_X1 U12299 ( .A1(n8424), .A2(n8443), .ZN(n8487) );
  BUF_X1 U12300 ( .A(n8487), .Z(n29850) );
  AOI22_X1 U12301 ( .A1(n29851), .A2(\xmem_data[34][5] ), .B1(n29850), .B2(
        \xmem_data[35][5] ), .ZN(n8427) );
  NAND2_X1 U12302 ( .A1(n8423), .A2(n8421), .ZN(n8444) );
  NOR2_X1 U12303 ( .A1(n8424), .A2(n8444), .ZN(n8488) );
  BUF_X1 U12304 ( .A(n8488), .Z(n29853) );
  NAND3_X1 U12305 ( .A1(n8423), .A2(n3248), .A3(n37198), .ZN(n8445) );
  NOR2_X1 U12306 ( .A1(n8424), .A2(n8445), .ZN(n11699) );
  BUF_X1 U12307 ( .A(n11699), .Z(n29852) );
  AOI22_X1 U12308 ( .A1(n29853), .A2(\xmem_data[36][5] ), .B1(n29852), .B2(
        \xmem_data[37][5] ), .ZN(n8426) );
  NAND3_X1 U12309 ( .A1(n8422), .A2(n8423), .A3(n6173), .ZN(n8447) );
  NOR2_X1 U12310 ( .A1(n8424), .A2(n8447), .ZN(n8489) );
  NAND3_X1 U12311 ( .A1(n8423), .A2(n8422), .A3(n3248), .ZN(n8449) );
  NOR2_X1 U12312 ( .A1(n8424), .A2(n8449), .ZN(n11700) );
  AOI22_X1 U12313 ( .A1(n29855), .A2(\xmem_data[38][5] ), .B1(n29854), .B2(
        \xmem_data[39][5] ), .ZN(n8425) );
  NAND4_X1 U12314 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n8425), .ZN(n8459)
         );
  NOR2_X1 U12315 ( .A1(n8440), .A2(n8430), .ZN(n8494) );
  BUF_X1 U12316 ( .A(n8494), .Z(n29860) );
  NOR2_X1 U12317 ( .A1(n8441), .A2(n8430), .ZN(n8464) );
  BUF_X1 U12318 ( .A(n8464), .Z(n29942) );
  AOI22_X1 U12319 ( .A1(n29860), .A2(\xmem_data[40][5] ), .B1(n29942), .B2(
        \xmem_data[41][5] ), .ZN(n8434) );
  NOR2_X1 U12320 ( .A1(n8442), .A2(n8430), .ZN(n8495) );
  BUF_X1 U12321 ( .A(n8495), .Z(n29943) );
  NOR2_X1 U12322 ( .A1(n8443), .A2(n8430), .ZN(n8558) );
  AOI22_X1 U12323 ( .A1(n29943), .A2(\xmem_data[42][5] ), .B1(n3195), .B2(
        \xmem_data[43][5] ), .ZN(n8433) );
  NOR2_X1 U12324 ( .A1(n8444), .A2(n8430), .ZN(n8496) );
  BUF_X1 U12325 ( .A(n8496), .Z(n29945) );
  NOR2_X1 U12326 ( .A1(n8445), .A2(n8430), .ZN(n8601) );
  BUF_X1 U12327 ( .A(n8601), .Z(n29979) );
  AOI22_X1 U12328 ( .A1(n29945), .A2(\xmem_data[44][5] ), .B1(n29979), .B2(
        \xmem_data[45][5] ), .ZN(n8432) );
  NOR2_X1 U12329 ( .A1(n8447), .A2(n8430), .ZN(n8497) );
  BUF_X1 U12330 ( .A(n8497), .Z(n29947) );
  NOR2_X1 U12331 ( .A1(n8449), .A2(n8430), .ZN(n8622) );
  BUF_X1 U12332 ( .A(n8622), .Z(n29981) );
  AOI22_X1 U12333 ( .A1(n29947), .A2(\xmem_data[46][5] ), .B1(n29981), .B2(
        \xmem_data[47][5] ), .ZN(n8431) );
  NAND4_X1 U12334 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n8458)
         );
  NOR2_X1 U12335 ( .A1(n8440), .A2(n8435), .ZN(n8502) );
  BUF_X1 U12336 ( .A(n8502), .Z(n29866) );
  NOR2_X1 U12337 ( .A1(n8441), .A2(n8435), .ZN(n8503) );
  AOI22_X1 U12338 ( .A1(n29866), .A2(\xmem_data[48][5] ), .B1(n29865), .B2(
        \xmem_data[49][5] ), .ZN(n8439) );
  NOR2_X1 U12339 ( .A1(n8442), .A2(n8435), .ZN(n8504) );
  BUF_X1 U12340 ( .A(n8504), .Z(n29868) );
  NOR2_X1 U12341 ( .A1(n8443), .A2(n8435), .ZN(n8505) );
  BUF_X1 U12342 ( .A(n8505), .Z(n29867) );
  AOI22_X1 U12343 ( .A1(n29868), .A2(\xmem_data[50][5] ), .B1(n29867), .B2(
        \xmem_data[51][5] ), .ZN(n8438) );
  NOR2_X1 U12344 ( .A1(n8444), .A2(n8435), .ZN(n8506) );
  BUF_X1 U12345 ( .A(n8506), .Z(n29870) );
  NOR2_X1 U12346 ( .A1(n8445), .A2(n8435), .ZN(n8507) );
  AOI22_X1 U12347 ( .A1(n29870), .A2(\xmem_data[52][5] ), .B1(n29869), .B2(
        \xmem_data[53][5] ), .ZN(n8437) );
  NOR2_X1 U12348 ( .A1(n8447), .A2(n8435), .ZN(n8508) );
  BUF_X1 U12349 ( .A(n8508), .Z(n29871) );
  NOR2_X1 U12350 ( .A1(n8449), .A2(n8435), .ZN(n8537) );
  BUF_X1 U12351 ( .A(n8537), .Z(n29993) );
  AOI22_X1 U12352 ( .A1(n29871), .A2(\xmem_data[54][5] ), .B1(n29993), .B2(
        \xmem_data[55][5] ), .ZN(n8436) );
  NAND4_X1 U12353 ( .A1(n8439), .A2(n8438), .A3(n8437), .A4(n8436), .ZN(n8457)
         );
  NAND2_X1 U12354 ( .A1(n8448), .A2(n8429), .ZN(n8446) );
  NOR2_X1 U12355 ( .A1(n8440), .A2(n8446), .ZN(n8513) );
  BUF_X1 U12356 ( .A(n8513), .Z(n29877) );
  NOR2_X1 U12357 ( .A1(n8441), .A2(n8446), .ZN(n8514) );
  BUF_X1 U12358 ( .A(n8514), .Z(n29876) );
  AOI22_X1 U12359 ( .A1(n29877), .A2(\xmem_data[56][5] ), .B1(n29876), .B2(
        \xmem_data[57][5] ), .ZN(n8455) );
  NOR2_X1 U12360 ( .A1(n8442), .A2(n8446), .ZN(n8515) );
  BUF_X1 U12361 ( .A(n8515), .Z(n29879) );
  NOR2_X1 U12362 ( .A1(n8443), .A2(n8446), .ZN(n8516) );
  BUF_X1 U12363 ( .A(n8516), .Z(n29878) );
  AOI22_X1 U12364 ( .A1(n29879), .A2(\xmem_data[58][5] ), .B1(n29878), .B2(
        \xmem_data[59][5] ), .ZN(n8454) );
  NOR2_X1 U12365 ( .A1(n8444), .A2(n8446), .ZN(n8517) );
  BUF_X1 U12366 ( .A(n8517), .Z(n29881) );
  NOR2_X1 U12367 ( .A1(n8445), .A2(n8446), .ZN(n8518) );
  AOI22_X1 U12368 ( .A1(n29881), .A2(\xmem_data[60][5] ), .B1(n29880), .B2(
        \xmem_data[61][5] ), .ZN(n8453) );
  NOR2_X1 U12369 ( .A1(n8447), .A2(n8446), .ZN(n8519) );
  BUF_X1 U12370 ( .A(n8519), .Z(n29883) );
  INV_X1 U12371 ( .A(n8448), .ZN(n38991) );
  INV_X1 U12372 ( .A(n8449), .ZN(n8450) );
  NAND2_X1 U12373 ( .A1(n8429), .A2(n8450), .ZN(n8451) );
  NOR2_X1 U12374 ( .A1(n38991), .A2(n8451), .ZN(n8520) );
  BUF_X1 U12375 ( .A(n8520), .Z(n29882) );
  AOI22_X1 U12376 ( .A1(n29883), .A2(\xmem_data[62][5] ), .B1(n29882), .B2(
        \xmem_data[63][5] ), .ZN(n8452) );
  NAND4_X1 U12377 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n8456)
         );
  OR4_X1 U12378 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n8482)
         );
  NOR2_X1 U12379 ( .A1(n38992), .A2(n8483), .ZN(n29935) );
  BUF_X1 U12380 ( .A(n8484), .Z(n29893) );
  BUF_X1 U12381 ( .A(n8485), .Z(n29892) );
  AOI22_X1 U12382 ( .A1(n29893), .A2(\xmem_data[0][5] ), .B1(n29892), .B2(
        \xmem_data[1][5] ), .ZN(n8463) );
  BUF_X1 U12383 ( .A(n8486), .Z(n29895) );
  BUF_X1 U12384 ( .A(n8487), .Z(n29894) );
  AOI22_X1 U12385 ( .A1(n29895), .A2(\xmem_data[2][5] ), .B1(n29894), .B2(
        \xmem_data[3][5] ), .ZN(n8462) );
  BUF_X1 U12386 ( .A(n8488), .Z(n29897) );
  BUF_X2 U12387 ( .A(n11699), .Z(n29896) );
  AOI22_X1 U12388 ( .A1(n29897), .A2(\xmem_data[4][5] ), .B1(n29896), .B2(
        \xmem_data[5][5] ), .ZN(n8461) );
  BUF_X1 U12389 ( .A(n8489), .Z(n29899) );
  BUF_X1 U12390 ( .A(n11700), .Z(n29898) );
  AOI22_X1 U12391 ( .A1(n29899), .A2(\xmem_data[6][5] ), .B1(n29898), .B2(
        \xmem_data[7][5] ), .ZN(n8460) );
  NAND4_X1 U12392 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(n8480)
         );
  BUF_X1 U12393 ( .A(n8494), .Z(n29904) );
  AOI22_X1 U12394 ( .A1(n29904), .A2(\xmem_data[8][5] ), .B1(n29976), .B2(
        \xmem_data[9][5] ), .ZN(n8468) );
  BUF_X1 U12395 ( .A(n8495), .Z(n29905) );
  AOI22_X1 U12396 ( .A1(n29905), .A2(\xmem_data[10][5] ), .B1(n3196), .B2(
        \xmem_data[11][5] ), .ZN(n8467) );
  BUF_X1 U12397 ( .A(n8496), .Z(n29907) );
  AOI22_X1 U12398 ( .A1(n29907), .A2(\xmem_data[12][5] ), .B1(n29979), .B2(
        \xmem_data[13][5] ), .ZN(n8466) );
  BUF_X1 U12399 ( .A(n8497), .Z(n29909) );
  BUF_X1 U12400 ( .A(n8622), .Z(n29908) );
  AOI22_X1 U12401 ( .A1(n29909), .A2(\xmem_data[14][5] ), .B1(n29908), .B2(
        \xmem_data[15][5] ), .ZN(n8465) );
  NAND4_X1 U12402 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n8479)
         );
  BUF_X1 U12403 ( .A(n8502), .Z(n29915) );
  BUF_X1 U12404 ( .A(n8503), .Z(n29914) );
  AOI22_X1 U12405 ( .A1(n29915), .A2(\xmem_data[16][5] ), .B1(n29914), .B2(
        \xmem_data[17][5] ), .ZN(n8472) );
  BUF_X1 U12406 ( .A(n8504), .Z(n29917) );
  BUF_X1 U12407 ( .A(n8505), .Z(n29916) );
  AOI22_X1 U12408 ( .A1(n29917), .A2(\xmem_data[18][5] ), .B1(n29916), .B2(
        \xmem_data[19][5] ), .ZN(n8471) );
  BUF_X1 U12409 ( .A(n8507), .Z(n29918) );
  AOI22_X1 U12410 ( .A1(n29919), .A2(\xmem_data[20][5] ), .B1(n29918), .B2(
        \xmem_data[21][5] ), .ZN(n8470) );
  BUF_X1 U12411 ( .A(n8508), .Z(n29921) );
  AOI22_X1 U12412 ( .A1(n29921), .A2(\xmem_data[22][5] ), .B1(n29993), .B2(
        \xmem_data[23][5] ), .ZN(n8469) );
  NAND4_X1 U12413 ( .A1(n8472), .A2(n8471), .A3(n8470), .A4(n8469), .ZN(n8478)
         );
  AOI22_X1 U12414 ( .A1(n3243), .A2(\xmem_data[24][5] ), .B1(n3242), .B2(
        \xmem_data[25][5] ), .ZN(n8476) );
  AOI22_X1 U12415 ( .A1(n3235), .A2(\xmem_data[26][5] ), .B1(n3238), .B2(
        \xmem_data[27][5] ), .ZN(n8475) );
  AOI22_X1 U12416 ( .A1(n3236), .A2(\xmem_data[28][5] ), .B1(n3225), .B2(
        \xmem_data[29][5] ), .ZN(n8474) );
  AOI22_X1 U12417 ( .A1(n3237), .A2(\xmem_data[30][5] ), .B1(n3234), .B2(
        \xmem_data[31][5] ), .ZN(n8473) );
  NAND4_X1 U12418 ( .A1(n8476), .A2(n8475), .A3(n8474), .A4(n8473), .ZN(n8477)
         );
  OR4_X1 U12419 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8477), .ZN(n8481)
         );
  AOI22_X1 U12420 ( .A1(n29937), .A2(n8482), .B1(n29935), .B2(n8481), .ZN(
        n8553) );
  AND2_X1 U12421 ( .A1(n38992), .A2(n8483), .ZN(n30007) );
  BUF_X1 U12422 ( .A(n8484), .Z(n29966) );
  BUF_X1 U12423 ( .A(n8485), .Z(n29965) );
  AOI22_X1 U12424 ( .A1(n29966), .A2(\xmem_data[96][5] ), .B1(n29965), .B2(
        \xmem_data[97][5] ), .ZN(n8493) );
  BUF_X1 U12425 ( .A(n8486), .Z(n29968) );
  BUF_X1 U12426 ( .A(n8487), .Z(n29967) );
  AOI22_X1 U12427 ( .A1(n29968), .A2(\xmem_data[98][5] ), .B1(n29967), .B2(
        \xmem_data[99][5] ), .ZN(n8492) );
  BUF_X1 U12428 ( .A(n8488), .Z(n29969) );
  AOI22_X1 U12429 ( .A1(n29969), .A2(\xmem_data[100][5] ), .B1(n29896), .B2(
        \xmem_data[101][5] ), .ZN(n8491) );
  BUF_X1 U12430 ( .A(n8489), .Z(n29971) );
  BUF_X1 U12431 ( .A(n11700), .Z(n29970) );
  AOI22_X1 U12432 ( .A1(n29971), .A2(\xmem_data[102][5] ), .B1(n29970), .B2(
        \xmem_data[103][5] ), .ZN(n8490) );
  NAND4_X1 U12433 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(n8528)
         );
  BUF_X1 U12434 ( .A(n8494), .Z(n29977) );
  AOI22_X1 U12435 ( .A1(n29977), .A2(\xmem_data[104][5] ), .B1(n29976), .B2(
        \xmem_data[105][5] ), .ZN(n8501) );
  BUF_X1 U12436 ( .A(n8495), .Z(n29978) );
  AOI22_X1 U12437 ( .A1(n29978), .A2(\xmem_data[106][5] ), .B1(n3194), .B2(
        \xmem_data[107][5] ), .ZN(n8500) );
  BUF_X1 U12438 ( .A(n8601), .Z(n29906) );
  AOI22_X1 U12439 ( .A1(n29980), .A2(\xmem_data[108][5] ), .B1(n29906), .B2(
        \xmem_data[109][5] ), .ZN(n8499) );
  AOI22_X1 U12440 ( .A1(n29982), .A2(\xmem_data[110][5] ), .B1(n29908), .B2(
        \xmem_data[111][5] ), .ZN(n8498) );
  NAND4_X1 U12441 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n8527)
         );
  BUF_X1 U12442 ( .A(n8502), .Z(n29988) );
  BUF_X1 U12443 ( .A(n8503), .Z(n29987) );
  AOI22_X1 U12444 ( .A1(n29988), .A2(\xmem_data[112][5] ), .B1(n29987), .B2(
        \xmem_data[113][5] ), .ZN(n8512) );
  BUF_X1 U12445 ( .A(n8504), .Z(n29990) );
  BUF_X1 U12446 ( .A(n8505), .Z(n29989) );
  AOI22_X1 U12447 ( .A1(n29990), .A2(\xmem_data[114][5] ), .B1(n29989), .B2(
        \xmem_data[115][5] ), .ZN(n8511) );
  BUF_X1 U12448 ( .A(n8506), .Z(n29992) );
  AOI22_X1 U12449 ( .A1(n29992), .A2(\xmem_data[116][5] ), .B1(n29991), .B2(
        \xmem_data[117][5] ), .ZN(n8510) );
  BUF_X1 U12450 ( .A(n8508), .Z(n29994) );
  BUF_X1 U12451 ( .A(n8537), .Z(n29952) );
  AOI22_X1 U12452 ( .A1(n29994), .A2(\xmem_data[118][5] ), .B1(n29952), .B2(
        \xmem_data[119][5] ), .ZN(n8509) );
  NAND4_X1 U12453 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n8526)
         );
  AOI22_X1 U12454 ( .A1(n3243), .A2(\xmem_data[120][5] ), .B1(n3242), .B2(
        \xmem_data[121][5] ), .ZN(n8524) );
  AOI22_X1 U12455 ( .A1(n3235), .A2(\xmem_data[122][5] ), .B1(n3238), .B2(
        \xmem_data[123][5] ), .ZN(n8523) );
  AOI22_X1 U12456 ( .A1(n3236), .A2(\xmem_data[124][5] ), .B1(n3225), .B2(
        \xmem_data[125][5] ), .ZN(n8522) );
  AOI22_X1 U12457 ( .A1(n3237), .A2(\xmem_data[126][5] ), .B1(n3234), .B2(
        \xmem_data[127][5] ), .ZN(n8521) );
  NAND4_X1 U12458 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n8525)
         );
  OR4_X1 U12459 ( .A1(n8528), .A2(n8527), .A3(n8526), .A4(n8525), .ZN(n8551)
         );
  NOR2_X1 U12460 ( .A1(n38992), .A2(n37315), .ZN(n30009) );
  AOI22_X1 U12461 ( .A1(n29849), .A2(\xmem_data[64][5] ), .B1(n29848), .B2(
        \xmem_data[65][5] ), .ZN(n8532) );
  AOI22_X1 U12462 ( .A1(n29851), .A2(\xmem_data[66][5] ), .B1(n29850), .B2(
        \xmem_data[67][5] ), .ZN(n8531) );
  AOI22_X1 U12463 ( .A1(n29853), .A2(\xmem_data[68][5] ), .B1(n29852), .B2(
        \xmem_data[69][5] ), .ZN(n8530) );
  AOI22_X1 U12464 ( .A1(n29855), .A2(\xmem_data[70][5] ), .B1(n29854), .B2(
        \xmem_data[71][5] ), .ZN(n8529) );
  NAND4_X1 U12465 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n8549)
         );
  AOI22_X1 U12466 ( .A1(n29860), .A2(\xmem_data[72][5] ), .B1(n29942), .B2(
        \xmem_data[73][5] ), .ZN(n8536) );
  AOI22_X1 U12467 ( .A1(n29943), .A2(\xmem_data[74][5] ), .B1(n3195), .B2(
        \xmem_data[75][5] ), .ZN(n8535) );
  AOI22_X1 U12468 ( .A1(n29945), .A2(\xmem_data[76][5] ), .B1(n29906), .B2(
        \xmem_data[77][5] ), .ZN(n8534) );
  AOI22_X1 U12469 ( .A1(n29947), .A2(\xmem_data[78][5] ), .B1(n29981), .B2(
        \xmem_data[79][5] ), .ZN(n8533) );
  NAND4_X1 U12470 ( .A1(n8536), .A2(n8535), .A3(n8534), .A4(n8533), .ZN(n8548)
         );
  AOI22_X1 U12471 ( .A1(n29866), .A2(\xmem_data[80][5] ), .B1(n29865), .B2(
        \xmem_data[81][5] ), .ZN(n8541) );
  AOI22_X1 U12472 ( .A1(n29868), .A2(\xmem_data[82][5] ), .B1(n29867), .B2(
        \xmem_data[83][5] ), .ZN(n8540) );
  AOI22_X1 U12473 ( .A1(n29870), .A2(\xmem_data[84][5] ), .B1(n29869), .B2(
        \xmem_data[85][5] ), .ZN(n8539) );
  AOI22_X1 U12474 ( .A1(n29871), .A2(\xmem_data[86][5] ), .B1(n29920), .B2(
        \xmem_data[87][5] ), .ZN(n8538) );
  NAND4_X1 U12475 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n8547)
         );
  AOI22_X1 U12476 ( .A1(n29877), .A2(\xmem_data[88][5] ), .B1(n29876), .B2(
        \xmem_data[89][5] ), .ZN(n8545) );
  AOI22_X1 U12477 ( .A1(n29879), .A2(\xmem_data[90][5] ), .B1(n29878), .B2(
        \xmem_data[91][5] ), .ZN(n8544) );
  AOI22_X1 U12478 ( .A1(n29881), .A2(\xmem_data[92][5] ), .B1(n29880), .B2(
        \xmem_data[93][5] ), .ZN(n8543) );
  AOI22_X1 U12479 ( .A1(n29883), .A2(\xmem_data[94][5] ), .B1(n29882), .B2(
        \xmem_data[95][5] ), .ZN(n8542) );
  NAND4_X1 U12480 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n8546)
         );
  OR4_X1 U12481 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n8550)
         );
  AOI22_X1 U12482 ( .A1(n30007), .A2(n8551), .B1(n30009), .B2(n8550), .ZN(
        n8552) );
  AOI22_X1 U12483 ( .A1(n29849), .A2(\xmem_data[32][4] ), .B1(n29848), .B2(
        \xmem_data[33][4] ), .ZN(n8557) );
  AOI22_X1 U12484 ( .A1(n29851), .A2(\xmem_data[34][4] ), .B1(n29850), .B2(
        \xmem_data[35][4] ), .ZN(n8556) );
  AOI22_X1 U12485 ( .A1(n29853), .A2(\xmem_data[36][4] ), .B1(n29852), .B2(
        \xmem_data[37][4] ), .ZN(n8555) );
  AOI22_X1 U12486 ( .A1(n29855), .A2(\xmem_data[38][4] ), .B1(n29854), .B2(
        \xmem_data[39][4] ), .ZN(n8554) );
  NAND4_X1 U12487 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n8574)
         );
  AOI22_X1 U12488 ( .A1(n29860), .A2(\xmem_data[40][4] ), .B1(n29976), .B2(
        \xmem_data[41][4] ), .ZN(n8562) );
  AOI22_X1 U12489 ( .A1(n29943), .A2(\xmem_data[42][4] ), .B1(n3196), .B2(
        \xmem_data[43][4] ), .ZN(n8561) );
  AOI22_X1 U12490 ( .A1(n29907), .A2(\xmem_data[44][4] ), .B1(n29979), .B2(
        \xmem_data[45][4] ), .ZN(n8560) );
  AOI22_X1 U12491 ( .A1(n29909), .A2(\xmem_data[46][4] ), .B1(n29981), .B2(
        \xmem_data[47][4] ), .ZN(n8559) );
  NAND4_X1 U12492 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n8573)
         );
  AOI22_X1 U12493 ( .A1(n29866), .A2(\xmem_data[48][4] ), .B1(n29865), .B2(
        \xmem_data[49][4] ), .ZN(n8566) );
  AOI22_X1 U12494 ( .A1(n29868), .A2(\xmem_data[50][4] ), .B1(n29867), .B2(
        \xmem_data[51][4] ), .ZN(n8565) );
  AOI22_X1 U12495 ( .A1(n29870), .A2(\xmem_data[52][4] ), .B1(n29869), .B2(
        \xmem_data[53][4] ), .ZN(n8564) );
  AOI22_X1 U12496 ( .A1(n29871), .A2(\xmem_data[54][4] ), .B1(n29952), .B2(
        \xmem_data[55][4] ), .ZN(n8563) );
  NAND4_X1 U12497 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n8572)
         );
  AOI22_X1 U12498 ( .A1(n29877), .A2(\xmem_data[56][4] ), .B1(n29876), .B2(
        \xmem_data[57][4] ), .ZN(n8570) );
  AOI22_X1 U12499 ( .A1(n29879), .A2(\xmem_data[58][4] ), .B1(n29878), .B2(
        \xmem_data[59][4] ), .ZN(n8569) );
  AOI22_X1 U12500 ( .A1(n29881), .A2(\xmem_data[60][4] ), .B1(n29880), .B2(
        \xmem_data[61][4] ), .ZN(n8568) );
  AOI22_X1 U12501 ( .A1(n29883), .A2(\xmem_data[62][4] ), .B1(n29882), .B2(
        \xmem_data[63][4] ), .ZN(n8567) );
  NAND4_X1 U12502 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n8571)
         );
  OR4_X1 U12503 ( .A1(n8574), .A2(n8573), .A3(n8572), .A4(n8571), .ZN(n8596)
         );
  AOI22_X1 U12504 ( .A1(n29893), .A2(\xmem_data[0][4] ), .B1(n29892), .B2(
        \xmem_data[1][4] ), .ZN(n8578) );
  AOI22_X1 U12505 ( .A1(n29895), .A2(\xmem_data[2][4] ), .B1(n29894), .B2(
        \xmem_data[3][4] ), .ZN(n8577) );
  AOI22_X1 U12506 ( .A1(n29897), .A2(\xmem_data[4][4] ), .B1(n29896), .B2(
        \xmem_data[5][4] ), .ZN(n8576) );
  AOI22_X1 U12507 ( .A1(n29899), .A2(\xmem_data[6][4] ), .B1(n29898), .B2(
        \xmem_data[7][4] ), .ZN(n8575) );
  NAND4_X1 U12508 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n8594)
         );
  AOI22_X1 U12509 ( .A1(n29904), .A2(\xmem_data[8][4] ), .B1(n29976), .B2(
        \xmem_data[9][4] ), .ZN(n8582) );
  AOI22_X1 U12510 ( .A1(n29943), .A2(\xmem_data[10][4] ), .B1(n3196), .B2(
        \xmem_data[11][4] ), .ZN(n8581) );
  AOI22_X1 U12511 ( .A1(n29945), .A2(\xmem_data[12][4] ), .B1(n29906), .B2(
        \xmem_data[13][4] ), .ZN(n8580) );
  AOI22_X1 U12512 ( .A1(n29947), .A2(\xmem_data[14][4] ), .B1(n29908), .B2(
        \xmem_data[15][4] ), .ZN(n8579) );
  NAND4_X1 U12513 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n8593)
         );
  AOI22_X1 U12514 ( .A1(n29915), .A2(\xmem_data[16][4] ), .B1(n29914), .B2(
        \xmem_data[17][4] ), .ZN(n8586) );
  AOI22_X1 U12515 ( .A1(n29917), .A2(\xmem_data[18][4] ), .B1(n29916), .B2(
        \xmem_data[19][4] ), .ZN(n8585) );
  AOI22_X1 U12516 ( .A1(n29919), .A2(\xmem_data[20][4] ), .B1(n29918), .B2(
        \xmem_data[21][4] ), .ZN(n8584) );
  AOI22_X1 U12517 ( .A1(n29921), .A2(\xmem_data[22][4] ), .B1(n29952), .B2(
        \xmem_data[23][4] ), .ZN(n8583) );
  NAND4_X1 U12518 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n8592)
         );
  AOI22_X1 U12519 ( .A1(n3243), .A2(\xmem_data[24][4] ), .B1(n3242), .B2(
        \xmem_data[25][4] ), .ZN(n8590) );
  AOI22_X1 U12520 ( .A1(n3235), .A2(\xmem_data[26][4] ), .B1(n3238), .B2(
        \xmem_data[27][4] ), .ZN(n8589) );
  AOI22_X1 U12521 ( .A1(n3236), .A2(\xmem_data[28][4] ), .B1(n3225), .B2(
        \xmem_data[29][4] ), .ZN(n8588) );
  AOI22_X1 U12522 ( .A1(n3237), .A2(\xmem_data[30][4] ), .B1(n3234), .B2(
        \xmem_data[31][4] ), .ZN(n8587) );
  NAND4_X1 U12523 ( .A1(n8590), .A2(n8589), .A3(n8588), .A4(n8587), .ZN(n8591)
         );
  OR4_X1 U12524 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(n8595)
         );
  AOI22_X1 U12525 ( .A1(n29937), .A2(n8596), .B1(n29935), .B2(n8595), .ZN(
        n8642) );
  AOI22_X1 U12526 ( .A1(n29966), .A2(\xmem_data[96][4] ), .B1(n29965), .B2(
        \xmem_data[97][4] ), .ZN(n8600) );
  AOI22_X1 U12527 ( .A1(n29968), .A2(\xmem_data[98][4] ), .B1(n29967), .B2(
        \xmem_data[99][4] ), .ZN(n8599) );
  AOI22_X1 U12528 ( .A1(n29969), .A2(\xmem_data[100][4] ), .B1(n29896), .B2(
        \xmem_data[101][4] ), .ZN(n8598) );
  AOI22_X1 U12529 ( .A1(n29971), .A2(\xmem_data[102][4] ), .B1(n29970), .B2(
        \xmem_data[103][4] ), .ZN(n8597) );
  NAND4_X1 U12530 ( .A1(n8600), .A2(n8599), .A3(n8598), .A4(n8597), .ZN(n8617)
         );
  AOI22_X1 U12531 ( .A1(n29977), .A2(\xmem_data[104][4] ), .B1(n29942), .B2(
        \xmem_data[105][4] ), .ZN(n8605) );
  AOI22_X1 U12532 ( .A1(n29978), .A2(\xmem_data[106][4] ), .B1(n3195), .B2(
        \xmem_data[107][4] ), .ZN(n8604) );
  BUF_X1 U12533 ( .A(n8601), .Z(n29944) );
  AOI22_X1 U12534 ( .A1(n29945), .A2(\xmem_data[108][4] ), .B1(n29944), .B2(
        \xmem_data[109][4] ), .ZN(n8603) );
  AOI22_X1 U12535 ( .A1(n29947), .A2(\xmem_data[110][4] ), .B1(n29908), .B2(
        \xmem_data[111][4] ), .ZN(n8602) );
  NAND4_X1 U12536 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n8616)
         );
  AOI22_X1 U12537 ( .A1(n29988), .A2(\xmem_data[112][4] ), .B1(n29987), .B2(
        \xmem_data[113][4] ), .ZN(n8609) );
  AOI22_X1 U12538 ( .A1(n29990), .A2(\xmem_data[114][4] ), .B1(n29989), .B2(
        \xmem_data[115][4] ), .ZN(n8608) );
  AOI22_X1 U12539 ( .A1(n29992), .A2(\xmem_data[116][4] ), .B1(n29991), .B2(
        \xmem_data[117][4] ), .ZN(n8607) );
  AOI22_X1 U12540 ( .A1(n29994), .A2(\xmem_data[118][4] ), .B1(n29920), .B2(
        \xmem_data[119][4] ), .ZN(n8606) );
  NAND4_X1 U12541 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n8615)
         );
  AOI22_X1 U12542 ( .A1(n3243), .A2(\xmem_data[120][4] ), .B1(n3242), .B2(
        \xmem_data[121][4] ), .ZN(n8613) );
  AOI22_X1 U12543 ( .A1(n3235), .A2(\xmem_data[122][4] ), .B1(n3238), .B2(
        \xmem_data[123][4] ), .ZN(n8612) );
  AOI22_X1 U12544 ( .A1(n3236), .A2(\xmem_data[124][4] ), .B1(n3225), .B2(
        \xmem_data[125][4] ), .ZN(n8611) );
  AOI22_X1 U12545 ( .A1(n3237), .A2(\xmem_data[126][4] ), .B1(n3234), .B2(
        \xmem_data[127][4] ), .ZN(n8610) );
  NAND4_X1 U12546 ( .A1(n8613), .A2(n8612), .A3(n8611), .A4(n8610), .ZN(n8614)
         );
  OR4_X1 U12547 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n8640)
         );
  AOI22_X1 U12548 ( .A1(n29849), .A2(\xmem_data[64][4] ), .B1(n29848), .B2(
        \xmem_data[65][4] ), .ZN(n8621) );
  AOI22_X1 U12549 ( .A1(n29851), .A2(\xmem_data[66][4] ), .B1(n29850), .B2(
        \xmem_data[67][4] ), .ZN(n8620) );
  AOI22_X1 U12550 ( .A1(n29853), .A2(\xmem_data[68][4] ), .B1(n29852), .B2(
        \xmem_data[69][4] ), .ZN(n8619) );
  AOI22_X1 U12551 ( .A1(n29855), .A2(\xmem_data[70][4] ), .B1(n29854), .B2(
        \xmem_data[71][4] ), .ZN(n8618) );
  NAND4_X1 U12552 ( .A1(n8621), .A2(n8620), .A3(n8619), .A4(n8618), .ZN(n8638)
         );
  AOI22_X1 U12553 ( .A1(n29860), .A2(\xmem_data[72][4] ), .B1(n29942), .B2(
        \xmem_data[73][4] ), .ZN(n8626) );
  AOI22_X1 U12554 ( .A1(n29943), .A2(\xmem_data[74][4] ), .B1(n3195), .B2(
        \xmem_data[75][4] ), .ZN(n8625) );
  AOI22_X1 U12555 ( .A1(n29945), .A2(\xmem_data[76][4] ), .B1(n29944), .B2(
        \xmem_data[77][4] ), .ZN(n8624) );
  BUF_X1 U12556 ( .A(n8622), .Z(n29946) );
  AOI22_X1 U12557 ( .A1(n29947), .A2(\xmem_data[78][4] ), .B1(n29946), .B2(
        \xmem_data[79][4] ), .ZN(n8623) );
  NAND4_X1 U12558 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(n8637)
         );
  AOI22_X1 U12559 ( .A1(n29866), .A2(\xmem_data[80][4] ), .B1(n29865), .B2(
        \xmem_data[81][4] ), .ZN(n8630) );
  AOI22_X1 U12560 ( .A1(n29868), .A2(\xmem_data[82][4] ), .B1(n29867), .B2(
        \xmem_data[83][4] ), .ZN(n8629) );
  AOI22_X1 U12561 ( .A1(n29870), .A2(\xmem_data[84][4] ), .B1(n29869), .B2(
        \xmem_data[85][4] ), .ZN(n8628) );
  AOI22_X1 U12562 ( .A1(n29871), .A2(\xmem_data[86][4] ), .B1(n29993), .B2(
        \xmem_data[87][4] ), .ZN(n8627) );
  NAND4_X1 U12563 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n8636)
         );
  AOI22_X1 U12564 ( .A1(n29877), .A2(\xmem_data[88][4] ), .B1(n29876), .B2(
        \xmem_data[89][4] ), .ZN(n8634) );
  AOI22_X1 U12565 ( .A1(n29879), .A2(\xmem_data[90][4] ), .B1(n29878), .B2(
        \xmem_data[91][4] ), .ZN(n8633) );
  AOI22_X1 U12566 ( .A1(n29881), .A2(\xmem_data[92][4] ), .B1(n29880), .B2(
        \xmem_data[93][4] ), .ZN(n8632) );
  AOI22_X1 U12567 ( .A1(n29883), .A2(\xmem_data[94][4] ), .B1(n29882), .B2(
        \xmem_data[95][4] ), .ZN(n8631) );
  NAND4_X1 U12568 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), .ZN(n8635)
         );
  AOI22_X1 U12569 ( .A1(n30007), .A2(n8640), .B1(n30009), .B2(n8639), .ZN(
        n8641) );
  NAND2_X1 U12570 ( .A1(n8642), .A2(n8641), .ZN(n32176) );
  XOR2_X1 U12571 ( .A(\fmem_data[1][4] ), .B(\fmem_data[1][5] ), .Z(n8643) );
  AOI22_X1 U12572 ( .A1(n30743), .A2(\xmem_data[88][3] ), .B1(n29589), .B2(
        \xmem_data[89][3] ), .ZN(n8654) );
  AOI22_X1 U12573 ( .A1(n30635), .A2(\xmem_data[92][3] ), .B1(n30237), .B2(
        \xmem_data[93][3] ), .ZN(n8653) );
  AOI22_X1 U12574 ( .A1(n28240), .A2(\xmem_data[72][3] ), .B1(n28239), .B2(
        \xmem_data[73][3] ), .ZN(n8647) );
  AOI22_X1 U12575 ( .A1(n28242), .A2(\xmem_data[74][3] ), .B1(n28241), .B2(
        \xmem_data[75][3] ), .ZN(n8646) );
  AOI22_X1 U12576 ( .A1(n28244), .A2(\xmem_data[76][3] ), .B1(n28243), .B2(
        \xmem_data[77][3] ), .ZN(n8645) );
  AOI22_X1 U12577 ( .A1(n28246), .A2(\xmem_data[78][3] ), .B1(n28245), .B2(
        \xmem_data[79][3] ), .ZN(n8644) );
  NAND4_X1 U12578 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .ZN(n8651)
         );
  AOI22_X1 U12579 ( .A1(n3240), .A2(\xmem_data[94][3] ), .B1(n28231), .B2(
        \xmem_data[95][3] ), .ZN(n8649) );
  AOI22_X1 U12580 ( .A1(n3241), .A2(\xmem_data[90][3] ), .B1(n28233), .B2(
        \xmem_data[91][3] ), .ZN(n8648) );
  NAND2_X1 U12581 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  NOR2_X1 U12582 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  NAND3_X1 U12583 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n8665) );
  AOI22_X1 U12584 ( .A1(n30279), .A2(\xmem_data[82][3] ), .B1(n28218), .B2(
        \xmem_data[83][3] ), .ZN(n8658) );
  AOI22_X1 U12585 ( .A1(n29433), .A2(\xmem_data[80][3] ), .B1(n27832), .B2(
        \xmem_data[81][3] ), .ZN(n8657) );
  AOI22_X1 U12586 ( .A1(n28219), .A2(\xmem_data[84][3] ), .B1(n28786), .B2(
        \xmem_data[85][3] ), .ZN(n8656) );
  AOI22_X1 U12587 ( .A1(n28220), .A2(\xmem_data[86][3] ), .B1(n25417), .B2(
        \xmem_data[87][3] ), .ZN(n8655) );
  NAND4_X1 U12588 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n8664)
         );
  AOI22_X1 U12589 ( .A1(n3164), .A2(\xmem_data[64][3] ), .B1(n3185), .B2(
        \xmem_data[65][3] ), .ZN(n8662) );
  AOI22_X1 U12590 ( .A1(n30684), .A2(\xmem_data[66][3] ), .B1(n28232), .B2(
        \xmem_data[67][3] ), .ZN(n8661) );
  AOI22_X1 U12591 ( .A1(n28173), .A2(\xmem_data[68][3] ), .B1(n30716), .B2(
        \xmem_data[69][3] ), .ZN(n8660) );
  AOI22_X1 U12592 ( .A1(n3233), .A2(\xmem_data[70][3] ), .B1(n28226), .B2(
        \xmem_data[71][3] ), .ZN(n8659) );
  NAND4_X1 U12593 ( .A1(n8662), .A2(n8661), .A3(n8660), .A4(n8659), .ZN(n8663)
         );
  OR3_X1 U12594 ( .A1(n8665), .A2(n8664), .A3(n8663), .ZN(n8687) );
  AOI22_X1 U12595 ( .A1(n30633), .A2(\xmem_data[120][3] ), .B1(n28665), .B2(
        \xmem_data[121][3] ), .ZN(n8669) );
  AOI22_X1 U12596 ( .A1(n3241), .A2(\xmem_data[122][3] ), .B1(n28233), .B2(
        \xmem_data[123][3] ), .ZN(n8668) );
  AOI22_X1 U12597 ( .A1(n29769), .A2(\xmem_data[124][3] ), .B1(n27753), .B2(
        \xmem_data[125][3] ), .ZN(n8667) );
  AOI22_X1 U12598 ( .A1(n3240), .A2(\xmem_data[126][3] ), .B1(n28231), .B2(
        \xmem_data[127][3] ), .ZN(n8666) );
  NAND4_X1 U12599 ( .A1(n8669), .A2(n8668), .A3(n8667), .A4(n8666), .ZN(n8685)
         );
  AOI22_X1 U12600 ( .A1(n29788), .A2(\xmem_data[112][3] ), .B1(n27013), .B2(
        \xmem_data[113][3] ), .ZN(n8673) );
  AOI22_X1 U12601 ( .A1(n3392), .A2(\xmem_data[114][3] ), .B1(n28218), .B2(
        \xmem_data[115][3] ), .ZN(n8672) );
  AOI22_X1 U12602 ( .A1(n28219), .A2(\xmem_data[116][3] ), .B1(n30293), .B2(
        \xmem_data[117][3] ), .ZN(n8671) );
  AOI22_X1 U12603 ( .A1(n28220), .A2(\xmem_data[118][3] ), .B1(n28308), .B2(
        \xmem_data[119][3] ), .ZN(n8670) );
  NAND4_X1 U12604 ( .A1(n8673), .A2(n8672), .A3(n8671), .A4(n8670), .ZN(n8684)
         );
  AOI22_X1 U12605 ( .A1(n3165), .A2(\xmem_data[96][3] ), .B1(n3183), .B2(
        \xmem_data[97][3] ), .ZN(n8677) );
  AOI22_X1 U12606 ( .A1(n29476), .A2(\xmem_data[98][3] ), .B1(n28232), .B2(
        \xmem_data[99][3] ), .ZN(n8676) );
  AOI22_X1 U12607 ( .A1(n28173), .A2(\xmem_data[100][3] ), .B1(n30716), .B2(
        \xmem_data[101][3] ), .ZN(n8675) );
  AOI22_X1 U12608 ( .A1(n3233), .A2(\xmem_data[102][3] ), .B1(n28226), .B2(
        \xmem_data[103][3] ), .ZN(n8674) );
  NAND4_X1 U12609 ( .A1(n8677), .A2(n8676), .A3(n8675), .A4(n8674), .ZN(n8683)
         );
  AOI22_X1 U12610 ( .A1(n28240), .A2(\xmem_data[104][3] ), .B1(n28239), .B2(
        \xmem_data[105][3] ), .ZN(n8681) );
  AOI22_X1 U12611 ( .A1(n28242), .A2(\xmem_data[106][3] ), .B1(n28241), .B2(
        \xmem_data[107][3] ), .ZN(n8680) );
  AOI22_X1 U12612 ( .A1(n28244), .A2(\xmem_data[108][3] ), .B1(n28243), .B2(
        \xmem_data[109][3] ), .ZN(n8679) );
  AOI22_X1 U12613 ( .A1(n28246), .A2(\xmem_data[110][3] ), .B1(n28245), .B2(
        \xmem_data[111][3] ), .ZN(n8678) );
  NAND4_X1 U12614 ( .A1(n8681), .A2(n8680), .A3(n8679), .A4(n8678), .ZN(n8682)
         );
  AOI22_X1 U12615 ( .A1(n8687), .A2(n28258), .B1(n8686), .B2(n28133), .ZN(
        n8732) );
  AOI22_X1 U12616 ( .A1(n3161), .A2(\xmem_data[32][3] ), .B1(n3184), .B2(
        \xmem_data[33][3] ), .ZN(n8691) );
  AOI22_X1 U12617 ( .A1(n30715), .A2(\xmem_data[34][3] ), .B1(n28147), .B2(
        \xmem_data[35][3] ), .ZN(n8690) );
  AOI22_X1 U12618 ( .A1(n30717), .A2(\xmem_data[36][3] ), .B1(n29640), .B2(
        \xmem_data[37][3] ), .ZN(n8689) );
  AOI22_X1 U12619 ( .A1(n28151), .A2(\xmem_data[38][3] ), .B1(n28461), .B2(
        \xmem_data[39][3] ), .ZN(n8688) );
  NAND4_X1 U12620 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n8708)
         );
  AOI22_X1 U12621 ( .A1(n28160), .A2(\xmem_data[40][3] ), .B1(n28159), .B2(
        \xmem_data[41][3] ), .ZN(n8695) );
  AOI22_X1 U12622 ( .A1(n28161), .A2(\xmem_data[42][3] ), .B1(n13420), .B2(
        \xmem_data[43][3] ), .ZN(n8694) );
  AOI22_X1 U12623 ( .A1(n28163), .A2(\xmem_data[44][3] ), .B1(n28162), .B2(
        \xmem_data[45][3] ), .ZN(n8693) );
  AOI22_X1 U12624 ( .A1(n28165), .A2(\xmem_data[46][3] ), .B1(n28164), .B2(
        \xmem_data[47][3] ), .ZN(n8692) );
  NAND4_X1 U12625 ( .A1(n8695), .A2(n8694), .A3(n8693), .A4(n8692), .ZN(n8707)
         );
  AOI22_X1 U12626 ( .A1(n29421), .A2(\xmem_data[48][3] ), .B1(n29432), .B2(
        \xmem_data[49][3] ), .ZN(n8699) );
  AOI22_X1 U12627 ( .A1(n29699), .A2(\xmem_data[50][3] ), .B1(n28137), .B2(
        \xmem_data[51][3] ), .ZN(n8698) );
  AOI22_X1 U12628 ( .A1(n28139), .A2(\xmem_data[52][3] ), .B1(n28786), .B2(
        \xmem_data[53][3] ), .ZN(n8697) );
  AOI22_X1 U12629 ( .A1(n28140), .A2(\xmem_data[54][3] ), .B1(n25377), .B2(
        \xmem_data[55][3] ), .ZN(n8696) );
  NAND4_X1 U12630 ( .A1(n8699), .A2(n8698), .A3(n8697), .A4(n8696), .ZN(n8706)
         );
  AOI22_X1 U12631 ( .A1(n29602), .A2(\xmem_data[56][3] ), .B1(n28738), .B2(
        \xmem_data[57][3] ), .ZN(n8704) );
  AOI22_X1 U12632 ( .A1(n28153), .A2(\xmem_data[58][3] ), .B1(n28152), .B2(
        \xmem_data[59][3] ), .ZN(n8703) );
  BUF_X1 U12633 ( .A(n8700), .Z(n28684) );
  AOI22_X1 U12634 ( .A1(n28685), .A2(\xmem_data[60][3] ), .B1(n27753), .B2(
        \xmem_data[61][3] ), .ZN(n8702) );
  AOI22_X1 U12635 ( .A1(n28155), .A2(\xmem_data[62][3] ), .B1(n28154), .B2(
        \xmem_data[63][3] ), .ZN(n8701) );
  NAND4_X1 U12636 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n8705)
         );
  OR4_X1 U12637 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n8730)
         );
  AOI22_X1 U12638 ( .A1(n3165), .A2(\xmem_data[0][3] ), .B1(n3186), .B2(
        \xmem_data[1][3] ), .ZN(n8712) );
  AOI22_X1 U12639 ( .A1(n30062), .A2(\xmem_data[2][3] ), .B1(n28232), .B2(
        \xmem_data[3][3] ), .ZN(n8711) );
  AOI22_X1 U12640 ( .A1(n30076), .A2(\xmem_data[4][3] ), .B1(n29640), .B2(
        \xmem_data[5][3] ), .ZN(n8710) );
  AOI22_X1 U12641 ( .A1(n3233), .A2(\xmem_data[6][3] ), .B1(n28202), .B2(
        \xmem_data[7][3] ), .ZN(n8709) );
  NAND4_X1 U12642 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n8728)
         );
  AOI22_X1 U12643 ( .A1(n28191), .A2(\xmem_data[8][3] ), .B1(n28190), .B2(
        \xmem_data[9][3] ), .ZN(n8716) );
  AOI22_X1 U12644 ( .A1(n28193), .A2(\xmem_data[10][3] ), .B1(n28192), .B2(
        \xmem_data[11][3] ), .ZN(n8715) );
  AOI22_X1 U12645 ( .A1(n28195), .A2(\xmem_data[12][3] ), .B1(n28194), .B2(
        \xmem_data[13][3] ), .ZN(n8714) );
  AOI22_X1 U12646 ( .A1(n28196), .A2(\xmem_data[14][3] ), .B1(n3149), .B2(
        \xmem_data[15][3] ), .ZN(n8713) );
  NAND4_X1 U12647 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n8727)
         );
  AOI22_X1 U12648 ( .A1(n27740), .A2(\xmem_data[18][3] ), .B1(n27708), .B2(
        \xmem_data[19][3] ), .ZN(n8720) );
  AOI22_X1 U12649 ( .A1(n30708), .A2(\xmem_data[16][3] ), .B1(n30695), .B2(
        \xmem_data[17][3] ), .ZN(n8719) );
  AOI22_X1 U12650 ( .A1(n28209), .A2(\xmem_data[20][3] ), .B1(n30217), .B2(
        \xmem_data[21][3] ), .ZN(n8718) );
  AOI22_X1 U12651 ( .A1(n28210), .A2(\xmem_data[22][3] ), .B1(n30295), .B2(
        \xmem_data[23][3] ), .ZN(n8717) );
  NAND4_X1 U12652 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n8726)
         );
  AOI22_X1 U12653 ( .A1(n29705), .A2(\xmem_data[24][3] ), .B1(n29482), .B2(
        \xmem_data[25][3] ), .ZN(n8724) );
  AOI22_X1 U12654 ( .A1(n3241), .A2(\xmem_data[26][3] ), .B1(n30663), .B2(
        \xmem_data[27][3] ), .ZN(n8723) );
  AOI22_X1 U12655 ( .A1(n29436), .A2(\xmem_data[28][3] ), .B1(n29648), .B2(
        \xmem_data[29][3] ), .ZN(n8722) );
  AOI22_X1 U12656 ( .A1(n3240), .A2(\xmem_data[30][3] ), .B1(n28091), .B2(
        \xmem_data[31][3] ), .ZN(n8721) );
  NAND4_X1 U12657 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8721), .ZN(n8725)
         );
  AOI22_X1 U12658 ( .A1(n28177), .A2(n8730), .B1(n28215), .B2(n8729), .ZN(
        n8731) );
  XNOR2_X1 U12659 ( .A(n3303), .B(\fmem_data[31][7] ), .ZN(n31975) );
  AOI22_X1 U12660 ( .A1(n28139), .A2(\xmem_data[52][2] ), .B1(n3198), .B2(
        \xmem_data[53][2] ), .ZN(n8733) );
  INV_X1 U12661 ( .A(n8733), .ZN(n8736) );
  AOI22_X1 U12662 ( .A1(n30248), .A2(\xmem_data[56][2] ), .B1(n3368), .B2(
        \xmem_data[57][2] ), .ZN(n8734) );
  INV_X1 U12663 ( .A(n8734), .ZN(n8735) );
  AOI22_X1 U12664 ( .A1(n30215), .A2(\xmem_data[50][2] ), .B1(n28137), .B2(
        \xmem_data[51][2] ), .ZN(n8738) );
  AOI22_X1 U12665 ( .A1(n29421), .A2(\xmem_data[48][2] ), .B1(n30695), .B2(
        \xmem_data[49][2] ), .ZN(n8737) );
  AOI22_X1 U12666 ( .A1(n29395), .A2(\xmem_data[60][2] ), .B1(n30084), .B2(
        \xmem_data[61][2] ), .ZN(n8739) );
  INV_X1 U12667 ( .A(n8739), .ZN(n8749) );
  AOI22_X1 U12668 ( .A1(n28160), .A2(\xmem_data[40][2] ), .B1(n28159), .B2(
        \xmem_data[41][2] ), .ZN(n8743) );
  AOI22_X1 U12669 ( .A1(n28161), .A2(\xmem_data[42][2] ), .B1(n20952), .B2(
        \xmem_data[43][2] ), .ZN(n8742) );
  AOI22_X1 U12670 ( .A1(n28163), .A2(\xmem_data[44][2] ), .B1(n28162), .B2(
        \xmem_data[45][2] ), .ZN(n8741) );
  AOI22_X1 U12671 ( .A1(n28165), .A2(\xmem_data[46][2] ), .B1(n28164), .B2(
        \xmem_data[47][2] ), .ZN(n8740) );
  NAND4_X1 U12672 ( .A1(n8743), .A2(n8742), .A3(n8741), .A4(n8740), .ZN(n8748)
         );
  AOI22_X1 U12673 ( .A1(n28153), .A2(\xmem_data[58][2] ), .B1(n28152), .B2(
        \xmem_data[59][2] ), .ZN(n8746) );
  AOI22_X1 U12674 ( .A1(n28140), .A2(\xmem_data[54][2] ), .B1(n20808), .B2(
        \xmem_data[55][2] ), .ZN(n8745) );
  AOI22_X1 U12675 ( .A1(n28155), .A2(\xmem_data[62][2] ), .B1(n28154), .B2(
        \xmem_data[63][2] ), .ZN(n8744) );
  NOR3_X1 U12676 ( .A1(n8749), .A2(n8748), .A3(n8747), .ZN(n8754) );
  AOI22_X1 U12677 ( .A1(n3162), .A2(\xmem_data[32][2] ), .B1(n3183), .B2(
        \xmem_data[33][2] ), .ZN(n8753) );
  AOI22_X1 U12678 ( .A1(n30070), .A2(\xmem_data[34][2] ), .B1(n28147), .B2(
        \xmem_data[35][2] ), .ZN(n8752) );
  AOI22_X1 U12679 ( .A1(n28680), .A2(\xmem_data[36][2] ), .B1(n30716), .B2(
        \xmem_data[37][2] ), .ZN(n8751) );
  AOI22_X1 U12680 ( .A1(n28151), .A2(\xmem_data[38][2] ), .B1(n24571), .B2(
        \xmem_data[39][2] ), .ZN(n8750) );
  NAND3_X1 U12681 ( .A1(n8755), .A2(n8754), .A3(n3753), .ZN(n8756) );
  OAI21_X1 U12682 ( .B1(n3992), .B2(n8756), .A(n28177), .ZN(n8832) );
  AOI22_X1 U12683 ( .A1(n29628), .A2(\xmem_data[82][2] ), .B1(n28218), .B2(
        \xmem_data[83][2] ), .ZN(n8757) );
  INV_X1 U12684 ( .A(n8757), .ZN(n8761) );
  AOI22_X1 U12685 ( .A1(n28219), .A2(\xmem_data[84][2] ), .B1(n30696), .B2(
        \xmem_data[85][2] ), .ZN(n8759) );
  AOI22_X1 U12686 ( .A1(n30191), .A2(\xmem_data[88][2] ), .B1(n28738), .B2(
        \xmem_data[89][2] ), .ZN(n8758) );
  NAND2_X1 U12687 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  AOI22_X1 U12688 ( .A1(n28240), .A2(\xmem_data[72][2] ), .B1(n28239), .B2(
        \xmem_data[73][2] ), .ZN(n8765) );
  AOI22_X1 U12689 ( .A1(n28242), .A2(\xmem_data[74][2] ), .B1(n28241), .B2(
        \xmem_data[75][2] ), .ZN(n8764) );
  AOI22_X1 U12690 ( .A1(n28244), .A2(\xmem_data[76][2] ), .B1(n28243), .B2(
        \xmem_data[77][2] ), .ZN(n8763) );
  AOI22_X1 U12691 ( .A1(n28246), .A2(\xmem_data[78][2] ), .B1(n28245), .B2(
        \xmem_data[79][2] ), .ZN(n8762) );
  NAND4_X1 U12692 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n8772)
         );
  AOI22_X1 U12693 ( .A1(n27811), .A2(\xmem_data[92][2] ), .B1(n29768), .B2(
        \xmem_data[93][2] ), .ZN(n8766) );
  INV_X1 U12694 ( .A(n8766), .ZN(n8771) );
  AOI22_X1 U12695 ( .A1(n3241), .A2(\xmem_data[90][2] ), .B1(n28233), .B2(
        \xmem_data[91][2] ), .ZN(n8769) );
  AOI22_X1 U12696 ( .A1(n28220), .A2(\xmem_data[86][2] ), .B1(n3128), .B2(
        \xmem_data[87][2] ), .ZN(n8768) );
  AOI22_X1 U12697 ( .A1(n3240), .A2(\xmem_data[94][2] ), .B1(n28231), .B2(
        \xmem_data[95][2] ), .ZN(n8767) );
  NOR3_X1 U12698 ( .A1(n8772), .A2(n8771), .A3(n8770), .ZN(n8778) );
  AOI22_X1 U12699 ( .A1(n3166), .A2(\xmem_data[64][2] ), .B1(n3186), .B2(
        \xmem_data[65][2] ), .ZN(n8776) );
  AOI22_X1 U12700 ( .A1(n30715), .A2(\xmem_data[66][2] ), .B1(n28232), .B2(
        \xmem_data[67][2] ), .ZN(n8775) );
  AOI22_X1 U12701 ( .A1(n29815), .A2(\xmem_data[68][2] ), .B1(n29640), .B2(
        \xmem_data[69][2] ), .ZN(n8774) );
  AOI22_X1 U12702 ( .A1(n3233), .A2(\xmem_data[70][2] ), .B1(n28226), .B2(
        \xmem_data[71][2] ), .ZN(n8773) );
  AOI22_X1 U12703 ( .A1(n29421), .A2(\xmem_data[80][2] ), .B1(n29432), .B2(
        \xmem_data[81][2] ), .ZN(n8777) );
  NAND3_X1 U12704 ( .A1(n8778), .A2(n3766), .A3(n8777), .ZN(n8779) );
  OAI21_X1 U12705 ( .B1(n8780), .B2(n8779), .A(n28258), .ZN(n8831) );
  AOI22_X1 U12706 ( .A1(\xmem_data[117][2] ), .A2(n30776), .B1(n29602), .B2(
        \xmem_data[120][2] ), .ZN(n8785) );
  AND2_X1 U12707 ( .A1(n28218), .A2(\xmem_data[115][2] ), .ZN(n8781) );
  AOI21_X1 U12708 ( .B1(n28219), .B2(\xmem_data[116][2] ), .A(n8781), .ZN(
        n8784) );
  NAND2_X1 U12709 ( .A1(n28145), .A2(\xmem_data[121][2] ), .ZN(n8783) );
  NAND2_X1 U12710 ( .A1(n28700), .A2(\xmem_data[114][2] ), .ZN(n8782) );
  NAND4_X1 U12711 ( .A1(n8785), .A2(n8784), .A3(n8783), .A4(n8782), .ZN(n8804)
         );
  AOI22_X1 U12712 ( .A1(n28240), .A2(\xmem_data[104][2] ), .B1(n28239), .B2(
        \xmem_data[105][2] ), .ZN(n8789) );
  AOI22_X1 U12713 ( .A1(n28242), .A2(\xmem_data[106][2] ), .B1(n28241), .B2(
        \xmem_data[107][2] ), .ZN(n8788) );
  AOI22_X1 U12714 ( .A1(n28244), .A2(\xmem_data[108][2] ), .B1(n28243), .B2(
        \xmem_data[109][2] ), .ZN(n8787) );
  AOI22_X1 U12715 ( .A1(n28246), .A2(\xmem_data[110][2] ), .B1(n28245), .B2(
        \xmem_data[111][2] ), .ZN(n8786) );
  NAND4_X1 U12716 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8796)
         );
  AOI22_X1 U12717 ( .A1(n30302), .A2(\xmem_data[124][2] ), .B1(n28110), .B2(
        \xmem_data[125][2] ), .ZN(n8790) );
  INV_X1 U12718 ( .A(n8790), .ZN(n8795) );
  AOI22_X1 U12719 ( .A1(n3241), .A2(\xmem_data[122][2] ), .B1(n28233), .B2(
        \xmem_data[123][2] ), .ZN(n8793) );
  AOI22_X1 U12720 ( .A1(n28220), .A2(\xmem_data[118][2] ), .B1(n28084), .B2(
        \xmem_data[119][2] ), .ZN(n8792) );
  AOI22_X1 U12721 ( .A1(n3240), .A2(\xmem_data[126][2] ), .B1(n28231), .B2(
        \xmem_data[127][2] ), .ZN(n8791) );
  NOR3_X1 U12722 ( .A1(n8796), .A2(n8795), .A3(n8794), .ZN(n8802) );
  AOI22_X1 U12723 ( .A1(n3163), .A2(\xmem_data[96][2] ), .B1(n3187), .B2(
        \xmem_data[97][2] ), .ZN(n8800) );
  AOI22_X1 U12724 ( .A1(n29610), .A2(\xmem_data[98][2] ), .B1(n28232), .B2(
        \xmem_data[99][2] ), .ZN(n8799) );
  AOI22_X1 U12725 ( .A1(n29722), .A2(\xmem_data[100][2] ), .B1(n30170), .B2(
        \xmem_data[101][2] ), .ZN(n8798) );
  AOI22_X1 U12726 ( .A1(n3233), .A2(\xmem_data[102][2] ), .B1(n28226), .B2(
        \xmem_data[103][2] ), .ZN(n8797) );
  AOI22_X1 U12727 ( .A1(n29626), .A2(\xmem_data[112][2] ), .B1(n30222), .B2(
        \xmem_data[113][2] ), .ZN(n8801) );
  NAND3_X1 U12728 ( .A1(n8802), .A2(n3759), .A3(n8801), .ZN(n8803) );
  OAI21_X1 U12729 ( .B1(n8804), .B2(n8803), .A(n28133), .ZN(n8830) );
  AOI22_X1 U12730 ( .A1(n30279), .A2(\xmem_data[18][2] ), .B1(n30278), .B2(
        \xmem_data[19][2] ), .ZN(n8806) );
  AOI22_X1 U12731 ( .A1(n28136), .A2(\xmem_data[16][2] ), .B1(n30222), .B2(
        \xmem_data[17][2] ), .ZN(n8805) );
  NAND2_X1 U12732 ( .A1(n8806), .A2(n8805), .ZN(n8812) );
  AOI22_X1 U12733 ( .A1(n3161), .A2(\xmem_data[0][2] ), .B1(n3190), .B2(
        \xmem_data[1][2] ), .ZN(n8810) );
  AOI22_X1 U12734 ( .A1(n29610), .A2(\xmem_data[2][2] ), .B1(n25400), .B2(
        \xmem_data[3][2] ), .ZN(n8809) );
  AOI22_X1 U12735 ( .A1(n30766), .A2(\xmem_data[4][2] ), .B1(n29721), .B2(
        \xmem_data[5][2] ), .ZN(n8808) );
  AOI22_X1 U12736 ( .A1(n3233), .A2(\xmem_data[6][2] ), .B1(n28202), .B2(
        \xmem_data[7][2] ), .ZN(n8807) );
  NAND4_X1 U12737 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n8811)
         );
  OR2_X1 U12738 ( .A1(n8812), .A2(n8811), .ZN(n8828) );
  AOI22_X1 U12739 ( .A1(n29705), .A2(\xmem_data[24][2] ), .B1(n27761), .B2(
        \xmem_data[25][2] ), .ZN(n8816) );
  AOI22_X1 U12740 ( .A1(n3241), .A2(\xmem_data[26][2] ), .B1(n28089), .B2(
        \xmem_data[27][2] ), .ZN(n8815) );
  AOI22_X1 U12741 ( .A1(n3174), .A2(\xmem_data[28][2] ), .B1(n29592), .B2(
        \xmem_data[29][2] ), .ZN(n8814) );
  AOI22_X1 U12742 ( .A1(n3240), .A2(\xmem_data[30][2] ), .B1(n23795), .B2(
        \xmem_data[31][2] ), .ZN(n8813) );
  AOI22_X1 U12743 ( .A1(n28209), .A2(\xmem_data[20][2] ), .B1(n28667), .B2(
        \xmem_data[21][2] ), .ZN(n8817) );
  INV_X1 U12744 ( .A(n8817), .ZN(n8825) );
  AOI22_X1 U12745 ( .A1(n28191), .A2(\xmem_data[8][2] ), .B1(n28190), .B2(
        \xmem_data[9][2] ), .ZN(n8821) );
  AOI22_X1 U12746 ( .A1(n28193), .A2(\xmem_data[10][2] ), .B1(n28192), .B2(
        \xmem_data[11][2] ), .ZN(n8820) );
  AOI22_X1 U12747 ( .A1(n28195), .A2(\xmem_data[12][2] ), .B1(n28194), .B2(
        \xmem_data[13][2] ), .ZN(n8819) );
  AOI22_X1 U12748 ( .A1(n28196), .A2(\xmem_data[14][2] ), .B1(n3333), .B2(
        \xmem_data[15][2] ), .ZN(n8818) );
  NAND4_X1 U12749 ( .A1(n8821), .A2(n8820), .A3(n8819), .A4(n8818), .ZN(n8824)
         );
  AOI22_X1 U12750 ( .A1(n28210), .A2(\xmem_data[22][2] ), .B1(n3138), .B2(
        \xmem_data[23][2] ), .ZN(n8822) );
  INV_X1 U12751 ( .A(n8822), .ZN(n8823) );
  NOR3_X1 U12752 ( .A1(n8825), .A2(n8824), .A3(n8823), .ZN(n8826) );
  NAND2_X1 U12753 ( .A1(n3791), .A2(n8826), .ZN(n8827) );
  OAI21_X1 U12754 ( .B1(n8828), .B2(n8827), .A(n28215), .ZN(n8829) );
  XOR2_X1 U12755 ( .A(\fmem_data[31][6] ), .B(\fmem_data[31][7] ), .Z(n8833)
         );
  OAI22_X1 U12756 ( .A1(n31975), .A2(n35663), .B1(n26148), .B2(n35662), .ZN(
        n34271) );
  OAI21_X1 U12757 ( .B1(n12727), .B2(n12725), .A(n12724), .ZN(n8835) );
  NAND2_X1 U12758 ( .A1(n12727), .A2(n12725), .ZN(n8834) );
  NAND2_X1 U12759 ( .A1(n8835), .A2(n8834), .ZN(n35158) );
  BUF_X1 U12760 ( .A(n14882), .Z(n30598) );
  AOI22_X1 U12761 ( .A1(n30899), .A2(\xmem_data[96][7] ), .B1(n21009), .B2(
        \xmem_data[97][7] ), .ZN(n8839) );
  BUF_X1 U12762 ( .A(n14974), .Z(n30600) );
  BUF_X1 U12763 ( .A(n14914), .Z(n30599) );
  AOI22_X1 U12764 ( .A1(n30600), .A2(\xmem_data[98][7] ), .B1(n30599), .B2(
        \xmem_data[99][7] ), .ZN(n8838) );
  AOI22_X1 U12765 ( .A1(n22684), .A2(\xmem_data[100][7] ), .B1(n25359), .B2(
        \xmem_data[101][7] ), .ZN(n8837) );
  BUF_X1 U12766 ( .A(n13457), .Z(n30601) );
  AOI22_X1 U12767 ( .A1(n30674), .A2(\xmem_data[102][7] ), .B1(n30601), .B2(
        \xmem_data[103][7] ), .ZN(n8836) );
  NAND4_X1 U12768 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n8855)
         );
  BUF_X1 U12769 ( .A(n29064), .Z(n30592) );
  AOI22_X1 U12770 ( .A1(n30592), .A2(\xmem_data[108][7] ), .B1(n3219), .B2(
        \xmem_data[109][7] ), .ZN(n8843) );
  AOI22_X1 U12771 ( .A1(n3229), .A2(\xmem_data[106][7] ), .B1(n30589), .B2(
        \xmem_data[107][7] ), .ZN(n8842) );
  BUF_X1 U12772 ( .A(n31263), .Z(n30588) );
  AOI22_X1 U12773 ( .A1(n30588), .A2(\xmem_data[104][7] ), .B1(n28317), .B2(
        \xmem_data[105][7] ), .ZN(n8841) );
  BUF_X1 U12774 ( .A(n14988), .Z(n30593) );
  AOI22_X1 U12775 ( .A1(n30593), .A2(\xmem_data[110][7] ), .B1(n20723), .B2(
        \xmem_data[111][7] ), .ZN(n8840) );
  NAND4_X1 U12776 ( .A1(n8843), .A2(n8842), .A3(n8841), .A4(n8840), .ZN(n8854)
         );
  BUF_X1 U12777 ( .A(n14990), .Z(n30606) );
  AOI22_X1 U12778 ( .A1(n30606), .A2(\xmem_data[112][7] ), .B1(n23811), .B2(
        \xmem_data[113][7] ), .ZN(n8847) );
  AOI22_X1 U12779 ( .A1(n28084), .A2(\xmem_data[114][7] ), .B1(n31252), .B2(
        \xmem_data[115][7] ), .ZN(n8846) );
  BUF_X1 U12780 ( .A(n31276), .Z(n30607) );
  AOI22_X1 U12781 ( .A1(n30607), .A2(\xmem_data[116][7] ), .B1(n28481), .B2(
        \xmem_data[117][7] ), .ZN(n8845) );
  BUF_X1 U12782 ( .A(n14997), .Z(n30608) );
  AOI22_X1 U12783 ( .A1(n30608), .A2(\xmem_data[118][7] ), .B1(n24516), .B2(
        \xmem_data[119][7] ), .ZN(n8844) );
  NAND4_X1 U12784 ( .A1(n8847), .A2(n8846), .A3(n8845), .A4(n8844), .ZN(n8853)
         );
  BUF_X1 U12785 ( .A(n14935), .Z(n30613) );
  AOI22_X1 U12786 ( .A1(n30614), .A2(\xmem_data[120][7] ), .B1(n30613), .B2(
        \xmem_data[121][7] ), .ZN(n8851) );
  AOI22_X1 U12787 ( .A1(n29770), .A2(\xmem_data[122][7] ), .B1(n30615), .B2(
        \xmem_data[123][7] ), .ZN(n8850) );
  AOI22_X1 U12788 ( .A1(n23717), .A2(\xmem_data[124][7] ), .B1(n24459), .B2(
        \xmem_data[125][7] ), .ZN(n8849) );
  BUF_X1 U12789 ( .A(n14971), .Z(n30617) );
  BUF_X1 U12790 ( .A(n14913), .Z(n30616) );
  AOI22_X1 U12791 ( .A1(n30617), .A2(\xmem_data[126][7] ), .B1(n30616), .B2(
        \xmem_data[127][7] ), .ZN(n8848) );
  NAND4_X1 U12792 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(n8852)
         );
  OR4_X1 U12793 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n8881)
         );
  NAND2_X1 U12794 ( .A1(n8856), .A2(n37190), .ZN(n8857) );
  INV_X1 U12795 ( .A(n8857), .ZN(n8858) );
  AOI22_X1 U12796 ( .A1(load_xaddr_val[5]), .A2(n8857), .B1(n8858), .B2(n4499), 
        .ZN(n8924) );
  AOI22_X1 U12797 ( .A1(n8858), .A2(n39040), .B1(n14909), .B2(n8857), .ZN(
        n8923) );
  INV_X1 U12798 ( .A(n8923), .ZN(n8902) );
  BUF_X1 U12799 ( .A(n29064), .Z(n30503) );
  AND2_X1 U12800 ( .A1(n3217), .A2(\xmem_data[77][7] ), .ZN(n8859) );
  AOI21_X1 U12801 ( .B1(n30503), .B2(\xmem_data[76][7] ), .A(n8859), .ZN(n8863) );
  AOI22_X1 U12802 ( .A1(n3382), .A2(\xmem_data[74][7] ), .B1(n29286), .B2(
        \xmem_data[75][7] ), .ZN(n8862) );
  BUF_X1 U12803 ( .A(n28974), .Z(n30571) );
  AOI22_X1 U12804 ( .A1(n25724), .A2(\xmem_data[72][7] ), .B1(n30571), .B2(
        \xmem_data[73][7] ), .ZN(n8861) );
  AOI22_X1 U12805 ( .A1(n29256), .A2(\xmem_data[78][7] ), .B1(n31367), .B2(
        \xmem_data[79][7] ), .ZN(n8860) );
  NAND4_X1 U12806 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n8879)
         );
  BUF_X1 U12807 ( .A(n14973), .Z(n30495) );
  AOI22_X1 U12808 ( .A1(n24615), .A2(\xmem_data[64][7] ), .B1(n30495), .B2(
        \xmem_data[65][7] ), .ZN(n8867) );
  AOI22_X1 U12809 ( .A1(n28202), .A2(\xmem_data[66][7] ), .B1(n24167), .B2(
        \xmem_data[67][7] ), .ZN(n8866) );
  BUF_X1 U12810 ( .A(n13486), .Z(n30497) );
  BUF_X1 U12811 ( .A(n14919), .Z(n30496) );
  AOI22_X1 U12812 ( .A1(n30497), .A2(\xmem_data[68][7] ), .B1(n30496), .B2(
        \xmem_data[69][7] ), .ZN(n8865) );
  BUF_X1 U12813 ( .A(n13457), .Z(n30498) );
  AOI22_X1 U12814 ( .A1(n28192), .A2(\xmem_data[70][7] ), .B1(n30498), .B2(
        \xmem_data[71][7] ), .ZN(n8864) );
  NAND4_X1 U12815 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n8878)
         );
  AOI22_X1 U12816 ( .A1(n24565), .A2(\xmem_data[80][7] ), .B1(n3255), .B2(
        \xmem_data[81][7] ), .ZN(n8871) );
  AOI22_X1 U12817 ( .A1(n3126), .A2(\xmem_data[82][7] ), .B1(n23771), .B2(
        \xmem_data[83][7] ), .ZN(n8870) );
  AOI22_X1 U12818 ( .A1(n25670), .A2(\xmem_data[84][7] ), .B1(n29307), .B2(
        \xmem_data[85][7] ), .ZN(n8869) );
  BUF_X1 U12819 ( .A(n14997), .Z(n30508) );
  AOI22_X1 U12820 ( .A1(n30508), .A2(\xmem_data[86][7] ), .B1(n20775), .B2(
        \xmem_data[87][7] ), .ZN(n8868) );
  NAND4_X1 U12821 ( .A1(n8871), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(n8877)
         );
  AOI22_X1 U12822 ( .A1(n29237), .A2(\xmem_data[90][7] ), .B1(n27516), .B2(
        \xmem_data[91][7] ), .ZN(n8875) );
  BUF_X1 U12823 ( .A(n14935), .Z(n30513) );
  AOI22_X1 U12824 ( .A1(n30514), .A2(\xmem_data[88][7] ), .B1(n30513), .B2(
        \xmem_data[89][7] ), .ZN(n8874) );
  AOI22_X1 U12825 ( .A1(n21007), .A2(\xmem_data[92][7] ), .B1(n28492), .B2(
        \xmem_data[93][7] ), .ZN(n8873) );
  BUF_X1 U12826 ( .A(n14913), .Z(n30515) );
  AOI22_X1 U12827 ( .A1(n17044), .A2(\xmem_data[94][7] ), .B1(n30515), .B2(
        \xmem_data[95][7] ), .ZN(n8872) );
  NAND4_X1 U12828 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n8876)
         );
  AOI22_X1 U12829 ( .A1(n8881), .A2(n30626), .B1(n30628), .B2(n8880), .ZN(
        n8928) );
  AOI22_X1 U12830 ( .A1(n28428), .A2(\xmem_data[32][7] ), .B1(n30495), .B2(
        \xmem_data[33][7] ), .ZN(n8886) );
  AOI22_X1 U12831 ( .A1(n29054), .A2(\xmem_data[34][7] ), .B1(n23779), .B2(
        \xmem_data[35][7] ), .ZN(n8885) );
  AOI22_X1 U12832 ( .A1(n30497), .A2(\xmem_data[36][7] ), .B1(n30496), .B2(
        \xmem_data[37][7] ), .ZN(n8884) );
  AND2_X1 U12833 ( .A1(n30498), .A2(\xmem_data[39][7] ), .ZN(n8882) );
  AOI21_X1 U12834 ( .B1(n25584), .B2(\xmem_data[38][7] ), .A(n8882), .ZN(n8883) );
  AOI22_X1 U12835 ( .A1(n30503), .A2(\xmem_data[44][7] ), .B1(n3219), .B2(
        \xmem_data[45][7] ), .ZN(n8901) );
  AOI22_X1 U12836 ( .A1(n22709), .A2(\xmem_data[48][7] ), .B1(n3256), .B2(
        \xmem_data[49][7] ), .ZN(n8890) );
  AOI22_X1 U12837 ( .A1(n28308), .A2(\xmem_data[50][7] ), .B1(n29306), .B2(
        \xmem_data[51][7] ), .ZN(n8889) );
  AOI22_X1 U12838 ( .A1(n27447), .A2(\xmem_data[52][7] ), .B1(n25481), .B2(
        \xmem_data[53][7] ), .ZN(n8888) );
  AOI22_X1 U12839 ( .A1(n30508), .A2(\xmem_data[54][7] ), .B1(n27513), .B2(
        \xmem_data[55][7] ), .ZN(n8887) );
  NAND4_X1 U12840 ( .A1(n8890), .A2(n8889), .A3(n8888), .A4(n8887), .ZN(n8895)
         );
  AOI22_X1 U12841 ( .A1(n21061), .A2(\xmem_data[40][7] ), .B1(n28317), .B2(
        \xmem_data[41][7] ), .ZN(n8893) );
  AOI22_X1 U12842 ( .A1(n20724), .A2(\xmem_data[46][7] ), .B1(n28476), .B2(
        \xmem_data[47][7] ), .ZN(n8892) );
  AOI22_X1 U12843 ( .A1(n3434), .A2(\xmem_data[42][7] ), .B1(n14875), .B2(
        \xmem_data[43][7] ), .ZN(n8891) );
  NOR2_X1 U12844 ( .A1(n8895), .A2(n8894), .ZN(n8900) );
  AOI22_X1 U12845 ( .A1(n30514), .A2(\xmem_data[56][7] ), .B1(n30513), .B2(
        \xmem_data[57][7] ), .ZN(n8899) );
  AOI22_X1 U12846 ( .A1(n28994), .A2(\xmem_data[62][7] ), .B1(n30515), .B2(
        \xmem_data[63][7] ), .ZN(n8898) );
  AOI22_X1 U12847 ( .A1(n25635), .A2(\xmem_data[60][7] ), .B1(n14912), .B2(
        \xmem_data[61][7] ), .ZN(n8897) );
  AOI22_X1 U12848 ( .A1(n3212), .A2(\xmem_data[59][7] ), .B1(
        \xmem_data[58][7] ), .B2(n29807), .ZN(n8896) );
  NAND4_X1 U12849 ( .A1(n3827), .A2(n8901), .A3(n8900), .A4(n3501), .ZN(n8926)
         );
  AND2_X1 U12850 ( .A1(n8902), .A2(n8924), .ZN(n30565) );
  BUF_X1 U12851 ( .A(n14881), .Z(n30557) );
  AOI22_X1 U12852 ( .A1(n30557), .A2(\xmem_data[0][7] ), .B1(n28327), .B2(
        \xmem_data[1][7] ), .ZN(n8906) );
  AOI22_X1 U12853 ( .A1(n29816), .A2(\xmem_data[2][7] ), .B1(n27525), .B2(
        \xmem_data[3][7] ), .ZN(n8905) );
  AOI22_X1 U12854 ( .A1(n3171), .A2(\xmem_data[4][7] ), .B1(n20733), .B2(
        \xmem_data[5][7] ), .ZN(n8904) );
  BUF_X1 U12855 ( .A(n10456), .Z(n30524) );
  AOI22_X1 U12856 ( .A1(n20985), .A2(\xmem_data[6][7] ), .B1(n30524), .B2(
        \xmem_data[7][7] ), .ZN(n8903) );
  NAND4_X1 U12857 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n8922)
         );
  AOI22_X1 U12858 ( .A1(n28076), .A2(\xmem_data[8][7] ), .B1(n27563), .B2(
        \xmem_data[9][7] ), .ZN(n8910) );
  AOI22_X1 U12859 ( .A1(n29661), .A2(\xmem_data[10][7] ), .B1(n24172), .B2(
        \xmem_data[11][7] ), .ZN(n8909) );
  AOI22_X1 U12860 ( .A1(n28503), .A2(\xmem_data[12][7] ), .B1(n3221), .B2(
        \xmem_data[13][7] ), .ZN(n8908) );
  BUF_X1 U12861 ( .A(n14925), .Z(n30534) );
  AOI22_X1 U12862 ( .A1(n24696), .A2(\xmem_data[14][7] ), .B1(n30534), .B2(
        \xmem_data[15][7] ), .ZN(n8907) );
  NAND4_X1 U12863 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n8921)
         );
  BUF_X1 U12864 ( .A(n14890), .Z(n30550) );
  AOI22_X1 U12865 ( .A1(n24697), .A2(\xmem_data[16][7] ), .B1(n30550), .B2(
        \xmem_data[17][7] ), .ZN(n8914) );
  AOI22_X1 U12866 ( .A1(n29706), .A2(\xmem_data[18][7] ), .B1(n27446), .B2(
        \xmem_data[19][7] ), .ZN(n8913) );
  AOI22_X1 U12867 ( .A1(n30551), .A2(\xmem_data[20][7] ), .B1(n30884), .B2(
        \xmem_data[21][7] ), .ZN(n8912) );
  BUF_X1 U12868 ( .A(n13435), .Z(n30552) );
  AOI22_X1 U12869 ( .A1(n23792), .A2(\xmem_data[22][7] ), .B1(n30552), .B2(
        \xmem_data[23][7] ), .ZN(n8911) );
  NAND4_X1 U12870 ( .A1(n8914), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n8920)
         );
  BUF_X1 U12871 ( .A(n14898), .Z(n30541) );
  AOI22_X1 U12872 ( .A1(n28980), .A2(\xmem_data[24][7] ), .B1(n30541), .B2(
        \xmem_data[25][7] ), .ZN(n8918) );
  BUF_X1 U12873 ( .A(n29187), .Z(n30543) );
  BUF_X1 U12874 ( .A(n13188), .Z(n30542) );
  AOI22_X1 U12875 ( .A1(n23795), .A2(\xmem_data[26][7] ), .B1(n30542), .B2(
        \xmem_data[27][7] ), .ZN(n8917) );
  BUF_X1 U12876 ( .A(n14912), .Z(n30544) );
  AOI22_X1 U12877 ( .A1(n31330), .A2(\xmem_data[28][7] ), .B1(n30544), .B2(
        \xmem_data[29][7] ), .ZN(n8916) );
  BUF_X1 U12878 ( .A(n13452), .Z(n30545) );
  AOI22_X1 U12879 ( .A1(n17021), .A2(\xmem_data[30][7] ), .B1(n30545), .B2(
        \xmem_data[31][7] ), .ZN(n8915) );
  NAND4_X1 U12880 ( .A1(n8918), .A2(n8917), .A3(n8916), .A4(n8915), .ZN(n8919)
         );
  OR4_X1 U12881 ( .A1(n8922), .A2(n8921), .A3(n8920), .A4(n8919), .ZN(n8925)
         );
  NOR2_X1 U12882 ( .A1(n8924), .A2(n8923), .ZN(n30563) );
  AOI22_X1 U12883 ( .A1(n8926), .A2(n30565), .B1(n8925), .B2(n30563), .ZN(
        n8927) );
  NAND2_X1 U12884 ( .A1(n8928), .A2(n8927), .ZN(n35106) );
  XNOR2_X1 U12885 ( .A(n35106), .B(\fmem_data[26][5] ), .ZN(n35032) );
  AOI22_X1 U12886 ( .A1(n30514), .A2(\xmem_data[88][6] ), .B1(n30513), .B2(
        \xmem_data[89][6] ), .ZN(n8932) );
  AOI22_X1 U12887 ( .A1(n25461), .A2(\xmem_data[90][6] ), .B1(n3208), .B2(
        \xmem_data[91][6] ), .ZN(n8931) );
  AOI22_X1 U12888 ( .A1(n24509), .A2(\xmem_data[92][6] ), .B1(n21006), .B2(
        \xmem_data[93][6] ), .ZN(n8930) );
  AOI22_X1 U12889 ( .A1(n30950), .A2(\xmem_data[94][6] ), .B1(n30515), .B2(
        \xmem_data[95][6] ), .ZN(n8929) );
  NAND4_X1 U12890 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n8938)
         );
  AOI22_X1 U12891 ( .A1(n25630), .A2(\xmem_data[72][6] ), .B1(n30571), .B2(
        \xmem_data[73][6] ), .ZN(n8936) );
  AOI22_X1 U12892 ( .A1(n29065), .A2(\xmem_data[78][6] ), .B1(n20500), .B2(
        \xmem_data[79][6] ), .ZN(n8934) );
  AOI22_X1 U12893 ( .A1(n3229), .A2(\xmem_data[74][6] ), .B1(n27437), .B2(
        \xmem_data[75][6] ), .ZN(n8933) );
  NAND2_X1 U12894 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  NOR2_X1 U12895 ( .A1(n8938), .A2(n8937), .ZN(n8949) );
  AOI22_X1 U12896 ( .A1(n30557), .A2(\xmem_data[64][6] ), .B1(n30495), .B2(
        \xmem_data[65][6] ), .ZN(n8942) );
  AOI22_X1 U12897 ( .A1(n14974), .A2(n20682), .B1(n29245), .B2(
        \xmem_data[67][6] ), .ZN(n8941) );
  AOI22_X1 U12898 ( .A1(n30497), .A2(\xmem_data[68][6] ), .B1(n30496), .B2(
        \xmem_data[69][6] ), .ZN(n8940) );
  AOI22_X1 U12899 ( .A1(n30901), .A2(\xmem_data[70][6] ), .B1(n30498), .B2(
        \xmem_data[71][6] ), .ZN(n8939) );
  AND2_X1 U12900 ( .A1(n3222), .A2(\xmem_data[77][6] ), .ZN(n8943) );
  AOI22_X1 U12901 ( .A1(n25617), .A2(\xmem_data[80][6] ), .B1(n3255), .B2(
        \xmem_data[81][6] ), .ZN(n8947) );
  AOI22_X1 U12902 ( .A1(n3280), .A2(\xmem_data[82][6] ), .B1(n29306), .B2(
        \xmem_data[83][6] ), .ZN(n8946) );
  AOI22_X1 U12903 ( .A1(n25707), .A2(\xmem_data[84][6] ), .B1(n24130), .B2(
        \xmem_data[85][6] ), .ZN(n8945) );
  AOI22_X1 U12904 ( .A1(n30508), .A2(\xmem_data[86][6] ), .B1(n13168), .B2(
        \xmem_data[87][6] ), .ZN(n8944) );
  NAND2_X1 U12905 ( .A1(n8950), .A2(n30628), .ZN(n9025) );
  AOI22_X1 U12906 ( .A1(n3178), .A2(\xmem_data[32][6] ), .B1(n30495), .B2(
        \xmem_data[33][6] ), .ZN(n8954) );
  AOI22_X1 U12907 ( .A1(n28955), .A2(\xmem_data[34][6] ), .B1(n22685), .B2(
        \xmem_data[35][6] ), .ZN(n8953) );
  AOI22_X1 U12908 ( .A1(n30497), .A2(\xmem_data[36][6] ), .B1(n30496), .B2(
        \xmem_data[37][6] ), .ZN(n8952) );
  AOI22_X1 U12909 ( .A1(n30674), .A2(\xmem_data[38][6] ), .B1(n30498), .B2(
        \xmem_data[39][6] ), .ZN(n8951) );
  AOI22_X1 U12910 ( .A1(n21061), .A2(\xmem_data[40][6] ), .B1(n30908), .B2(
        \xmem_data[41][6] ), .ZN(n8957) );
  AOI22_X1 U12911 ( .A1(n24139), .A2(\xmem_data[46][6] ), .B1(n22667), .B2(
        \xmem_data[47][6] ), .ZN(n8956) );
  AOI22_X1 U12912 ( .A1(n3414), .A2(\xmem_data[42][6] ), .B1(n27437), .B2(
        \xmem_data[43][6] ), .ZN(n8955) );
  AOI22_X1 U12913 ( .A1(n25449), .A2(\xmem_data[48][6] ), .B1(n3256), .B2(
        \xmem_data[49][6] ), .ZN(n8961) );
  AOI22_X1 U12914 ( .A1(n29157), .A2(\xmem_data[50][6] ), .B1(n3231), .B2(
        \xmem_data[51][6] ), .ZN(n8960) );
  AOI22_X1 U12915 ( .A1(n20961), .A2(\xmem_data[52][6] ), .B1(n3357), .B2(
        \xmem_data[53][6] ), .ZN(n8959) );
  AOI22_X1 U12916 ( .A1(n30508), .A2(\xmem_data[54][6] ), .B1(n24159), .B2(
        \xmem_data[55][6] ), .ZN(n8958) );
  NAND4_X1 U12917 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n8962)
         );
  NOR2_X1 U12918 ( .A1(n8963), .A2(n8962), .ZN(n8964) );
  NAND2_X1 U12919 ( .A1(n3773), .A2(n8964), .ZN(n8971) );
  AOI22_X1 U12920 ( .A1(n30514), .A2(\xmem_data[56][6] ), .B1(n30513), .B2(
        \xmem_data[57][6] ), .ZN(n8968) );
  AOI22_X1 U12921 ( .A1(n29010), .A2(\xmem_data[60][6] ), .B1(n20505), .B2(
        \xmem_data[61][6] ), .ZN(n8966) );
  AOI22_X1 U12922 ( .A1(n28302), .A2(\xmem_data[62][6] ), .B1(n30515), .B2(
        \xmem_data[63][6] ), .ZN(n8965) );
  AOI22_X1 U12923 ( .A1(n30503), .A2(\xmem_data[44][6] ), .B1(n3222), .B2(
        \xmem_data[45][6] ), .ZN(n8969) );
  NAND2_X1 U12924 ( .A1(n3774), .A2(n8969), .ZN(n8970) );
  OAI21_X1 U12925 ( .B1(n8971), .B2(n8970), .A(n30565), .ZN(n9024) );
  AOI22_X1 U12926 ( .A1(n3205), .A2(\xmem_data[96][6] ), .B1(n20506), .B2(
        \xmem_data[97][6] ), .ZN(n8975) );
  AOI22_X1 U12927 ( .A1(n30600), .A2(\xmem_data[98][6] ), .B1(n30599), .B2(
        \xmem_data[99][6] ), .ZN(n8974) );
  AOI22_X1 U12928 ( .A1(n24572), .A2(\xmem_data[100][6] ), .B1(n20488), .B2(
        \xmem_data[101][6] ), .ZN(n8973) );
  AOI22_X1 U12929 ( .A1(n29383), .A2(\xmem_data[102][6] ), .B1(n30601), .B2(
        \xmem_data[103][6] ), .ZN(n8972) );
  NAND4_X1 U12930 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n8987)
         );
  AOI22_X1 U12931 ( .A1(n30606), .A2(\xmem_data[112][6] ), .B1(n25415), .B2(
        \xmem_data[113][6] ), .ZN(n8979) );
  AOI22_X1 U12932 ( .A1(n29762), .A2(\xmem_data[114][6] ), .B1(n28343), .B2(
        \xmem_data[115][6] ), .ZN(n8978) );
  AOI22_X1 U12933 ( .A1(n30607), .A2(\xmem_data[116][6] ), .B1(n22739), .B2(
        \xmem_data[117][6] ), .ZN(n8977) );
  AOI22_X1 U12934 ( .A1(n30608), .A2(\xmem_data[118][6] ), .B1(n24639), .B2(
        \xmem_data[119][6] ), .ZN(n8976) );
  NAND4_X1 U12935 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(n8985)
         );
  AOI22_X1 U12936 ( .A1(n30614), .A2(\xmem_data[120][6] ), .B1(n30613), .B2(
        \xmem_data[121][6] ), .ZN(n8983) );
  AOI22_X1 U12937 ( .A1(n20939), .A2(\xmem_data[122][6] ), .B1(n30615), .B2(
        \xmem_data[123][6] ), .ZN(n8982) );
  AOI22_X1 U12938 ( .A1(n24593), .A2(\xmem_data[124][6] ), .B1(n25715), .B2(
        \xmem_data[125][6] ), .ZN(n8981) );
  AOI22_X1 U12939 ( .A1(n30617), .A2(\xmem_data[126][6] ), .B1(n30616), .B2(
        \xmem_data[127][6] ), .ZN(n8980) );
  NAND4_X1 U12940 ( .A1(n8983), .A2(n8982), .A3(n8981), .A4(n8980), .ZN(n8984)
         );
  OR2_X1 U12941 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  OR2_X1 U12942 ( .A1(n8987), .A2(n8986), .ZN(n8996) );
  AOI22_X1 U12943 ( .A1(n30592), .A2(\xmem_data[108][6] ), .B1(n3220), .B2(
        \xmem_data[109][6] ), .ZN(n8994) );
  AOI22_X1 U12944 ( .A1(n30588), .A2(\xmem_data[104][6] ), .B1(n12471), .B2(
        \xmem_data[105][6] ), .ZN(n8988) );
  INV_X1 U12945 ( .A(n8988), .ZN(n8992) );
  AOI22_X1 U12946 ( .A1(n30593), .A2(\xmem_data[110][6] ), .B1(n25562), .B2(
        \xmem_data[111][6] ), .ZN(n8990) );
  AOI22_X1 U12947 ( .A1(n3348), .A2(\xmem_data[106][6] ), .B1(n30589), .B2(
        \xmem_data[107][6] ), .ZN(n8989) );
  NAND2_X1 U12948 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NOR2_X1 U12949 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U12950 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  OAI21_X1 U12951 ( .B1(n8996), .B2(n8995), .A(n30626), .ZN(n9023) );
  AOI22_X1 U12952 ( .A1(n27502), .A2(\xmem_data[12][6] ), .B1(n3217), .B2(
        \xmem_data[13][6] ), .ZN(n8998) );
  AOI22_X1 U12953 ( .A1(n30674), .A2(\xmem_data[6][6] ), .B1(n30524), .B2(
        \xmem_data[7][6] ), .ZN(n8997) );
  AOI22_X1 U12954 ( .A1(n20541), .A2(\xmem_data[24][6] ), .B1(n30541), .B2(
        \xmem_data[25][6] ), .ZN(n9002) );
  AOI22_X1 U12955 ( .A1(n27818), .A2(\xmem_data[26][6] ), .B1(n30542), .B2(
        \xmem_data[27][6] ), .ZN(n9001) );
  AOI22_X1 U12956 ( .A1(n30949), .A2(\xmem_data[28][6] ), .B1(n30544), .B2(
        \xmem_data[29][6] ), .ZN(n9000) );
  AOI22_X1 U12957 ( .A1(n28781), .A2(\xmem_data[30][6] ), .B1(n30545), .B2(
        \xmem_data[31][6] ), .ZN(n8999) );
  AOI22_X1 U12958 ( .A1(n25686), .A2(\xmem_data[8][6] ), .B1(n30571), .B2(
        \xmem_data[9][6] ), .ZN(n9019) );
  AOI22_X1 U12959 ( .A1(n27904), .A2(\xmem_data[16][6] ), .B1(n30550), .B2(
        \xmem_data[17][6] ), .ZN(n9006) );
  AOI22_X1 U12960 ( .A1(n3126), .A2(\xmem_data[18][6] ), .B1(n3231), .B2(
        \xmem_data[19][6] ), .ZN(n9005) );
  AOI22_X1 U12961 ( .A1(n30551), .A2(\xmem_data[20][6] ), .B1(n30884), .B2(
        \xmem_data[21][6] ), .ZN(n9004) );
  AOI22_X1 U12962 ( .A1(n28671), .A2(\xmem_data[22][6] ), .B1(n30552), .B2(
        \xmem_data[23][6] ), .ZN(n9003) );
  NAND4_X1 U12963 ( .A1(n9006), .A2(n9005), .A3(n9004), .A4(n9003), .ZN(n9017)
         );
  AOI22_X1 U12964 ( .A1(n30557), .A2(\xmem_data[0][6] ), .B1(n27461), .B2(
        \xmem_data[1][6] ), .ZN(n9015) );
  AOI22_X1 U12965 ( .A1(n29151), .A2(\xmem_data[4][6] ), .B1(n28979), .B2(
        \xmem_data[5][6] ), .ZN(n9007) );
  INV_X1 U12966 ( .A(n9007), .ZN(n9013) );
  AOI22_X1 U12967 ( .A1(n29026), .A2(\xmem_data[14][6] ), .B1(n30534), .B2(
        \xmem_data[15][6] ), .ZN(n9008) );
  INV_X1 U12968 ( .A(n9008), .ZN(n9012) );
  AOI22_X1 U12969 ( .A1(n20984), .A2(\xmem_data[2][6] ), .B1(n14975), .B2(
        \xmem_data[3][6] ), .ZN(n9010) );
  AOI22_X1 U12970 ( .A1(n30907), .A2(\xmem_data[10][6] ), .B1(n3247), .B2(
        \xmem_data[11][6] ), .ZN(n9009) );
  NAND2_X1 U12971 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  NOR3_X1 U12972 ( .A1(n9013), .A2(n9012), .A3(n9011), .ZN(n9014) );
  NAND2_X1 U12973 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  NOR2_X1 U12974 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  NAND4_X1 U12975 ( .A1(n9018), .A2(n3779), .A3(n9019), .A4(n9020), .ZN(n9021)
         );
  NAND2_X1 U12976 ( .A1(n9021), .A2(n30563), .ZN(n9022) );
  XNOR2_X1 U12977 ( .A(n31670), .B(\fmem_data[26][5] ), .ZN(n24436) );
  OAI22_X1 U12978 ( .A1(n35032), .A2(n35034), .B1(n24436), .B2(n35033), .ZN(
        n31830) );
  AOI22_X1 U12979 ( .A1(n27959), .A2(\xmem_data[40][5] ), .B1(n20489), .B2(
        \xmem_data[41][5] ), .ZN(n9030) );
  AOI22_X1 U12980 ( .A1(n23732), .A2(\xmem_data[42][5] ), .B1(n3247), .B2(
        \xmem_data[43][5] ), .ZN(n9029) );
  AOI22_X1 U12981 ( .A1(n30503), .A2(\xmem_data[44][5] ), .B1(n3221), .B2(
        \xmem_data[45][5] ), .ZN(n9028) );
  AOI22_X1 U12982 ( .A1(n29698), .A2(\xmem_data[46][5] ), .B1(n25562), .B2(
        \xmem_data[47][5] ), .ZN(n9027) );
  NAND4_X1 U12983 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n9046)
         );
  AOI22_X1 U12984 ( .A1(n27524), .A2(\xmem_data[32][5] ), .B1(n30495), .B2(
        \xmem_data[33][5] ), .ZN(n9034) );
  AOI22_X1 U12985 ( .A1(n24571), .A2(\xmem_data[34][5] ), .B1(n29126), .B2(
        \xmem_data[35][5] ), .ZN(n9033) );
  AOI22_X1 U12986 ( .A1(n30497), .A2(\xmem_data[36][5] ), .B1(n30496), .B2(
        \xmem_data[37][5] ), .ZN(n9032) );
  AOI22_X1 U12987 ( .A1(n30754), .A2(\xmem_data[38][5] ), .B1(n30498), .B2(
        \xmem_data[39][5] ), .ZN(n9031) );
  NAND4_X1 U12988 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(n9045)
         );
  AOI22_X1 U12989 ( .A1(n30606), .A2(\xmem_data[48][5] ), .B1(n3256), .B2(
        \xmem_data[49][5] ), .ZN(n9038) );
  AOI22_X1 U12990 ( .A1(n3140), .A2(\xmem_data[50][5] ), .B1(n28007), .B2(
        \xmem_data[51][5] ), .ZN(n9037) );
  AOI22_X1 U12991 ( .A1(n27447), .A2(\xmem_data[52][5] ), .B1(n27988), .B2(
        \xmem_data[53][5] ), .ZN(n9036) );
  AOI22_X1 U12992 ( .A1(n30508), .A2(\xmem_data[54][5] ), .B1(n22702), .B2(
        \xmem_data[55][5] ), .ZN(n9035) );
  NAND4_X1 U12993 ( .A1(n9038), .A2(n9037), .A3(n9036), .A4(n9035), .ZN(n9044)
         );
  AOI22_X1 U12994 ( .A1(n30514), .A2(\xmem_data[56][5] ), .B1(n30513), .B2(
        \xmem_data[57][5] ), .ZN(n9042) );
  AOI22_X1 U12995 ( .A1(n28231), .A2(\xmem_data[58][5] ), .B1(n29162), .B2(
        \xmem_data[59][5] ), .ZN(n9041) );
  AOI22_X1 U12996 ( .A1(n20585), .A2(\xmem_data[60][5] ), .B1(n28492), .B2(
        \xmem_data[61][5] ), .ZN(n9040) );
  AOI22_X1 U12997 ( .A1(n28302), .A2(\xmem_data[62][5] ), .B1(n30515), .B2(
        \xmem_data[63][5] ), .ZN(n9039) );
  NAND4_X1 U12998 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n9043)
         );
  OR4_X1 U12999 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(n9068)
         );
  AOI22_X1 U13000 ( .A1(n30557), .A2(\xmem_data[0][5] ), .B1(n30898), .B2(
        \xmem_data[1][5] ), .ZN(n9050) );
  AOI22_X1 U13001 ( .A1(n28226), .A2(\xmem_data[2][5] ), .B1(n24622), .B2(
        \xmem_data[3][5] ), .ZN(n9049) );
  AOI22_X1 U13002 ( .A1(n3172), .A2(\xmem_data[4][5] ), .B1(n27463), .B2(
        \xmem_data[5][5] ), .ZN(n9048) );
  AOI22_X1 U13003 ( .A1(n20952), .A2(\xmem_data[6][5] ), .B1(n30524), .B2(
        \xmem_data[7][5] ), .ZN(n9047) );
  NAND4_X1 U13004 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n9066)
         );
  AOI22_X1 U13005 ( .A1(n27436), .A2(\xmem_data[8][5] ), .B1(n30571), .B2(
        \xmem_data[9][5] ), .ZN(n9054) );
  AOI22_X1 U13006 ( .A1(n20828), .A2(\xmem_data[10][5] ), .B1(n23731), .B2(
        \xmem_data[11][5] ), .ZN(n9053) );
  AOI22_X1 U13007 ( .A1(n28044), .A2(\xmem_data[12][5] ), .B1(n3222), .B2(
        \xmem_data[13][5] ), .ZN(n9052) );
  AOI22_X1 U13008 ( .A1(n30593), .A2(\xmem_data[14][5] ), .B1(n30534), .B2(
        \xmem_data[15][5] ), .ZN(n9051) );
  NAND4_X1 U13009 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n9065)
         );
  AOI22_X1 U13010 ( .A1(n3340), .A2(\xmem_data[16][5] ), .B1(n30550), .B2(
        \xmem_data[17][5] ), .ZN(n9058) );
  AOI22_X1 U13011 ( .A1(n3134), .A2(\xmem_data[18][5] ), .B1(n29306), .B2(
        \xmem_data[19][5] ), .ZN(n9057) );
  AOI22_X1 U13012 ( .A1(n30551), .A2(\xmem_data[20][5] ), .B1(n20546), .B2(
        \xmem_data[21][5] ), .ZN(n9056) );
  AOI22_X1 U13013 ( .A1(n28309), .A2(\xmem_data[22][5] ), .B1(n30552), .B2(
        \xmem_data[23][5] ), .ZN(n9055) );
  NAND4_X1 U13014 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n9064)
         );
  AOI22_X1 U13015 ( .A1(n3175), .A2(\xmem_data[24][5] ), .B1(n30541), .B2(
        \xmem_data[25][5] ), .ZN(n9062) );
  AOI22_X1 U13016 ( .A1(n27517), .A2(\xmem_data[26][5] ), .B1(n30542), .B2(
        \xmem_data[27][5] ), .ZN(n9061) );
  AOI22_X1 U13017 ( .A1(n24509), .A2(\xmem_data[28][5] ), .B1(n30544), .B2(
        \xmem_data[29][5] ), .ZN(n9060) );
  AOI22_X1 U13018 ( .A1(n30872), .A2(\xmem_data[30][5] ), .B1(n30545), .B2(
        \xmem_data[31][5] ), .ZN(n9059) );
  NAND4_X1 U13019 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n9063)
         );
  OR4_X1 U13020 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n9067)
         );
  AOI22_X1 U13021 ( .A1(n9068), .A2(n30565), .B1(n9067), .B2(n30563), .ZN(
        n9113) );
  AOI22_X1 U13022 ( .A1(n29240), .A2(\xmem_data[96][5] ), .B1(n20816), .B2(
        \xmem_data[97][5] ), .ZN(n9072) );
  AOI22_X1 U13023 ( .A1(n30600), .A2(\xmem_data[98][5] ), .B1(n30599), .B2(
        \xmem_data[99][5] ), .ZN(n9071) );
  AOI22_X1 U13024 ( .A1(n20818), .A2(\xmem_data[100][5] ), .B1(n29086), .B2(
        \xmem_data[101][5] ), .ZN(n9070) );
  AOI22_X1 U13025 ( .A1(n29820), .A2(\xmem_data[102][5] ), .B1(n30601), .B2(
        \xmem_data[103][5] ), .ZN(n9069) );
  NAND4_X1 U13026 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n9088)
         );
  AOI22_X1 U13027 ( .A1(n30592), .A2(\xmem_data[108][5] ), .B1(n3222), .B2(
        \xmem_data[109][5] ), .ZN(n9076) );
  AOI22_X1 U13028 ( .A1(n3229), .A2(\xmem_data[106][5] ), .B1(n30589), .B2(
        \xmem_data[107][5] ), .ZN(n9075) );
  AOI22_X1 U13029 ( .A1(n30588), .A2(\xmem_data[104][5] ), .B1(n30571), .B2(
        \xmem_data[105][5] ), .ZN(n9074) );
  AOI22_X1 U13030 ( .A1(n30593), .A2(\xmem_data[110][5] ), .B1(n22710), .B2(
        \xmem_data[111][5] ), .ZN(n9073) );
  NAND4_X1 U13031 ( .A1(n9076), .A2(n9075), .A3(n9074), .A4(n9073), .ZN(n9087)
         );
  AOI22_X1 U13032 ( .A1(n30606), .A2(\xmem_data[112][5] ), .B1(n22669), .B2(
        \xmem_data[113][5] ), .ZN(n9080) );
  AOI22_X1 U13033 ( .A1(n3135), .A2(\xmem_data[114][5] ), .B1(n29306), .B2(
        \xmem_data[115][5] ), .ZN(n9079) );
  AOI22_X1 U13034 ( .A1(n30607), .A2(\xmem_data[116][5] ), .B1(n22701), .B2(
        \xmem_data[117][5] ), .ZN(n9078) );
  AOI22_X1 U13035 ( .A1(n30608), .A2(\xmem_data[118][5] ), .B1(n25605), .B2(
        \xmem_data[119][5] ), .ZN(n9077) );
  NAND4_X1 U13036 ( .A1(n9080), .A2(n9079), .A3(n9078), .A4(n9077), .ZN(n9086)
         );
  AOI22_X1 U13037 ( .A1(n30614), .A2(\xmem_data[120][5] ), .B1(n30613), .B2(
        \xmem_data[121][5] ), .ZN(n9084) );
  AOI22_X1 U13038 ( .A1(n30303), .A2(\xmem_data[122][5] ), .B1(n30615), .B2(
        \xmem_data[123][5] ), .ZN(n9083) );
  AOI22_X1 U13039 ( .A1(n29317), .A2(\xmem_data[124][5] ), .B1(n17043), .B2(
        \xmem_data[125][5] ), .ZN(n9082) );
  AOI22_X1 U13040 ( .A1(n30617), .A2(\xmem_data[126][5] ), .B1(n30616), .B2(
        \xmem_data[127][5] ), .ZN(n9081) );
  NAND4_X1 U13041 ( .A1(n9084), .A2(n9083), .A3(n9082), .A4(n9081), .ZN(n9085)
         );
  OR4_X1 U13042 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n9111)
         );
  AND2_X1 U13043 ( .A1(n3221), .A2(\xmem_data[77][5] ), .ZN(n9089) );
  AOI21_X1 U13044 ( .B1(n30503), .B2(\xmem_data[76][5] ), .A(n9089), .ZN(n9093) );
  AOI22_X1 U13045 ( .A1(n27813), .A2(\xmem_data[74][5] ), .B1(n29286), .B2(
        \xmem_data[75][5] ), .ZN(n9092) );
  AOI22_X1 U13046 ( .A1(n27500), .A2(\xmem_data[72][5] ), .B1(n30571), .B2(
        \xmem_data[73][5] ), .ZN(n9091) );
  AOI22_X1 U13047 ( .A1(n22708), .A2(\xmem_data[78][5] ), .B1(n27507), .B2(
        \xmem_data[79][5] ), .ZN(n9090) );
  NAND4_X1 U13048 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n9109)
         );
  AOI22_X1 U13049 ( .A1(n28428), .A2(\xmem_data[64][5] ), .B1(n30495), .B2(
        \xmem_data[65][5] ), .ZN(n9097) );
  AOI22_X1 U13050 ( .A1(n30269), .A2(\xmem_data[66][5] ), .B1(n24622), .B2(
        \xmem_data[67][5] ), .ZN(n9096) );
  AOI22_X1 U13051 ( .A1(n30497), .A2(\xmem_data[68][5] ), .B1(n30496), .B2(
        \xmem_data[69][5] ), .ZN(n9095) );
  AOI22_X1 U13052 ( .A1(n29298), .A2(\xmem_data[70][5] ), .B1(n30498), .B2(
        \xmem_data[71][5] ), .ZN(n9094) );
  NAND4_X1 U13053 ( .A1(n9097), .A2(n9096), .A3(n9095), .A4(n9094), .ZN(n9108)
         );
  AOI22_X1 U13054 ( .A1(n23741), .A2(\xmem_data[80][5] ), .B1(n3255), .B2(
        \xmem_data[81][5] ), .ZN(n9101) );
  AOI22_X1 U13055 ( .A1(n29350), .A2(\xmem_data[82][5] ), .B1(n23771), .B2(
        \xmem_data[83][5] ), .ZN(n9100) );
  AOI22_X1 U13056 ( .A1(n20961), .A2(\xmem_data[84][5] ), .B1(n27943), .B2(
        \xmem_data[85][5] ), .ZN(n9099) );
  AOI22_X1 U13057 ( .A1(n30508), .A2(\xmem_data[86][5] ), .B1(n13168), .B2(
        \xmem_data[87][5] ), .ZN(n9098) );
  NAND4_X1 U13058 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n9107)
         );
  AOI22_X1 U13059 ( .A1(n30514), .A2(\xmem_data[88][5] ), .B1(n30513), .B2(
        \xmem_data[89][5] ), .ZN(n9105) );
  AOI22_X1 U13060 ( .A1(n21005), .A2(\xmem_data[90][5] ), .B1(n27516), .B2(
        \xmem_data[91][5] ), .ZN(n9104) );
  AOI22_X1 U13061 ( .A1(n22676), .A2(\xmem_data[92][5] ), .B1(n28492), .B2(
        \xmem_data[93][5] ), .ZN(n9103) );
  AOI22_X1 U13062 ( .A1(n31255), .A2(\xmem_data[94][5] ), .B1(n30515), .B2(
        \xmem_data[95][5] ), .ZN(n9102) );
  NAND4_X1 U13063 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n9106)
         );
  OR4_X1 U13064 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n9110)
         );
  AOI22_X1 U13065 ( .A1(n9111), .A2(n30626), .B1(n30628), .B2(n9110), .ZN(
        n9112) );
  XNOR2_X1 U13066 ( .A(n32163), .B(\fmem_data[26][7] ), .ZN(n31671) );
  XOR2_X1 U13067 ( .A(\fmem_data[26][6] ), .B(\fmem_data[26][7] ), .Z(n9114)
         );
  AOI22_X1 U13068 ( .A1(n29100), .A2(\xmem_data[64][4] ), .B1(n30495), .B2(
        \xmem_data[65][4] ), .ZN(n9118) );
  AOI22_X1 U13069 ( .A1(n20732), .A2(\xmem_data[66][4] ), .B1(n24622), .B2(
        \xmem_data[67][4] ), .ZN(n9117) );
  AOI22_X1 U13070 ( .A1(n30497), .A2(\xmem_data[68][4] ), .B1(n30496), .B2(
        \xmem_data[69][4] ), .ZN(n9116) );
  AOI22_X1 U13071 ( .A1(n29725), .A2(\xmem_data[70][4] ), .B1(n30498), .B2(
        \xmem_data[71][4] ), .ZN(n9115) );
  NAND4_X1 U13072 ( .A1(n9118), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n9138)
         );
  AOI22_X1 U13073 ( .A1(n30503), .A2(\xmem_data[76][4] ), .B1(n3219), .B2(
        \xmem_data[77][4] ), .ZN(n9126) );
  NAND2_X1 U13074 ( .A1(n24470), .A2(\xmem_data[73][4] ), .ZN(n9120) );
  NAND2_X1 U13075 ( .A1(n20953), .A2(\xmem_data[72][4] ), .ZN(n9119) );
  NAND2_X1 U13076 ( .A1(n9120), .A2(n9119), .ZN(n9124) );
  AOI22_X1 U13077 ( .A1(n25612), .A2(\xmem_data[78][4] ), .B1(n30534), .B2(
        \xmem_data[79][4] ), .ZN(n9122) );
  AOI22_X1 U13078 ( .A1(n3335), .A2(\xmem_data[74][4] ), .B1(n14983), .B2(
        \xmem_data[75][4] ), .ZN(n9121) );
  NAND2_X1 U13079 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  NOR2_X1 U13080 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  NAND2_X1 U13081 ( .A1(n9126), .A2(n9125), .ZN(n9137) );
  AOI22_X1 U13082 ( .A1(n20969), .A2(\xmem_data[80][4] ), .B1(n3256), .B2(
        \xmem_data[81][4] ), .ZN(n9130) );
  AOI22_X1 U13083 ( .A1(n3140), .A2(\xmem_data[82][4] ), .B1(n28045), .B2(
        \xmem_data[83][4] ), .ZN(n9129) );
  AOI22_X1 U13084 ( .A1(n25422), .A2(\xmem_data[84][4] ), .B1(n22739), .B2(
        \xmem_data[85][4] ), .ZN(n9128) );
  AOI22_X1 U13085 ( .A1(n30508), .A2(\xmem_data[86][4] ), .B1(n13168), .B2(
        \xmem_data[87][4] ), .ZN(n9127) );
  NAND4_X1 U13086 ( .A1(n9130), .A2(n9129), .A3(n9128), .A4(n9127), .ZN(n9136)
         );
  AOI22_X1 U13087 ( .A1(n30514), .A2(\xmem_data[88][4] ), .B1(n30513), .B2(
        \xmem_data[89][4] ), .ZN(n9134) );
  AOI22_X1 U13088 ( .A1(n27755), .A2(\xmem_data[90][4] ), .B1(n27516), .B2(
        \xmem_data[91][4] ), .ZN(n9133) );
  AOI22_X1 U13089 ( .A1(n25573), .A2(\xmem_data[92][4] ), .B1(n28492), .B2(
        \xmem_data[93][4] ), .ZN(n9132) );
  AOI22_X1 U13090 ( .A1(n24710), .A2(\xmem_data[94][4] ), .B1(n30515), .B2(
        \xmem_data[95][4] ), .ZN(n9131) );
  NAND4_X1 U13091 ( .A1(n9134), .A2(n9133), .A3(n9132), .A4(n9131), .ZN(n9135)
         );
  OR4_X1 U13092 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9135), .ZN(n9139)
         );
  NAND2_X1 U13093 ( .A1(n9139), .A2(n30628), .ZN(n9207) );
  AND2_X1 U13094 ( .A1(n3218), .A2(\xmem_data[45][4] ), .ZN(n9140) );
  AOI21_X1 U13095 ( .B1(n30503), .B2(\xmem_data[44][4] ), .A(n9140), .ZN(n9144) );
  AOI22_X1 U13096 ( .A1(n3351), .A2(\xmem_data[42][4] ), .B1(n23731), .B2(
        \xmem_data[43][4] ), .ZN(n9143) );
  AOI22_X1 U13097 ( .A1(n27564), .A2(\xmem_data[40][4] ), .B1(n30571), .B2(
        \xmem_data[41][4] ), .ZN(n9142) );
  AOI22_X1 U13098 ( .A1(n22708), .A2(\xmem_data[46][4] ), .B1(n29028), .B2(
        \xmem_data[47][4] ), .ZN(n9141) );
  NAND4_X1 U13099 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n9160)
         );
  AOI22_X1 U13100 ( .A1(n25521), .A2(\xmem_data[32][4] ), .B1(n30495), .B2(
        \xmem_data[33][4] ), .ZN(n9148) );
  AOI22_X1 U13101 ( .A1(n29246), .A2(\xmem_data[34][4] ), .B1(n24622), .B2(
        \xmem_data[35][4] ), .ZN(n9147) );
  AOI22_X1 U13102 ( .A1(n30497), .A2(\xmem_data[36][4] ), .B1(n30496), .B2(
        \xmem_data[37][4] ), .ZN(n9146) );
  AOI22_X1 U13103 ( .A1(n31345), .A2(\xmem_data[38][4] ), .B1(n30498), .B2(
        \xmem_data[39][4] ), .ZN(n9145) );
  NAND4_X1 U13104 ( .A1(n9148), .A2(n9147), .A3(n9146), .A4(n9145), .ZN(n9159)
         );
  AOI22_X1 U13105 ( .A1(n24438), .A2(\xmem_data[48][4] ), .B1(n3256), .B2(
        \xmem_data[49][4] ), .ZN(n9152) );
  AOI22_X1 U13106 ( .A1(n20808), .A2(\xmem_data[50][4] ), .B1(n28007), .B2(
        \xmem_data[51][4] ), .ZN(n9151) );
  AOI22_X1 U13107 ( .A1(n27447), .A2(\xmem_data[52][4] ), .B1(n24130), .B2(
        \xmem_data[53][4] ), .ZN(n9150) );
  AOI22_X1 U13108 ( .A1(n30508), .A2(\xmem_data[54][4] ), .B1(n22675), .B2(
        \xmem_data[55][4] ), .ZN(n9149) );
  NAND4_X1 U13109 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n9158)
         );
  AOI22_X1 U13110 ( .A1(n30514), .A2(\xmem_data[56][4] ), .B1(n30513), .B2(
        \xmem_data[57][4] ), .ZN(n9156) );
  AOI22_X1 U13111 ( .A1(n28091), .A2(\xmem_data[58][4] ), .B1(n27516), .B2(
        \xmem_data[59][4] ), .ZN(n9155) );
  AOI22_X1 U13112 ( .A1(n25635), .A2(\xmem_data[60][4] ), .B1(n28492), .B2(
        \xmem_data[61][4] ), .ZN(n9154) );
  AOI22_X1 U13113 ( .A1(n21050), .A2(\xmem_data[62][4] ), .B1(n30515), .B2(
        \xmem_data[63][4] ), .ZN(n9153) );
  NAND4_X1 U13114 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n9157)
         );
  OR4_X1 U13115 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n9161)
         );
  NAND2_X1 U13116 ( .A1(n9161), .A2(n30565), .ZN(n9206) );
  AOI22_X1 U13117 ( .A1(n14972), .A2(\xmem_data[96][4] ), .B1(n21051), .B2(
        \xmem_data[97][4] ), .ZN(n9166) );
  AOI22_X1 U13118 ( .A1(n30600), .A2(\xmem_data[98][4] ), .B1(n30599), .B2(
        \xmem_data[99][4] ), .ZN(n9165) );
  AOI22_X1 U13119 ( .A1(n24685), .A2(\xmem_data[100][4] ), .B1(n29247), .B2(
        \xmem_data[101][4] ), .ZN(n9164) );
  AND2_X1 U13120 ( .A1(n30601), .A2(\xmem_data[103][4] ), .ZN(n9162) );
  AOI21_X1 U13121 ( .B1(n28241), .B2(\xmem_data[102][4] ), .A(n9162), .ZN(
        n9163) );
  AOI22_X1 U13122 ( .A1(n30592), .A2(\xmem_data[108][4] ), .B1(n3217), .B2(
        \xmem_data[109][4] ), .ZN(n9181) );
  AOI22_X1 U13123 ( .A1(n30606), .A2(\xmem_data[112][4] ), .B1(n13444), .B2(
        \xmem_data[113][4] ), .ZN(n9170) );
  AOI22_X1 U13124 ( .A1(n29157), .A2(\xmem_data[114][4] ), .B1(n29306), .B2(
        \xmem_data[115][4] ), .ZN(n9169) );
  AOI22_X1 U13125 ( .A1(n30607), .A2(\xmem_data[116][4] ), .B1(n28481), .B2(
        \xmem_data[117][4] ), .ZN(n9168) );
  AOI22_X1 U13126 ( .A1(n30608), .A2(\xmem_data[118][4] ), .B1(n24555), .B2(
        \xmem_data[119][4] ), .ZN(n9167) );
  NAND4_X1 U13127 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n9175)
         );
  AOI22_X1 U13128 ( .A1(n30588), .A2(\xmem_data[104][4] ), .B1(n28037), .B2(
        \xmem_data[105][4] ), .ZN(n9173) );
  AOI22_X1 U13129 ( .A1(n30593), .A2(\xmem_data[110][4] ), .B1(n25491), .B2(
        \xmem_data[111][4] ), .ZN(n9172) );
  AOI22_X1 U13130 ( .A1(n3348), .A2(\xmem_data[106][4] ), .B1(n30589), .B2(
        \xmem_data[107][4] ), .ZN(n9171) );
  NOR2_X1 U13131 ( .A1(n9175), .A2(n9174), .ZN(n9180) );
  AOI22_X1 U13132 ( .A1(n30614), .A2(\xmem_data[120][4] ), .B1(n30613), .B2(
        \xmem_data[121][4] ), .ZN(n9179) );
  AOI22_X1 U13133 ( .A1(n28154), .A2(\xmem_data[122][4] ), .B1(n30615), .B2(
        \xmem_data[123][4] ), .ZN(n9178) );
  AOI22_X1 U13134 ( .A1(n24509), .A2(\xmem_data[124][4] ), .B1(n23796), .B2(
        \xmem_data[125][4] ), .ZN(n9177) );
  AOI22_X1 U13135 ( .A1(n30617), .A2(\xmem_data[126][4] ), .B1(n30616), .B2(
        \xmem_data[127][4] ), .ZN(n9176) );
  NAND4_X1 U13136 ( .A1(n3864), .A2(n9181), .A3(n9180), .A4(n3530), .ZN(n9182)
         );
  NAND2_X1 U13137 ( .A1(n9182), .A2(n30626), .ZN(n9205) );
  AOI22_X1 U13138 ( .A1(n30557), .A2(\xmem_data[0][4] ), .B1(n20506), .B2(
        \xmem_data[1][4] ), .ZN(n9186) );
  AOI22_X1 U13139 ( .A1(n25401), .A2(\xmem_data[2][4] ), .B1(n23779), .B2(
        \xmem_data[3][4] ), .ZN(n9185) );
  AOI22_X1 U13140 ( .A1(n3171), .A2(\xmem_data[4][4] ), .B1(n25723), .B2(
        \xmem_data[5][4] ), .ZN(n9184) );
  AOI22_X1 U13141 ( .A1(n30674), .A2(\xmem_data[6][4] ), .B1(n30524), .B2(
        \xmem_data[7][4] ), .ZN(n9183) );
  NAND4_X1 U13142 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n9202)
         );
  AOI22_X1 U13143 ( .A1(n27564), .A2(\xmem_data[8][4] ), .B1(n22752), .B2(
        \xmem_data[9][4] ), .ZN(n9190) );
  AOI22_X1 U13144 ( .A1(n3228), .A2(\xmem_data[10][4] ), .B1(n27437), .B2(
        \xmem_data[11][4] ), .ZN(n9189) );
  AOI22_X1 U13145 ( .A1(n29254), .A2(\xmem_data[12][4] ), .B1(n3217), .B2(
        \xmem_data[13][4] ), .ZN(n9188) );
  AOI22_X1 U13146 ( .A1(n25448), .A2(\xmem_data[14][4] ), .B1(n30534), .B2(
        \xmem_data[15][4] ), .ZN(n9187) );
  NAND4_X1 U13147 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9187), .ZN(n9201)
         );
  AOI22_X1 U13148 ( .A1(n28475), .A2(\xmem_data[16][4] ), .B1(n30550), .B2(
        \xmem_data[17][4] ), .ZN(n9194) );
  AOI22_X1 U13149 ( .A1(n24702), .A2(\xmem_data[18][4] ), .B1(n25514), .B2(
        \xmem_data[19][4] ), .ZN(n9193) );
  AOI22_X1 U13150 ( .A1(n30551), .A2(\xmem_data[20][4] ), .B1(n13475), .B2(
        \xmem_data[21][4] ), .ZN(n9192) );
  AOI22_X1 U13151 ( .A1(n20545), .A2(\xmem_data[22][4] ), .B1(n30552), .B2(
        \xmem_data[23][4] ), .ZN(n9191) );
  NAND4_X1 U13152 ( .A1(n9194), .A2(n9193), .A3(n9192), .A4(n9191), .ZN(n9200)
         );
  AOI22_X1 U13153 ( .A1(n16986), .A2(\xmem_data[24][4] ), .B1(n30541), .B2(
        \xmem_data[25][4] ), .ZN(n9198) );
  AOI22_X1 U13154 ( .A1(n17018), .A2(\xmem_data[26][4] ), .B1(n30542), .B2(
        \xmem_data[27][4] ), .ZN(n9197) );
  AOI22_X1 U13155 ( .A1(n29010), .A2(\xmem_data[28][4] ), .B1(n30544), .B2(
        \xmem_data[29][4] ), .ZN(n9196) );
  AOI22_X1 U13156 ( .A1(n31255), .A2(\xmem_data[30][4] ), .B1(n30545), .B2(
        \xmem_data[31][4] ), .ZN(n9195) );
  NAND4_X1 U13157 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), .ZN(n9199)
         );
  OR4_X1 U13158 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), .ZN(n9203)
         );
  NAND2_X1 U13159 ( .A1(n9203), .A2(n30563), .ZN(n9204) );
  XNOR2_X1 U13160 ( .A(n31220), .B(\fmem_data[26][7] ), .ZN(n25146) );
  AOI22_X1 U13161 ( .A1(n16986), .A2(\xmem_data[96][7] ), .B1(n24597), .B2(
        \xmem_data[97][7] ), .ZN(n9211) );
  AOI22_X1 U13162 ( .A1(n16988), .A2(\xmem_data[98][7] ), .B1(n17019), .B2(
        \xmem_data[99][7] ), .ZN(n9210) );
  AOI22_X1 U13163 ( .A1(n20542), .A2(\xmem_data[100][7] ), .B1(n16989), .B2(
        \xmem_data[101][7] ), .ZN(n9209) );
  AOI22_X1 U13164 ( .A1(n16990), .A2(\xmem_data[102][7] ), .B1(n25399), .B2(
        \xmem_data[103][7] ), .ZN(n9208) );
  NAND4_X1 U13165 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n9229)
         );
  AOI22_X1 U13166 ( .A1(n30956), .A2(\xmem_data[104][7] ), .B1(n30955), .B2(
        \xmem_data[105][7] ), .ZN(n9215) );
  AOI22_X1 U13167 ( .A1(n3271), .A2(\xmem_data[106][7] ), .B1(n3200), .B2(
        \xmem_data[107][7] ), .ZN(n9214) );
  AOI22_X1 U13168 ( .A1(n20782), .A2(\xmem_data[108][7] ), .B1(n29136), .B2(
        \xmem_data[109][7] ), .ZN(n9213) );
  AOI22_X1 U13169 ( .A1(n30901), .A2(\xmem_data[110][7] ), .B1(n22727), .B2(
        \xmem_data[111][7] ), .ZN(n9212) );
  NAND4_X1 U13170 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n9228)
         );
  AND2_X1 U13171 ( .A1(n3222), .A2(\xmem_data[117][7] ), .ZN(n9216) );
  AOI21_X1 U13172 ( .B1(n25692), .B2(\xmem_data[116][7] ), .A(n9216), .ZN(
        n9221) );
  AOI22_X1 U13173 ( .A1(n16980), .A2(\xmem_data[114][7] ), .B1(n16979), .B2(
        \xmem_data[115][7] ), .ZN(n9220) );
  AND2_X1 U13174 ( .A1(n20986), .A2(\xmem_data[112][7] ), .ZN(n9217) );
  AOI21_X1 U13175 ( .B1(n25561), .B2(\xmem_data[113][7] ), .A(n9217), .ZN(
        n9219) );
  AOI22_X1 U13176 ( .A1(n25414), .A2(\xmem_data[118][7] ), .B1(n24695), .B2(
        \xmem_data[119][7] ), .ZN(n9218) );
  NAND4_X1 U13177 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(n9227)
         );
  AOI22_X1 U13178 ( .A1(n29174), .A2(\xmem_data[120][7] ), .B1(n3256), .B2(
        \xmem_data[121][7] ), .ZN(n9225) );
  AOI22_X1 U13179 ( .A1(n16973), .A2(\xmem_data[122][7] ), .B1(n16972), .B2(
        \xmem_data[123][7] ), .ZN(n9224) );
  AOI22_X1 U13180 ( .A1(n16974), .A2(\xmem_data[124][7] ), .B1(n29180), .B2(
        \xmem_data[125][7] ), .ZN(n9223) );
  AOI22_X1 U13181 ( .A1(n30943), .A2(\xmem_data[126][7] ), .B1(n25423), .B2(
        \xmem_data[127][7] ), .ZN(n9222) );
  NAND4_X1 U13182 ( .A1(n9225), .A2(n9224), .A3(n9223), .A4(n9222), .ZN(n9226)
         );
  OR4_X1 U13183 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(n9230)
         );
  NAND2_X1 U13184 ( .A1(n9230), .A2(n16997), .ZN(n9297) );
  AOI22_X1 U13185 ( .A1(n28298), .A2(\xmem_data[64][7] ), .B1(n24160), .B2(
        \xmem_data[65][7] ), .ZN(n9234) );
  AOI22_X1 U13186 ( .A1(n20776), .A2(\xmem_data[66][7] ), .B1(n3202), .B2(
        \xmem_data[67][7] ), .ZN(n9233) );
  AOI22_X1 U13187 ( .A1(n17020), .A2(\xmem_data[68][7] ), .B1(n28427), .B2(
        \xmem_data[69][7] ), .ZN(n9232) );
  AOI22_X1 U13188 ( .A1(n17021), .A2(\xmem_data[70][7] ), .B1(n29238), .B2(
        \xmem_data[71][7] ), .ZN(n9231) );
  NAND4_X1 U13189 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n9250)
         );
  AOI22_X1 U13190 ( .A1(n3326), .A2(\xmem_data[72][7] ), .B1(n17001), .B2(
        \xmem_data[73][7] ), .ZN(n9238) );
  AOI22_X1 U13191 ( .A1(n17004), .A2(\xmem_data[74][7] ), .B1(n3201), .B2(
        \xmem_data[75][7] ), .ZN(n9237) );
  AOI22_X1 U13192 ( .A1(n20552), .A2(\xmem_data[76][7] ), .B1(n17003), .B2(
        \xmem_data[77][7] ), .ZN(n9236) );
  AOI22_X1 U13193 ( .A1(n23730), .A2(\xmem_data[78][7] ), .B1(n16999), .B2(
        \xmem_data[79][7] ), .ZN(n9235) );
  NAND4_X1 U13194 ( .A1(n9238), .A2(n9237), .A3(n9236), .A4(n9235), .ZN(n9249)
         );
  AOI22_X1 U13195 ( .A1(n17030), .A2(\xmem_data[80][7] ), .B1(n20709), .B2(
        \xmem_data[81][7] ), .ZN(n9242) );
  AOI22_X1 U13196 ( .A1(n3388), .A2(\xmem_data[82][7] ), .B1(n17031), .B2(
        \xmem_data[83][7] ), .ZN(n9241) );
  AOI22_X1 U13197 ( .A1(n24562), .A2(\xmem_data[84][7] ), .B1(n3219), .B2(
        \xmem_data[85][7] ), .ZN(n9240) );
  AOI22_X1 U13198 ( .A1(n17033), .A2(\xmem_data[86][7] ), .B1(n29255), .B2(
        \xmem_data[87][7] ), .ZN(n9239) );
  NAND4_X1 U13199 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n9248)
         );
  AOI22_X1 U13200 ( .A1(n17010), .A2(\xmem_data[88][7] ), .B1(n22669), .B2(
        \xmem_data[89][7] ), .ZN(n9246) );
  AOI22_X1 U13201 ( .A1(n20808), .A2(\xmem_data[90][7] ), .B1(n17011), .B2(
        \xmem_data[91][7] ), .ZN(n9245) );
  AOI22_X1 U13202 ( .A1(n25422), .A2(\xmem_data[92][7] ), .B1(n13475), .B2(
        \xmem_data[93][7] ), .ZN(n9244) );
  AOI22_X1 U13203 ( .A1(n17013), .A2(\xmem_data[94][7] ), .B1(n17012), .B2(
        \xmem_data[95][7] ), .ZN(n9243) );
  NAND4_X1 U13204 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n9247)
         );
  OR4_X1 U13205 ( .A1(n9250), .A2(n9249), .A3(n9248), .A4(n9247), .ZN(n9251)
         );
  NAND2_X1 U13206 ( .A1(n9251), .A2(n16966), .ZN(n9296) );
  AOI22_X1 U13207 ( .A1(n30891), .A2(\xmem_data[32][7] ), .B1(n20717), .B2(
        \xmem_data[33][7] ), .ZN(n9255) );
  AOI22_X1 U13208 ( .A1(n30746), .A2(\xmem_data[34][7] ), .B1(n17019), .B2(
        \xmem_data[35][7] ), .ZN(n9254) );
  AOI22_X1 U13209 ( .A1(n17020), .A2(\xmem_data[36][7] ), .B1(n24219), .B2(
        \xmem_data[37][7] ), .ZN(n9253) );
  AOI22_X1 U13210 ( .A1(n17021), .A2(\xmem_data[38][7] ), .B1(n30515), .B2(
        \xmem_data[39][7] ), .ZN(n9252) );
  NAND4_X1 U13211 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n9271)
         );
  AOI22_X1 U13212 ( .A1(n3326), .A2(\xmem_data[40][7] ), .B1(n17001), .B2(
        \xmem_data[41][7] ), .ZN(n9259) );
  AOI22_X1 U13213 ( .A1(n17004), .A2(\xmem_data[42][7] ), .B1(n3199), .B2(
        \xmem_data[43][7] ), .ZN(n9258) );
  AOI22_X1 U13214 ( .A1(n3172), .A2(\xmem_data[44][7] ), .B1(n17003), .B2(
        \xmem_data[45][7] ), .ZN(n9257) );
  AOI22_X1 U13215 ( .A1(n20770), .A2(\xmem_data[46][7] ), .B1(n16999), .B2(
        \xmem_data[47][7] ), .ZN(n9256) );
  NAND4_X1 U13216 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n9270)
         );
  AOI22_X1 U13217 ( .A1(n17030), .A2(\xmem_data[48][7] ), .B1(n12471), .B2(
        \xmem_data[49][7] ), .ZN(n9263) );
  AOI22_X1 U13218 ( .A1(n3388), .A2(\xmem_data[50][7] ), .B1(n17031), .B2(
        \xmem_data[51][7] ), .ZN(n9262) );
  AOI22_X1 U13219 ( .A1(n30962), .A2(\xmem_data[52][7] ), .B1(n3218), .B2(
        \xmem_data[53][7] ), .ZN(n9261) );
  AOI22_X1 U13220 ( .A1(n17033), .A2(\xmem_data[54][7] ), .B1(n22667), .B2(
        \xmem_data[55][7] ), .ZN(n9260) );
  NAND4_X1 U13221 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n9269)
         );
  AOI22_X1 U13222 ( .A1(n17010), .A2(\xmem_data[56][7] ), .B1(n30550), .B2(
        \xmem_data[57][7] ), .ZN(n9267) );
  AOI22_X1 U13223 ( .A1(n29350), .A2(\xmem_data[58][7] ), .B1(n17011), .B2(
        \xmem_data[59][7] ), .ZN(n9266) );
  AOI22_X1 U13224 ( .A1(n25422), .A2(\xmem_data[60][7] ), .B1(n27863), .B2(
        \xmem_data[61][7] ), .ZN(n9265) );
  AOI22_X1 U13225 ( .A1(n17013), .A2(\xmem_data[62][7] ), .B1(n17012), .B2(
        \xmem_data[63][7] ), .ZN(n9264) );
  NAND4_X1 U13226 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n9268)
         );
  OR4_X1 U13227 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9272)
         );
  NAND2_X1 U13228 ( .A1(n9272), .A2(n17038), .ZN(n9295) );
  AOI22_X1 U13229 ( .A1(n17041), .A2(\xmem_data[0][7] ), .B1(n24160), .B2(
        \xmem_data[1][7] ), .ZN(n9276) );
  AOI22_X1 U13230 ( .A1(n3465), .A2(\xmem_data[2][7] ), .B1(n3202), .B2(
        \xmem_data[3][7] ), .ZN(n9275) );
  AOI22_X1 U13231 ( .A1(n24708), .A2(\xmem_data[4][7] ), .B1(n17043), .B2(
        \xmem_data[5][7] ), .ZN(n9274) );
  AOI22_X1 U13232 ( .A1(n17044), .A2(\xmem_data[6][7] ), .B1(n28301), .B2(
        \xmem_data[7][7] ), .ZN(n9273) );
  NAND4_X1 U13233 ( .A1(n9276), .A2(n9275), .A3(n9274), .A4(n9273), .ZN(n9292)
         );
  AOI22_X1 U13234 ( .A1(n3205), .A2(\xmem_data[8][7] ), .B1(n20816), .B2(
        \xmem_data[9][7] ), .ZN(n9280) );
  AOI22_X1 U13235 ( .A1(n28461), .A2(\xmem_data[10][7] ), .B1(n3200), .B2(
        \xmem_data[11][7] ), .ZN(n9279) );
  AOI22_X1 U13236 ( .A1(n21058), .A2(\xmem_data[12][7] ), .B1(n17049), .B2(
        \xmem_data[13][7] ), .ZN(n9278) );
  AOI22_X1 U13237 ( .A1(n17051), .A2(\xmem_data[14][7] ), .B1(n17050), .B2(
        \xmem_data[15][7] ), .ZN(n9277) );
  NAND4_X1 U13238 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n9291)
         );
  AOI22_X1 U13239 ( .A1(n17056), .A2(\xmem_data[16][7] ), .B1(n28037), .B2(
        \xmem_data[17][7] ), .ZN(n9284) );
  AOI22_X1 U13240 ( .A1(n20828), .A2(\xmem_data[18][7] ), .B1(n16979), .B2(
        \xmem_data[19][7] ), .ZN(n9283) );
  AOI22_X1 U13241 ( .A1(n23756), .A2(\xmem_data[20][7] ), .B1(n3220), .B2(
        \xmem_data[21][7] ), .ZN(n9282) );
  AOI22_X1 U13242 ( .A1(n20724), .A2(\xmem_data[22][7] ), .B1(n23739), .B2(
        \xmem_data[23][7] ), .ZN(n9281) );
  NAND4_X1 U13243 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n9290)
         );
  AOI22_X1 U13244 ( .A1(n25617), .A2(\xmem_data[24][7] ), .B1(n17061), .B2(
        \xmem_data[25][7] ), .ZN(n9288) );
  AOI22_X1 U13245 ( .A1(n17063), .A2(\xmem_data[26][7] ), .B1(n17062), .B2(
        \xmem_data[27][7] ), .ZN(n9287) );
  AOI22_X1 U13246 ( .A1(n27447), .A2(\xmem_data[28][7] ), .B1(n14996), .B2(
        \xmem_data[29][7] ), .ZN(n9286) );
  AOI22_X1 U13247 ( .A1(n17064), .A2(\xmem_data[30][7] ), .B1(n21015), .B2(
        \xmem_data[31][7] ), .ZN(n9285) );
  NAND4_X1 U13248 ( .A1(n9288), .A2(n9287), .A3(n9286), .A4(n9285), .ZN(n9289)
         );
  OR4_X1 U13249 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n9293)
         );
  NAND2_X1 U13250 ( .A1(n9293), .A2(n17073), .ZN(n9294) );
  XNOR2_X1 U13251 ( .A(n35336), .B(\fmem_data[2][5] ), .ZN(n35017) );
  AOI22_X1 U13252 ( .A1(n16986), .A2(\xmem_data[96][6] ), .B1(n29009), .B2(
        \xmem_data[97][6] ), .ZN(n9301) );
  AOI22_X1 U13253 ( .A1(n16988), .A2(\xmem_data[98][6] ), .B1(n16987), .B2(
        \xmem_data[99][6] ), .ZN(n9300) );
  AOI22_X1 U13254 ( .A1(n23717), .A2(\xmem_data[100][6] ), .B1(n16989), .B2(
        \xmem_data[101][6] ), .ZN(n9299) );
  AOI22_X1 U13255 ( .A1(n16990), .A2(\xmem_data[102][6] ), .B1(n31254), .B2(
        \xmem_data[103][6] ), .ZN(n9298) );
  NAND4_X1 U13256 ( .A1(n9301), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(n9317)
         );
  AOI22_X1 U13257 ( .A1(n24647), .A2(\xmem_data[104][6] ), .B1(n21051), .B2(
        \xmem_data[105][6] ), .ZN(n9305) );
  AOI22_X1 U13258 ( .A1(n3271), .A2(\xmem_data[106][6] ), .B1(n3199), .B2(
        \xmem_data[107][6] ), .ZN(n9304) );
  AOI22_X1 U13259 ( .A1(n24467), .A2(\xmem_data[108][6] ), .B1(n17003), .B2(
        \xmem_data[109][6] ), .ZN(n9303) );
  AOI22_X1 U13260 ( .A1(n25407), .A2(\xmem_data[110][6] ), .B1(n31344), .B2(
        \xmem_data[111][6] ), .ZN(n9302) );
  NAND4_X1 U13261 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n9316)
         );
  AOI22_X1 U13262 ( .A1(n24532), .A2(\xmem_data[116][6] ), .B1(n3219), .B2(
        \xmem_data[117][6] ), .ZN(n9309) );
  AOI22_X1 U13263 ( .A1(n16980), .A2(\xmem_data[114][6] ), .B1(n16979), .B2(
        \xmem_data[115][6] ), .ZN(n9308) );
  AOI22_X1 U13264 ( .A1(n20953), .A2(\xmem_data[112][6] ), .B1(n25685), .B2(
        \xmem_data[113][6] ), .ZN(n9307) );
  AOI22_X1 U13265 ( .A1(n25448), .A2(\xmem_data[118][6] ), .B1(n24695), .B2(
        \xmem_data[119][6] ), .ZN(n9306) );
  NAND4_X1 U13266 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n9315)
         );
  AOI22_X1 U13267 ( .A1(n20725), .A2(\xmem_data[120][6] ), .B1(n27550), .B2(
        \xmem_data[121][6] ), .ZN(n9313) );
  AOI22_X1 U13268 ( .A1(n16973), .A2(\xmem_data[122][6] ), .B1(n16972), .B2(
        \xmem_data[123][6] ), .ZN(n9312) );
  AOI22_X1 U13269 ( .A1(n16974), .A2(\xmem_data[124][6] ), .B1(n29180), .B2(
        \xmem_data[125][6] ), .ZN(n9311) );
  AOI22_X1 U13270 ( .A1(n31327), .A2(\xmem_data[126][6] ), .B1(n13168), .B2(
        \xmem_data[127][6] ), .ZN(n9310) );
  NAND4_X1 U13271 ( .A1(n9313), .A2(n9312), .A3(n9311), .A4(n9310), .ZN(n9314)
         );
  OR4_X1 U13272 ( .A1(n9317), .A2(n9316), .A3(n9315), .A4(n9314), .ZN(n9318)
         );
  NAND2_X1 U13273 ( .A1(n9318), .A2(n16997), .ZN(n9385) );
  AOI22_X1 U13274 ( .A1(n17041), .A2(\xmem_data[0][6] ), .B1(n20717), .B2(
        \xmem_data[1][6] ), .ZN(n9322) );
  AOI22_X1 U13275 ( .A1(n24458), .A2(\xmem_data[2][6] ), .B1(n16987), .B2(
        \xmem_data[3][6] ), .ZN(n9321) );
  AOI22_X1 U13276 ( .A1(n24133), .A2(\xmem_data[4][6] ), .B1(n17043), .B2(
        \xmem_data[5][6] ), .ZN(n9320) );
  AOI22_X1 U13277 ( .A1(n17044), .A2(\xmem_data[6][6] ), .B1(n24709), .B2(
        \xmem_data[7][6] ), .ZN(n9319) );
  NAND4_X1 U13278 ( .A1(n9322), .A2(n9321), .A3(n9320), .A4(n9319), .ZN(n9338)
         );
  AOI22_X1 U13279 ( .A1(n24190), .A2(\xmem_data[8][6] ), .B1(n29281), .B2(
        \xmem_data[9][6] ), .ZN(n9326) );
  AOI22_X1 U13280 ( .A1(n25636), .A2(\xmem_data[10][6] ), .B1(n3201), .B2(
        \xmem_data[11][6] ), .ZN(n9325) );
  AOI22_X1 U13281 ( .A1(n29325), .A2(\xmem_data[12][6] ), .B1(n17049), .B2(
        \xmem_data[13][6] ), .ZN(n9324) );
  AOI22_X1 U13282 ( .A1(n17051), .A2(\xmem_data[14][6] ), .B1(n17050), .B2(
        \xmem_data[15][6] ), .ZN(n9323) );
  NAND4_X1 U13283 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9323), .ZN(n9337)
         );
  AOI22_X1 U13284 ( .A1(n17056), .A2(\xmem_data[16][6] ), .B1(n12471), .B2(
        \xmem_data[17][6] ), .ZN(n9330) );
  AOI22_X1 U13285 ( .A1(n3245), .A2(\xmem_data[18][6] ), .B1(n16979), .B2(
        \xmem_data[19][6] ), .ZN(n9329) );
  AOI22_X1 U13286 ( .A1(n25692), .A2(\xmem_data[20][6] ), .B1(n3222), .B2(
        \xmem_data[21][6] ), .ZN(n9328) );
  AOI22_X1 U13287 ( .A1(n25731), .A2(\xmem_data[22][6] ), .B1(n23739), .B2(
        \xmem_data[23][6] ), .ZN(n9327) );
  NAND4_X1 U13288 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(n9336)
         );
  AOI22_X1 U13289 ( .A1(n24565), .A2(\xmem_data[24][6] ), .B1(n17061), .B2(
        \xmem_data[25][6] ), .ZN(n9334) );
  AOI22_X1 U13290 ( .A1(n17063), .A2(\xmem_data[26][6] ), .B1(n17062), .B2(
        \xmem_data[27][6] ), .ZN(n9333) );
  AOI22_X1 U13291 ( .A1(n25422), .A2(\xmem_data[28][6] ), .B1(n24590), .B2(
        \xmem_data[29][6] ), .ZN(n9332) );
  AOI22_X1 U13292 ( .A1(n17064), .A2(\xmem_data[30][6] ), .B1(n28416), .B2(
        \xmem_data[31][6] ), .ZN(n9331) );
  NAND4_X1 U13293 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n9335)
         );
  OR4_X1 U13294 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n9339)
         );
  NAND2_X1 U13295 ( .A1(n9339), .A2(n17073), .ZN(n9384) );
  AOI22_X1 U13296 ( .A1(n16986), .A2(\xmem_data[32][6] ), .B1(n30541), .B2(
        \xmem_data[33][6] ), .ZN(n9343) );
  AOI22_X1 U13297 ( .A1(n31354), .A2(\xmem_data[34][6] ), .B1(n16987), .B2(
        \xmem_data[35][6] ), .ZN(n9342) );
  AOI22_X1 U13298 ( .A1(n17020), .A2(\xmem_data[36][6] ), .B1(n31270), .B2(
        \xmem_data[37][6] ), .ZN(n9341) );
  AOI22_X1 U13299 ( .A1(n17021), .A2(\xmem_data[38][6] ), .B1(n27920), .B2(
        \xmem_data[39][6] ), .ZN(n9340) );
  NAND4_X1 U13300 ( .A1(n9343), .A2(n9342), .A3(n9341), .A4(n9340), .ZN(n9359)
         );
  AOI22_X1 U13301 ( .A1(n28460), .A2(\xmem_data[40][6] ), .B1(n17001), .B2(
        \xmem_data[41][6] ), .ZN(n9347) );
  AOI22_X1 U13302 ( .A1(n17004), .A2(\xmem_data[42][6] ), .B1(n3201), .B2(
        \xmem_data[43][6] ), .ZN(n9346) );
  AOI22_X1 U13303 ( .A1(n25526), .A2(\xmem_data[44][6] ), .B1(n17003), .B2(
        \xmem_data[45][6] ), .ZN(n9345) );
  AOI22_X1 U13304 ( .A1(n14982), .A2(\xmem_data[46][6] ), .B1(n16999), .B2(
        \xmem_data[47][6] ), .ZN(n9344) );
  NAND4_X1 U13305 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9358)
         );
  AOI22_X1 U13306 ( .A1(n17030), .A2(\xmem_data[48][6] ), .B1(n29118), .B2(
        \xmem_data[49][6] ), .ZN(n9351) );
  AOI22_X1 U13307 ( .A1(n3387), .A2(\xmem_data[50][6] ), .B1(n17031), .B2(
        \xmem_data[51][6] ), .ZN(n9350) );
  AOI22_X1 U13308 ( .A1(n28364), .A2(\xmem_data[52][6] ), .B1(n3221), .B2(
        \xmem_data[53][6] ), .ZN(n9349) );
  AOI22_X1 U13309 ( .A1(n17033), .A2(\xmem_data[54][6] ), .B1(n23769), .B2(
        \xmem_data[55][6] ), .ZN(n9348) );
  NAND4_X1 U13310 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n9357)
         );
  AOI22_X1 U13311 ( .A1(n17010), .A2(\xmem_data[56][6] ), .B1(n22711), .B2(
        \xmem_data[57][6] ), .ZN(n9355) );
  AOI22_X1 U13312 ( .A1(n25377), .A2(\xmem_data[58][6] ), .B1(n17011), .B2(
        \xmem_data[59][6] ), .ZN(n9354) );
  AOI22_X1 U13313 ( .A1(n25707), .A2(\xmem_data[60][6] ), .B1(n25481), .B2(
        \xmem_data[61][6] ), .ZN(n9353) );
  AOI22_X1 U13314 ( .A1(n17013), .A2(\xmem_data[62][6] ), .B1(n17012), .B2(
        \xmem_data[63][6] ), .ZN(n9352) );
  NAND4_X1 U13315 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9356)
         );
  OR4_X1 U13316 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n9360)
         );
  NAND2_X1 U13317 ( .A1(n9360), .A2(n17038), .ZN(n9383) );
  AOI22_X1 U13318 ( .A1(n16986), .A2(\xmem_data[64][6] ), .B1(n20544), .B2(
        \xmem_data[65][6] ), .ZN(n9364) );
  AOI22_X1 U13319 ( .A1(n23795), .A2(n20682), .B1(n3202), .B2(
        \xmem_data[67][6] ), .ZN(n9363) );
  AOI22_X1 U13320 ( .A1(n17020), .A2(\xmem_data[68][6] ), .B1(n23796), .B2(
        \xmem_data[69][6] ), .ZN(n9362) );
  AOI22_X1 U13321 ( .A1(n17021), .A2(\xmem_data[70][6] ), .B1(n27523), .B2(
        \xmem_data[71][6] ), .ZN(n9361) );
  NAND4_X1 U13322 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9380)
         );
  AOI22_X1 U13323 ( .A1(n24615), .A2(\xmem_data[72][6] ), .B1(n17001), .B2(
        \xmem_data[73][6] ), .ZN(n9368) );
  AOI22_X1 U13324 ( .A1(n17004), .A2(\xmem_data[74][6] ), .B1(n3199), .B2(
        \xmem_data[75][6] ), .ZN(n9367) );
  AOI22_X1 U13325 ( .A1(n20782), .A2(\xmem_data[76][6] ), .B1(n17003), .B2(
        \xmem_data[77][6] ), .ZN(n9366) );
  AOI22_X1 U13326 ( .A1(n25628), .A2(\xmem_data[78][6] ), .B1(n16999), .B2(
        \xmem_data[79][6] ), .ZN(n9365) );
  NAND4_X1 U13327 ( .A1(n9368), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n9379)
         );
  AOI22_X1 U13328 ( .A1(n17030), .A2(\xmem_data[80][6] ), .B1(n25685), .B2(
        \xmem_data[81][6] ), .ZN(n9372) );
  AOI22_X1 U13329 ( .A1(n3387), .A2(\xmem_data[82][6] ), .B1(n17031), .B2(
        \xmem_data[83][6] ), .ZN(n9371) );
  AOI22_X1 U13330 ( .A1(n25730), .A2(\xmem_data[84][6] ), .B1(n3222), .B2(
        \xmem_data[85][6] ), .ZN(n9370) );
  AOI22_X1 U13331 ( .A1(n17033), .A2(\xmem_data[86][6] ), .B1(n29028), .B2(
        \xmem_data[87][6] ), .ZN(n9369) );
  NAND4_X1 U13332 ( .A1(n9372), .A2(n9371), .A3(n9370), .A4(n9369), .ZN(n9378)
         );
  AOI22_X1 U13333 ( .A1(n17010), .A2(\xmem_data[88][6] ), .B1(n29181), .B2(
        \xmem_data[89][6] ), .ZN(n9376) );
  AOI22_X1 U13334 ( .A1(n16973), .A2(\xmem_data[90][6] ), .B1(n17011), .B2(
        \xmem_data[91][6] ), .ZN(n9375) );
  AOI22_X1 U13335 ( .A1(n30551), .A2(\xmem_data[92][6] ), .B1(n24130), .B2(
        \xmem_data[93][6] ), .ZN(n9374) );
  AOI22_X1 U13336 ( .A1(n17013), .A2(\xmem_data[94][6] ), .B1(n17012), .B2(
        \xmem_data[95][6] ), .ZN(n9373) );
  NAND4_X1 U13337 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n9377)
         );
  OR4_X1 U13338 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n9381)
         );
  NAND2_X1 U13339 ( .A1(n9381), .A2(n16966), .ZN(n9382) );
  XNOR2_X1 U13340 ( .A(n32014), .B(\fmem_data[2][5] ), .ZN(n12809) );
  XOR2_X1 U13341 ( .A(\fmem_data[2][4] ), .B(\fmem_data[2][5] ), .Z(n9386) );
  BUF_X1 U13342 ( .A(n14919), .Z(n25359) );
  AOI22_X1 U13343 ( .A1(n24606), .A2(\xmem_data[8][5] ), .B1(n25359), .B2(
        \xmem_data[9][5] ), .ZN(n9390) );
  BUF_X1 U13344 ( .A(n13487), .Z(n25388) );
  AOI22_X1 U13345 ( .A1(n28772), .A2(\xmem_data[10][5] ), .B1(n25388), .B2(
        \xmem_data[11][5] ), .ZN(n9389) );
  BUF_X1 U13346 ( .A(n31263), .Z(n25358) );
  AOI22_X1 U13347 ( .A1(n25358), .A2(\xmem_data[12][5] ), .B1(n25357), .B2(
        \xmem_data[13][5] ), .ZN(n9388) );
  AOI22_X1 U13348 ( .A1(n27813), .A2(\xmem_data[14][5] ), .B1(n25360), .B2(
        \xmem_data[15][5] ), .ZN(n9387) );
  NAND4_X1 U13349 ( .A1(n9390), .A2(n9389), .A3(n9388), .A4(n9387), .ZN(n9397)
         );
  AOI22_X1 U13350 ( .A1(n28152), .A2(\xmem_data[26][5] ), .B1(n20958), .B2(
        \xmem_data[27][5] ), .ZN(n9395) );
  BUF_X1 U13351 ( .A(n14898), .Z(n25382) );
  NAND2_X1 U13352 ( .A1(n25456), .A2(\xmem_data[25][5] ), .ZN(n9392) );
  NAND2_X1 U13353 ( .A1(n3465), .A2(\xmem_data[30][5] ), .ZN(n9391) );
  NAND2_X1 U13354 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  AOI21_X1 U13355 ( .B1(\xmem_data[29][5] ), .B2(n25382), .A(n9393), .ZN(n9394) );
  NAND2_X1 U13356 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  OR3_X1 U13357 ( .A1(n9397), .A2(n9396), .A3(n4016), .ZN(n9416) );
  BUF_X1 U13358 ( .A(n29064), .Z(n25354) );
  AOI22_X1 U13359 ( .A1(n25354), .A2(\xmem_data[16][5] ), .B1(n3219), .B2(
        \xmem_data[17][5] ), .ZN(n9398) );
  INV_X1 U13360 ( .A(n9398), .ZN(n9405) );
  NAND2_X1 U13361 ( .A1(n28374), .A2(\xmem_data[24][5] ), .ZN(n9400) );
  NAND2_X1 U13362 ( .A1(n17041), .A2(\xmem_data[28][5] ), .ZN(n9399) );
  AND2_X1 U13363 ( .A1(n9400), .A2(n9399), .ZN(n9403) );
  AOI22_X1 U13364 ( .A1(n29257), .A2(\xmem_data[20][5] ), .B1(n20993), .B2(
        \xmem_data[21][5] ), .ZN(n9402) );
  BUF_X1 U13365 ( .A(n14991), .Z(n25377) );
  NAND2_X1 U13366 ( .A1(n25377), .A2(\xmem_data[22][5] ), .ZN(n9401) );
  NAND3_X1 U13367 ( .A1(n9403), .A2(n9402), .A3(n9401), .ZN(n9404) );
  NOR2_X1 U13368 ( .A1(n9405), .A2(n9404), .ZN(n9414) );
  AOI22_X1 U13369 ( .A1(n30949), .A2(\xmem_data[0][5] ), .B1(n24645), .B2(
        \xmem_data[1][5] ), .ZN(n9409) );
  BUF_X1 U13370 ( .A(n13452), .Z(n25367) );
  AOI22_X1 U13371 ( .A1(n17021), .A2(\xmem_data[2][5] ), .B1(n25367), .B2(
        \xmem_data[3][5] ), .ZN(n9408) );
  BUF_X1 U13372 ( .A(n14973), .Z(n25364) );
  AOI22_X1 U13373 ( .A1(n3178), .A2(\xmem_data[4][5] ), .B1(n25364), .B2(
        \xmem_data[5][5] ), .ZN(n9407) );
  AOI22_X1 U13374 ( .A1(n20817), .A2(\xmem_data[6][5] ), .B1(n29126), .B2(
        \xmem_data[7][5] ), .ZN(n9406) );
  NAND4_X1 U13375 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n9412)
         );
  AOI22_X1 U13376 ( .A1(n29431), .A2(\xmem_data[18][5] ), .B1(n29028), .B2(
        \xmem_data[19][5] ), .ZN(n9410) );
  NAND2_X1 U13377 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  OR2_X1 U13378 ( .A1(n9416), .A2(n9415), .ZN(n9422) );
  AND2_X1 U13379 ( .A1(n23771), .A2(\xmem_data[23][5] ), .ZN(n9421) );
  INV_X1 U13380 ( .A(n9420), .ZN(n9419) );
  AOI21_X1 U13381 ( .B1(load_xaddr_val[5]), .B2(n9419), .A(n9418), .ZN(n9466)
         );
  AOI22_X1 U13382 ( .A1(n9420), .A2(n39040), .B1(n14909), .B2(n9419), .ZN(
        n9444) );
  NOR2_X1 U13383 ( .A1(n9466), .A2(n9444), .ZN(n16443) );
  OAI21_X1 U13384 ( .B1(n9422), .B2(n9421), .A(n16443), .ZN(n9491) );
  BUF_X1 U13385 ( .A(n14937), .Z(n25434) );
  AOI22_X1 U13386 ( .A1(n25434), .A2(\xmem_data[32][5] ), .B1(n31329), .B2(
        \xmem_data[33][5] ), .ZN(n9426) );
  AOI22_X1 U13387 ( .A1(n30617), .A2(\xmem_data[34][5] ), .B1(n25435), .B2(
        \xmem_data[35][5] ), .ZN(n9425) );
  AOI22_X1 U13388 ( .A1(n24461), .A2(\xmem_data[36][5] ), .B1(n27856), .B2(
        \xmem_data[37][5] ), .ZN(n9424) );
  AOI22_X1 U13389 ( .A1(n3308), .A2(\xmem_data[38][5] ), .B1(n28495), .B2(
        \xmem_data[39][5] ), .ZN(n9423) );
  NAND4_X1 U13390 ( .A1(n9426), .A2(n9425), .A3(n9424), .A4(n9423), .ZN(n9442)
         );
  AOI22_X1 U13391 ( .A1(n13486), .A2(\xmem_data[40][5] ), .B1(n30496), .B2(
        \xmem_data[41][5] ), .ZN(n9430) );
  BUF_X1 U13392 ( .A(n13487), .Z(n25440) );
  AOI22_X1 U13393 ( .A1(n28192), .A2(\xmem_data[42][5] ), .B1(n25440), .B2(
        \xmem_data[43][5] ), .ZN(n9429) );
  BUF_X1 U13394 ( .A(n31263), .Z(n25441) );
  AOI22_X1 U13395 ( .A1(n25441), .A2(\xmem_data[44][5] ), .B1(n25629), .B2(
        \xmem_data[45][5] ), .ZN(n9428) );
  BUF_X1 U13396 ( .A(n28973), .Z(n25443) );
  BUF_X1 U13397 ( .A(n13468), .Z(n25442) );
  AOI22_X1 U13398 ( .A1(n25443), .A2(\xmem_data[46][5] ), .B1(n25442), .B2(
        \xmem_data[47][5] ), .ZN(n9427) );
  NAND4_X1 U13399 ( .A1(n9430), .A2(n9429), .A3(n9428), .A4(n9427), .ZN(n9441)
         );
  AOI22_X1 U13400 ( .A1(n30906), .A2(\xmem_data[48][5] ), .B1(n3222), .B2(
        \xmem_data[49][5] ), .ZN(n9434) );
  BUF_X1 U13401 ( .A(n14988), .Z(n25448) );
  AOI22_X1 U13402 ( .A1(n25448), .A2(\xmem_data[50][5] ), .B1(n31367), .B2(
        \xmem_data[51][5] ), .ZN(n9433) );
  BUF_X1 U13403 ( .A(n14990), .Z(n25449) );
  AOI22_X1 U13404 ( .A1(n25449), .A2(\xmem_data[52][5] ), .B1(n24140), .B2(
        \xmem_data[53][5] ), .ZN(n9432) );
  BUF_X1 U13405 ( .A(n14991), .Z(n25451) );
  AOI22_X1 U13406 ( .A1(n25451), .A2(\xmem_data[54][5] ), .B1(n24553), .B2(
        \xmem_data[55][5] ), .ZN(n9431) );
  NAND4_X1 U13407 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(n9440)
         );
  BUF_X1 U13408 ( .A(n14933), .Z(n25456) );
  AOI22_X1 U13409 ( .A1(n20809), .A2(\xmem_data[56][5] ), .B1(n3358), .B2(
        \xmem_data[57][5] ), .ZN(n9438) );
  BUF_X1 U13410 ( .A(n14997), .Z(n25457) );
  AOI22_X1 U13411 ( .A1(n25457), .A2(\xmem_data[58][5] ), .B1(n24132), .B2(
        \xmem_data[59][5] ), .ZN(n9437) );
  BUF_X1 U13412 ( .A(n13476), .Z(n25459) );
  BUF_X1 U13413 ( .A(n14999), .Z(n25458) );
  AOI22_X1 U13414 ( .A1(n25459), .A2(\xmem_data[60][5] ), .B1(n25458), .B2(
        \xmem_data[61][5] ), .ZN(n9436) );
  BUF_X1 U13415 ( .A(n29187), .Z(n25461) );
  BUF_X1 U13416 ( .A(n15000), .Z(n25460) );
  AOI22_X1 U13417 ( .A1(n3466), .A2(\xmem_data[62][5] ), .B1(n25460), .B2(
        \xmem_data[63][5] ), .ZN(n9435) );
  NAND4_X1 U13418 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(n9439)
         );
  OR4_X1 U13419 ( .A1(n9442), .A2(n9441), .A3(n9440), .A4(n9439), .ZN(n9443)
         );
  INV_X1 U13420 ( .A(n9444), .ZN(n9465) );
  AND2_X1 U13421 ( .A1(n9465), .A2(n9466), .ZN(n25396) );
  NAND2_X1 U13422 ( .A1(n9443), .A2(n25396), .ZN(n9490) );
  AND2_X1 U13423 ( .A1(n9466), .A2(n9444), .ZN(n25473) );
  AOI22_X1 U13424 ( .A1(n23717), .A2(\xmem_data[96][5] ), .B1(n25398), .B2(
        \xmem_data[97][5] ), .ZN(n9448) );
  BUF_X1 U13425 ( .A(n14971), .Z(n25400) );
  BUF_X1 U13426 ( .A(n13452), .Z(n25399) );
  AOI22_X1 U13427 ( .A1(n25400), .A2(\xmem_data[98][5] ), .B1(n25399), .B2(
        \xmem_data[99][5] ), .ZN(n9447) );
  AOI22_X1 U13428 ( .A1(n3178), .A2(\xmem_data[100][5] ), .B1(n29281), .B2(
        \xmem_data[101][5] ), .ZN(n9446) );
  BUF_X1 U13429 ( .A(n14974), .Z(n25401) );
  AOI22_X1 U13430 ( .A1(n25401), .A2(\xmem_data[102][5] ), .B1(n14975), .B2(
        \xmem_data[103][5] ), .ZN(n9445) );
  NAND4_X1 U13431 ( .A1(n9448), .A2(n9447), .A3(n9446), .A4(n9445), .ZN(n9464)
         );
  BUF_X1 U13432 ( .A(n14919), .Z(n25406) );
  AOI22_X1 U13433 ( .A1(n29325), .A2(\xmem_data[104][5] ), .B1(n25406), .B2(
        \xmem_data[105][5] ), .ZN(n9452) );
  BUF_X1 U13434 ( .A(n13127), .Z(n25407) );
  AOI22_X1 U13435 ( .A1(n25407), .A2(\xmem_data[106][5] ), .B1(n27435), .B2(
        \xmem_data[107][5] ), .ZN(n9451) );
  BUF_X1 U13436 ( .A(n31263), .Z(n25408) );
  AOI22_X1 U13437 ( .A1(n25408), .A2(\xmem_data[108][5] ), .B1(n30571), .B2(
        \xmem_data[109][5] ), .ZN(n9450) );
  AOI22_X1 U13438 ( .A1(n3318), .A2(\xmem_data[110][5] ), .B1(n20711), .B2(
        \xmem_data[111][5] ), .ZN(n9449) );
  NAND4_X1 U13439 ( .A1(n9452), .A2(n9451), .A3(n9450), .A4(n9449), .ZN(n9463)
         );
  BUF_X1 U13440 ( .A(n29064), .Z(n25413) );
  AOI22_X1 U13441 ( .A1(n25413), .A2(\xmem_data[112][5] ), .B1(n3220), .B2(
        \xmem_data[113][5] ), .ZN(n9456) );
  BUF_X1 U13442 ( .A(n14988), .Z(n25414) );
  AOI22_X1 U13443 ( .A1(n25414), .A2(\xmem_data[114][5] ), .B1(n20787), .B2(
        \xmem_data[115][5] ), .ZN(n9455) );
  BUF_X1 U13444 ( .A(n14990), .Z(n25416) );
  BUF_X1 U13445 ( .A(n14890), .Z(n25415) );
  AOI22_X1 U13446 ( .A1(n25416), .A2(\xmem_data[116][5] ), .B1(n25415), .B2(
        \xmem_data[117][5] ), .ZN(n9454) );
  BUF_X1 U13447 ( .A(n14991), .Z(n25417) );
  AOI22_X1 U13448 ( .A1(n25417), .A2(\xmem_data[118][5] ), .B1(n25514), .B2(
        \xmem_data[119][5] ), .ZN(n9453) );
  NAND4_X1 U13449 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n9462)
         );
  AOI22_X1 U13450 ( .A1(n25422), .A2(\xmem_data[120][5] ), .B1(n24158), .B2(
        \xmem_data[121][5] ), .ZN(n9460) );
  BUF_X1 U13451 ( .A(n14997), .Z(n25424) );
  BUF_X1 U13452 ( .A(n14934), .Z(n25423) );
  AOI22_X1 U13453 ( .A1(n25424), .A2(\xmem_data[122][5] ), .B1(n25423), .B2(
        \xmem_data[123][5] ), .ZN(n9459) );
  AOI22_X1 U13454 ( .A1(n25425), .A2(\xmem_data[124][5] ), .B1(n22674), .B2(
        \xmem_data[125][5] ), .ZN(n9458) );
  AOI22_X1 U13455 ( .A1(n28336), .A2(\xmem_data[126][5] ), .B1(n27454), .B2(
        \xmem_data[127][5] ), .ZN(n9457) );
  NAND4_X1 U13456 ( .A1(n9460), .A2(n9459), .A3(n9458), .A4(n9457), .ZN(n9461)
         );
  OR4_X1 U13457 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9461), .ZN(n9488)
         );
  NOR2_X1 U13458 ( .A1(n9466), .A2(n9465), .ZN(n25471) );
  AOI22_X1 U13459 ( .A1(n25434), .A2(\xmem_data[64][5] ), .B1(n25398), .B2(
        \xmem_data[65][5] ), .ZN(n9470) );
  AOI22_X1 U13460 ( .A1(n24710), .A2(\xmem_data[66][5] ), .B1(n25435), .B2(
        \xmem_data[67][5] ), .ZN(n9469) );
  AOI22_X1 U13461 ( .A1(n28493), .A2(\xmem_data[68][5] ), .B1(n30898), .B2(
        \xmem_data[69][5] ), .ZN(n9468) );
  AOI22_X1 U13462 ( .A1(n3308), .A2(\xmem_data[70][5] ), .B1(n27975), .B2(
        \xmem_data[71][5] ), .ZN(n9467) );
  NAND4_X1 U13463 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n9486)
         );
  AOI22_X1 U13464 ( .A1(n3172), .A2(\xmem_data[72][5] ), .B1(n22751), .B2(
        \xmem_data[73][5] ), .ZN(n9474) );
  AOI22_X1 U13465 ( .A1(n28036), .A2(\xmem_data[74][5] ), .B1(n25440), .B2(
        \xmem_data[75][5] ), .ZN(n9473) );
  AOI22_X1 U13466 ( .A1(n25441), .A2(\xmem_data[76][5] ), .B1(n28366), .B2(
        \xmem_data[77][5] ), .ZN(n9472) );
  AOI22_X1 U13467 ( .A1(n25443), .A2(\xmem_data[78][5] ), .B1(n25442), .B2(
        \xmem_data[79][5] ), .ZN(n9471) );
  NAND4_X1 U13468 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n9485)
         );
  AOI22_X1 U13469 ( .A1(n28470), .A2(\xmem_data[80][5] ), .B1(n3220), .B2(
        \xmem_data[81][5] ), .ZN(n9478) );
  AOI22_X1 U13470 ( .A1(n25448), .A2(\xmem_data[82][5] ), .B1(n24695), .B2(
        \xmem_data[83][5] ), .ZN(n9477) );
  AOI22_X1 U13471 ( .A1(n25449), .A2(\xmem_data[84][5] ), .B1(n21068), .B2(
        \xmem_data[85][5] ), .ZN(n9476) );
  AOI22_X1 U13472 ( .A1(n25451), .A2(\xmem_data[86][5] ), .B1(n23771), .B2(
        \xmem_data[87][5] ), .ZN(n9475) );
  NAND4_X1 U13473 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(n9484)
         );
  AOI22_X1 U13474 ( .A1(n27447), .A2(\xmem_data[88][5] ), .B1(n28373), .B2(
        \xmem_data[89][5] ), .ZN(n9482) );
  AOI22_X1 U13475 ( .A1(n25457), .A2(\xmem_data[90][5] ), .B1(n24448), .B2(
        \xmem_data[91][5] ), .ZN(n9481) );
  AOI22_X1 U13476 ( .A1(n25459), .A2(\xmem_data[92][5] ), .B1(n25458), .B2(
        \xmem_data[93][5] ), .ZN(n9480) );
  AOI22_X1 U13477 ( .A1(n3466), .A2(\xmem_data[94][5] ), .B1(n25460), .B2(
        \xmem_data[95][5] ), .ZN(n9479) );
  NAND4_X1 U13478 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9483)
         );
  OR4_X1 U13479 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n9487)
         );
  AOI22_X1 U13480 ( .A1(n25473), .A2(n9488), .B1(n25471), .B2(n9487), .ZN(
        n9489) );
  XOR2_X1 U13481 ( .A(\fmem_data[30][5] ), .B(\fmem_data[30][4] ), .Z(n9492)
         );
  AOI22_X1 U13482 ( .A1(n25358), .A2(\xmem_data[12][6] ), .B1(n25357), .B2(
        \xmem_data[13][6] ), .ZN(n9506) );
  AOI22_X1 U13483 ( .A1(n3177), .A2(\xmem_data[4][6] ), .B1(n25364), .B2(
        \xmem_data[5][6] ), .ZN(n9493) );
  INV_X1 U13484 ( .A(n9493), .ZN(n9498) );
  AOI22_X1 U13485 ( .A1(n30893), .A2(\xmem_data[2][6] ), .B1(n25367), .B2(
        \xmem_data[3][6] ), .ZN(n9496) );
  AOI22_X1 U13486 ( .A1(n24509), .A2(\xmem_data[0][6] ), .B1(n14970), .B2(
        \xmem_data[1][6] ), .ZN(n9495) );
  AOI22_X1 U13487 ( .A1(n21056), .A2(\xmem_data[6][6] ), .B1(n20949), .B2(
        \xmem_data[7][6] ), .ZN(n9494) );
  NOR2_X1 U13488 ( .A1(n9498), .A2(n9497), .ZN(n9505) );
  AOI22_X1 U13489 ( .A1(n28467), .A2(\xmem_data[10][6] ), .B1(n25388), .B2(
        \xmem_data[11][6] ), .ZN(n9504) );
  AOI22_X1 U13490 ( .A1(n28293), .A2(\xmem_data[8][6] ), .B1(n25359), .B2(
        \xmem_data[9][6] ), .ZN(n9499) );
  INV_X1 U13491 ( .A(n9499), .ZN(n9502) );
  AOI22_X1 U13492 ( .A1(n3306), .A2(\xmem_data[14][6] ), .B1(n25360), .B2(
        \xmem_data[15][6] ), .ZN(n9500) );
  INV_X1 U13493 ( .A(n9500), .ZN(n9501) );
  NOR2_X1 U13494 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  NAND4_X1 U13495 ( .A1(n9506), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(n9519)
         );
  AOI22_X1 U13496 ( .A1(n28374), .A2(\xmem_data[24][6] ), .B1(n13475), .B2(
        \xmem_data[25][6] ), .ZN(n9510) );
  AOI22_X1 U13497 ( .A1(n30886), .A2(\xmem_data[26][6] ), .B1(n21075), .B2(
        \xmem_data[27][6] ), .ZN(n9509) );
  AOI22_X1 U13498 ( .A1(n30514), .A2(\xmem_data[28][6] ), .B1(n25382), .B2(
        \xmem_data[29][6] ), .ZN(n9508) );
  AOI22_X1 U13499 ( .A1(n31328), .A2(\xmem_data[30][6] ), .B1(n25383), .B2(
        \xmem_data[31][6] ), .ZN(n9507) );
  AOI22_X1 U13500 ( .A1(n25354), .A2(\xmem_data[16][6] ), .B1(n3220), .B2(
        \xmem_data[17][6] ), .ZN(n9517) );
  AOI22_X1 U13501 ( .A1(n24697), .A2(\xmem_data[20][6] ), .B1(n20559), .B2(
        \xmem_data[21][6] ), .ZN(n9511) );
  INV_X1 U13502 ( .A(n9511), .ZN(n9515) );
  AOI22_X1 U13503 ( .A1(n28733), .A2(\xmem_data[18][6] ), .B1(n28356), .B2(
        \xmem_data[19][6] ), .ZN(n9513) );
  NAND2_X1 U13504 ( .A1(n25377), .A2(\xmem_data[22][6] ), .ZN(n9512) );
  NAND2_X1 U13505 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  NOR2_X1 U13506 ( .A1(n9515), .A2(n9514), .ZN(n9516) );
  NAND3_X1 U13507 ( .A1(n3784), .A2(n9517), .A3(n9516), .ZN(n9518) );
  NOR2_X1 U13508 ( .A1(n9519), .A2(n9518), .ZN(n9521) );
  NAND2_X1 U13509 ( .A1(n25450), .A2(\xmem_data[23][6] ), .ZN(n9520) );
  INV_X1 U13510 ( .A(n16443), .ZN(n25392) );
  AOI21_X1 U13511 ( .B1(n9521), .B2(n9520), .A(n25392), .ZN(n9522) );
  INV_X1 U13512 ( .A(n9522), .ZN(n9588) );
  AOI22_X1 U13513 ( .A1(n17020), .A2(\xmem_data[96][6] ), .B1(n25398), .B2(
        \xmem_data[97][6] ), .ZN(n9526) );
  AOI22_X1 U13514 ( .A1(n25400), .A2(\xmem_data[98][6] ), .B1(n25399), .B2(
        \xmem_data[99][6] ), .ZN(n9525) );
  AOI22_X1 U13515 ( .A1(n3177), .A2(\xmem_data[100][6] ), .B1(n30598), .B2(
        \xmem_data[101][6] ), .ZN(n9524) );
  AOI22_X1 U13516 ( .A1(n25401), .A2(\xmem_data[102][6] ), .B1(n14975), .B2(
        \xmem_data[103][6] ), .ZN(n9523) );
  NAND4_X1 U13517 ( .A1(n9526), .A2(n9525), .A3(n9524), .A4(n9523), .ZN(n9542)
         );
  AOI22_X1 U13518 ( .A1(n29325), .A2(\xmem_data[104][6] ), .B1(n25406), .B2(
        \xmem_data[105][6] ), .ZN(n9530) );
  AOI22_X1 U13519 ( .A1(n25407), .A2(\xmem_data[106][6] ), .B1(n20579), .B2(
        \xmem_data[107][6] ), .ZN(n9529) );
  AOI22_X1 U13520 ( .A1(n25408), .A2(\xmem_data[108][6] ), .B1(n3203), .B2(
        \xmem_data[109][6] ), .ZN(n9528) );
  AOI22_X1 U13521 ( .A1(n3318), .A2(\xmem_data[110][6] ), .B1(n29173), .B2(
        \xmem_data[111][6] ), .ZN(n9527) );
  NAND4_X1 U13522 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n9541)
         );
  AOI22_X1 U13523 ( .A1(n25413), .A2(\xmem_data[112][6] ), .B1(n3222), .B2(
        \xmem_data[113][6] ), .ZN(n9534) );
  AOI22_X1 U13524 ( .A1(n25414), .A2(\xmem_data[114][6] ), .B1(n23739), .B2(
        \xmem_data[115][6] ), .ZN(n9533) );
  AOI22_X1 U13525 ( .A1(n25416), .A2(\xmem_data[116][6] ), .B1(n25415), .B2(
        \xmem_data[117][6] ), .ZN(n9532) );
  AOI22_X1 U13526 ( .A1(n25417), .A2(\xmem_data[118][6] ), .B1(n25492), .B2(
        \xmem_data[119][6] ), .ZN(n9531) );
  NAND4_X1 U13527 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n9540)
         );
  AOI22_X1 U13528 ( .A1(n25422), .A2(\xmem_data[120][6] ), .B1(n13475), .B2(
        \xmem_data[121][6] ), .ZN(n9538) );
  AOI22_X1 U13529 ( .A1(n25424), .A2(\xmem_data[122][6] ), .B1(n25423), .B2(
        \xmem_data[123][6] ), .ZN(n9537) );
  AOI22_X1 U13530 ( .A1(n25425), .A2(\xmem_data[124][6] ), .B1(n25671), .B2(
        \xmem_data[125][6] ), .ZN(n9536) );
  AOI22_X1 U13531 ( .A1(n29605), .A2(\xmem_data[126][6] ), .B1(n25460), .B2(
        \xmem_data[127][6] ), .ZN(n9535) );
  NAND4_X1 U13532 ( .A1(n9538), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(n9539)
         );
  OR4_X1 U13533 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(n9564)
         );
  AOI22_X1 U13534 ( .A1(n25434), .A2(\xmem_data[64][6] ), .B1(n23796), .B2(
        \xmem_data[65][6] ), .ZN(n9546) );
  AOI22_X1 U13535 ( .A1(n22717), .A2(n20682), .B1(n25435), .B2(
        \xmem_data[67][6] ), .ZN(n9545) );
  AOI22_X1 U13536 ( .A1(n28428), .A2(\xmem_data[68][6] ), .B1(n30955), .B2(
        \xmem_data[69][6] ), .ZN(n9544) );
  AOI22_X1 U13537 ( .A1(n3308), .A2(\xmem_data[70][6] ), .B1(n28098), .B2(
        \xmem_data[71][6] ), .ZN(n9543) );
  NAND4_X1 U13538 ( .A1(n9546), .A2(n9545), .A3(n9544), .A4(n9543), .ZN(n9562)
         );
  AOI22_X1 U13539 ( .A1(n24685), .A2(\xmem_data[72][6] ), .B1(n31256), .B2(
        \xmem_data[73][6] ), .ZN(n9550) );
  AOI22_X1 U13540 ( .A1(n29725), .A2(\xmem_data[74][6] ), .B1(n25440), .B2(
        \xmem_data[75][6] ), .ZN(n9549) );
  AOI22_X1 U13541 ( .A1(n25441), .A2(\xmem_data[76][6] ), .B1(n24525), .B2(
        \xmem_data[77][6] ), .ZN(n9548) );
  AOI22_X1 U13542 ( .A1(n25443), .A2(\xmem_data[78][6] ), .B1(n25442), .B2(
        \xmem_data[79][6] ), .ZN(n9547) );
  NAND4_X1 U13543 ( .A1(n9550), .A2(n9549), .A3(n9548), .A4(n9547), .ZN(n9561)
         );
  AOI22_X1 U13544 ( .A1(n31348), .A2(\xmem_data[80][6] ), .B1(n3220), .B2(
        \xmem_data[81][6] ), .ZN(n9554) );
  AOI22_X1 U13545 ( .A1(n25448), .A2(\xmem_data[82][6] ), .B1(n20500), .B2(
        \xmem_data[83][6] ), .ZN(n9553) );
  AOI22_X1 U13546 ( .A1(n25449), .A2(\xmem_data[84][6] ), .B1(n31275), .B2(
        \xmem_data[85][6] ), .ZN(n9552) );
  AOI22_X1 U13547 ( .A1(n25451), .A2(\xmem_data[86][6] ), .B1(n3231), .B2(
        \xmem_data[87][6] ), .ZN(n9551) );
  NAND4_X1 U13548 ( .A1(n9554), .A2(n9553), .A3(n9552), .A4(n9551), .ZN(n9560)
         );
  AOI22_X1 U13549 ( .A1(n31321), .A2(\xmem_data[88][6] ), .B1(n3358), .B2(
        \xmem_data[89][6] ), .ZN(n9558) );
  AOI22_X1 U13550 ( .A1(n25457), .A2(\xmem_data[90][6] ), .B1(n14998), .B2(
        \xmem_data[91][6] ), .ZN(n9557) );
  AOI22_X1 U13551 ( .A1(n25459), .A2(\xmem_data[92][6] ), .B1(n25458), .B2(
        \xmem_data[93][6] ), .ZN(n9556) );
  AOI22_X1 U13552 ( .A1(n3466), .A2(\xmem_data[94][6] ), .B1(n25460), .B2(
        \xmem_data[95][6] ), .ZN(n9555) );
  NAND4_X1 U13553 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9559)
         );
  OR4_X1 U13554 ( .A1(n9562), .A2(n9561), .A3(n9560), .A4(n9559), .ZN(n9563)
         );
  AOI22_X1 U13555 ( .A1(n25473), .A2(n9564), .B1(n25471), .B2(n9563), .ZN(
        n9587) );
  AOI22_X1 U13556 ( .A1(n25434), .A2(\xmem_data[32][6] ), .B1(n28492), .B2(
        \xmem_data[33][6] ), .ZN(n9568) );
  AOI22_X1 U13557 ( .A1(n17021), .A2(\xmem_data[34][6] ), .B1(n25435), .B2(
        \xmem_data[35][6] ), .ZN(n9567) );
  AOI22_X1 U13558 ( .A1(n28428), .A2(\xmem_data[36][6] ), .B1(n17001), .B2(
        \xmem_data[37][6] ), .ZN(n9566) );
  AOI22_X1 U13559 ( .A1(n3308), .A2(\xmem_data[38][6] ), .B1(n24223), .B2(
        \xmem_data[39][6] ), .ZN(n9565) );
  NAND4_X1 U13560 ( .A1(n9568), .A2(n9567), .A3(n9566), .A4(n9565), .ZN(n9584)
         );
  AOI22_X1 U13561 ( .A1(n3172), .A2(\xmem_data[40][6] ), .B1(n27526), .B2(
        \xmem_data[41][6] ), .ZN(n9572) );
  AOI22_X1 U13562 ( .A1(n28241), .A2(\xmem_data[42][6] ), .B1(n25440), .B2(
        \xmem_data[43][6] ), .ZN(n9571) );
  AOI22_X1 U13563 ( .A1(n25441), .A2(\xmem_data[44][6] ), .B1(n28075), .B2(
        \xmem_data[45][6] ), .ZN(n9570) );
  AOI22_X1 U13564 ( .A1(n25443), .A2(\xmem_data[46][6] ), .B1(n25442), .B2(
        \xmem_data[47][6] ), .ZN(n9569) );
  NAND4_X1 U13565 ( .A1(n9572), .A2(n9571), .A3(n9570), .A4(n9569), .ZN(n9583)
         );
  AOI22_X1 U13566 ( .A1(n28318), .A2(\xmem_data[48][6] ), .B1(n3220), .B2(
        \xmem_data[49][6] ), .ZN(n9576) );
  AOI22_X1 U13567 ( .A1(n25448), .A2(\xmem_data[50][6] ), .B1(n28319), .B2(
        \xmem_data[51][6] ), .ZN(n9575) );
  AOI22_X1 U13568 ( .A1(n25449), .A2(\xmem_data[52][6] ), .B1(n3255), .B2(
        \xmem_data[53][6] ), .ZN(n9574) );
  AOI22_X1 U13569 ( .A1(n25451), .A2(\xmem_data[54][6] ), .B1(n3231), .B2(
        \xmem_data[55][6] ), .ZN(n9573) );
  NAND4_X1 U13570 ( .A1(n9576), .A2(n9575), .A3(n9574), .A4(n9573), .ZN(n9582)
         );
  AOI22_X1 U13571 ( .A1(n24554), .A2(\xmem_data[56][6] ), .B1(n20546), .B2(
        \xmem_data[57][6] ), .ZN(n9580) );
  AOI22_X1 U13572 ( .A1(n25457), .A2(\xmem_data[58][6] ), .B1(n24555), .B2(
        \xmem_data[59][6] ), .ZN(n9579) );
  AOI22_X1 U13573 ( .A1(n25459), .A2(\xmem_data[60][6] ), .B1(n25458), .B2(
        \xmem_data[61][6] ), .ZN(n9578) );
  AOI22_X1 U13574 ( .A1(n30303), .A2(\xmem_data[62][6] ), .B1(n25460), .B2(
        \xmem_data[63][6] ), .ZN(n9577) );
  NAND4_X1 U13575 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n9581)
         );
  OR4_X1 U13576 ( .A1(n9584), .A2(n9583), .A3(n9582), .A4(n9581), .ZN(n9585)
         );
  NAND2_X1 U13577 ( .A1(n9585), .A2(n25396), .ZN(n9586) );
  XNOR2_X1 U13578 ( .A(n31659), .B(\fmem_data[30][5] ), .ZN(n33104) );
  OAI22_X1 U13579 ( .A1(n30420), .A2(n33103), .B1(n33104), .B2(n33105), .ZN(
        n23597) );
  AOI22_X1 U13580 ( .A1(n20730), .A2(\xmem_data[96][5] ), .B1(n24510), .B2(
        \xmem_data[97][5] ), .ZN(n9592) );
  AOI22_X1 U13581 ( .A1(n20731), .A2(\xmem_data[98][5] ), .B1(n29281), .B2(
        \xmem_data[99][5] ), .ZN(n9591) );
  AOI22_X1 U13582 ( .A1(n20732), .A2(\xmem_data[100][5] ), .B1(n30599), .B2(
        \xmem_data[101][5] ), .ZN(n9590) );
  AOI22_X1 U13583 ( .A1(n20734), .A2(\xmem_data[102][5] ), .B1(n20733), .B2(
        \xmem_data[103][5] ), .ZN(n9589) );
  NAND4_X1 U13584 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n9608)
         );
  AOI22_X1 U13585 ( .A1(n20708), .A2(\xmem_data[104][5] ), .B1(n20707), .B2(
        \xmem_data[105][5] ), .ZN(n9596) );
  AOI22_X1 U13586 ( .A1(n20710), .A2(\xmem_data[106][5] ), .B1(n20709), .B2(
        \xmem_data[107][5] ), .ZN(n9595) );
  AOI22_X1 U13587 ( .A1(n3305), .A2(\xmem_data[108][5] ), .B1(n20711), .B2(
        \xmem_data[109][5] ), .ZN(n9594) );
  AOI22_X1 U13588 ( .A1(n29254), .A2(\xmem_data[110][5] ), .B1(n3220), .B2(
        \xmem_data[111][5] ), .ZN(n9593) );
  NAND4_X1 U13589 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9607)
         );
  AOI22_X1 U13590 ( .A1(n20724), .A2(\xmem_data[112][5] ), .B1(n20723), .B2(
        \xmem_data[113][5] ), .ZN(n9600) );
  AOI22_X1 U13591 ( .A1(n20725), .A2(\xmem_data[114][5] ), .B1(n3256), .B2(
        \xmem_data[115][5] ), .ZN(n9599) );
  AOI22_X1 U13592 ( .A1(n3344), .A2(\xmem_data[116][5] ), .B1(n25514), .B2(
        \xmem_data[117][5] ), .ZN(n9598) );
  AOI22_X1 U13593 ( .A1(n28050), .A2(\xmem_data[118][5] ), .B1(n27863), .B2(
        \xmem_data[119][5] ), .ZN(n9597) );
  NAND4_X1 U13594 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9606)
         );
  AOI22_X1 U13595 ( .A1(n20716), .A2(\xmem_data[120][5] ), .B1(n27535), .B2(
        \xmem_data[121][5] ), .ZN(n9604) );
  AOI22_X1 U13596 ( .A1(n25567), .A2(\xmem_data[122][5] ), .B1(n20717), .B2(
        \xmem_data[123][5] ), .ZN(n9603) );
  AOI22_X1 U13597 ( .A1(n27455), .A2(\xmem_data[124][5] ), .B1(n29188), .B2(
        \xmem_data[125][5] ), .ZN(n9602) );
  AOI22_X1 U13598 ( .A1(n24547), .A2(\xmem_data[126][5] ), .B1(n27518), .B2(
        \xmem_data[127][5] ), .ZN(n9601) );
  NAND4_X1 U13599 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n9605)
         );
  OR4_X1 U13600 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9631)
         );
  AOI22_X1 U13601 ( .A1(n20826), .A2(\xmem_data[72][5] ), .B1(n20769), .B2(
        \xmem_data[73][5] ), .ZN(n9613) );
  AOI22_X1 U13602 ( .A1(n20827), .A2(\xmem_data[74][5] ), .B1(n25685), .B2(
        \xmem_data[75][5] ), .ZN(n9612) );
  AOI22_X1 U13603 ( .A1(n20828), .A2(\xmem_data[76][5] ), .B1(n30589), .B2(
        \xmem_data[77][5] ), .ZN(n9611) );
  AND2_X1 U13604 ( .A1(n3222), .A2(\xmem_data[79][5] ), .ZN(n9609) );
  AOI21_X1 U13605 ( .B1(n24443), .B2(\xmem_data[78][5] ), .A(n9609), .ZN(n9610) );
  NAND4_X1 U13606 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), .ZN(n9629)
         );
  AOI22_X1 U13607 ( .A1(n20799), .A2(\xmem_data[88][5] ), .B1(n25605), .B2(
        \xmem_data[89][5] ), .ZN(n9617) );
  AOI22_X1 U13608 ( .A1(n25425), .A2(\xmem_data[90][5] ), .B1(n20798), .B2(
        \xmem_data[91][5] ), .ZN(n9616) );
  AOI22_X1 U13609 ( .A1(n28231), .A2(\xmem_data[92][5] ), .B1(n24134), .B2(
        \xmem_data[93][5] ), .ZN(n9615) );
  AOI22_X1 U13610 ( .A1(n20800), .A2(\xmem_data[94][5] ), .B1(n25398), .B2(
        \xmem_data[95][5] ), .ZN(n9614) );
  NAND4_X1 U13611 ( .A1(n9617), .A2(n9616), .A3(n9615), .A4(n9614), .ZN(n9628)
         );
  AOI22_X1 U13612 ( .A1(n20805), .A2(\xmem_data[80][5] ), .B1(n20598), .B2(
        \xmem_data[81][5] ), .ZN(n9621) );
  AOI22_X1 U13613 ( .A1(n20807), .A2(\xmem_data[82][5] ), .B1(n20806), .B2(
        \xmem_data[83][5] ), .ZN(n9620) );
  AOI22_X1 U13614 ( .A1(n20808), .A2(\xmem_data[84][5] ), .B1(n15011), .B2(
        \xmem_data[85][5] ), .ZN(n9619) );
  AOI22_X1 U13615 ( .A1(n20809), .A2(\xmem_data[86][5] ), .B1(n3357), .B2(
        \xmem_data[87][5] ), .ZN(n9618) );
  NAND4_X1 U13616 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n9627)
         );
  AOI22_X1 U13617 ( .A1(n20815), .A2(\xmem_data[64][5] ), .B1(n20814), .B2(
        \xmem_data[65][5] ), .ZN(n9625) );
  AOI22_X1 U13618 ( .A1(n28385), .A2(\xmem_data[66][5] ), .B1(n28327), .B2(
        \xmem_data[67][5] ), .ZN(n9624) );
  AOI22_X1 U13619 ( .A1(n20817), .A2(\xmem_data[68][5] ), .B1(n28098), .B2(
        \xmem_data[69][5] ), .ZN(n9623) );
  AOI22_X1 U13620 ( .A1(n20818), .A2(\xmem_data[70][5] ), .B1(n27526), .B2(
        \xmem_data[71][5] ), .ZN(n9622) );
  NAND4_X1 U13621 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), .ZN(n9626)
         );
  OR4_X1 U13622 ( .A1(n9629), .A2(n9628), .A3(n9627), .A4(n9626), .ZN(n9630)
         );
  AOI22_X1 U13623 ( .A1(n9631), .A2(n20742), .B1(n20833), .B2(n9630), .ZN(
        n9685) );
  AOI22_X1 U13624 ( .A1(n27708), .A2(\xmem_data[16][5] ), .B1(n20787), .B2(
        \xmem_data[17][5] ), .ZN(n9638) );
  AOI22_X1 U13625 ( .A1(n3322), .A2(\xmem_data[18][5] ), .B1(n21068), .B2(
        \xmem_data[19][5] ), .ZN(n9632) );
  INV_X1 U13626 ( .A(n9632), .ZN(n9636) );
  AOI22_X1 U13627 ( .A1(n25422), .A2(\xmem_data[22][5] ), .B1(n3358), .B2(
        \xmem_data[23][5] ), .ZN(n9634) );
  NAND2_X1 U13628 ( .A1(n17063), .A2(\xmem_data[20][5] ), .ZN(n9633) );
  NAND2_X1 U13629 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  NOR2_X1 U13630 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NAND2_X1 U13631 ( .A1(n9638), .A2(n9637), .ZN(n9644) );
  AOI22_X1 U13632 ( .A1(n30744), .A2(\xmem_data[24][5] ), .B1(n20775), .B2(
        \xmem_data[25][5] ), .ZN(n9642) );
  AOI22_X1 U13633 ( .A1(n27537), .A2(\xmem_data[26][5] ), .B1(n20717), .B2(
        \xmem_data[27][5] ), .ZN(n9641) );
  AOI22_X1 U13634 ( .A1(n3158), .A2(\xmem_data[28][5] ), .B1(n27864), .B2(
        \xmem_data[29][5] ), .ZN(n9640) );
  AOI22_X1 U13635 ( .A1(n23717), .A2(\xmem_data[30][5] ), .B1(n28427), .B2(
        \xmem_data[31][5] ), .ZN(n9639) );
  NAND4_X1 U13636 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(n9643)
         );
  OR2_X1 U13637 ( .A1(n9644), .A2(n9643), .ZN(n9659) );
  AOI22_X1 U13638 ( .A1(n3317), .A2(\xmem_data[12][5] ), .B1(n20711), .B2(
        \xmem_data[13][5] ), .ZN(n9645) );
  INV_X1 U13639 ( .A(n9645), .ZN(n9653) );
  AOI22_X1 U13640 ( .A1(n20782), .A2(\xmem_data[6][5] ), .B1(n28328), .B2(
        \xmem_data[7][5] ), .ZN(n9647) );
  AOI22_X1 U13641 ( .A1(n3300), .A2(\xmem_data[4][5] ), .B1(n20781), .B2(
        \xmem_data[5][5] ), .ZN(n9646) );
  NAND2_X1 U13642 ( .A1(n9647), .A2(n9646), .ZN(n9652) );
  AOI22_X1 U13643 ( .A1(n20731), .A2(\xmem_data[2][5] ), .B1(n28327), .B2(
        \xmem_data[3][5] ), .ZN(n9648) );
  INV_X1 U13644 ( .A(n9648), .ZN(n9651) );
  AOI22_X1 U13645 ( .A1(n21008), .A2(\xmem_data[0][5] ), .B1(n27523), .B2(
        \xmem_data[1][5] ), .ZN(n9649) );
  INV_X1 U13646 ( .A(n9649), .ZN(n9650) );
  NOR4_X1 U13647 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n9657)
         );
  AOI22_X1 U13648 ( .A1(n30592), .A2(\xmem_data[14][5] ), .B1(n3219), .B2(
        \xmem_data[15][5] ), .ZN(n9656) );
  AOI22_X1 U13649 ( .A1(n20770), .A2(\xmem_data[8][5] ), .B1(n20769), .B2(
        \xmem_data[9][5] ), .ZN(n9655) );
  AOI22_X1 U13650 ( .A1(n30862), .A2(\xmem_data[10][5] ), .B1(n29118), .B2(
        \xmem_data[11][5] ), .ZN(n9654) );
  NAND4_X1 U13651 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9658)
         );
  NOR2_X1 U13652 ( .A1(n9659), .A2(n9658), .ZN(n9660) );
  AOI22_X1 U13653 ( .A1(n20815), .A2(\xmem_data[32][5] ), .B1(n20814), .B2(
        \xmem_data[33][5] ), .ZN(n9664) );
  AOI22_X1 U13654 ( .A1(n27974), .A2(\xmem_data[34][5] ), .B1(n29281), .B2(
        \xmem_data[35][5] ), .ZN(n9663) );
  AOI22_X1 U13655 ( .A1(n20817), .A2(\xmem_data[36][5] ), .B1(n25583), .B2(
        \xmem_data[37][5] ), .ZN(n9662) );
  AOI22_X1 U13656 ( .A1(n20818), .A2(\xmem_data[38][5] ), .B1(n27981), .B2(
        \xmem_data[39][5] ), .ZN(n9661) );
  NAND4_X1 U13657 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9680)
         );
  AOI22_X1 U13658 ( .A1(n20826), .A2(\xmem_data[40][5] ), .B1(n24686), .B2(
        \xmem_data[41][5] ), .ZN(n9668) );
  AOI22_X1 U13659 ( .A1(n20827), .A2(\xmem_data[42][5] ), .B1(n21309), .B2(
        \xmem_data[43][5] ), .ZN(n9667) );
  AOI22_X1 U13660 ( .A1(n20828), .A2(\xmem_data[44][5] ), .B1(n27437), .B2(
        \xmem_data[45][5] ), .ZN(n9666) );
  AOI22_X1 U13661 ( .A1(n24694), .A2(\xmem_data[46][5] ), .B1(n3217), .B2(
        \xmem_data[47][5] ), .ZN(n9665) );
  NAND4_X1 U13662 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n9679)
         );
  AOI22_X1 U13663 ( .A1(n20805), .A2(\xmem_data[48][5] ), .B1(n20500), .B2(
        \xmem_data[49][5] ), .ZN(n9672) );
  AOI22_X1 U13664 ( .A1(n20807), .A2(\xmem_data[50][5] ), .B1(n20806), .B2(
        \xmem_data[51][5] ), .ZN(n9671) );
  AOI22_X1 U13665 ( .A1(n20808), .A2(\xmem_data[52][5] ), .B1(n27547), .B2(
        \xmem_data[53][5] ), .ZN(n9670) );
  AOI22_X1 U13666 ( .A1(n20809), .A2(\xmem_data[54][5] ), .B1(n3358), .B2(
        \xmem_data[55][5] ), .ZN(n9669) );
  NAND4_X1 U13667 ( .A1(n9672), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n9678)
         );
  AOI22_X1 U13668 ( .A1(n20799), .A2(\xmem_data[56][5] ), .B1(n28375), .B2(
        \xmem_data[57][5] ), .ZN(n9676) );
  AOI22_X1 U13669 ( .A1(n3175), .A2(\xmem_data[58][5] ), .B1(n20798), .B2(
        \xmem_data[59][5] ), .ZN(n9675) );
  AOI22_X1 U13670 ( .A1(n30948), .A2(\xmem_data[60][5] ), .B1(n29188), .B2(
        \xmem_data[61][5] ), .ZN(n9674) );
  AOI22_X1 U13671 ( .A1(n20800), .A2(\xmem_data[62][5] ), .B1(n27918), .B2(
        \xmem_data[63][5] ), .ZN(n9673) );
  NAND4_X1 U13672 ( .A1(n9676), .A2(n9675), .A3(n9674), .A4(n9673), .ZN(n9677)
         );
  OR4_X1 U13673 ( .A1(n9680), .A2(n9679), .A3(n9678), .A4(n9677), .ZN(n9682)
         );
  NOR2_X1 U13674 ( .A1(n20188), .A2(n39004), .ZN(n9681) );
  AOI21_X1 U13675 ( .B1(n9682), .B2(n20765), .A(n3895), .ZN(n9683) );
  XNOR2_X1 U13676 ( .A(n31656), .B(\fmem_data[28][5] ), .ZN(n30157) );
  XOR2_X1 U13677 ( .A(\fmem_data[28][4] ), .B(\fmem_data[28][5] ), .Z(n9686)
         );
  AOI22_X1 U13678 ( .A1(n29439), .A2(\xmem_data[0][6] ), .B1(n27920), .B2(
        \xmem_data[1][6] ), .ZN(n9690) );
  AOI22_X1 U13679 ( .A1(n30899), .A2(\xmem_data[2][6] ), .B1(n21009), .B2(
        \xmem_data[3][6] ), .ZN(n9689) );
  AOI22_X1 U13680 ( .A1(n28226), .A2(\xmem_data[4][6] ), .B1(n20781), .B2(
        \xmem_data[5][6] ), .ZN(n9688) );
  AOI22_X1 U13681 ( .A1(n20782), .A2(\xmem_data[6][6] ), .B1(n14981), .B2(
        \xmem_data[7][6] ), .ZN(n9687) );
  NAND4_X1 U13682 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n9706)
         );
  AOI22_X1 U13683 ( .A1(n20770), .A2(\xmem_data[8][6] ), .B1(n20769), .B2(
        \xmem_data[9][6] ), .ZN(n9694) );
  AOI22_X1 U13684 ( .A1(n17030), .A2(\xmem_data[10][6] ), .B1(n29118), .B2(
        \xmem_data[11][6] ), .ZN(n9693) );
  AOI22_X1 U13685 ( .A1(n3352), .A2(\xmem_data[12][6] ), .B1(n28501), .B2(
        \xmem_data[13][6] ), .ZN(n9692) );
  AOI22_X1 U13686 ( .A1(n28503), .A2(\xmem_data[14][6] ), .B1(n3217), .B2(
        \xmem_data[15][6] ), .ZN(n9691) );
  NAND4_X1 U13687 ( .A1(n9694), .A2(n9693), .A3(n9692), .A4(n9691), .ZN(n9705)
         );
  AOI22_X1 U13688 ( .A1(n29494), .A2(\xmem_data[16][6] ), .B1(n20787), .B2(
        \xmem_data[17][6] ), .ZN(n9698) );
  AOI22_X1 U13689 ( .A1(n20725), .A2(\xmem_data[18][6] ), .B1(n23811), .B2(
        \xmem_data[19][6] ), .ZN(n9697) );
  AOI22_X1 U13690 ( .A1(n30710), .A2(\xmem_data[20][6] ), .B1(n24657), .B2(
        \xmem_data[21][6] ), .ZN(n9696) );
  AOI22_X1 U13691 ( .A1(n25707), .A2(\xmem_data[22][6] ), .B1(n28373), .B2(
        \xmem_data[23][6] ), .ZN(n9695) );
  NAND4_X1 U13692 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9704)
         );
  AOI22_X1 U13693 ( .A1(n27763), .A2(\xmem_data[24][6] ), .B1(n20775), .B2(
        \xmem_data[25][6] ), .ZN(n9702) );
  AOI22_X1 U13694 ( .A1(n31268), .A2(\xmem_data[26][6] ), .B1(n21076), .B2(
        \xmem_data[27][6] ), .ZN(n9701) );
  AOI22_X1 U13695 ( .A1(n31328), .A2(\xmem_data[28][6] ), .B1(n23716), .B2(
        \xmem_data[29][6] ), .ZN(n9700) );
  AOI22_X1 U13696 ( .A1(n28059), .A2(\xmem_data[30][6] ), .B1(n31329), .B2(
        \xmem_data[31][6] ), .ZN(n9699) );
  NAND4_X1 U13697 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n9703)
         );
  OR4_X1 U13698 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n9707)
         );
  AOI22_X1 U13699 ( .A1(n20799), .A2(\xmem_data[88][6] ), .B1(n23761), .B2(
        \xmem_data[89][6] ), .ZN(n9711) );
  AOI22_X1 U13700 ( .A1(n3176), .A2(\xmem_data[90][6] ), .B1(n20798), .B2(
        \xmem_data[91][6] ), .ZN(n9710) );
  AOI22_X1 U13701 ( .A1(n30303), .A2(\xmem_data[92][6] ), .B1(n25460), .B2(
        \xmem_data[93][6] ), .ZN(n9709) );
  AOI22_X1 U13702 ( .A1(n20800), .A2(\xmem_data[94][6] ), .B1(n21006), .B2(
        \xmem_data[95][6] ), .ZN(n9708) );
  NAND4_X1 U13703 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n9722)
         );
  AOI22_X1 U13704 ( .A1(n20805), .A2(\xmem_data[80][6] ), .B1(n27507), .B2(
        \xmem_data[81][6] ), .ZN(n9715) );
  AOI22_X1 U13705 ( .A1(n20807), .A2(\xmem_data[82][6] ), .B1(n20806), .B2(
        \xmem_data[83][6] ), .ZN(n9714) );
  AOI22_X1 U13706 ( .A1(n20808), .A2(\xmem_data[84][6] ), .B1(n3231), .B2(
        \xmem_data[85][6] ), .ZN(n9713) );
  AOI22_X1 U13707 ( .A1(n20809), .A2(\xmem_data[86][6] ), .B1(n20982), .B2(
        \xmem_data[87][6] ), .ZN(n9712) );
  NAND4_X1 U13708 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n9721)
         );
  AOI22_X1 U13709 ( .A1(n20815), .A2(\xmem_data[64][6] ), .B1(n20814), .B2(
        \xmem_data[65][6] ), .ZN(n9719) );
  AOI22_X1 U13710 ( .A1(n28428), .A2(n20682), .B1(n27856), .B2(
        \xmem_data[67][6] ), .ZN(n9718) );
  AOI22_X1 U13711 ( .A1(n20817), .A2(\xmem_data[68][6] ), .B1(n27365), .B2(
        \xmem_data[69][6] ), .ZN(n9717) );
  AOI22_X1 U13712 ( .A1(n20818), .A2(\xmem_data[70][6] ), .B1(n25406), .B2(
        \xmem_data[71][6] ), .ZN(n9716) );
  NAND4_X1 U13713 ( .A1(n9719), .A2(n9718), .A3(n9717), .A4(n9716), .ZN(n9720)
         );
  OR3_X1 U13714 ( .A1(n9722), .A2(n9721), .A3(n9720), .ZN(n9728) );
  AOI22_X1 U13715 ( .A1(n20826), .A2(\xmem_data[72][6] ), .B1(n25528), .B2(
        \xmem_data[73][6] ), .ZN(n9726) );
  AOI22_X1 U13716 ( .A1(n20827), .A2(\xmem_data[74][6] ), .B1(n31346), .B2(
        \xmem_data[75][6] ), .ZN(n9725) );
  AOI22_X1 U13717 ( .A1(n20828), .A2(\xmem_data[76][6] ), .B1(n29286), .B2(
        \xmem_data[77][6] ), .ZN(n9724) );
  AOI22_X1 U13718 ( .A1(n25692), .A2(\xmem_data[78][6] ), .B1(n3217), .B2(
        \xmem_data[79][6] ), .ZN(n9723) );
  NAND4_X1 U13719 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n9727)
         );
  OAI21_X1 U13720 ( .B1(n9728), .B2(n9727), .A(n20833), .ZN(n9773) );
  AOI22_X1 U13721 ( .A1(n20716), .A2(\xmem_data[120][6] ), .B1(n21015), .B2(
        \xmem_data[121][6] ), .ZN(n9732) );
  AOI22_X1 U13722 ( .A1(n16986), .A2(\xmem_data[122][6] ), .B1(n20717), .B2(
        \xmem_data[123][6] ), .ZN(n9731) );
  AOI22_X1 U13723 ( .A1(n24213), .A2(\xmem_data[124][6] ), .B1(n29162), .B2(
        \xmem_data[125][6] ), .ZN(n9730) );
  AOI22_X1 U13724 ( .A1(n24593), .A2(\xmem_data[126][6] ), .B1(n24546), .B2(
        \xmem_data[127][6] ), .ZN(n9729) );
  NAND4_X1 U13725 ( .A1(n9732), .A2(n9731), .A3(n9730), .A4(n9729), .ZN(n9743)
         );
  AOI22_X1 U13726 ( .A1(n20724), .A2(\xmem_data[112][6] ), .B1(n20723), .B2(
        \xmem_data[113][6] ), .ZN(n9736) );
  AOI22_X1 U13727 ( .A1(n20725), .A2(\xmem_data[114][6] ), .B1(n20806), .B2(
        \xmem_data[115][6] ), .ZN(n9735) );
  AOI22_X1 U13728 ( .A1(n23742), .A2(\xmem_data[116][6] ), .B1(n27446), .B2(
        \xmem_data[117][6] ), .ZN(n9734) );
  AOI22_X1 U13729 ( .A1(n23813), .A2(\xmem_data[118][6] ), .B1(n13475), .B2(
        \xmem_data[119][6] ), .ZN(n9733) );
  NAND4_X1 U13730 ( .A1(n9736), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(n9742)
         );
  AOI22_X1 U13731 ( .A1(n20730), .A2(\xmem_data[96][6] ), .B1(n25435), .B2(
        \xmem_data[97][6] ), .ZN(n9740) );
  AOI22_X1 U13732 ( .A1(n20731), .A2(\xmem_data[98][6] ), .B1(n25679), .B2(
        \xmem_data[99][6] ), .ZN(n9739) );
  AOI22_X1 U13733 ( .A1(n20732), .A2(\xmem_data[100][6] ), .B1(n20949), .B2(
        \xmem_data[101][6] ), .ZN(n9738) );
  AOI22_X1 U13734 ( .A1(n20734), .A2(\xmem_data[102][6] ), .B1(n20733), .B2(
        \xmem_data[103][6] ), .ZN(n9737) );
  NAND4_X1 U13735 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n9741)
         );
  OR3_X1 U13736 ( .A1(n9743), .A2(n9742), .A3(n9741), .ZN(n9749) );
  AOI22_X1 U13737 ( .A1(n20708), .A2(\xmem_data[104][6] ), .B1(n20707), .B2(
        \xmem_data[105][6] ), .ZN(n9747) );
  AOI22_X1 U13738 ( .A1(n20710), .A2(\xmem_data[106][6] ), .B1(n20709), .B2(
        \xmem_data[107][6] ), .ZN(n9746) );
  AOI22_X1 U13739 ( .A1(n3228), .A2(\xmem_data[108][6] ), .B1(n20711), .B2(
        \xmem_data[109][6] ), .ZN(n9745) );
  AOI22_X1 U13740 ( .A1(n27502), .A2(\xmem_data[110][6] ), .B1(n3218), .B2(
        \xmem_data[111][6] ), .ZN(n9744) );
  NAND4_X1 U13741 ( .A1(n9747), .A2(n9746), .A3(n9745), .A4(n9744), .ZN(n9748)
         );
  OAI21_X1 U13742 ( .B1(n9749), .B2(n9748), .A(n20742), .ZN(n9772) );
  AOI22_X1 U13743 ( .A1(n20799), .A2(\xmem_data[56][6] ), .B1(n24516), .B2(
        \xmem_data[57][6] ), .ZN(n9753) );
  AOI22_X1 U13744 ( .A1(n28334), .A2(\xmem_data[58][6] ), .B1(n20798), .B2(
        \xmem_data[59][6] ), .ZN(n9752) );
  AOI22_X1 U13745 ( .A1(n28752), .A2(\xmem_data[60][6] ), .B1(n23716), .B2(
        \xmem_data[61][6] ), .ZN(n9751) );
  AOI22_X1 U13746 ( .A1(n20800), .A2(\xmem_data[62][6] ), .B1(n17043), .B2(
        \xmem_data[63][6] ), .ZN(n9750) );
  NAND4_X1 U13747 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n9764)
         );
  AOI22_X1 U13748 ( .A1(n20805), .A2(\xmem_data[48][6] ), .B1(n24695), .B2(
        \xmem_data[49][6] ), .ZN(n9757) );
  AOI22_X1 U13749 ( .A1(n20807), .A2(\xmem_data[50][6] ), .B1(n20806), .B2(
        \xmem_data[51][6] ), .ZN(n9756) );
  AOI22_X1 U13750 ( .A1(n20808), .A2(\xmem_data[52][6] ), .B1(n25450), .B2(
        \xmem_data[53][6] ), .ZN(n9755) );
  AOI22_X1 U13751 ( .A1(n20809), .A2(\xmem_data[54][6] ), .B1(n25456), .B2(
        \xmem_data[55][6] ), .ZN(n9754) );
  NAND4_X1 U13752 ( .A1(n9757), .A2(n9756), .A3(n9755), .A4(n9754), .ZN(n9763)
         );
  AOI22_X1 U13753 ( .A1(n20815), .A2(\xmem_data[32][6] ), .B1(n20814), .B2(
        \xmem_data[33][6] ), .ZN(n9761) );
  AOI22_X1 U13754 ( .A1(n21010), .A2(\xmem_data[34][6] ), .B1(n25716), .B2(
        \xmem_data[35][6] ), .ZN(n9760) );
  AOI22_X1 U13755 ( .A1(n20817), .A2(\xmem_data[36][6] ), .B1(n27365), .B2(
        \xmem_data[37][6] ), .ZN(n9759) );
  AOI22_X1 U13756 ( .A1(n20818), .A2(\xmem_data[38][6] ), .B1(n29136), .B2(
        \xmem_data[39][6] ), .ZN(n9758) );
  NAND4_X1 U13757 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n9762)
         );
  OR3_X1 U13758 ( .A1(n9764), .A2(n9763), .A3(n9762), .ZN(n9770) );
  AOI22_X1 U13759 ( .A1(n20826), .A2(\xmem_data[40][6] ), .B1(n20769), .B2(
        \xmem_data[41][6] ), .ZN(n9768) );
  AOI22_X1 U13760 ( .A1(n20827), .A2(\xmem_data[42][6] ), .B1(n24470), .B2(
        \xmem_data[43][6] ), .ZN(n9767) );
  AOI22_X1 U13761 ( .A1(n20828), .A2(\xmem_data[44][6] ), .B1(n25442), .B2(
        \xmem_data[45][6] ), .ZN(n9766) );
  AOI22_X1 U13762 ( .A1(n30962), .A2(\xmem_data[46][6] ), .B1(n3220), .B2(
        \xmem_data[47][6] ), .ZN(n9765) );
  NAND4_X1 U13763 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n9769)
         );
  OAI21_X1 U13764 ( .B1(n9770), .B2(n9769), .A(n20765), .ZN(n9771) );
  XNOR2_X1 U13765 ( .A(n31657), .B(\fmem_data[28][5] ), .ZN(n33322) );
  AOI22_X1 U13766 ( .A1(n27902), .A2(\xmem_data[96][5] ), .B1(n3218), .B2(
        \xmem_data[97][5] ), .ZN(n9778) );
  AOI22_X1 U13767 ( .A1(n20805), .A2(\xmem_data[98][5] ), .B1(n25509), .B2(
        \xmem_data[99][5] ), .ZN(n9777) );
  AOI22_X1 U13768 ( .A1(n27904), .A2(\xmem_data[100][5] ), .B1(n27903), .B2(
        \xmem_data[101][5] ), .ZN(n9776) );
  AOI22_X1 U13769 ( .A1(n27905), .A2(\xmem_data[102][5] ), .B1(n13474), .B2(
        \xmem_data[103][5] ), .ZN(n9775) );
  NAND4_X1 U13770 ( .A1(n9778), .A2(n9777), .A3(n9776), .A4(n9775), .ZN(n9794)
         );
  AOI22_X1 U13771 ( .A1(n25582), .A2(\xmem_data[120][5] ), .B1(n28328), .B2(
        \xmem_data[121][5] ), .ZN(n9782) );
  AOI22_X1 U13772 ( .A1(n30901), .A2(\xmem_data[122][5] ), .B1(n20769), .B2(
        \xmem_data[123][5] ), .ZN(n9781) );
  AOI22_X1 U13773 ( .A1(n27925), .A2(\xmem_data[124][5] ), .B1(n12471), .B2(
        \xmem_data[125][5] ), .ZN(n9780) );
  AOI22_X1 U13774 ( .A1(n23732), .A2(\xmem_data[126][5] ), .B1(n30589), .B2(
        \xmem_data[127][5] ), .ZN(n9779) );
  NAND4_X1 U13775 ( .A1(n9782), .A2(n9781), .A3(n9780), .A4(n9779), .ZN(n9793)
         );
  AOI22_X1 U13776 ( .A1(n27919), .A2(\xmem_data[112][5] ), .B1(n27918), .B2(
        \xmem_data[113][5] ), .ZN(n9786) );
  AOI22_X1 U13777 ( .A1(n27855), .A2(\xmem_data[114][5] ), .B1(n27920), .B2(
        \xmem_data[115][5] ), .ZN(n9785) );
  AOI22_X1 U13778 ( .A1(n3178), .A2(\xmem_data[116][5] ), .B1(n25679), .B2(
        \xmem_data[117][5] ), .ZN(n9784) );
  AOI22_X1 U13779 ( .A1(n29324), .A2(\xmem_data[118][5] ), .B1(n27525), .B2(
        \xmem_data[119][5] ), .ZN(n9783) );
  NAND4_X1 U13780 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(n9792)
         );
  AOI22_X1 U13781 ( .A1(n27910), .A2(\xmem_data[104][5] ), .B1(n28415), .B2(
        \xmem_data[105][5] ), .ZN(n9790) );
  AOI22_X1 U13782 ( .A1(n27911), .A2(\xmem_data[106][5] ), .B1(n24212), .B2(
        \xmem_data[107][5] ), .ZN(n9789) );
  AOI22_X1 U13783 ( .A1(n3176), .A2(\xmem_data[108][5] ), .B1(n27912), .B2(
        \xmem_data[109][5] ), .ZN(n9788) );
  AOI22_X1 U13784 ( .A1(n25519), .A2(\xmem_data[110][5] ), .B1(n22742), .B2(
        \xmem_data[111][5] ), .ZN(n9787) );
  NAND4_X1 U13785 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n9791)
         );
  AOI22_X1 U13786 ( .A1(n27439), .A2(\xmem_data[32][5] ), .B1(n3220), .B2(
        \xmem_data[33][5] ), .ZN(n9799) );
  AOI22_X1 U13787 ( .A1(n28733), .A2(\xmem_data[34][5] ), .B1(n20723), .B2(
        \xmem_data[35][5] ), .ZN(n9798) );
  AOI22_X1 U13788 ( .A1(n27938), .A2(\xmem_data[36][5] ), .B1(n22711), .B2(
        \xmem_data[37][5] ), .ZN(n9797) );
  AOI22_X1 U13789 ( .A1(n29706), .A2(\xmem_data[38][5] ), .B1(n25450), .B2(
        \xmem_data[39][5] ), .ZN(n9796) );
  NAND4_X1 U13790 ( .A1(n9799), .A2(n9798), .A3(n9797), .A4(n9796), .ZN(n9815)
         );
  AOI22_X1 U13791 ( .A1(n22684), .A2(\xmem_data[56][5] ), .B1(n28468), .B2(
        \xmem_data[57][5] ), .ZN(n9803) );
  AOI22_X1 U13792 ( .A1(n31345), .A2(\xmem_data[58][5] ), .B1(n27957), .B2(
        \xmem_data[59][5] ), .ZN(n9802) );
  AOI22_X1 U13793 ( .A1(n27959), .A2(\xmem_data[60][5] ), .B1(n27958), .B2(
        \xmem_data[61][5] ), .ZN(n9801) );
  AOI22_X1 U13794 ( .A1(n3352), .A2(\xmem_data[62][5] ), .B1(n20568), .B2(
        \xmem_data[63][5] ), .ZN(n9800) );
  NAND4_X1 U13795 ( .A1(n9803), .A2(n9802), .A3(n9801), .A4(n9800), .ZN(n9814)
         );
  AOI22_X1 U13796 ( .A1(n20585), .A2(\xmem_data[48][5] ), .B1(n29048), .B2(
        \xmem_data[49][5] ), .ZN(n9807) );
  AOI22_X1 U13797 ( .A1(n29047), .A2(\xmem_data[50][5] ), .B1(n27950), .B2(
        \xmem_data[51][5] ), .ZN(n9806) );
  AOI22_X1 U13798 ( .A1(n27952), .A2(\xmem_data[52][5] ), .B1(n27951), .B2(
        \xmem_data[53][5] ), .ZN(n9805) );
  AOI22_X1 U13799 ( .A1(n17004), .A2(\xmem_data[54][5] ), .B1(n31362), .B2(
        \xmem_data[55][5] ), .ZN(n9804) );
  NAND4_X1 U13800 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n9813)
         );
  AOI22_X1 U13801 ( .A1(n25422), .A2(\xmem_data[40][5] ), .B1(n3357), .B2(
        \xmem_data[41][5] ), .ZN(n9811) );
  AOI22_X1 U13802 ( .A1(n27944), .A2(\xmem_data[42][5] ), .B1(n20775), .B2(
        \xmem_data[43][5] ), .ZN(n9810) );
  AOI22_X1 U13803 ( .A1(n24131), .A2(\xmem_data[44][5] ), .B1(n23793), .B2(
        \xmem_data[45][5] ), .ZN(n9809) );
  AOI22_X1 U13804 ( .A1(n29437), .A2(\xmem_data[46][5] ), .B1(n27516), .B2(
        \xmem_data[47][5] ), .ZN(n9808) );
  NAND4_X1 U13805 ( .A1(n9811), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(n9812)
         );
  AOI22_X1 U13806 ( .A1(n31348), .A2(\xmem_data[64][5] ), .B1(n3221), .B2(
        \xmem_data[65][5] ), .ZN(n9823) );
  AOI22_X1 U13807 ( .A1(n27938), .A2(\xmem_data[68][5] ), .B1(n20559), .B2(
        \xmem_data[69][5] ), .ZN(n9817) );
  INV_X1 U13808 ( .A(n9817), .ZN(n9821) );
  AOI22_X1 U13809 ( .A1(n29026), .A2(\xmem_data[66][5] ), .B1(n25491), .B2(
        \xmem_data[67][5] ), .ZN(n9819) );
  AOI22_X1 U13810 ( .A1(n24702), .A2(\xmem_data[70][5] ), .B1(n28045), .B2(
        \xmem_data[71][5] ), .ZN(n9818) );
  NAND2_X1 U13811 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  NOR2_X1 U13812 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U13813 ( .A1(n9823), .A2(n9822), .ZN(n9842) );
  AOI22_X1 U13814 ( .A1(n28337), .A2(\xmem_data[80][5] ), .B1(n25677), .B2(
        \xmem_data[81][5] ), .ZN(n9827) );
  AOI22_X1 U13815 ( .A1(n31255), .A2(\xmem_data[82][5] ), .B1(n27950), .B2(
        \xmem_data[83][5] ), .ZN(n9826) );
  AOI22_X1 U13816 ( .A1(n27952), .A2(\xmem_data[84][5] ), .B1(n27951), .B2(
        \xmem_data[85][5] ), .ZN(n9825) );
  AOI22_X1 U13817 ( .A1(n3301), .A2(\xmem_data[86][5] ), .B1(n31314), .B2(
        \xmem_data[87][5] ), .ZN(n9824) );
  NAND4_X1 U13818 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9841)
         );
  AOI22_X1 U13819 ( .A1(n27447), .A2(\xmem_data[72][5] ), .B1(n28415), .B2(
        \xmem_data[73][5] ), .ZN(n9831) );
  AOI22_X1 U13820 ( .A1(n27944), .A2(\xmem_data[74][5] ), .B1(n24448), .B2(
        \xmem_data[75][5] ), .ZN(n9830) );
  AOI22_X1 U13821 ( .A1(n29272), .A2(\xmem_data[76][5] ), .B1(n22741), .B2(
        \xmem_data[77][5] ), .ZN(n9829) );
  AOI22_X1 U13822 ( .A1(n30746), .A2(\xmem_data[78][5] ), .B1(n29162), .B2(
        \xmem_data[79][5] ), .ZN(n9828) );
  NAND4_X1 U13823 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n9840)
         );
  AOI22_X1 U13824 ( .A1(n27498), .A2(\xmem_data[90][5] ), .B1(n27957), .B2(
        \xmem_data[91][5] ), .ZN(n9838) );
  AOI22_X1 U13825 ( .A1(n27959), .A2(\xmem_data[92][5] ), .B1(n27958), .B2(
        \xmem_data[93][5] ), .ZN(n9837) );
  AOI22_X1 U13826 ( .A1(n25582), .A2(\xmem_data[88][5] ), .B1(n25359), .B2(
        \xmem_data[89][5] ), .ZN(n9832) );
  INV_X1 U13827 ( .A(n9832), .ZN(n9835) );
  AOI22_X1 U13828 ( .A1(n3335), .A2(\xmem_data[94][5] ), .B1(n29286), .B2(
        \xmem_data[95][5] ), .ZN(n9833) );
  INV_X1 U13829 ( .A(n9833), .ZN(n9834) );
  NOR2_X1 U13830 ( .A1(n9835), .A2(n9834), .ZN(n9836) );
  NAND3_X1 U13831 ( .A1(n9838), .A2(n9837), .A3(n9836), .ZN(n9839) );
  AND2_X1 U13832 ( .A1(n25422), .A2(\xmem_data[8][5] ), .ZN(n9845) );
  AND2_X1 U13833 ( .A1(n29157), .A2(\xmem_data[6][5] ), .ZN(n9844) );
  OR2_X1 U13834 ( .A1(n9845), .A2(n9844), .ZN(n9848) );
  AOI22_X1 U13835 ( .A1(n23770), .A2(\xmem_data[2][5] ), .B1(n27869), .B2(
        \xmem_data[3][5] ), .ZN(n9846) );
  INV_X1 U13836 ( .A(n9846), .ZN(n9847) );
  NOR2_X1 U13837 ( .A1(n9848), .A2(n9847), .ZN(n9851) );
  AOI22_X1 U13838 ( .A1(n27502), .A2(\xmem_data[0][5] ), .B1(n3219), .B2(
        \xmem_data[1][5] ), .ZN(n9850) );
  AOI22_X1 U13839 ( .A1(n21069), .A2(\xmem_data[4][5] ), .B1(n30550), .B2(
        \xmem_data[5][5] ), .ZN(n9849) );
  AOI22_X1 U13840 ( .A1(n24133), .A2(\xmem_data[16][5] ), .B1(n31270), .B2(
        \xmem_data[17][5] ), .ZN(n9855) );
  AOI22_X1 U13841 ( .A1(n27855), .A2(\xmem_data[18][5] ), .B1(n29190), .B2(
        \xmem_data[19][5] ), .ZN(n9854) );
  AOI22_X1 U13842 ( .A1(n27462), .A2(\xmem_data[20][5] ), .B1(n25679), .B2(
        \xmem_data[21][5] ), .ZN(n9853) );
  AOI22_X1 U13843 ( .A1(n29573), .A2(\xmem_data[22][5] ), .B1(n20553), .B2(
        \xmem_data[23][5] ), .ZN(n9852) );
  NAND4_X1 U13844 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9856)
         );
  AOI22_X1 U13845 ( .A1(n22738), .A2(\xmem_data[10][5] ), .B1(n31326), .B2(
        \xmem_data[11][5] ), .ZN(n9861) );
  AOI22_X1 U13846 ( .A1(n28052), .A2(\xmem_data[13][5] ), .B1(
        \xmem_data[9][5] ), .B2(n27863), .ZN(n9859) );
  AOI22_X1 U13847 ( .A1(n27864), .A2(\xmem_data[15][5] ), .B1(
        \xmem_data[14][5] ), .B2(n3121), .ZN(n9858) );
  AND2_X1 U13848 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  NAND2_X1 U13849 ( .A1(n9861), .A2(n9860), .ZN(n9868) );
  AOI22_X1 U13850 ( .A1(n27847), .A2(\xmem_data[24][5] ), .B1(n28292), .B2(
        \xmem_data[25][5] ), .ZN(n9866) );
  AND2_X1 U13851 ( .A1(n25440), .A2(\xmem_data[27][5] ), .ZN(n9862) );
  AOI21_X1 U13852 ( .B1(n27852), .B2(\xmem_data[26][5] ), .A(n9862), .ZN(n9865) );
  AOI22_X1 U13853 ( .A1(n27564), .A2(\xmem_data[28][5] ), .B1(n31262), .B2(
        \xmem_data[29][5] ), .ZN(n9864) );
  AOI22_X1 U13854 ( .A1(n3413), .A2(\xmem_data[30][5] ), .B1(n20568), .B2(
        \xmem_data[31][5] ), .ZN(n9863) );
  NAND4_X1 U13855 ( .A1(n9866), .A2(n9865), .A3(n9864), .A4(n9863), .ZN(n9867)
         );
  XOR2_X1 U13856 ( .A(\fmem_data[14][5] ), .B(\fmem_data[14][4] ), .Z(n9875)
         );
  AOI22_X1 U13857 ( .A1(n3131), .A2(\xmem_data[6][6] ), .B1(n29045), .B2(
        \xmem_data[7][6] ), .ZN(n9876) );
  INV_X1 U13858 ( .A(n9876), .ZN(n9898) );
  AOI22_X1 U13859 ( .A1(n20518), .A2(\xmem_data[0][6] ), .B1(n3217), .B2(
        \xmem_data[1][6] ), .ZN(n9879) );
  AOI22_X1 U13860 ( .A1(n28475), .A2(\xmem_data[4][6] ), .B1(n27994), .B2(
        \xmem_data[5][6] ), .ZN(n9878) );
  AOI22_X1 U13861 ( .A1(n28733), .A2(\xmem_data[2][6] ), .B1(n27869), .B2(
        \xmem_data[3][6] ), .ZN(n9877) );
  NAND3_X1 U13862 ( .A1(n9879), .A2(n9878), .A3(n9877), .ZN(n9895) );
  AOI22_X1 U13863 ( .A1(n28050), .A2(\xmem_data[8][6] ), .B1(n27863), .B2(
        \xmem_data[9][6] ), .ZN(n9883) );
  AOI22_X1 U13864 ( .A1(n22738), .A2(\xmem_data[10][6] ), .B1(n25605), .B2(
        \xmem_data[11][6] ), .ZN(n9882) );
  AOI22_X1 U13865 ( .A1(n28298), .A2(\xmem_data[12][6] ), .B1(n25572), .B2(
        \xmem_data[13][6] ), .ZN(n9881) );
  AOI22_X1 U13866 ( .A1(n24545), .A2(\xmem_data[14][6] ), .B1(n27864), .B2(
        \xmem_data[15][6] ), .ZN(n9880) );
  NAND4_X1 U13867 ( .A1(n9883), .A2(n9882), .A3(n9881), .A4(n9880), .ZN(n9894)
         );
  AOI22_X1 U13868 ( .A1(n28337), .A2(\xmem_data[16][6] ), .B1(n22718), .B2(
        \xmem_data[17][6] ), .ZN(n9887) );
  AOI22_X1 U13869 ( .A1(n27855), .A2(\xmem_data[18][6] ), .B1(n28380), .B2(
        \xmem_data[19][6] ), .ZN(n9886) );
  AOI22_X1 U13870 ( .A1(n30899), .A2(\xmem_data[20][6] ), .B1(n27856), .B2(
        \xmem_data[21][6] ), .ZN(n9885) );
  AOI22_X1 U13871 ( .A1(n3337), .A2(\xmem_data[22][6] ), .B1(n29245), .B2(
        \xmem_data[23][6] ), .ZN(n9884) );
  NAND4_X1 U13872 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n9893)
         );
  AOI22_X1 U13873 ( .A1(n27847), .A2(\xmem_data[24][6] ), .B1(n20733), .B2(
        \xmem_data[25][6] ), .ZN(n9891) );
  AOI22_X1 U13874 ( .A1(n27852), .A2(\xmem_data[26][6] ), .B1(n24624), .B2(
        \xmem_data[27][6] ), .ZN(n9890) );
  AOI22_X1 U13875 ( .A1(n29124), .A2(\xmem_data[28][6] ), .B1(n22752), .B2(
        \xmem_data[29][6] ), .ZN(n9889) );
  AOI22_X1 U13876 ( .A1(n3384), .A2(\xmem_data[30][6] ), .B1(n27437), .B2(
        \xmem_data[31][6] ), .ZN(n9888) );
  NAND4_X1 U13877 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n9892)
         );
  OR4_X1 U13878 ( .A1(n9895), .A2(n9894), .A3(n9893), .A4(n9892), .ZN(n9897)
         );
  OAI21_X1 U13879 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9899) );
  AOI22_X1 U13880 ( .A1(n31348), .A2(\xmem_data[64][6] ), .B1(n3219), .B2(
        \xmem_data[65][6] ), .ZN(n9907) );
  AOI22_X1 U13881 ( .A1(n27938), .A2(\xmem_data[68][6] ), .B1(n3255), .B2(
        \xmem_data[69][6] ), .ZN(n9900) );
  INV_X1 U13882 ( .A(n9900), .ZN(n9905) );
  AOI22_X1 U13883 ( .A1(n17063), .A2(\xmem_data[70][6] ), .B1(n15011), .B2(
        \xmem_data[71][6] ), .ZN(n9901) );
  INV_X1 U13884 ( .A(n9901), .ZN(n9904) );
  AOI22_X1 U13885 ( .A1(n29698), .A2(n20682), .B1(n14989), .B2(
        \xmem_data[67][6] ), .ZN(n9902) );
  INV_X1 U13886 ( .A(n9902), .ZN(n9903) );
  NOR3_X1 U13887 ( .A1(n9905), .A2(n9904), .A3(n9903), .ZN(n9906) );
  NAND2_X1 U13888 ( .A1(n9907), .A2(n9906), .ZN(n9923) );
  AOI22_X1 U13889 ( .A1(n27447), .A2(\xmem_data[72][6] ), .B1(n25456), .B2(
        \xmem_data[73][6] ), .ZN(n9911) );
  AOI22_X1 U13890 ( .A1(n27944), .A2(\xmem_data[74][6] ), .B1(n20775), .B2(
        \xmem_data[75][6] ), .ZN(n9910) );
  AOI22_X1 U13891 ( .A1(n31268), .A2(\xmem_data[76][6] ), .B1(n24160), .B2(
        \xmem_data[77][6] ), .ZN(n9909) );
  AOI22_X1 U13892 ( .A1(n27818), .A2(\xmem_data[78][6] ), .B1(n27516), .B2(
        \xmem_data[79][6] ), .ZN(n9908) );
  NAND4_X1 U13893 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(n9922)
         );
  AOI22_X1 U13894 ( .A1(n21007), .A2(\xmem_data[80][6] ), .B1(n25398), .B2(
        \xmem_data[81][6] ), .ZN(n9915) );
  AOI22_X1 U13895 ( .A1(n29239), .A2(\xmem_data[82][6] ), .B1(n27950), .B2(
        \xmem_data[83][6] ), .ZN(n9914) );
  AOI22_X1 U13896 ( .A1(n27952), .A2(\xmem_data[84][6] ), .B1(n27951), .B2(
        \xmem_data[85][6] ), .ZN(n9913) );
  AOI22_X1 U13897 ( .A1(n20984), .A2(\xmem_data[86][6] ), .B1(n25583), .B2(
        \xmem_data[87][6] ), .ZN(n9912) );
  NAND4_X1 U13898 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n9921)
         );
  AOI22_X1 U13899 ( .A1(n25582), .A2(\xmem_data[88][6] ), .B1(n11008), .B2(
        \xmem_data[89][6] ), .ZN(n9919) );
  AOI22_X1 U13900 ( .A1(n25584), .A2(\xmem_data[90][6] ), .B1(n27957), .B2(
        \xmem_data[91][6] ), .ZN(n9918) );
  AOI22_X1 U13901 ( .A1(n27959), .A2(\xmem_data[92][6] ), .B1(n27958), .B2(
        \xmem_data[93][6] ), .ZN(n9917) );
  AOI22_X1 U13902 ( .A1(n3228), .A2(\xmem_data[94][6] ), .B1(n25485), .B2(
        \xmem_data[95][6] ), .ZN(n9916) );
  NAND4_X1 U13903 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n9920)
         );
  OR4_X1 U13904 ( .A1(n9923), .A2(n9922), .A3(n9921), .A4(n9920), .ZN(n9924)
         );
  NAND2_X1 U13905 ( .A1(n9924), .A2(n27935), .ZN(n9947) );
  AOI22_X1 U13906 ( .A1(n27902), .A2(\xmem_data[96][6] ), .B1(n3220), .B2(
        \xmem_data[97][6] ), .ZN(n9928) );
  AOI22_X1 U13907 ( .A1(n21067), .A2(\xmem_data[98][6] ), .B1(n20787), .B2(
        \xmem_data[99][6] ), .ZN(n9927) );
  AOI22_X1 U13908 ( .A1(n27904), .A2(\xmem_data[100][6] ), .B1(n27903), .B2(
        \xmem_data[101][6] ), .ZN(n9926) );
  AOI22_X1 U13909 ( .A1(n27905), .A2(\xmem_data[102][6] ), .B1(n23771), .B2(
        \xmem_data[103][6] ), .ZN(n9925) );
  NAND4_X1 U13910 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n9944)
         );
  AOI22_X1 U13911 ( .A1(n27910), .A2(\xmem_data[104][6] ), .B1(n28415), .B2(
        \xmem_data[105][6] ), .ZN(n9932) );
  AOI22_X1 U13912 ( .A1(n27911), .A2(\xmem_data[106][6] ), .B1(n24212), .B2(
        \xmem_data[107][6] ), .ZN(n9931) );
  AOI22_X1 U13913 ( .A1(n3175), .A2(\xmem_data[108][6] ), .B1(n27912), .B2(
        \xmem_data[109][6] ), .ZN(n9930) );
  AOI22_X1 U13914 ( .A1(n28053), .A2(\xmem_data[110][6] ), .B1(n25383), .B2(
        \xmem_data[111][6] ), .ZN(n9929) );
  NAND4_X1 U13915 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9943)
         );
  AOI22_X1 U13916 ( .A1(n27919), .A2(\xmem_data[112][6] ), .B1(n27918), .B2(
        \xmem_data[113][6] ), .ZN(n9936) );
  AOI22_X1 U13917 ( .A1(n28302), .A2(\xmem_data[114][6] ), .B1(n27920), .B2(
        \xmem_data[115][6] ), .ZN(n9935) );
  AOI22_X1 U13918 ( .A1(n21010), .A2(\xmem_data[116][6] ), .B1(n20943), .B2(
        \xmem_data[117][6] ), .ZN(n9934) );
  AOI22_X1 U13919 ( .A1(n3300), .A2(\xmem_data[118][6] ), .B1(n14883), .B2(
        \xmem_data[119][6] ), .ZN(n9933) );
  NAND4_X1 U13920 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(n9942)
         );
  AOI22_X1 U13921 ( .A1(n24467), .A2(\xmem_data[120][6] ), .B1(n27981), .B2(
        \xmem_data[121][6] ), .ZN(n9940) );
  AOI22_X1 U13922 ( .A1(n14982), .A2(\xmem_data[122][6] ), .B1(n28329), .B2(
        \xmem_data[123][6] ), .ZN(n9939) );
  AOI22_X1 U13923 ( .A1(n27925), .A2(\xmem_data[124][6] ), .B1(n22752), .B2(
        \xmem_data[125][6] ), .ZN(n9938) );
  AOI22_X1 U13924 ( .A1(n23754), .A2(\xmem_data[126][6] ), .B1(n25360), .B2(
        \xmem_data[127][6] ), .ZN(n9937) );
  NAND4_X1 U13925 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), .ZN(n9941)
         );
  OR4_X1 U13926 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9945)
         );
  NAND2_X1 U13927 ( .A1(n9945), .A2(n27937), .ZN(n9946) );
  NAND2_X1 U13928 ( .A1(n9947), .A2(n9946), .ZN(n9970) );
  AOI22_X1 U13929 ( .A1(n31348), .A2(\xmem_data[32][6] ), .B1(n3218), .B2(
        \xmem_data[33][6] ), .ZN(n9951) );
  AOI22_X1 U13930 ( .A1(n24563), .A2(\xmem_data[34][6] ), .B1(n29028), .B2(
        \xmem_data[35][6] ), .ZN(n9950) );
  AOI22_X1 U13931 ( .A1(n27938), .A2(\xmem_data[36][6] ), .B1(n28509), .B2(
        \xmem_data[37][6] ), .ZN(n9949) );
  AOI22_X1 U13932 ( .A1(n24702), .A2(\xmem_data[38][6] ), .B1(n28007), .B2(
        \xmem_data[39][6] ), .ZN(n9948) );
  NAND4_X1 U13933 ( .A1(n9951), .A2(n9950), .A3(n9949), .A4(n9948), .ZN(n9967)
         );
  AOI22_X1 U13934 ( .A1(n25422), .A2(\xmem_data[40][6] ), .B1(n27943), .B2(
        \xmem_data[41][6] ), .ZN(n9955) );
  AOI22_X1 U13935 ( .A1(n27944), .A2(\xmem_data[42][6] ), .B1(n24212), .B2(
        \xmem_data[43][6] ), .ZN(n9954) );
  AOI22_X1 U13936 ( .A1(n29023), .A2(\xmem_data[44][6] ), .B1(n23793), .B2(
        \xmem_data[45][6] ), .ZN(n9953) );
  AOI22_X1 U13937 ( .A1(n29605), .A2(\xmem_data[46][6] ), .B1(n27516), .B2(
        \xmem_data[47][6] ), .ZN(n9952) );
  NAND4_X1 U13938 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9966)
         );
  AOI22_X1 U13939 ( .A1(n23764), .A2(\xmem_data[48][6] ), .B1(n24707), .B2(
        \xmem_data[49][6] ), .ZN(n9959) );
  AOI22_X1 U13940 ( .A1(n30893), .A2(\xmem_data[50][6] ), .B1(n27950), .B2(
        \xmem_data[51][6] ), .ZN(n9958) );
  AOI22_X1 U13941 ( .A1(n27952), .A2(\xmem_data[52][6] ), .B1(n27951), .B2(
        \xmem_data[53][6] ), .ZN(n9957) );
  AOI22_X1 U13942 ( .A1(n29297), .A2(\xmem_data[54][6] ), .B1(n27975), .B2(
        \xmem_data[55][6] ), .ZN(n9956) );
  NAND4_X1 U13943 ( .A1(n9959), .A2(n9958), .A3(n9957), .A4(n9956), .ZN(n9965)
         );
  AOI22_X1 U13944 ( .A1(n25582), .A2(\xmem_data[56][6] ), .B1(n25406), .B2(
        \xmem_data[57][6] ), .ZN(n9963) );
  AOI22_X1 U13945 ( .A1(n28241), .A2(\xmem_data[58][6] ), .B1(n27957), .B2(
        \xmem_data[59][6] ), .ZN(n9962) );
  AOI22_X1 U13946 ( .A1(n27959), .A2(\xmem_data[60][6] ), .B1(n27958), .B2(
        \xmem_data[61][6] ), .ZN(n9961) );
  AOI22_X1 U13947 ( .A1(n25624), .A2(\xmem_data[62][6] ), .B1(n25442), .B2(
        \xmem_data[63][6] ), .ZN(n9960) );
  NAND4_X1 U13948 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9964)
         );
  OR4_X1 U13949 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n9968)
         );
  AND2_X1 U13950 ( .A1(n9968), .A2(n27968), .ZN(n9969) );
  XNOR2_X1 U13951 ( .A(n31799), .B(\fmem_data[14][5] ), .ZN(n33099) );
  XOR2_X1 U13952 ( .A(\fmem_data[21][2] ), .B(\fmem_data[21][3] ), .Z(n9972)
         );
  AOI22_X1 U13953 ( .A1(n20488), .A2(\xmem_data[32][7] ), .B1(n20577), .B2(
        \xmem_data[33][7] ), .ZN(n9977) );
  AOI22_X1 U13954 ( .A1(n20579), .A2(\xmem_data[34][7] ), .B1(n27436), .B2(
        \xmem_data[35][7] ), .ZN(n9976) );
  AOI22_X1 U13955 ( .A1(n20578), .A2(\xmem_data[36][7] ), .B1(n28677), .B2(
        \xmem_data[37][7] ), .ZN(n9975) );
  AND2_X1 U13956 ( .A1(n25442), .A2(\xmem_data[38][7] ), .ZN(n9973) );
  AOI21_X1 U13957 ( .B1(n20518), .B2(\xmem_data[39][7] ), .A(n9973), .ZN(n9974) );
  NAND4_X1 U13958 ( .A1(n9977), .A2(n9976), .A3(n9975), .A4(n9974), .ZN(n9994)
         );
  AOI22_X1 U13959 ( .A1(n20588), .A2(\xmem_data[48][7] ), .B1(n20587), .B2(
        \xmem_data[49][7] ), .ZN(n9981) );
  AOI22_X1 U13960 ( .A1(n25605), .A2(\xmem_data[50][7] ), .B1(n30514), .B2(
        \xmem_data[51][7] ), .ZN(n9980) );
  AOI22_X1 U13961 ( .A1(n20584), .A2(\xmem_data[52][7] ), .B1(n31354), .B2(
        \xmem_data[53][7] ), .ZN(n9979) );
  AOI22_X1 U13962 ( .A1(n20586), .A2(\xmem_data[54][7] ), .B1(n20585), .B2(
        \xmem_data[55][7] ), .ZN(n9978) );
  NAND4_X1 U13963 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n9992)
         );
  AOI22_X1 U13964 ( .A1(n31355), .A2(\xmem_data[56][7] ), .B1(n20730), .B2(
        \xmem_data[57][7] ), .ZN(n9985) );
  AOI22_X1 U13965 ( .A1(n25435), .A2(\xmem_data[58][7] ), .B1(n17002), .B2(
        \xmem_data[59][7] ), .ZN(n9984) );
  AOI22_X1 U13966 ( .A1(n27951), .A2(\xmem_data[60][7] ), .B1(n24571), .B2(
        \xmem_data[61][7] ), .ZN(n9983) );
  AOI22_X1 U13967 ( .A1(n14975), .A2(\xmem_data[62][7] ), .B1(n25526), .B2(
        \xmem_data[63][7] ), .ZN(n9982) );
  NAND4_X1 U13968 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n9991)
         );
  AOI22_X1 U13969 ( .A1(n3222), .A2(\xmem_data[40][7] ), .B1(n20724), .B2(
        \xmem_data[41][7] ), .ZN(n9989) );
  AOI22_X1 U13970 ( .A1(n20598), .A2(\xmem_data[42][7] ), .B1(n25694), .B2(
        \xmem_data[43][7] ), .ZN(n9988) );
  AOI22_X1 U13971 ( .A1(n13444), .A2(\xmem_data[44][7] ), .B1(n20962), .B2(
        \xmem_data[45][7] ), .ZN(n9987) );
  AOI22_X1 U13972 ( .A1(n28007), .A2(\xmem_data[46][7] ), .B1(n25422), .B2(
        \xmem_data[47][7] ), .ZN(n9986) );
  NAND4_X1 U13973 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n9990)
         );
  OR3_X1 U13974 ( .A1(n9992), .A2(n9991), .A3(n9990), .ZN(n9993) );
  OAI21_X1 U13975 ( .B1(n9994), .B2(n9993), .A(n20606), .ZN(n9995) );
  INV_X1 U13976 ( .A(n9995), .ZN(n10043) );
  AOI22_X1 U13977 ( .A1(n3222), .A2(\xmem_data[104][7] ), .B1(n27445), .B2(
        \xmem_data[105][7] ), .ZN(n9999) );
  AOI22_X1 U13978 ( .A1(n20558), .A2(\xmem_data[106][7] ), .B1(n20994), .B2(
        \xmem_data[107][7] ), .ZN(n9998) );
  AOI22_X1 U13979 ( .A1(n20559), .A2(\xmem_data[108][7] ), .B1(n25417), .B2(
        \xmem_data[109][7] ), .ZN(n9997) );
  AOI22_X1 U13980 ( .A1(n27446), .A2(\xmem_data[110][7] ), .B1(n25707), .B2(
        \xmem_data[111][7] ), .ZN(n9996) );
  NAND4_X1 U13981 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n10010) );
  AOI22_X1 U13982 ( .A1(n20546), .A2(\xmem_data[112][7] ), .B1(n20545), .B2(
        \xmem_data[113][7] ), .ZN(n10003) );
  AOI22_X1 U13983 ( .A1(n22675), .A2(\xmem_data[114][7] ), .B1(n28980), .B2(
        \xmem_data[115][7] ), .ZN(n10002) );
  AOI22_X1 U13984 ( .A1(n20544), .A2(\xmem_data[116][7] ), .B1(n28752), .B2(
        \xmem_data[117][7] ), .ZN(n10001) );
  AOI22_X1 U13985 ( .A1(n20543), .A2(\xmem_data[118][7] ), .B1(n20542), .B2(
        \xmem_data[119][7] ), .ZN(n10000) );
  NAND4_X1 U13986 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10009) );
  AOI22_X1 U13987 ( .A1(n25677), .A2(\xmem_data[120][7] ), .B1(n22717), .B2(
        \xmem_data[121][7] ), .ZN(n10007) );
  AOI22_X1 U13988 ( .A1(n27950), .A2(\xmem_data[122][7] ), .B1(n28428), .B2(
        \xmem_data[123][7] ), .ZN(n10006) );
  AOI22_X1 U13989 ( .A1(n20551), .A2(\xmem_data[124][7] ), .B1(n23780), .B2(
        \xmem_data[125][7] ), .ZN(n10005) );
  AOI22_X1 U13990 ( .A1(n20553), .A2(\xmem_data[126][7] ), .B1(n20552), .B2(
        \xmem_data[127][7] ), .ZN(n10004) );
  NAND4_X1 U13991 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n10008) );
  AOI22_X1 U13992 ( .A1(n29136), .A2(\xmem_data[96][7] ), .B1(n20567), .B2(
        \xmem_data[97][7] ), .ZN(n10014) );
  AOI22_X1 U13993 ( .A1(n17050), .A2(\xmem_data[98][7] ), .B1(n28038), .B2(
        \xmem_data[99][7] ), .ZN(n10013) );
  AOI22_X1 U13994 ( .A1(n29118), .A2(\xmem_data[100][7] ), .B1(n28718), .B2(
        \xmem_data[101][7] ), .ZN(n10012) );
  AOI22_X1 U13995 ( .A1(n20568), .A2(\xmem_data[102][7] ), .B1(n20518), .B2(
        \xmem_data[103][7] ), .ZN(n10011) );
  NAND4_X1 U13996 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10015) );
  OAI21_X1 U13997 ( .B1(n10016), .B2(n10015), .A(n20538), .ZN(n10041) );
  AND2_X1 U13998 ( .A1(n23725), .A2(\xmem_data[64][7] ), .ZN(n10017) );
  AOI21_X1 U13999 ( .B1(n20577), .B2(\xmem_data[65][7] ), .A(n10017), .ZN(
        n10022) );
  AOI22_X1 U14000 ( .A1(n20579), .A2(\xmem_data[66][7] ), .B1(n25630), .B2(
        \xmem_data[67][7] ), .ZN(n10021) );
  AOI22_X1 U14001 ( .A1(n20578), .A2(\xmem_data[68][7] ), .B1(n3434), .B2(
        \xmem_data[69][7] ), .ZN(n10020) );
  AND2_X1 U14002 ( .A1(n22753), .A2(\xmem_data[70][7] ), .ZN(n10018) );
  AOI21_X1 U14003 ( .B1(n20576), .B2(\xmem_data[71][7] ), .A(n10018), .ZN(
        n10019) );
  NAND4_X1 U14004 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10039) );
  AOI22_X1 U14005 ( .A1(n20584), .A2(\xmem_data[84][7] ), .B1(n25672), .B2(
        \xmem_data[85][7] ), .ZN(n10026) );
  AOI22_X1 U14006 ( .A1(n30552), .A2(\xmem_data[82][7] ), .B1(n28298), .B2(
        \xmem_data[83][7] ), .ZN(n10025) );
  AOI22_X1 U14007 ( .A1(n20588), .A2(\xmem_data[80][7] ), .B1(n20587), .B2(
        \xmem_data[81][7] ), .ZN(n10024) );
  AOI22_X1 U14008 ( .A1(n20586), .A2(\xmem_data[86][7] ), .B1(n20585), .B2(
        \xmem_data[87][7] ), .ZN(n10023) );
  NAND4_X1 U14009 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10037) );
  AOI22_X1 U14010 ( .A1(n31270), .A2(\xmem_data[88][7] ), .B1(n24710), .B2(
        \xmem_data[89][7] ), .ZN(n10030) );
  AOI22_X1 U14011 ( .A1(n30515), .A2(\xmem_data[90][7] ), .B1(n24190), .B2(
        \xmem_data[91][7] ), .ZN(n10029) );
  AOI22_X1 U14012 ( .A1(n20551), .A2(\xmem_data[92][7] ), .B1(n29324), .B2(
        \xmem_data[93][7] ), .ZN(n10028) );
  AOI22_X1 U14013 ( .A1(n24521), .A2(\xmem_data[94][7] ), .B1(n3179), .B2(
        \xmem_data[95][7] ), .ZN(n10027) );
  NAND4_X1 U14014 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n10036) );
  AOI22_X1 U14015 ( .A1(n3220), .A2(\xmem_data[72][7] ), .B1(n21067), .B2(
        \xmem_data[73][7] ), .ZN(n10034) );
  AOI22_X1 U14016 ( .A1(n20598), .A2(\xmem_data[74][7] ), .B1(n25617), .B2(
        \xmem_data[75][7] ), .ZN(n10033) );
  AOI22_X1 U14017 ( .A1(n25486), .A2(\xmem_data[76][7] ), .B1(n29157), .B2(
        \xmem_data[77][7] ), .ZN(n10032) );
  AOI22_X1 U14018 ( .A1(n3231), .A2(\xmem_data[78][7] ), .B1(n24450), .B2(
        \xmem_data[79][7] ), .ZN(n10031) );
  NAND4_X1 U14019 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10035) );
  OR3_X1 U14020 ( .A1(n10037), .A2(n10036), .A3(n10035), .ZN(n10038) );
  OAI21_X1 U14021 ( .B1(n10039), .B2(n10038), .A(n20573), .ZN(n10040) );
  NAND2_X1 U14022 ( .A1(n10041), .A2(n10040), .ZN(n10042) );
  NOR2_X1 U14023 ( .A1(n10043), .A2(n10042), .ZN(n10067) );
  AOI22_X1 U14024 ( .A1(n28045), .A2(\xmem_data[14][7] ), .B1(n25422), .B2(
        \xmem_data[15][7] ), .ZN(n10044) );
  INV_X1 U14025 ( .A(n10044), .ZN(n10065) );
  AOI22_X1 U14026 ( .A1(n20505), .A2(\xmem_data[24][7] ), .B1(n30309), .B2(
        \xmem_data[25][7] ), .ZN(n10048) );
  AOI22_X1 U14027 ( .A1(n13481), .A2(\xmem_data[26][7] ), .B1(n14972), .B2(
        \xmem_data[27][7] ), .ZN(n10047) );
  AOI22_X1 U14028 ( .A1(n28327), .A2(\xmem_data[28][7] ), .B1(n29816), .B2(
        \xmem_data[29][7] ), .ZN(n10046) );
  AOI22_X1 U14029 ( .A1(n20507), .A2(\xmem_data[30][7] ), .B1(n20734), .B2(
        \xmem_data[31][7] ), .ZN(n10045) );
  NAND4_X1 U14030 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10063) );
  AOI22_X1 U14031 ( .A1(n20546), .A2(\xmem_data[16][7] ), .B1(n20799), .B2(
        \xmem_data[17][7] ), .ZN(n10052) );
  AOI22_X1 U14032 ( .A1(n13168), .A2(\xmem_data[18][7] ), .B1(n29023), .B2(
        \xmem_data[19][7] ), .ZN(n10051) );
  AOI22_X1 U14033 ( .A1(n29046), .A2(\xmem_data[20][7] ), .B1(n3120), .B2(
        \xmem_data[21][7] ), .ZN(n10050) );
  AOI22_X1 U14034 ( .A1(n31269), .A2(\xmem_data[22][7] ), .B1(n28096), .B2(
        \xmem_data[23][7] ), .ZN(n10049) );
  NAND4_X1 U14035 ( .A1(n10052), .A2(n10051), .A3(n10050), .A4(n10049), .ZN(
        n10062) );
  AOI22_X1 U14036 ( .A1(n20488), .A2(\xmem_data[0][7] ), .B1(n20708), .B2(
        \xmem_data[1][7] ), .ZN(n10056) );
  AOI22_X1 U14037 ( .A1(n20707), .A2(\xmem_data[2][7] ), .B1(n24526), .B2(
        \xmem_data[3][7] ), .ZN(n10055) );
  AOI22_X1 U14038 ( .A1(n20489), .A2(\xmem_data[4][7] ), .B1(n3412), .B2(
        \xmem_data[5][7] ), .ZN(n10054) );
  AOI22_X1 U14039 ( .A1(n25360), .A2(\xmem_data[6][7] ), .B1(n20576), .B2(
        \xmem_data[7][7] ), .ZN(n10053) );
  NAND4_X1 U14040 ( .A1(n10056), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(
        n10061) );
  AOI22_X1 U14041 ( .A1(n25415), .A2(\xmem_data[12][7] ), .B1(n30295), .B2(
        \xmem_data[13][7] ), .ZN(n10059) );
  AOI22_X1 U14042 ( .A1(n20500), .A2(\xmem_data[10][7] ), .B1(n24697), .B2(
        \xmem_data[11][7] ), .ZN(n10058) );
  AOI22_X1 U14043 ( .A1(n3222), .A2(\xmem_data[8][7] ), .B1(n20805), .B2(
        \xmem_data[9][7] ), .ZN(n10057) );
  NAND3_X1 U14044 ( .A1(n10059), .A2(n10058), .A3(n10057), .ZN(n10060) );
  OR4_X1 U14045 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10064) );
  OAI21_X1 U14046 ( .B1(n10065), .B2(n10064), .A(n20515), .ZN(n10066) );
  XNOR2_X1 U14047 ( .A(n35403), .B(\fmem_data[21][3] ), .ZN(n30413) );
  AOI21_X1 U14048 ( .B1(n34201), .B2(n34199), .A(n30413), .ZN(n10068) );
  INV_X1 U14049 ( .A(n10068), .ZN(n11336) );
  NAND2_X1 U14050 ( .A1(n10069), .A2(n10589), .ZN(n10070) );
  INV_X1 U14051 ( .A(n10070), .ZN(n10071) );
  AOI22_X1 U14052 ( .A1(n37191), .A2(n10071), .B1(n10070), .B2(n4499), .ZN(
        n10162) );
  NAND2_X1 U14053 ( .A1(n37191), .A2(n10071), .ZN(n10072) );
  XOR2_X1 U14054 ( .A(n39040), .B(n10072), .Z(n10161) );
  AND2_X1 U14055 ( .A1(n10162), .A2(n10161), .ZN(n30976) );
  AOI22_X1 U14056 ( .A1(n20725), .A2(\xmem_data[96][5] ), .B1(n27994), .B2(
        \xmem_data[97][5] ), .ZN(n10076) );
  BUF_X1 U14057 ( .A(n14991), .Z(n30942) );
  AOI22_X1 U14058 ( .A1(n3129), .A2(\xmem_data[98][5] ), .B1(n24657), .B2(
        \xmem_data[99][5] ), .ZN(n10075) );
  AOI22_X1 U14059 ( .A1(n27551), .A2(\xmem_data[100][5] ), .B1(n27988), .B2(
        \xmem_data[101][5] ), .ZN(n10074) );
  BUF_X1 U14060 ( .A(n14997), .Z(n30943) );
  AOI22_X1 U14061 ( .A1(n30943), .A2(\xmem_data[102][5] ), .B1(n13168), .B2(
        \xmem_data[103][5] ), .ZN(n10073) );
  NAND4_X1 U14062 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10092) );
  AOI22_X1 U14063 ( .A1(n31268), .A2(\xmem_data[104][5] ), .B1(n14999), .B2(
        \xmem_data[105][5] ), .ZN(n10080) );
  BUF_X1 U14064 ( .A(n29187), .Z(n30948) );
  AOI22_X1 U14065 ( .A1(n28053), .A2(\xmem_data[106][5] ), .B1(n22677), .B2(
        \xmem_data[107][5] ), .ZN(n10079) );
  BUF_X1 U14066 ( .A(n14937), .Z(n30949) );
  AOI22_X1 U14067 ( .A1(n30949), .A2(\xmem_data[108][5] ), .B1(n25398), .B2(
        \xmem_data[109][5] ), .ZN(n10078) );
  BUF_X1 U14068 ( .A(n14971), .Z(n30950) );
  AOI22_X1 U14069 ( .A1(n30950), .A2(\xmem_data[110][5] ), .B1(n28380), .B2(
        \xmem_data[111][5] ), .ZN(n10077) );
  NAND4_X1 U14070 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10091) );
  BUF_X1 U14071 ( .A(n14881), .Z(n30956) );
  BUF_X1 U14072 ( .A(n14973), .Z(n30955) );
  AOI22_X1 U14073 ( .A1(n30956), .A2(\xmem_data[112][5] ), .B1(n30955), .B2(
        \xmem_data[113][5] ), .ZN(n10084) );
  AOI22_X1 U14074 ( .A1(n28226), .A2(\xmem_data[114][5] ), .B1(n28098), .B2(
        \xmem_data[115][5] ), .ZN(n10083) );
  AOI22_X1 U14075 ( .A1(n21058), .A2(\xmem_data[116][5] ), .B1(n28500), .B2(
        \xmem_data[117][5] ), .ZN(n10082) );
  AOI22_X1 U14076 ( .A1(n20567), .A2(\xmem_data[118][5] ), .B1(n29125), .B2(
        \xmem_data[119][5] ), .ZN(n10081) );
  NAND4_X1 U14077 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10090) );
  AOI22_X1 U14078 ( .A1(n31263), .A2(\xmem_data[120][5] ), .B1(n22729), .B2(
        \xmem_data[121][5] ), .ZN(n10088) );
  AOI22_X1 U14079 ( .A1(n3333), .A2(\xmem_data[122][5] ), .B1(n31347), .B2(
        \xmem_data[123][5] ), .ZN(n10087) );
  BUF_X1 U14080 ( .A(n29064), .Z(n30962) );
  AOI22_X1 U14081 ( .A1(n30962), .A2(\xmem_data[124][5] ), .B1(n3218), .B2(
        \xmem_data[125][5] ), .ZN(n10086) );
  BUF_X1 U14082 ( .A(n14988), .Z(n30964) );
  BUF_X1 U14083 ( .A(n14989), .Z(n30963) );
  AOI22_X1 U14084 ( .A1(n30964), .A2(\xmem_data[126][5] ), .B1(n30963), .B2(
        \xmem_data[127][5] ), .ZN(n10085) );
  NAND4_X1 U14085 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10089) );
  OR4_X1 U14086 ( .A1(n10092), .A2(n10091), .A3(n10090), .A4(n10089), .ZN(
        n10114) );
  INV_X1 U14087 ( .A(n10161), .ZN(n10135) );
  NOR2_X1 U14088 ( .A1(n10162), .A2(n10135), .ZN(n30974) );
  BUF_X1 U14089 ( .A(n14926), .Z(n30883) );
  AOI22_X1 U14090 ( .A1(n30883), .A2(\xmem_data[64][5] ), .B1(n30882), .B2(
        \xmem_data[65][5] ), .ZN(n10096) );
  AOI22_X1 U14091 ( .A1(n20962), .A2(\xmem_data[66][5] ), .B1(n29306), .B2(
        \xmem_data[67][5] ), .ZN(n10095) );
  BUF_X1 U14092 ( .A(n10999), .Z(n30884) );
  AOI22_X1 U14093 ( .A1(n30885), .A2(\xmem_data[68][5] ), .B1(n30884), .B2(
        \xmem_data[69][5] ), .ZN(n10094) );
  BUF_X1 U14094 ( .A(n14997), .Z(n30886) );
  AOI22_X1 U14095 ( .A1(n30886), .A2(\xmem_data[70][5] ), .B1(n24639), .B2(
        \xmem_data[71][5] ), .ZN(n10093) );
  NAND4_X1 U14096 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10112) );
  AOI22_X1 U14097 ( .A1(n27537), .A2(\xmem_data[72][5] ), .B1(n30613), .B2(
        \xmem_data[73][5] ), .ZN(n10100) );
  BUF_X1 U14098 ( .A(n29187), .Z(n30892) );
  AOI22_X1 U14099 ( .A1(n25461), .A2(\xmem_data[74][5] ), .B1(n28993), .B2(
        \xmem_data[75][5] ), .ZN(n10099) );
  AOI22_X1 U14100 ( .A1(n28337), .A2(\xmem_data[76][5] ), .B1(n27918), .B2(
        \xmem_data[77][5] ), .ZN(n10098) );
  BUF_X1 U14101 ( .A(n14971), .Z(n30893) );
  AOI22_X1 U14102 ( .A1(n30893), .A2(\xmem_data[78][5] ), .B1(n20941), .B2(
        \xmem_data[79][5] ), .ZN(n10097) );
  NAND4_X1 U14103 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10111) );
  BUF_X1 U14104 ( .A(n3324), .Z(n30899) );
  BUF_X1 U14105 ( .A(n14973), .Z(n30898) );
  AOI22_X1 U14106 ( .A1(n24220), .A2(\xmem_data[80][5] ), .B1(n30898), .B2(
        \xmem_data[81][5] ), .ZN(n10104) );
  AOI22_X1 U14107 ( .A1(n3301), .A2(\xmem_data[82][5] ), .B1(n28098), .B2(
        \xmem_data[83][5] ), .ZN(n10103) );
  AOI22_X1 U14108 ( .A1(n28293), .A2(\xmem_data[84][5] ), .B1(n11008), .B2(
        \xmem_data[85][5] ), .ZN(n10102) );
  BUF_X1 U14109 ( .A(n13457), .Z(n30900) );
  AOI22_X1 U14110 ( .A1(n30901), .A2(\xmem_data[86][5] ), .B1(n30900), .B2(
        \xmem_data[87][5] ), .ZN(n10101) );
  NAND4_X1 U14111 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10110) );
  BUF_X1 U14112 ( .A(n31263), .Z(n30909) );
  BUF_X1 U14113 ( .A(n28974), .Z(n30908) );
  AOI22_X1 U14114 ( .A1(n30909), .A2(\xmem_data[88][5] ), .B1(n30908), .B2(
        \xmem_data[89][5] ), .ZN(n10108) );
  AOI22_X1 U14115 ( .A1(n3350), .A2(\xmem_data[90][5] ), .B1(n27437), .B2(
        \xmem_data[91][5] ), .ZN(n10107) );
  BUF_X1 U14116 ( .A(n29064), .Z(n30906) );
  AOI22_X1 U14117 ( .A1(n30906), .A2(\xmem_data[92][5] ), .B1(n3222), .B2(
        \xmem_data[93][5] ), .ZN(n10106) );
  AOI22_X1 U14118 ( .A1(n31368), .A2(\xmem_data[94][5] ), .B1(n28356), .B2(
        \xmem_data[95][5] ), .ZN(n10105) );
  NAND4_X1 U14119 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10109) );
  OR4_X1 U14120 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10113) );
  AOI22_X1 U14121 ( .A1(n30976), .A2(n10114), .B1(n30974), .B2(n10113), .ZN(
        n10166) );
  AOI22_X1 U14122 ( .A1(n30883), .A2(\xmem_data[32][5] ), .B1(n30882), .B2(
        \xmem_data[33][5] ), .ZN(n10118) );
  AOI22_X1 U14123 ( .A1(n29350), .A2(\xmem_data[34][5] ), .B1(n30877), .B2(
        \xmem_data[35][5] ), .ZN(n10117) );
  AOI22_X1 U14124 ( .A1(n30885), .A2(\xmem_data[36][5] ), .B1(n30884), .B2(
        \xmem_data[37][5] ), .ZN(n10116) );
  AOI22_X1 U14125 ( .A1(n30886), .A2(\xmem_data[38][5] ), .B1(n17012), .B2(
        \xmem_data[39][5] ), .ZN(n10115) );
  NAND4_X1 U14126 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10134) );
  AOI22_X1 U14127 ( .A1(n28980), .A2(\xmem_data[40][5] ), .B1(n22674), .B2(
        \xmem_data[41][5] ), .ZN(n10122) );
  AOI22_X1 U14128 ( .A1(n31354), .A2(\xmem_data[42][5] ), .B1(n27516), .B2(
        \xmem_data[43][5] ), .ZN(n10121) );
  AOI22_X1 U14129 ( .A1(n21007), .A2(\xmem_data[44][5] ), .B1(n29048), .B2(
        \xmem_data[45][5] ), .ZN(n10120) );
  AOI22_X1 U14130 ( .A1(n30893), .A2(\xmem_data[46][5] ), .B1(n30515), .B2(
        \xmem_data[47][5] ), .ZN(n10119) );
  NAND4_X1 U14131 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10133) );
  AOI22_X1 U14132 ( .A1(n24615), .A2(\xmem_data[48][5] ), .B1(n30898), .B2(
        \xmem_data[49][5] ), .ZN(n10126) );
  AOI22_X1 U14133 ( .A1(n3302), .A2(\xmem_data[50][5] ), .B1(n28983), .B2(
        \xmem_data[51][5] ), .ZN(n10125) );
  AOI22_X1 U14134 ( .A1(n27847), .A2(\xmem_data[52][5] ), .B1(n22751), .B2(
        \xmem_data[53][5] ), .ZN(n10124) );
  AOI22_X1 U14135 ( .A1(n30901), .A2(\xmem_data[54][5] ), .B1(n30900), .B2(
        \xmem_data[55][5] ), .ZN(n10123) );
  NAND4_X1 U14136 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10132) );
  AOI22_X1 U14137 ( .A1(n30909), .A2(\xmem_data[56][5] ), .B1(n30908), .B2(
        \xmem_data[57][5] ), .ZN(n10130) );
  AOI22_X1 U14138 ( .A1(n3351), .A2(\xmem_data[58][5] ), .B1(n25360), .B2(
        \xmem_data[59][5] ), .ZN(n10129) );
  AOI22_X1 U14139 ( .A1(n30906), .A2(\xmem_data[60][5] ), .B1(n3220), .B2(
        \xmem_data[61][5] ), .ZN(n10128) );
  AOI22_X1 U14140 ( .A1(n29256), .A2(\xmem_data[62][5] ), .B1(n24695), .B2(
        \xmem_data[63][5] ), .ZN(n10127) );
  NAND4_X1 U14141 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10131) );
  OR4_X1 U14142 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10136) );
  NAND2_X1 U14143 ( .A1(n10136), .A2(n30918), .ZN(n10165) );
  AOI22_X1 U14144 ( .A1(n23756), .A2(\xmem_data[28][5] ), .B1(n3220), .B2(
        \xmem_data[29][5] ), .ZN(n10148) );
  AOI22_X1 U14145 ( .A1(n13436), .A2(\xmem_data[8][5] ), .B1(n25671), .B2(
        \xmem_data[9][5] ), .ZN(n10140) );
  AOI22_X1 U14146 ( .A1(n27455), .A2(\xmem_data[10][5] ), .B1(n3208), .B2(
        \xmem_data[11][5] ), .ZN(n10139) );
  AOI22_X1 U14147 ( .A1(n14937), .A2(\xmem_data[12][5] ), .B1(n20940), .B2(
        \xmem_data[13][5] ), .ZN(n10138) );
  BUF_X1 U14148 ( .A(n14971), .Z(n30872) );
  BUF_X1 U14149 ( .A(n13481), .Z(n30871) );
  AOI22_X1 U14150 ( .A1(n30872), .A2(\xmem_data[14][5] ), .B1(n30871), .B2(
        \xmem_data[15][5] ), .ZN(n10137) );
  AOI22_X1 U14151 ( .A1(n28367), .A2(\xmem_data[30][5] ), .B1(n20723), .B2(
        \xmem_data[31][5] ), .ZN(n10141) );
  INV_X1 U14152 ( .A(n10141), .ZN(n10144) );
  BUF_X1 U14153 ( .A(n28973), .Z(n30864) );
  BUF_X1 U14154 ( .A(n13468), .Z(n30863) );
  AOI22_X1 U14155 ( .A1(n30864), .A2(\xmem_data[26][5] ), .B1(n30863), .B2(
        \xmem_data[27][5] ), .ZN(n10142) );
  INV_X1 U14156 ( .A(n10142), .ZN(n10143) );
  NOR2_X1 U14157 ( .A1(n10144), .A2(n10143), .ZN(n10146) );
  BUF_X1 U14158 ( .A(n31263), .Z(n30862) );
  BUF_X1 U14159 ( .A(n28947), .Z(n30861) );
  AOI22_X1 U14160 ( .A1(n30862), .A2(\xmem_data[24][5] ), .B1(n30861), .B2(
        \xmem_data[25][5] ), .ZN(n10145) );
  NAND4_X1 U14161 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10160) );
  BUF_X1 U14162 ( .A(n14972), .Z(n30849) );
  AOI22_X1 U14163 ( .A1(n30849), .A2(\xmem_data[16][5] ), .B1(n28327), .B2(
        \xmem_data[17][5] ), .ZN(n10152) );
  AOI22_X1 U14164 ( .A1(n23724), .A2(\xmem_data[18][5] ), .B1(n14975), .B2(
        \xmem_data[19][5] ), .ZN(n10151) );
  AOI22_X1 U14165 ( .A1(n22684), .A2(\xmem_data[20][5] ), .B1(n29136), .B2(
        \xmem_data[21][5] ), .ZN(n10150) );
  AOI22_X1 U14166 ( .A1(n21060), .A2(\xmem_data[22][5] ), .B1(n28035), .B2(
        \xmem_data[23][5] ), .ZN(n10149) );
  NAND4_X1 U14167 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10159) );
  BUF_X1 U14168 ( .A(n14928), .Z(n30877) );
  NAND2_X1 U14169 ( .A1(n25450), .A2(\xmem_data[3][5] ), .ZN(n10153) );
  AOI22_X1 U14170 ( .A1(n25457), .A2(\xmem_data[6][5] ), .B1(n24212), .B2(
        \xmem_data[7][5] ), .ZN(n10156) );
  AOI22_X1 U14171 ( .A1(n23813), .A2(\xmem_data[4][5] ), .B1(n30854), .B2(
        \xmem_data[5][5] ), .ZN(n10155) );
  AOI22_X1 U14172 ( .A1(n29174), .A2(\xmem_data[0][5] ), .B1(n20993), .B2(
        \xmem_data[1][5] ), .ZN(n10154) );
  NAND3_X1 U14173 ( .A1(n10156), .A2(n10155), .A3(n10154), .ZN(n10157) );
  NOR2_X1 U14174 ( .A1(n10162), .A2(n10161), .ZN(n10213) );
  NAND2_X1 U14175 ( .A1(n10163), .A2(n10213), .ZN(n10164) );
  XOR2_X1 U14176 ( .A(\fmem_data[10][4] ), .B(\fmem_data[10][5] ), .Z(n10167)
         );
  AOI22_X1 U14177 ( .A1(n30883), .A2(\xmem_data[32][6] ), .B1(n30882), .B2(
        \xmem_data[33][6] ), .ZN(n10171) );
  AOI22_X1 U14178 ( .A1(n3345), .A2(\xmem_data[34][6] ), .B1(n25514), .B2(
        \xmem_data[35][6] ), .ZN(n10170) );
  AOI22_X1 U14179 ( .A1(n30885), .A2(\xmem_data[36][6] ), .B1(n30884), .B2(
        \xmem_data[37][6] ), .ZN(n10169) );
  AOI22_X1 U14180 ( .A1(n30886), .A2(\xmem_data[38][6] ), .B1(n22675), .B2(
        \xmem_data[39][6] ), .ZN(n10168) );
  NAND4_X1 U14181 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10187) );
  AOI22_X1 U14182 ( .A1(n29023), .A2(\xmem_data[40][6] ), .B1(n14999), .B2(
        \xmem_data[41][6] ), .ZN(n10175) );
  AOI22_X1 U14183 ( .A1(n29396), .A2(\xmem_data[42][6] ), .B1(n20938), .B2(
        \xmem_data[43][6] ), .ZN(n10174) );
  AOI22_X1 U14184 ( .A1(n24547), .A2(\xmem_data[44][6] ), .B1(n31270), .B2(
        \xmem_data[45][6] ), .ZN(n10173) );
  AOI22_X1 U14185 ( .A1(n30893), .A2(\xmem_data[46][6] ), .B1(n25435), .B2(
        \xmem_data[47][6] ), .ZN(n10172) );
  NAND4_X1 U14186 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10186) );
  AOI22_X1 U14187 ( .A1(n28460), .A2(\xmem_data[48][6] ), .B1(n30898), .B2(
        \xmem_data[49][6] ), .ZN(n10179) );
  AOI22_X1 U14188 ( .A1(n3302), .A2(\xmem_data[50][6] ), .B1(n24622), .B2(
        \xmem_data[51][6] ), .ZN(n10178) );
  AOI22_X1 U14189 ( .A1(n24685), .A2(\xmem_data[52][6] ), .B1(n21057), .B2(
        \xmem_data[53][6] ), .ZN(n10177) );
  AOI22_X1 U14190 ( .A1(n30901), .A2(\xmem_data[54][6] ), .B1(n30900), .B2(
        \xmem_data[55][6] ), .ZN(n10176) );
  NAND4_X1 U14191 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10185) );
  AOI22_X1 U14192 ( .A1(n30909), .A2(\xmem_data[56][6] ), .B1(n30908), .B2(
        \xmem_data[57][6] ), .ZN(n10183) );
  AOI22_X1 U14193 ( .A1(n3352), .A2(\xmem_data[58][6] ), .B1(n30863), .B2(
        \xmem_data[59][6] ), .ZN(n10182) );
  AOI22_X1 U14194 ( .A1(n30906), .A2(\xmem_data[60][6] ), .B1(n3218), .B2(
        \xmem_data[61][6] ), .ZN(n10181) );
  AOI22_X1 U14195 ( .A1(n29789), .A2(\xmem_data[62][6] ), .B1(n28356), .B2(
        \xmem_data[63][6] ), .ZN(n10180) );
  NAND4_X1 U14196 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10184) );
  OR4_X1 U14197 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10216) );
  AOI22_X1 U14198 ( .A1(n30862), .A2(\xmem_data[24][6] ), .B1(n30861), .B2(
        \xmem_data[25][6] ), .ZN(n10191) );
  AOI22_X1 U14199 ( .A1(n30864), .A2(\xmem_data[26][6] ), .B1(n30863), .B2(
        \xmem_data[27][6] ), .ZN(n10190) );
  AOI22_X1 U14200 ( .A1(n23734), .A2(\xmem_data[28][6] ), .B1(n3217), .B2(
        \xmem_data[29][6] ), .ZN(n10189) );
  AOI22_X1 U14201 ( .A1(n25693), .A2(\xmem_data[30][6] ), .B1(n29095), .B2(
        \xmem_data[31][6] ), .ZN(n10188) );
  AOI22_X1 U14202 ( .A1(n29310), .A2(\xmem_data[8][6] ), .B1(n28052), .B2(
        \xmem_data[9][6] ), .ZN(n10195) );
  AOI22_X1 U14203 ( .A1(n28154), .A2(\xmem_data[10][6] ), .B1(n20586), .B2(
        \xmem_data[11][6] ), .ZN(n10194) );
  AOI22_X1 U14204 ( .A1(n25434), .A2(\xmem_data[12][6] ), .B1(n31355), .B2(
        \xmem_data[13][6] ), .ZN(n10193) );
  AOI22_X1 U14205 ( .A1(n30872), .A2(\xmem_data[14][6] ), .B1(n30871), .B2(
        \xmem_data[15][6] ), .ZN(n10192) );
  NAND4_X1 U14206 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10212) );
  AOI22_X1 U14207 ( .A1(n3341), .A2(\xmem_data[0][6] ), .B1(n22759), .B2(
        \xmem_data[1][6] ), .ZN(n10196) );
  INV_X1 U14208 ( .A(n10196), .ZN(n10200) );
  AOI22_X1 U14209 ( .A1(n23813), .A2(\xmem_data[4][6] ), .B1(n30854), .B2(
        \xmem_data[5][6] ), .ZN(n10198) );
  NAND2_X1 U14210 ( .A1(n3374), .A2(\xmem_data[2][6] ), .ZN(n10197) );
  NAND2_X1 U14211 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  AOI22_X1 U14212 ( .A1(n14982), .A2(\xmem_data[22][6] ), .B1(n27435), .B2(
        \xmem_data[23][6] ), .ZN(n10210) );
  AOI22_X1 U14213 ( .A1(n30849), .A2(\xmem_data[16][6] ), .B1(n23778), .B2(
        \xmem_data[17][6] ), .ZN(n10201) );
  INV_X1 U14214 ( .A(n10201), .ZN(n10208) );
  AOI22_X1 U14215 ( .A1(n20545), .A2(\xmem_data[6][6] ), .B1(n28345), .B2(
        \xmem_data[7][6] ), .ZN(n10202) );
  INV_X1 U14216 ( .A(n10202), .ZN(n10207) );
  AOI22_X1 U14217 ( .A1(n30525), .A2(\xmem_data[20][6] ), .B1(n31256), .B2(
        \xmem_data[21][6] ), .ZN(n10205) );
  AOI22_X1 U14218 ( .A1(n21056), .A2(\xmem_data[18][6] ), .B1(n14975), .B2(
        \xmem_data[19][6] ), .ZN(n10204) );
  NAND2_X1 U14219 ( .A1(n31252), .A2(\xmem_data[3][6] ), .ZN(n10203) );
  NOR3_X1 U14220 ( .A1(n10208), .A2(n10207), .A3(n10206), .ZN(n10209) );
  NAND2_X1 U14221 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  NOR3_X1 U14222 ( .A1(n10212), .A2(n3986), .A3(n10211), .ZN(n10214) );
  INV_X1 U14223 ( .A(n10213), .ZN(n30879) );
  AOI21_X1 U14224 ( .B1(n3748), .B2(n10214), .A(n30879), .ZN(n10215) );
  AOI21_X1 U14225 ( .B1(n10216), .B2(n30918), .A(n10215), .ZN(n10260) );
  AOI22_X1 U14226 ( .A1(n3342), .A2(\xmem_data[96][6] ), .B1(n28342), .B2(
        \xmem_data[97][6] ), .ZN(n10220) );
  AOI22_X1 U14227 ( .A1(n3128), .A2(\xmem_data[98][6] ), .B1(n28343), .B2(
        \xmem_data[99][6] ), .ZN(n10219) );
  AOI22_X1 U14228 ( .A1(n27551), .A2(\xmem_data[100][6] ), .B1(n3357), .B2(
        \xmem_data[101][6] ), .ZN(n10218) );
  AOI22_X1 U14229 ( .A1(n30943), .A2(\xmem_data[102][6] ), .B1(n13168), .B2(
        \xmem_data[103][6] ), .ZN(n10217) );
  NAND4_X1 U14230 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10236) );
  AOI22_X1 U14231 ( .A1(n16986), .A2(\xmem_data[104][6] ), .B1(n22674), .B2(
        \xmem_data[105][6] ), .ZN(n10224) );
  AOI22_X1 U14232 ( .A1(n25519), .A2(\xmem_data[106][6] ), .B1(n25574), .B2(
        \xmem_data[107][6] ), .ZN(n10223) );
  AOI22_X1 U14233 ( .A1(n30949), .A2(\xmem_data[108][6] ), .B1(n23796), .B2(
        \xmem_data[109][6] ), .ZN(n10222) );
  AOI22_X1 U14234 ( .A1(n30950), .A2(\xmem_data[110][6] ), .B1(n29238), .B2(
        \xmem_data[111][6] ), .ZN(n10221) );
  NAND4_X1 U14235 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(
        n10235) );
  AOI22_X1 U14236 ( .A1(n30956), .A2(\xmem_data[112][6] ), .B1(n30955), .B2(
        \xmem_data[113][6] ), .ZN(n10228) );
  AOI22_X1 U14237 ( .A1(n24623), .A2(\xmem_data[114][6] ), .B1(n20553), .B2(
        \xmem_data[115][6] ), .ZN(n10227) );
  AOI22_X1 U14238 ( .A1(n3171), .A2(\xmem_data[116][6] ), .B1(n25406), .B2(
        \xmem_data[117][6] ), .ZN(n10226) );
  AOI22_X1 U14239 ( .A1(n28192), .A2(\xmem_data[118][6] ), .B1(n21059), .B2(
        \xmem_data[119][6] ), .ZN(n10225) );
  NAND4_X1 U14240 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(
        n10234) );
  AOI22_X1 U14241 ( .A1(n3380), .A2(\xmem_data[120][6] ), .B1(n25357), .B2(
        \xmem_data[121][6] ), .ZN(n10232) );
  AOI22_X1 U14242 ( .A1(n3333), .A2(\xmem_data[122][6] ), .B1(n14875), .B2(
        \xmem_data[123][6] ), .ZN(n10231) );
  AOI22_X1 U14243 ( .A1(n30962), .A2(\xmem_data[124][6] ), .B1(n3218), .B2(
        \xmem_data[125][6] ), .ZN(n10230) );
  AOI22_X1 U14244 ( .A1(n30964), .A2(\xmem_data[126][6] ), .B1(n30963), .B2(
        \xmem_data[127][6] ), .ZN(n10229) );
  NAND4_X1 U14245 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10233) );
  OR4_X1 U14246 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10258) );
  AOI22_X1 U14247 ( .A1(n30883), .A2(\xmem_data[64][6] ), .B1(n30882), .B2(
        \xmem_data[65][6] ), .ZN(n10240) );
  AOI22_X1 U14248 ( .A1(n28084), .A2(n20682), .B1(n24553), .B2(
        \xmem_data[67][6] ), .ZN(n10239) );
  AOI22_X1 U14249 ( .A1(n30885), .A2(\xmem_data[68][6] ), .B1(n30884), .B2(
        \xmem_data[69][6] ), .ZN(n10238) );
  AOI22_X1 U14250 ( .A1(n30886), .A2(\xmem_data[70][6] ), .B1(n27535), .B2(
        \xmem_data[71][6] ), .ZN(n10237) );
  NAND4_X1 U14251 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10256) );
  AOI22_X1 U14252 ( .A1(n20495), .A2(\xmem_data[72][6] ), .B1(n27912), .B2(
        \xmem_data[73][6] ), .ZN(n10244) );
  AOI22_X1 U14253 ( .A1(n29396), .A2(\xmem_data[74][6] ), .B1(n25383), .B2(
        \xmem_data[75][6] ), .ZN(n10243) );
  AOI22_X1 U14254 ( .A1(n27919), .A2(\xmem_data[76][6] ), .B1(n24707), .B2(
        \xmem_data[77][6] ), .ZN(n10242) );
  AOI22_X1 U14255 ( .A1(n30893), .A2(\xmem_data[78][6] ), .B1(n28380), .B2(
        \xmem_data[79][6] ), .ZN(n10241) );
  NAND4_X1 U14256 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10255) );
  AOI22_X1 U14257 ( .A1(n3326), .A2(\xmem_data[80][6] ), .B1(n30898), .B2(
        \xmem_data[81][6] ), .ZN(n10248) );
  AOI22_X1 U14258 ( .A1(n3301), .A2(\xmem_data[82][6] ), .B1(n28098), .B2(
        \xmem_data[83][6] ), .ZN(n10247) );
  AOI22_X1 U14259 ( .A1(n25526), .A2(\xmem_data[84][6] ), .B1(n11008), .B2(
        \xmem_data[85][6] ), .ZN(n10246) );
  AOI22_X1 U14260 ( .A1(n30901), .A2(\xmem_data[86][6] ), .B1(n30900), .B2(
        \xmem_data[87][6] ), .ZN(n10245) );
  NAND4_X1 U14261 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10254) );
  AOI22_X1 U14262 ( .A1(n30906), .A2(\xmem_data[92][6] ), .B1(n3222), .B2(
        \xmem_data[93][6] ), .ZN(n10252) );
  AOI22_X1 U14263 ( .A1(n3352), .A2(\xmem_data[90][6] ), .B1(n31347), .B2(
        \xmem_data[91][6] ), .ZN(n10251) );
  AOI22_X1 U14264 ( .A1(n30909), .A2(\xmem_data[88][6] ), .B1(n30908), .B2(
        \xmem_data[89][6] ), .ZN(n10250) );
  AOI22_X1 U14265 ( .A1(n30964), .A2(\xmem_data[94][6] ), .B1(n20558), .B2(
        \xmem_data[95][6] ), .ZN(n10249) );
  NAND4_X1 U14266 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10253) );
  OR4_X1 U14267 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10257) );
  AOI22_X1 U14268 ( .A1(n30976), .A2(n10258), .B1(n30974), .B2(n10257), .ZN(
        n10259) );
  AOI22_X1 U14269 ( .A1(n14997), .A2(\xmem_data[20][7] ), .B1(n13168), .B2(
        \xmem_data[21][7] ), .ZN(n10261) );
  INV_X1 U14270 ( .A(n10261), .ZN(n10268) );
  BUF_X1 U14271 ( .A(n10999), .Z(n24590) );
  AOI22_X1 U14272 ( .A1(n25422), .A2(\xmem_data[18][7] ), .B1(n24590), .B2(
        \xmem_data[19][7] ), .ZN(n10263) );
  NAND2_X1 U14273 ( .A1(n3374), .A2(\xmem_data[16][7] ), .ZN(n10262) );
  NAND2_X1 U14274 ( .A1(n10263), .A2(n10262), .ZN(n10267) );
  BUF_X1 U14275 ( .A(n14898), .Z(n24597) );
  NAND2_X1 U14276 ( .A1(n10265), .A2(n10264), .ZN(n10266) );
  OR3_X1 U14277 ( .A1(n10268), .A2(n10267), .A3(n10266), .ZN(n10274) );
  AOI22_X1 U14278 ( .A1(n28231), .A2(\xmem_data[24][7] ), .B1(n20543), .B2(
        \xmem_data[25][7] ), .ZN(n10272) );
  BUF_X1 U14279 ( .A(n14937), .Z(n24593) );
  AOI22_X1 U14280 ( .A1(n24593), .A2(\xmem_data[26][7] ), .B1(n29048), .B2(
        \xmem_data[27][7] ), .ZN(n10271) );
  BUF_X1 U14281 ( .A(n14913), .Z(n24592) );
  AOI22_X1 U14282 ( .A1(n16990), .A2(\xmem_data[28][7] ), .B1(n24592), .B2(
        \xmem_data[29][7] ), .ZN(n10270) );
  BUF_X1 U14283 ( .A(n3324), .Z(n24615) );
  AOI22_X1 U14284 ( .A1(n24615), .A2(\xmem_data[30][7] ), .B1(n31361), .B2(
        \xmem_data[31][7] ), .ZN(n10269) );
  NAND4_X1 U14285 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  OR2_X1 U14286 ( .A1(n10274), .A2(n10273), .ZN(n10281) );
  AOI22_X1 U14287 ( .A1(n28718), .A2(\xmem_data[8][7] ), .B1(n3247), .B2(
        \xmem_data[9][7] ), .ZN(n10279) );
  AND2_X1 U14288 ( .A1(n3219), .A2(\xmem_data[11][7] ), .ZN(n10275) );
  AOI21_X1 U14289 ( .B1(n24631), .B2(\xmem_data[10][7] ), .A(n10275), .ZN(
        n10278) );
  AOI22_X1 U14290 ( .A1(n29627), .A2(\xmem_data[12][7] ), .B1(n25509), .B2(
        \xmem_data[13][7] ), .ZN(n10277) );
  AOI22_X1 U14291 ( .A1(n23741), .A2(\xmem_data[14][7] ), .B1(n27903), .B2(
        \xmem_data[15][7] ), .ZN(n10276) );
  NAND4_X1 U14292 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  NOR2_X1 U14293 ( .A1(n10281), .A2(n10280), .ZN(n10290) );
  AOI22_X1 U14294 ( .A1(n29573), .A2(\xmem_data[0][7] ), .B1(n22685), .B2(
        \xmem_data[1][7] ), .ZN(n10285) );
  BUF_X1 U14295 ( .A(n13486), .Z(n24606) );
  AOI22_X1 U14296 ( .A1(n24606), .A2(\xmem_data[2][7] ), .B1(n28468), .B2(
        \xmem_data[3][7] ), .ZN(n10284) );
  AOI22_X1 U14297 ( .A1(n28772), .A2(\xmem_data[4][7] ), .B1(n24686), .B2(
        \xmem_data[5][7] ), .ZN(n10283) );
  BUF_X1 U14298 ( .A(n31263), .Z(n24607) );
  AOI22_X1 U14299 ( .A1(n24607), .A2(\xmem_data[6][7] ), .B1(n27563), .B2(
        \xmem_data[7][7] ), .ZN(n10282) );
  NAND4_X1 U14300 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  BUF_X1 U14301 ( .A(n14928), .Z(n24657) );
  NOR2_X1 U14302 ( .A1(n10286), .A2(n3873), .ZN(n10289) );
  OAI21_X1 U14303 ( .B1(load_xaddr_val[5]), .B2(n37190), .A(n10287), .ZN(
        n10356) );
  AOI22_X1 U14304 ( .A1(n37190), .A2(n39040), .B1(n14909), .B2(n10288), .ZN(
        n10333) );
  NOR2_X1 U14305 ( .A1(n10356), .A2(n10333), .ZN(n21278) );
  AOI21_X1 U14306 ( .B1(n10290), .B2(n10289), .A(n24662), .ZN(n10291) );
  INV_X1 U14307 ( .A(n10291), .ZN(n10362) );
  BUF_X1 U14308 ( .A(n28973), .Z(n24630) );
  AOI22_X1 U14309 ( .A1(n24630), .A2(\xmem_data[72][7] ), .B1(n3247), .B2(
        \xmem_data[73][7] ), .ZN(n10295) );
  BUF_X1 U14310 ( .A(n29064), .Z(n24631) );
  AOI22_X1 U14311 ( .A1(n24631), .A2(\xmem_data[74][7] ), .B1(n3222), .B2(
        \xmem_data[75][7] ), .ZN(n10294) );
  BUF_X1 U14312 ( .A(n14988), .Z(n24632) );
  AOI22_X1 U14313 ( .A1(n24632), .A2(\xmem_data[76][7] ), .B1(n27444), .B2(
        \xmem_data[77][7] ), .ZN(n10293) );
  BUF_X1 U14314 ( .A(n14890), .Z(n24633) );
  AOI22_X1 U14315 ( .A1(n3342), .A2(\xmem_data[78][7] ), .B1(n24633), .B2(
        \xmem_data[79][7] ), .ZN(n10292) );
  NAND4_X1 U14316 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10311) );
  BUF_X1 U14317 ( .A(n14974), .Z(n24623) );
  AOI22_X1 U14318 ( .A1(n24623), .A2(\xmem_data[64][7] ), .B1(n24622), .B2(
        \xmem_data[65][7] ), .ZN(n10299) );
  AOI22_X1 U14319 ( .A1(n29325), .A2(\xmem_data[66][7] ), .B1(n28468), .B2(
        \xmem_data[67][7] ), .ZN(n10298) );
  BUF_X1 U14320 ( .A(n10456), .Z(n24624) );
  AOI22_X1 U14321 ( .A1(n29298), .A2(\xmem_data[68][7] ), .B1(n24624), .B2(
        \xmem_data[69][7] ), .ZN(n10297) );
  BUF_X1 U14322 ( .A(n28974), .Z(n24625) );
  AOI22_X1 U14323 ( .A1(n20953), .A2(\xmem_data[70][7] ), .B1(n3203), .B2(
        \xmem_data[71][7] ), .ZN(n10296) );
  NAND4_X1 U14324 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10310) );
  AOI22_X1 U14325 ( .A1(n3281), .A2(\xmem_data[80][7] ), .B1(n28343), .B2(
        \xmem_data[81][7] ), .ZN(n10303) );
  BUF_X1 U14326 ( .A(n4478), .Z(n24638) );
  AOI22_X1 U14327 ( .A1(n24638), .A2(\xmem_data[82][7] ), .B1(n27943), .B2(
        \xmem_data[83][7] ), .ZN(n10302) );
  BUF_X1 U14328 ( .A(n14997), .Z(n24640) );
  BUF_X1 U14329 ( .A(n13435), .Z(n24639) );
  AOI22_X1 U14330 ( .A1(n24640), .A2(\xmem_data[84][7] ), .B1(n24639), .B2(
        \xmem_data[85][7] ), .ZN(n10301) );
  AOI22_X1 U14331 ( .A1(n25425), .A2(\xmem_data[86][7] ), .B1(n30613), .B2(
        \xmem_data[87][7] ), .ZN(n10300) );
  NAND4_X1 U14332 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10309) );
  AOI22_X1 U14333 ( .A1(n20718), .A2(\xmem_data[88][7] ), .B1(n23716), .B2(
        \xmem_data[89][7] ), .ZN(n10307) );
  BUF_X1 U14334 ( .A(n14912), .Z(n24645) );
  AOI22_X1 U14335 ( .A1(n23717), .A2(\xmem_data[90][7] ), .B1(n24645), .B2(
        \xmem_data[91][7] ), .ZN(n10306) );
  BUF_X1 U14336 ( .A(n13452), .Z(n24646) );
  AOI22_X1 U14337 ( .A1(n20942), .A2(\xmem_data[92][7] ), .B1(n24646), .B2(
        \xmem_data[93][7] ), .ZN(n10305) );
  BUF_X2 U14338 ( .A(n14881), .Z(n24647) );
  AOI22_X1 U14339 ( .A1(n24647), .A2(\xmem_data[94][7] ), .B1(n25679), .B2(
        \xmem_data[95][7] ), .ZN(n10304) );
  NAND4_X1 U14340 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  OR4_X1 U14341 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  INV_X1 U14342 ( .A(n10333), .ZN(n10357) );
  NOR2_X1 U14343 ( .A1(n10356), .A2(n10357), .ZN(n24720) );
  NAND2_X1 U14344 ( .A1(n10312), .A2(n24720), .ZN(n10361) );
  BUF_X1 U14345 ( .A(n28973), .Z(n24693) );
  AOI22_X1 U14346 ( .A1(n24693), .A2(\xmem_data[104][7] ), .B1(n3247), .B2(
        \xmem_data[105][7] ), .ZN(n10316) );
  BUF_X1 U14347 ( .A(n29064), .Z(n24694) );
  AOI22_X1 U14348 ( .A1(n24694), .A2(\xmem_data[106][7] ), .B1(n3222), .B2(
        \xmem_data[107][7] ), .ZN(n10315) );
  BUF_X1 U14349 ( .A(n14988), .Z(n24696) );
  AOI22_X1 U14350 ( .A1(n24696), .A2(\xmem_data[108][7] ), .B1(n24695), .B2(
        \xmem_data[109][7] ), .ZN(n10314) );
  AOI22_X1 U14351 ( .A1(n24697), .A2(\xmem_data[110][7] ), .B1(n25616), .B2(
        \xmem_data[111][7] ), .ZN(n10313) );
  NAND4_X1 U14352 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10332) );
  AOI22_X1 U14353 ( .A1(n25636), .A2(\xmem_data[96][7] ), .B1(n24622), .B2(
        \xmem_data[97][7] ), .ZN(n10320) );
  AOI22_X1 U14354 ( .A1(n24685), .A2(\xmem_data[98][7] ), .B1(n25359), .B2(
        \xmem_data[99][7] ), .ZN(n10319) );
  BUF_X1 U14355 ( .A(n13127), .Z(n24687) );
  BUF_X1 U14356 ( .A(n13487), .Z(n24686) );
  AOI22_X1 U14357 ( .A1(n24687), .A2(\xmem_data[100][7] ), .B1(n24686), .B2(
        \xmem_data[101][7] ), .ZN(n10318) );
  BUF_X1 U14358 ( .A(n31263), .Z(n24688) );
  AOI22_X1 U14359 ( .A1(n24688), .A2(\xmem_data[102][7] ), .B1(n30908), .B2(
        \xmem_data[103][7] ), .ZN(n10317) );
  NAND4_X1 U14360 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10331) );
  BUF_X1 U14361 ( .A(n14991), .Z(n24702) );
  AOI22_X1 U14362 ( .A1(n24702), .A2(\xmem_data[112][7] ), .B1(n29103), .B2(
        \xmem_data[113][7] ), .ZN(n10324) );
  AOI22_X1 U14363 ( .A1(n25422), .A2(\xmem_data[114][7] ), .B1(n3357), .B2(
        \xmem_data[115][7] ), .ZN(n10323) );
  AOI22_X1 U14364 ( .A1(n27944), .A2(\xmem_data[116][7] ), .B1(n13168), .B2(
        \xmem_data[117][7] ), .ZN(n10322) );
  AOI22_X1 U14365 ( .A1(n28298), .A2(\xmem_data[118][7] ), .B1(n27536), .B2(
        \xmem_data[119][7] ), .ZN(n10321) );
  NAND4_X1 U14366 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10330) );
  AOI22_X1 U14367 ( .A1(n27455), .A2(\xmem_data[120][7] ), .B1(n24457), .B2(
        \xmem_data[121][7] ), .ZN(n10328) );
  BUF_X1 U14368 ( .A(n14937), .Z(n24708) );
  BUF_X1 U14369 ( .A(n14912), .Z(n24707) );
  AOI22_X1 U14370 ( .A1(n24708), .A2(\xmem_data[122][7] ), .B1(n24707), .B2(
        \xmem_data[123][7] ), .ZN(n10327) );
  BUF_X1 U14371 ( .A(n14971), .Z(n24710) );
  BUF_X1 U14372 ( .A(n13452), .Z(n24709) );
  AOI22_X1 U14373 ( .A1(n24710), .A2(\xmem_data[124][7] ), .B1(n24709), .B2(
        \xmem_data[125][7] ), .ZN(n10326) );
  AOI22_X1 U14374 ( .A1(n3206), .A2(\xmem_data[126][7] ), .B1(n24117), .B2(
        \xmem_data[127][7] ), .ZN(n10325) );
  NAND4_X1 U14375 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  OR4_X1 U14376 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10334) );
  AND2_X1 U14377 ( .A1(n10356), .A2(n10333), .ZN(n24722) );
  NAND2_X1 U14378 ( .A1(n10334), .A2(n24722), .ZN(n10360) );
  AOI22_X1 U14379 ( .A1(n24630), .A2(\xmem_data[40][7] ), .B1(n3247), .B2(
        \xmem_data[41][7] ), .ZN(n10339) );
  AND2_X1 U14380 ( .A1(n3222), .A2(\xmem_data[43][7] ), .ZN(n10335) );
  AOI21_X1 U14381 ( .B1(n24631), .B2(\xmem_data[42][7] ), .A(n10335), .ZN(
        n10338) );
  AOI22_X1 U14382 ( .A1(n24632), .A2(\xmem_data[44][7] ), .B1(n22710), .B2(
        \xmem_data[45][7] ), .ZN(n10337) );
  AOI22_X1 U14383 ( .A1(n3322), .A2(\xmem_data[46][7] ), .B1(n24633), .B2(
        \xmem_data[47][7] ), .ZN(n10336) );
  NAND4_X1 U14384 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10355) );
  AOI22_X1 U14385 ( .A1(n24623), .A2(\xmem_data[32][7] ), .B1(n24622), .B2(
        \xmem_data[33][7] ), .ZN(n10343) );
  AOI22_X1 U14386 ( .A1(n31316), .A2(\xmem_data[34][7] ), .B1(n17049), .B2(
        \xmem_data[35][7] ), .ZN(n10342) );
  AOI22_X1 U14387 ( .A1(n29298), .A2(\xmem_data[36][7] ), .B1(n24624), .B2(
        \xmem_data[37][7] ), .ZN(n10341) );
  AOI22_X1 U14388 ( .A1(n25441), .A2(\xmem_data[38][7] ), .B1(n3203), .B2(
        \xmem_data[39][7] ), .ZN(n10340) );
  NAND4_X1 U14389 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10354) );
  AOI22_X1 U14390 ( .A1(n3281), .A2(\xmem_data[48][7] ), .B1(n30877), .B2(
        \xmem_data[49][7] ), .ZN(n10347) );
  AOI22_X1 U14391 ( .A1(n24638), .A2(\xmem_data[50][7] ), .B1(n3357), .B2(
        \xmem_data[51][7] ), .ZN(n10346) );
  AOI22_X1 U14392 ( .A1(n24640), .A2(\xmem_data[52][7] ), .B1(n24639), .B2(
        \xmem_data[53][7] ), .ZN(n10345) );
  AOI22_X1 U14393 ( .A1(n17041), .A2(\xmem_data[54][7] ), .B1(n20717), .B2(
        \xmem_data[55][7] ), .ZN(n10344) );
  NAND4_X1 U14394 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10353) );
  AOI22_X1 U14395 ( .A1(n29008), .A2(\xmem_data[56][7] ), .B1(n30615), .B2(
        \xmem_data[57][7] ), .ZN(n10351) );
  AOI22_X1 U14396 ( .A1(n24133), .A2(\xmem_data[58][7] ), .B1(n24645), .B2(
        \xmem_data[59][7] ), .ZN(n10350) );
  AOI22_X1 U14397 ( .A1(n21050), .A2(\xmem_data[60][7] ), .B1(n24646), .B2(
        \xmem_data[61][7] ), .ZN(n10349) );
  AOI22_X1 U14398 ( .A1(n24647), .A2(\xmem_data[62][7] ), .B1(n23778), .B2(
        \xmem_data[63][7] ), .ZN(n10348) );
  NAND4_X1 U14399 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  OR4_X1 U14400 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10358) );
  AND2_X1 U14401 ( .A1(n10357), .A2(n10356), .ZN(n24659) );
  NAND2_X1 U14402 ( .A1(n10358), .A2(n24659), .ZN(n10359) );
  NAND4_X1 U14403 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n35395) );
  XNOR2_X1 U14404 ( .A(n35395), .B(\fmem_data[24][3] ), .ZN(n30471) );
  XOR2_X1 U14405 ( .A(\fmem_data[24][3] ), .B(\fmem_data[24][2] ), .Z(n10363)
         );
  AND2_X1 U14406 ( .A1(n34433), .A2(n34431), .ZN(n10364) );
  BUF_X1 U14407 ( .A(n3464), .Z(n20939) );
  BUF_X1 U14408 ( .A(n13188), .Z(n20938) );
  AOI22_X1 U14409 ( .A1(n20939), .A2(\xmem_data[64][5] ), .B1(n20938), .B2(
        \xmem_data[65][5] ), .ZN(n10368) );
  BUF_X1 U14410 ( .A(n13415), .Z(n20940) );
  AOI22_X1 U14411 ( .A1(n23764), .A2(\xmem_data[66][5] ), .B1(n20940), .B2(
        \xmem_data[67][5] ), .ZN(n10367) );
  BUF_X1 U14412 ( .A(n14971), .Z(n20942) );
  BUF_X1 U14413 ( .A(n14913), .Z(n20941) );
  AOI22_X1 U14414 ( .A1(n20942), .A2(\xmem_data[68][5] ), .B1(n20941), .B2(
        \xmem_data[69][5] ), .ZN(n10366) );
  BUF_X1 U14415 ( .A(n14973), .Z(n20943) );
  AOI22_X1 U14416 ( .A1(n24511), .A2(\xmem_data[70][5] ), .B1(n20943), .B2(
        \xmem_data[71][5] ), .ZN(n10365) );
  NAND4_X1 U14417 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10384) );
  BUF_X1 U14418 ( .A(n14974), .Z(n20950) );
  BUF_X1 U14419 ( .A(n14883), .Z(n20949) );
  AOI22_X1 U14420 ( .A1(n20950), .A2(\xmem_data[72][5] ), .B1(n20949), .B2(
        \xmem_data[73][5] ), .ZN(n10372) );
  AOI22_X1 U14421 ( .A1(n20818), .A2(\xmem_data[74][5] ), .B1(n20733), .B2(
        \xmem_data[75][5] ), .ZN(n10371) );
  BUF_X1 U14422 ( .A(n13127), .Z(n20952) );
  BUF_X1 U14423 ( .A(n13487), .Z(n20951) );
  AOI22_X1 U14424 ( .A1(n20952), .A2(\xmem_data[76][5] ), .B1(n20951), .B2(
        \xmem_data[77][5] ), .ZN(n10370) );
  BUF_X1 U14425 ( .A(n31263), .Z(n20953) );
  AOI22_X1 U14426 ( .A1(n20953), .A2(\xmem_data[78][5] ), .B1(n28317), .B2(
        \xmem_data[79][5] ), .ZN(n10369) );
  NAND4_X1 U14427 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10383) );
  AOI22_X1 U14428 ( .A1(n3414), .A2(\xmem_data[80][5] ), .B1(n29173), .B2(
        \xmem_data[81][5] ), .ZN(n10376) );
  AOI22_X1 U14429 ( .A1(n20518), .A2(\xmem_data[82][5] ), .B1(n3219), .B2(
        \xmem_data[83][5] ), .ZN(n10375) );
  AOI22_X1 U14430 ( .A1(n29698), .A2(\xmem_data[84][5] ), .B1(n27444), .B2(
        \xmem_data[85][5] ), .ZN(n10374) );
  BUF_X1 U14431 ( .A(n14926), .Z(n20969) );
  AOI22_X1 U14432 ( .A1(n20969), .A2(\xmem_data[86][5] ), .B1(n28342), .B2(
        \xmem_data[87][5] ), .ZN(n10373) );
  NAND4_X1 U14433 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10382) );
  BUF_X1 U14434 ( .A(n14991), .Z(n20962) );
  AOI22_X1 U14435 ( .A1(n20962), .A2(\xmem_data[88][5] ), .B1(n31252), .B2(
        \xmem_data[89][5] ), .ZN(n10380) );
  BUF_X1 U14436 ( .A(n31276), .Z(n20961) );
  AOI22_X1 U14437 ( .A1(n20961), .A2(\xmem_data[90][5] ), .B1(n24130), .B2(
        \xmem_data[91][5] ), .ZN(n10379) );
  BUF_X1 U14438 ( .A(n14934), .Z(n20958) );
  AOI22_X1 U14439 ( .A1(n23792), .A2(\xmem_data[92][5] ), .B1(n20958), .B2(
        \xmem_data[93][5] ), .ZN(n10378) );
  BUF_X1 U14440 ( .A(n13476), .Z(n20959) );
  AOI22_X1 U14441 ( .A1(n20959), .A2(\xmem_data[94][5] ), .B1(n25709), .B2(
        \xmem_data[95][5] ), .ZN(n10377) );
  NAND4_X1 U14442 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  OR4_X1 U14443 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  NOR2_X1 U14444 ( .A1(n37191), .A2(n39040), .ZN(n21086) );
  NAND2_X1 U14445 ( .A1(n10385), .A2(n21086), .ZN(n10408) );
  BUF_X1 U14446 ( .A(n3464), .Z(n21048) );
  AOI22_X1 U14447 ( .A1(n21048), .A2(\xmem_data[96][5] ), .B1(n20586), .B2(
        \xmem_data[97][5] ), .ZN(n10389) );
  AOI22_X1 U14448 ( .A1(n20542), .A2(\xmem_data[98][5] ), .B1(n24707), .B2(
        \xmem_data[99][5] ), .ZN(n10388) );
  BUF_X1 U14449 ( .A(n14971), .Z(n21050) );
  BUF_X1 U14450 ( .A(n13452), .Z(n21049) );
  AOI22_X1 U14451 ( .A1(n21050), .A2(\xmem_data[100][5] ), .B1(n21049), .B2(
        \xmem_data[101][5] ), .ZN(n10387) );
  BUF_X1 U14452 ( .A(n14882), .Z(n21051) );
  AOI22_X1 U14453 ( .A1(n27974), .A2(\xmem_data[102][5] ), .B1(n25679), .B2(
        \xmem_data[103][5] ), .ZN(n10386) );
  NAND4_X1 U14454 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10405) );
  BUF_X1 U14455 ( .A(n14974), .Z(n21056) );
  AOI22_X1 U14456 ( .A1(n21056), .A2(\xmem_data[104][5] ), .B1(n28098), .B2(
        \xmem_data[105][5] ), .ZN(n10393) );
  BUF_X1 U14457 ( .A(n14976), .Z(n21058) );
  BUF_X1 U14458 ( .A(n14919), .Z(n21057) );
  AOI22_X1 U14459 ( .A1(n21058), .A2(\xmem_data[106][5] ), .B1(n21057), .B2(
        \xmem_data[107][5] ), .ZN(n10392) );
  BUF_X1 U14460 ( .A(n13487), .Z(n21059) );
  AOI22_X1 U14461 ( .A1(n21060), .A2(\xmem_data[108][5] ), .B1(n21059), .B2(
        \xmem_data[109][5] ), .ZN(n10391) );
  BUF_X1 U14462 ( .A(n31263), .Z(n21061) );
  AOI22_X1 U14463 ( .A1(n21061), .A2(\xmem_data[110][5] ), .B1(n20709), .B2(
        \xmem_data[111][5] ), .ZN(n10390) );
  NAND4_X1 U14464 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10404) );
  AOI22_X1 U14465 ( .A1(n3449), .A2(\xmem_data[112][5] ), .B1(n29173), .B2(
        \xmem_data[113][5] ), .ZN(n10397) );
  BUF_X1 U14466 ( .A(n29064), .Z(n21066) );
  AOI22_X1 U14467 ( .A1(n21066), .A2(\xmem_data[114][5] ), .B1(n3218), .B2(
        \xmem_data[115][5] ), .ZN(n10396) );
  BUF_X1 U14468 ( .A(n14988), .Z(n21067) );
  AOI22_X1 U14469 ( .A1(n21067), .A2(\xmem_data[116][5] ), .B1(n30534), .B2(
        \xmem_data[117][5] ), .ZN(n10395) );
  BUF_X1 U14470 ( .A(n14990), .Z(n21069) );
  BUF_X1 U14471 ( .A(n14927), .Z(n21068) );
  AOI22_X1 U14472 ( .A1(n21069), .A2(\xmem_data[118][5] ), .B1(n21068), .B2(
        \xmem_data[119][5] ), .ZN(n10394) );
  NAND4_X1 U14473 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n10403) );
  BUF_X1 U14474 ( .A(n14991), .Z(n21074) );
  AOI22_X1 U14475 ( .A1(n21074), .A2(\xmem_data[120][5] ), .B1(n28007), .B2(
        \xmem_data[121][5] ), .ZN(n10401) );
  AOI22_X1 U14476 ( .A1(n27910), .A2(\xmem_data[122][5] ), .B1(n24130), .B2(
        \xmem_data[123][5] ), .ZN(n10400) );
  BUF_X1 U14477 ( .A(n14934), .Z(n21075) );
  AOI22_X1 U14478 ( .A1(n17013), .A2(\xmem_data[124][5] ), .B1(n21075), .B2(
        \xmem_data[125][5] ), .ZN(n10399) );
  BUF_X1 U14479 ( .A(n14935), .Z(n21076) );
  AOI22_X1 U14480 ( .A1(n24131), .A2(\xmem_data[126][5] ), .B1(n21076), .B2(
        \xmem_data[127][5] ), .ZN(n10398) );
  NAND4_X1 U14481 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  OR4_X1 U14482 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10406) );
  AND2_X1 U14483 ( .A1(n37191), .A2(load_xaddr_val[6]), .ZN(n21088) );
  NAND2_X1 U14484 ( .A1(n10406), .A2(n21088), .ZN(n10407) );
  NAND2_X1 U14485 ( .A1(n10408), .A2(n10407), .ZN(n10431) );
  AOI22_X1 U14486 ( .A1(n20939), .A2(\xmem_data[32][5] ), .B1(n20938), .B2(
        \xmem_data[33][5] ), .ZN(n10412) );
  AOI22_X1 U14487 ( .A1(n20800), .A2(\xmem_data[34][5] ), .B1(n20940), .B2(
        \xmem_data[35][5] ), .ZN(n10411) );
  AOI22_X1 U14488 ( .A1(n20942), .A2(\xmem_data[36][5] ), .B1(n20941), .B2(
        \xmem_data[37][5] ), .ZN(n10410) );
  AOI22_X1 U14489 ( .A1(n30899), .A2(\xmem_data[38][5] ), .B1(n20943), .B2(
        \xmem_data[39][5] ), .ZN(n10409) );
  NAND4_X1 U14490 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n10428) );
  AOI22_X1 U14491 ( .A1(n20950), .A2(\xmem_data[40][5] ), .B1(n20949), .B2(
        \xmem_data[41][5] ), .ZN(n10416) );
  AOI22_X1 U14492 ( .A1(n24166), .A2(\xmem_data[42][5] ), .B1(n14981), .B2(
        \xmem_data[43][5] ), .ZN(n10415) );
  AOI22_X1 U14493 ( .A1(n20952), .A2(\xmem_data[44][5] ), .B1(n20951), .B2(
        \xmem_data[45][5] ), .ZN(n10414) );
  AOI22_X1 U14494 ( .A1(n20953), .A2(\xmem_data[46][5] ), .B1(n27563), .B2(
        \xmem_data[47][5] ), .ZN(n10413) );
  NAND4_X1 U14495 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10427) );
  AOI22_X1 U14496 ( .A1(n16980), .A2(\xmem_data[48][5] ), .B1(n30589), .B2(
        \xmem_data[49][5] ), .ZN(n10420) );
  AOI22_X1 U14497 ( .A1(n24631), .A2(\xmem_data[50][5] ), .B1(n3222), .B2(
        \xmem_data[51][5] ), .ZN(n10419) );
  AOI22_X1 U14498 ( .A1(n29026), .A2(\xmem_data[52][5] ), .B1(n27444), .B2(
        \xmem_data[53][5] ), .ZN(n10418) );
  AOI22_X1 U14499 ( .A1(n20969), .A2(\xmem_data[54][5] ), .B1(n22759), .B2(
        \xmem_data[55][5] ), .ZN(n10417) );
  NAND4_X1 U14500 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10426) );
  AOI22_X1 U14501 ( .A1(n20962), .A2(\xmem_data[56][5] ), .B1(n29103), .B2(
        \xmem_data[57][5] ), .ZN(n10424) );
  AOI22_X1 U14502 ( .A1(n20961), .A2(\xmem_data[58][5] ), .B1(n27943), .B2(
        \xmem_data[59][5] ), .ZN(n10423) );
  AOI22_X1 U14503 ( .A1(n20799), .A2(\xmem_data[60][5] ), .B1(n20958), .B2(
        \xmem_data[61][5] ), .ZN(n10422) );
  AOI22_X1 U14504 ( .A1(n20959), .A2(\xmem_data[62][5] ), .B1(n25606), .B2(
        \xmem_data[63][5] ), .ZN(n10421) );
  NAND4_X1 U14505 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  OR4_X1 U14506 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10429) );
  NOR2_X1 U14507 ( .A1(n10431), .A2(n10430), .ZN(n10467) );
  NAND2_X1 U14508 ( .A1(n24131), .A2(\xmem_data[30][5] ), .ZN(n10433) );
  BUF_X1 U14509 ( .A(n14972), .Z(n21010) );
  AOI22_X1 U14510 ( .A1(n25422), .A2(\xmem_data[26][5] ), .B1(n20982), .B2(
        \xmem_data[27][5] ), .ZN(n10434) );
  BUF_X1 U14511 ( .A(n14926), .Z(n20994) );
  BUF_X1 U14512 ( .A(n14890), .Z(n20993) );
  AOI22_X1 U14513 ( .A1(n20994), .A2(\xmem_data[22][5] ), .B1(n20993), .B2(
        \xmem_data[23][5] ), .ZN(n10435) );
  BUF_X1 U14514 ( .A(n14989), .Z(n20992) );
  AOI22_X1 U14515 ( .A1(n25612), .A2(\xmem_data[20][5] ), .B1(n20992), .B2(
        \xmem_data[21][5] ), .ZN(n10436) );
  AOI22_X1 U14516 ( .A1(n3142), .A2(\xmem_data[16][5] ), .B1(n27437), .B2(
        \xmem_data[17][5] ), .ZN(n10438) );
  BUF_X1 U14517 ( .A(n14974), .Z(n20984) );
  BUF_X1 U14518 ( .A(n14914), .Z(n20983) );
  AOI22_X1 U14519 ( .A1(n20984), .A2(\xmem_data[8][5] ), .B1(n20983), .B2(
        \xmem_data[9][5] ), .ZN(n10437) );
  AOI22_X1 U14520 ( .A1(n29325), .A2(\xmem_data[10][5] ), .B1(n29086), .B2(
        \xmem_data[11][5] ), .ZN(n10440) );
  AOI22_X1 U14521 ( .A1(n25732), .A2(\xmem_data[24][5] ), .B1(n13474), .B2(
        \xmem_data[25][5] ), .ZN(n10439) );
  BUF_X1 U14522 ( .A(n14934), .Z(n21015) );
  AOI22_X1 U14523 ( .A1(n31327), .A2(\xmem_data[28][5] ), .B1(n21015), .B2(
        \xmem_data[29][5] ), .ZN(n10448) );
  INV_X1 U14524 ( .A(n10448), .ZN(n10451) );
  BUF_X1 U14525 ( .A(n14971), .Z(n21008) );
  AOI22_X1 U14526 ( .A1(n21008), .A2(\xmem_data[4][5] ), .B1(n29238), .B2(
        \xmem_data[5][5] ), .ZN(n10449) );
  INV_X1 U14527 ( .A(n10449), .ZN(n10450) );
  BUF_X1 U14528 ( .A(n29064), .Z(n20991) );
  AOI22_X1 U14529 ( .A1(n20991), .A2(\xmem_data[18][5] ), .B1(n3222), .B2(
        \xmem_data[19][5] ), .ZN(n10452) );
  BUF_X1 U14530 ( .A(n3464), .Z(n21005) );
  AOI22_X1 U14531 ( .A1(n21005), .A2(\xmem_data[0][5] ), .B1(n20543), .B2(
        \xmem_data[1][5] ), .ZN(n10455) );
  BUF_X1 U14532 ( .A(n14882), .Z(n21009) );
  AOI22_X1 U14533 ( .A1(n14935), .A2(\xmem_data[31][5] ), .B1(n20816), .B2(
        \xmem_data[7][5] ), .ZN(n10454) );
  BUF_X1 U14534 ( .A(n13420), .Z(n20985) );
  AOI22_X1 U14535 ( .A1(n20985), .A2(\xmem_data[12][5] ), .B1(n24686), .B2(
        \xmem_data[13][5] ), .ZN(n10457) );
  BUF_X1 U14536 ( .A(n31263), .Z(n20986) );
  AOI22_X1 U14537 ( .A1(n20986), .A2(\xmem_data[14][5] ), .B1(n20578), .B2(
        \xmem_data[15][5] ), .ZN(n10459) );
  BUF_X1 U14538 ( .A(n14912), .Z(n21006) );
  AOI22_X1 U14539 ( .A1(n21007), .A2(\xmem_data[2][5] ), .B1(n21006), .B2(
        \xmem_data[3][5] ), .ZN(n10458) );
  NOR2_X1 U14540 ( .A1(n37191), .A2(load_xaddr_val[6]), .ZN(n20980) );
  AOI22_X1 U14541 ( .A1(n31268), .A2(\xmem_data[30][4] ), .B1(n29309), .B2(
        \xmem_data[31][4] ), .ZN(n10468) );
  INV_X1 U14542 ( .A(n10468), .ZN(n10471) );
  AOI22_X1 U14543 ( .A1(n29179), .A2(\xmem_data[28][4] ), .B1(n21015), .B2(
        \xmem_data[29][4] ), .ZN(n10469) );
  INV_X1 U14544 ( .A(n10469), .ZN(n10470) );
  NOR2_X1 U14545 ( .A1(n10471), .A2(n10470), .ZN(n10474) );
  AOI22_X1 U14546 ( .A1(n23813), .A2(\xmem_data[26][4] ), .B1(n20982), .B2(
        \xmem_data[27][4] ), .ZN(n10473) );
  NAND2_X1 U14547 ( .A1(n17063), .A2(\xmem_data[24][4] ), .ZN(n10472) );
  NAND2_X1 U14548 ( .A1(n10474), .A2(n3925), .ZN(n10486) );
  AOI22_X1 U14549 ( .A1(n21005), .A2(\xmem_data[0][4] ), .B1(n3212), .B2(
        \xmem_data[1][4] ), .ZN(n10478) );
  AOI22_X1 U14550 ( .A1(n21007), .A2(\xmem_data[2][4] ), .B1(n21006), .B2(
        \xmem_data[3][4] ), .ZN(n10477) );
  AOI22_X1 U14551 ( .A1(n21008), .A2(\xmem_data[4][4] ), .B1(n29238), .B2(
        \xmem_data[5][4] ), .ZN(n10476) );
  AOI22_X1 U14552 ( .A1(n21010), .A2(\xmem_data[6][4] ), .B1(n28327), .B2(
        \xmem_data[7][4] ), .ZN(n10475) );
  NAND4_X1 U14553 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n10485) );
  AOI22_X1 U14554 ( .A1(n3332), .A2(\xmem_data[16][4] ), .B1(n25442), .B2(
        \xmem_data[17][4] ), .ZN(n10483) );
  AND2_X1 U14555 ( .A1(n3217), .A2(\xmem_data[19][4] ), .ZN(n10479) );
  AOI21_X1 U14556 ( .B1(n20991), .B2(\xmem_data[18][4] ), .A(n10479), .ZN(
        n10482) );
  AOI22_X1 U14557 ( .A1(n27708), .A2(\xmem_data[20][4] ), .B1(n20992), .B2(
        \xmem_data[21][4] ), .ZN(n10481) );
  AOI22_X1 U14558 ( .A1(n20994), .A2(\xmem_data[22][4] ), .B1(n20993), .B2(
        \xmem_data[23][4] ), .ZN(n10480) );
  NAND4_X1 U14559 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10484) );
  AOI22_X1 U14560 ( .A1(n20984), .A2(\xmem_data[8][4] ), .B1(n20983), .B2(
        \xmem_data[9][4] ), .ZN(n10490) );
  AOI22_X1 U14561 ( .A1(n31316), .A2(\xmem_data[10][4] ), .B1(n28328), .B2(
        \xmem_data[11][4] ), .ZN(n10489) );
  AOI22_X1 U14562 ( .A1(n20985), .A2(\xmem_data[12][4] ), .B1(n20769), .B2(
        \xmem_data[13][4] ), .ZN(n10488) );
  AOI22_X1 U14563 ( .A1(n20986), .A2(\xmem_data[14][4] ), .B1(n29118), .B2(
        \xmem_data[15][4] ), .ZN(n10487) );
  NAND4_X1 U14564 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  NOR2_X1 U14565 ( .A1(n10491), .A2(n3877), .ZN(n10492) );
  INV_X1 U14566 ( .A(n20980), .ZN(n20386) );
  AOI21_X1 U14567 ( .B1(n10493), .B2(n10492), .A(n20386), .ZN(n10494) );
  INV_X1 U14568 ( .A(n10494), .ZN(n10561) );
  AOI22_X1 U14569 ( .A1(n20939), .A2(\xmem_data[32][4] ), .B1(n20938), .B2(
        \xmem_data[33][4] ), .ZN(n10498) );
  AOI22_X1 U14570 ( .A1(n20585), .A2(\xmem_data[34][4] ), .B1(n20940), .B2(
        \xmem_data[35][4] ), .ZN(n10497) );
  AOI22_X1 U14571 ( .A1(n20942), .A2(\xmem_data[36][4] ), .B1(n20941), .B2(
        \xmem_data[37][4] ), .ZN(n10496) );
  AOI22_X1 U14572 ( .A1(n29240), .A2(\xmem_data[38][4] ), .B1(n20943), .B2(
        \xmem_data[39][4] ), .ZN(n10495) );
  NAND4_X1 U14573 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10514) );
  AOI22_X1 U14574 ( .A1(n20950), .A2(\xmem_data[40][4] ), .B1(n20949), .B2(
        \xmem_data[41][4] ), .ZN(n10502) );
  AOI22_X1 U14575 ( .A1(n29325), .A2(\xmem_data[42][4] ), .B1(n29136), .B2(
        \xmem_data[43][4] ), .ZN(n10501) );
  AOI22_X1 U14576 ( .A1(n20952), .A2(\xmem_data[44][4] ), .B1(n20951), .B2(
        \xmem_data[45][4] ), .ZN(n10500) );
  AOI22_X1 U14577 ( .A1(n20953), .A2(\xmem_data[46][4] ), .B1(n27499), .B2(
        \xmem_data[47][4] ), .ZN(n10499) );
  NAND4_X1 U14578 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10513) );
  AOI22_X1 U14579 ( .A1(n3348), .A2(\xmem_data[48][4] ), .B1(n29173), .B2(
        \xmem_data[49][4] ), .ZN(n10506) );
  AOI22_X1 U14580 ( .A1(n27502), .A2(\xmem_data[50][4] ), .B1(n3219), .B2(
        \xmem_data[51][4] ), .ZN(n10505) );
  AOI22_X1 U14581 ( .A1(n25448), .A2(\xmem_data[52][4] ), .B1(n22667), .B2(
        \xmem_data[53][4] ), .ZN(n10504) );
  AOI22_X1 U14582 ( .A1(n20969), .A2(\xmem_data[54][4] ), .B1(n13444), .B2(
        \xmem_data[55][4] ), .ZN(n10503) );
  NAND4_X1 U14583 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10512) );
  AOI22_X1 U14584 ( .A1(n20962), .A2(\xmem_data[56][4] ), .B1(n28343), .B2(
        \xmem_data[57][4] ), .ZN(n10510) );
  AOI22_X1 U14585 ( .A1(n20961), .A2(\xmem_data[58][4] ), .B1(n24130), .B2(
        \xmem_data[59][4] ), .ZN(n10509) );
  AOI22_X1 U14586 ( .A1(n28743), .A2(\xmem_data[60][4] ), .B1(n20958), .B2(
        \xmem_data[61][4] ), .ZN(n10508) );
  AOI22_X1 U14587 ( .A1(n20959), .A2(\xmem_data[62][4] ), .B1(n30541), .B2(
        \xmem_data[63][4] ), .ZN(n10507) );
  NAND4_X1 U14588 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10511) );
  OR4_X1 U14589 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10515) );
  NAND2_X1 U14590 ( .A1(n10515), .A2(n20311), .ZN(n10560) );
  AOI22_X1 U14591 ( .A1(n21048), .A2(\xmem_data[96][4] ), .B1(n28299), .B2(
        \xmem_data[97][4] ), .ZN(n10519) );
  AOI22_X1 U14592 ( .A1(n22676), .A2(\xmem_data[98][4] ), .B1(n28492), .B2(
        \xmem_data[99][4] ), .ZN(n10518) );
  AOI22_X1 U14593 ( .A1(n21050), .A2(\xmem_data[100][4] ), .B1(n21049), .B2(
        \xmem_data[101][4] ), .ZN(n10517) );
  AOI22_X1 U14594 ( .A1(n25632), .A2(\xmem_data[102][4] ), .B1(n28429), .B2(
        \xmem_data[103][4] ), .ZN(n10516) );
  NAND4_X1 U14595 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10535) );
  AOI22_X1 U14596 ( .A1(n21056), .A2(\xmem_data[104][4] ), .B1(n28098), .B2(
        \xmem_data[105][4] ), .ZN(n10523) );
  AOI22_X1 U14597 ( .A1(n21058), .A2(\xmem_data[106][4] ), .B1(n21057), .B2(
        \xmem_data[107][4] ), .ZN(n10522) );
  AOI22_X1 U14598 ( .A1(n21060), .A2(\xmem_data[108][4] ), .B1(n21059), .B2(
        \xmem_data[109][4] ), .ZN(n10521) );
  AOI22_X1 U14599 ( .A1(n21061), .A2(\xmem_data[110][4] ), .B1(n24470), .B2(
        \xmem_data[111][4] ), .ZN(n10520) );
  NAND4_X1 U14600 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10534) );
  AOI22_X1 U14601 ( .A1(n3144), .A2(\xmem_data[112][4] ), .B1(n28501), .B2(
        \xmem_data[113][4] ), .ZN(n10527) );
  AOI22_X1 U14602 ( .A1(n21066), .A2(\xmem_data[114][4] ), .B1(n3218), .B2(
        \xmem_data[115][4] ), .ZN(n10526) );
  AOI22_X1 U14603 ( .A1(n21067), .A2(\xmem_data[116][4] ), .B1(n25509), .B2(
        \xmem_data[117][4] ), .ZN(n10525) );
  AOI22_X1 U14604 ( .A1(n21069), .A2(\xmem_data[118][4] ), .B1(n21068), .B2(
        \xmem_data[119][4] ), .ZN(n10524) );
  NAND4_X1 U14605 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10533) );
  AOI22_X1 U14606 ( .A1(n21074), .A2(\xmem_data[120][4] ), .B1(n25450), .B2(
        \xmem_data[121][4] ), .ZN(n10531) );
  AOI22_X1 U14607 ( .A1(n28050), .A2(\xmem_data[122][4] ), .B1(n3358), .B2(
        \xmem_data[123][4] ), .ZN(n10530) );
  AOI22_X1 U14608 ( .A1(n27911), .A2(\xmem_data[124][4] ), .B1(n21075), .B2(
        \xmem_data[125][4] ), .ZN(n10529) );
  AOI22_X1 U14609 ( .A1(n25459), .A2(\xmem_data[126][4] ), .B1(n21076), .B2(
        \xmem_data[127][4] ), .ZN(n10528) );
  NAND4_X1 U14610 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  OR4_X1 U14611 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10536) );
  NAND2_X1 U14612 ( .A1(n10536), .A2(n21088), .ZN(n10559) );
  AOI22_X1 U14613 ( .A1(n20939), .A2(\xmem_data[64][4] ), .B1(n20938), .B2(
        \xmem_data[65][4] ), .ZN(n10540) );
  AOI22_X1 U14614 ( .A1(n23717), .A2(\xmem_data[66][4] ), .B1(n20940), .B2(
        \xmem_data[67][4] ), .ZN(n10539) );
  AOI22_X1 U14615 ( .A1(n20942), .A2(\xmem_data[68][4] ), .B1(n20941), .B2(
        \xmem_data[69][4] ), .ZN(n10538) );
  AOI22_X1 U14616 ( .A1(n24647), .A2(\xmem_data[70][4] ), .B1(n20943), .B2(
        \xmem_data[71][4] ), .ZN(n10537) );
  NAND4_X1 U14617 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .ZN(
        n10556) );
  AOI22_X1 U14618 ( .A1(n20950), .A2(\xmem_data[72][4] ), .B1(n20949), .B2(
        \xmem_data[73][4] ), .ZN(n10544) );
  AOI22_X1 U14619 ( .A1(n20734), .A2(\xmem_data[74][4] ), .B1(n28468), .B2(
        \xmem_data[75][4] ), .ZN(n10543) );
  AOI22_X1 U14620 ( .A1(n20952), .A2(\xmem_data[76][4] ), .B1(n20951), .B2(
        \xmem_data[77][4] ), .ZN(n10542) );
  AOI22_X1 U14621 ( .A1(n20953), .A2(\xmem_data[78][4] ), .B1(n28317), .B2(
        \xmem_data[79][4] ), .ZN(n10541) );
  NAND4_X1 U14622 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10555) );
  AOI22_X1 U14623 ( .A1(n3228), .A2(\xmem_data[80][4] ), .B1(n20711), .B2(
        \xmem_data[81][4] ), .ZN(n10548) );
  AOI22_X1 U14624 ( .A1(n28503), .A2(\xmem_data[82][4] ), .B1(n3219), .B2(
        \xmem_data[83][4] ), .ZN(n10547) );
  AOI22_X1 U14625 ( .A1(n21067), .A2(\xmem_data[84][4] ), .B1(n22667), .B2(
        \xmem_data[85][4] ), .ZN(n10546) );
  AOI22_X1 U14626 ( .A1(n20969), .A2(\xmem_data[86][4] ), .B1(n24564), .B2(
        \xmem_data[87][4] ), .ZN(n10545) );
  NAND4_X1 U14627 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10554) );
  AOI22_X1 U14628 ( .A1(n20962), .A2(\xmem_data[88][4] ), .B1(n25450), .B2(
        \xmem_data[89][4] ), .ZN(n10552) );
  AOI22_X1 U14629 ( .A1(n20961), .A2(\xmem_data[90][4] ), .B1(n27863), .B2(
        \xmem_data[91][4] ), .ZN(n10551) );
  AOI22_X1 U14630 ( .A1(n20587), .A2(\xmem_data[92][4] ), .B1(n20958), .B2(
        \xmem_data[93][4] ), .ZN(n10550) );
  AOI22_X1 U14631 ( .A1(n20959), .A2(\xmem_data[94][4] ), .B1(n20584), .B2(
        \xmem_data[95][4] ), .ZN(n10549) );
  NAND4_X1 U14632 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10553) );
  OR4_X1 U14633 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10557) );
  NAND2_X1 U14634 ( .A1(n10557), .A2(n21086), .ZN(n10558) );
  XOR2_X1 U14635 ( .A(\fmem_data[0][5] ), .B(\fmem_data[0][4] ), .Z(n10562) );
  NAND2_X1 U14636 ( .A1(n27568), .A2(\xmem_data[0][5] ), .ZN(n10564) );
  BUF_X1 U14637 ( .A(n13457), .Z(n27567) );
  NAND2_X1 U14638 ( .A1(n27567), .A2(\xmem_data[1][5] ), .ZN(n10563) );
  NAND2_X1 U14639 ( .A1(n10564), .A2(n10563), .ZN(n10571) );
  AOI22_X1 U14640 ( .A1(n17020), .A2(\xmem_data[22][5] ), .B1(n21006), .B2(
        \xmem_data[23][5] ), .ZN(n10566) );
  NAND2_X1 U14641 ( .A1(n27551), .A2(\xmem_data[14][5] ), .ZN(n10565) );
  NAND2_X1 U14642 ( .A1(n10566), .A2(n10565), .ZN(n10570) );
  BUF_X1 U14643 ( .A(n13435), .Z(n27535) );
  AOI22_X1 U14644 ( .A1(n23762), .A2(\xmem_data[16][5] ), .B1(n27535), .B2(
        \xmem_data[17][5] ), .ZN(n10568) );
  AOI22_X1 U14645 ( .A1(n30292), .A2(\xmem_data[8][5] ), .B1(n20992), .B2(
        \xmem_data[9][5] ), .ZN(n10567) );
  AOI22_X1 U14646 ( .A1(n25354), .A2(\xmem_data[6][5] ), .B1(n3220), .B2(
        \xmem_data[7][5] ), .ZN(n10572) );
  INV_X1 U14647 ( .A(n10572), .ZN(n10585) );
  BUF_X1 U14648 ( .A(n31263), .Z(n27564) );
  BUF_X1 U14649 ( .A(n28974), .Z(n27563) );
  AOI22_X1 U14650 ( .A1(n27564), .A2(\xmem_data[2][5] ), .B1(n27563), .B2(
        \xmem_data[3][5] ), .ZN(n10573) );
  INV_X1 U14651 ( .A(n10573), .ZN(n10584) );
  BUF_X1 U14652 ( .A(n14890), .Z(n27550) );
  AOI22_X1 U14653 ( .A1(n27904), .A2(\xmem_data[10][5] ), .B1(n27550), .B2(
        \xmem_data[11][5] ), .ZN(n10574) );
  INV_X1 U14654 ( .A(n10574), .ZN(n10578) );
  AOI22_X1 U14655 ( .A1(n25607), .A2(\xmem_data[20][5] ), .B1(n30542), .B2(
        \xmem_data[21][5] ), .ZN(n10576) );
  BUF_X1 U14656 ( .A(n14999), .Z(n27536) );
  AOI22_X1 U14657 ( .A1(n27536), .A2(\xmem_data[19][5] ), .B1(
        \xmem_data[15][5] ), .B2(n28415), .ZN(n10575) );
  NAND2_X1 U14658 ( .A1(n10576), .A2(n10575), .ZN(n10577) );
  NOR2_X1 U14659 ( .A1(n10578), .A2(n10577), .ZN(n10582) );
  BUF_X1 U14660 ( .A(n10977), .Z(n27537) );
  AOI22_X1 U14661 ( .A1(n28677), .A2(\xmem_data[4][5] ), .B1(n25360), .B2(
        \xmem_data[5][5] ), .ZN(n10579) );
  INV_X1 U14662 ( .A(n10579), .ZN(n10580) );
  NOR2_X1 U14663 ( .A1(n3880), .A2(n10580), .ZN(n10581) );
  NAND2_X1 U14664 ( .A1(n10582), .A2(n10581), .ZN(n10583) );
  NOR3_X1 U14665 ( .A1(n10585), .A2(n10584), .A3(n10583), .ZN(n10587) );
  BUF_X1 U14666 ( .A(n14928), .Z(n27547) );
  AOI22_X1 U14667 ( .A1(n3132), .A2(\xmem_data[12][5] ), .B1(n3231), .B2(
        \xmem_data[13][5] ), .ZN(n10586) );
  NAND3_X1 U14668 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n10594) );
  NOR2_X1 U14669 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  INV_X1 U14670 ( .A(n10591), .ZN(n10592) );
  AOI22_X1 U14671 ( .A1(n37191), .A2(n10592), .B1(n10591), .B2(n4499), .ZN(
        n10650) );
  NAND2_X1 U14672 ( .A1(load_xaddr_val[5]), .A2(n10592), .ZN(n10593) );
  XOR2_X1 U14673 ( .A(n39040), .B(n10593), .Z(n10628) );
  NOR2_X1 U14674 ( .A1(n10650), .A2(n10628), .ZN(n19410) );
  NAND2_X1 U14675 ( .A1(n10594), .A2(n19410), .ZN(n10675) );
  BUF_X1 U14676 ( .A(n14997), .Z(n27514) );
  BUF_X1 U14677 ( .A(n13435), .Z(n27513) );
  AOI22_X1 U14678 ( .A1(n27514), .A2(\xmem_data[48][5] ), .B1(n27513), .B2(
        \xmem_data[49][5] ), .ZN(n10598) );
  BUF_X1 U14679 ( .A(n13476), .Z(n27515) );
  AOI22_X1 U14680 ( .A1(n27515), .A2(\xmem_data[50][5] ), .B1(n20798), .B2(
        \xmem_data[51][5] ), .ZN(n10597) );
  BUF_X1 U14681 ( .A(n29187), .Z(n27517) );
  AOI22_X1 U14682 ( .A1(n28091), .A2(\xmem_data[52][5] ), .B1(n27516), .B2(
        \xmem_data[53][5] ), .ZN(n10596) );
  BUF_X1 U14683 ( .A(n14912), .Z(n27518) );
  AOI22_X1 U14684 ( .A1(n24708), .A2(\xmem_data[54][5] ), .B1(n27518), .B2(
        \xmem_data[55][5] ), .ZN(n10595) );
  NAND4_X1 U14685 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10604) );
  BUF_X1 U14686 ( .A(n14913), .Z(n27523) );
  AOI22_X1 U14687 ( .A1(n30617), .A2(\xmem_data[56][5] ), .B1(n27523), .B2(
        \xmem_data[57][5] ), .ZN(n10602) );
  BUF_X1 U14688 ( .A(n14881), .Z(n27524) );
  AOI22_X1 U14689 ( .A1(n27524), .A2(\xmem_data[58][5] ), .B1(n30495), .B2(
        \xmem_data[59][5] ), .ZN(n10601) );
  BUF_X1 U14690 ( .A(n14914), .Z(n27525) );
  AOI22_X1 U14691 ( .A1(n30645), .A2(\xmem_data[60][5] ), .B1(n27525), .B2(
        \xmem_data[61][5] ), .ZN(n10600) );
  AOI22_X1 U14692 ( .A1(n22719), .A2(\xmem_data[62][5] ), .B1(n27526), .B2(
        \xmem_data[63][5] ), .ZN(n10599) );
  NAND4_X1 U14693 ( .A1(n10602), .A2(n10601), .A3(n10600), .A4(n10599), .ZN(
        n10603) );
  OR3_X1 U14694 ( .A1(n10604), .A2(n10603), .A3(n3932), .ZN(n10613) );
  BUF_X1 U14695 ( .A(n13469), .Z(n27507) );
  AOI22_X1 U14696 ( .A1(n29065), .A2(\xmem_data[40][5] ), .B1(n27507), .B2(
        \xmem_data[41][5] ), .ZN(n10605) );
  INV_X1 U14697 ( .A(n10605), .ZN(n10609) );
  BUF_X1 U14698 ( .A(n31276), .Z(n27508) );
  AOI22_X1 U14699 ( .A1(n27508), .A2(\xmem_data[46][5] ), .B1(n28373), .B2(
        \xmem_data[47][5] ), .ZN(n10606) );
  INV_X1 U14700 ( .A(n10606), .ZN(n10608) );
  AND2_X1 U14701 ( .A1(n3147), .A2(\xmem_data[44][5] ), .ZN(n10607) );
  NOR3_X1 U14702 ( .A1(n10609), .A2(n10608), .A3(n10607), .ZN(n10611) );
  AOI22_X1 U14703 ( .A1(n30606), .A2(\xmem_data[42][5] ), .B1(n13444), .B2(
        \xmem_data[43][5] ), .ZN(n10610) );
  NAND2_X1 U14704 ( .A1(n10611), .A2(n10610), .ZN(n10612) );
  NOR2_X1 U14705 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  INV_X1 U14706 ( .A(n10628), .ZN(n10649) );
  AND2_X1 U14707 ( .A1(n10649), .A2(n10650), .ZN(n27577) );
  INV_X1 U14708 ( .A(n27577), .ZN(n19406) );
  NOR2_X1 U14709 ( .A1(n10614), .A2(n19406), .ZN(n10627) );
  BUF_X1 U14710 ( .A(n13127), .Z(n27498) );
  AOI22_X1 U14711 ( .A1(n27498), .A2(\xmem_data[32][5] ), .B1(n24468), .B2(
        \xmem_data[33][5] ), .ZN(n10619) );
  BUF_X1 U14712 ( .A(n31263), .Z(n27500) );
  BUF_X1 U14713 ( .A(n28947), .Z(n27499) );
  AOI22_X1 U14714 ( .A1(n27500), .A2(\xmem_data[34][5] ), .B1(n27499), .B2(
        \xmem_data[35][5] ), .ZN(n10618) );
  BUF_X1 U14715 ( .A(n13468), .Z(n27501) );
  AOI22_X1 U14716 ( .A1(n22728), .A2(\xmem_data[36][5] ), .B1(n27501), .B2(
        \xmem_data[37][5] ), .ZN(n10617) );
  BUF_X1 U14717 ( .A(n29064), .Z(n27502) );
  AND2_X1 U14718 ( .A1(n3218), .A2(\xmem_data[39][5] ), .ZN(n10615) );
  AOI21_X1 U14719 ( .B1(n27502), .B2(\xmem_data[38][5] ), .A(n10615), .ZN(
        n10616) );
  AOI22_X1 U14720 ( .A1(n27855), .A2(\xmem_data[24][5] ), .B1(n13452), .B2(
        \xmem_data[25][5] ), .ZN(n10623) );
  AOI22_X1 U14721 ( .A1(n29240), .A2(\xmem_data[26][5] ), .B1(n27461), .B2(
        \xmem_data[27][5] ), .ZN(n10622) );
  AOI22_X1 U14722 ( .A1(n28701), .A2(\xmem_data[28][5] ), .B1(n28098), .B2(
        \xmem_data[29][5] ), .ZN(n10621) );
  BUF_X1 U14723 ( .A(n14976), .Z(n27542) );
  AOI22_X1 U14724 ( .A1(n27542), .A2(\xmem_data[30][5] ), .B1(n17049), .B2(
        \xmem_data[31][5] ), .ZN(n10620) );
  NAND4_X1 U14725 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10624) );
  NAND2_X1 U14726 ( .A1(n10624), .A2(n19410), .ZN(n10625) );
  OAI21_X1 U14727 ( .B1(n3754), .B2(n19406), .A(n10625), .ZN(n10626) );
  NOR2_X1 U14728 ( .A1(n10627), .A2(n10626), .ZN(n10674) );
  AND2_X1 U14729 ( .A1(n10650), .A2(n10628), .ZN(n27496) );
  BUF_X1 U14730 ( .A(n13487), .Z(n27435) );
  AOI22_X1 U14731 ( .A1(n25684), .A2(\xmem_data[96][5] ), .B1(n27435), .B2(
        \xmem_data[97][5] ), .ZN(n10632) );
  BUF_X1 U14732 ( .A(n31263), .Z(n27436) );
  AOI22_X1 U14733 ( .A1(n27436), .A2(\xmem_data[98][5] ), .B1(n28037), .B2(
        \xmem_data[99][5] ), .ZN(n10631) );
  AOI22_X1 U14734 ( .A1(n3334), .A2(\xmem_data[100][5] ), .B1(n27437), .B2(
        \xmem_data[101][5] ), .ZN(n10630) );
  BUF_X1 U14735 ( .A(n29064), .Z(n27439) );
  AOI22_X1 U14736 ( .A1(n27439), .A2(\xmem_data[102][5] ), .B1(n3218), .B2(
        \xmem_data[103][5] ), .ZN(n10629) );
  NAND4_X1 U14737 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10648) );
  BUF_X1 U14738 ( .A(n14988), .Z(n27445) );
  BUF_X1 U14739 ( .A(n14925), .Z(n27444) );
  AOI22_X1 U14740 ( .A1(n27445), .A2(\xmem_data[104][5] ), .B1(n27444), .B2(
        \xmem_data[105][5] ), .ZN(n10636) );
  AOI22_X1 U14741 ( .A1(n27938), .A2(\xmem_data[106][5] ), .B1(n24564), .B2(
        \xmem_data[107][5] ), .ZN(n10635) );
  BUF_X1 U14742 ( .A(n13474), .Z(n27446) );
  AOI22_X1 U14743 ( .A1(n3126), .A2(\xmem_data[108][5] ), .B1(n27446), .B2(
        \xmem_data[109][5] ), .ZN(n10634) );
  AOI22_X1 U14744 ( .A1(n27447), .A2(\xmem_data[110][5] ), .B1(n28481), .B2(
        \xmem_data[111][5] ), .ZN(n10633) );
  NAND4_X1 U14745 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n10647) );
  BUF_X1 U14746 ( .A(n14997), .Z(n27453) );
  BUF_X1 U14747 ( .A(n14998), .Z(n27452) );
  AOI22_X1 U14748 ( .A1(n27453), .A2(\xmem_data[112][5] ), .B1(n27452), .B2(
        \xmem_data[113][5] ), .ZN(n10640) );
  AOI22_X1 U14749 ( .A1(n16986), .A2(\xmem_data[114][5] ), .B1(n24160), .B2(
        \xmem_data[115][5] ), .ZN(n10639) );
  BUF_X1 U14750 ( .A(n3464), .Z(n27455) );
  BUF_X1 U14751 ( .A(n14936), .Z(n27454) );
  AOI22_X1 U14752 ( .A1(n3466), .A2(\xmem_data[116][5] ), .B1(n27454), .B2(
        \xmem_data[117][5] ), .ZN(n10638) );
  AOI22_X1 U14753 ( .A1(n20542), .A2(\xmem_data[118][5] ), .B1(n22718), .B2(
        \xmem_data[119][5] ), .ZN(n10637) );
  NAND4_X1 U14754 ( .A1(n10640), .A2(n10639), .A3(n10638), .A4(n10637), .ZN(
        n10646) );
  BUF_X1 U14755 ( .A(n13452), .Z(n27460) );
  AOI22_X1 U14756 ( .A1(n20730), .A2(\xmem_data[120][5] ), .B1(n27460), .B2(
        \xmem_data[121][5] ), .ZN(n10644) );
  BUF_X1 U14757 ( .A(n14881), .Z(n27462) );
  BUF_X1 U14758 ( .A(n14973), .Z(n27461) );
  AOI22_X1 U14759 ( .A1(n27462), .A2(\xmem_data[122][5] ), .B1(n27461), .B2(
        \xmem_data[123][5] ), .ZN(n10643) );
  AOI22_X1 U14760 ( .A1(n28202), .A2(\xmem_data[124][5] ), .B1(n28983), .B2(
        \xmem_data[125][5] ), .ZN(n10642) );
  BUF_X1 U14761 ( .A(n14919), .Z(n27463) );
  AOI22_X1 U14762 ( .A1(n22719), .A2(\xmem_data[126][5] ), .B1(n27463), .B2(
        \xmem_data[127][5] ), .ZN(n10641) );
  NAND4_X1 U14763 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        n10645) );
  OR4_X1 U14764 ( .A1(n10648), .A2(n10647), .A3(n10646), .A4(n10645), .ZN(
        n10672) );
  NOR2_X1 U14765 ( .A1(n10650), .A2(n10649), .ZN(n27494) );
  AOI22_X1 U14766 ( .A1(n27498), .A2(\xmem_data[64][5] ), .B1(n20951), .B2(
        \xmem_data[65][5] ), .ZN(n10654) );
  AOI22_X1 U14767 ( .A1(n27500), .A2(\xmem_data[66][5] ), .B1(n27499), .B2(
        \xmem_data[67][5] ), .ZN(n10653) );
  AOI22_X1 U14768 ( .A1(n30864), .A2(\xmem_data[68][5] ), .B1(n27501), .B2(
        \xmem_data[69][5] ), .ZN(n10652) );
  AOI22_X1 U14769 ( .A1(n27502), .A2(\xmem_data[70][5] ), .B1(n3217), .B2(
        \xmem_data[71][5] ), .ZN(n10651) );
  NAND4_X1 U14770 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10670) );
  AOI22_X1 U14771 ( .A1(n24632), .A2(\xmem_data[72][5] ), .B1(n27507), .B2(
        \xmem_data[73][5] ), .ZN(n10658) );
  AOI22_X1 U14772 ( .A1(n24534), .A2(\xmem_data[74][5] ), .B1(n13444), .B2(
        \xmem_data[75][5] ), .ZN(n10657) );
  AOI22_X1 U14773 ( .A1(n3140), .A2(\xmem_data[76][5] ), .B1(n27547), .B2(
        \xmem_data[77][5] ), .ZN(n10656) );
  AOI22_X1 U14774 ( .A1(n27508), .A2(\xmem_data[78][5] ), .B1(n25456), .B2(
        \xmem_data[79][5] ), .ZN(n10655) );
  NAND4_X1 U14775 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10669) );
  AOI22_X1 U14776 ( .A1(n27514), .A2(\xmem_data[80][5] ), .B1(n27513), .B2(
        \xmem_data[81][5] ), .ZN(n10662) );
  AOI22_X1 U14777 ( .A1(n27515), .A2(\xmem_data[82][5] ), .B1(n22674), .B2(
        \xmem_data[83][5] ), .ZN(n10661) );
  AOI22_X1 U14778 ( .A1(n28752), .A2(\xmem_data[84][5] ), .B1(n27516), .B2(
        \xmem_data[85][5] ), .ZN(n10660) );
  AOI22_X1 U14779 ( .A1(n20585), .A2(\xmem_data[86][5] ), .B1(n27518), .B2(
        \xmem_data[87][5] ), .ZN(n10659) );
  NAND4_X1 U14780 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10668) );
  AOI22_X1 U14781 ( .A1(n23802), .A2(\xmem_data[88][5] ), .B1(n27523), .B2(
        \xmem_data[89][5] ), .ZN(n10666) );
  AOI22_X1 U14782 ( .A1(n27524), .A2(\xmem_data[90][5] ), .B1(n30955), .B2(
        \xmem_data[91][5] ), .ZN(n10665) );
  AOI22_X1 U14783 ( .A1(n29573), .A2(\xmem_data[92][5] ), .B1(n27525), .B2(
        \xmem_data[93][5] ), .ZN(n10664) );
  AOI22_X1 U14784 ( .A1(n20734), .A2(\xmem_data[94][5] ), .B1(n27526), .B2(
        \xmem_data[95][5] ), .ZN(n10663) );
  NAND4_X1 U14785 ( .A1(n10666), .A2(n10665), .A3(n10664), .A4(n10663), .ZN(
        n10667) );
  OR4_X1 U14786 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10671) );
  AOI22_X1 U14787 ( .A1(n27496), .A2(n10672), .B1(n27494), .B2(n10671), .ZN(
        n10673) );
  XNOR2_X1 U14788 ( .A(n31642), .B(\fmem_data[20][5] ), .ZN(n33253) );
  AOI22_X1 U14789 ( .A1(n27498), .A2(\xmem_data[32][4] ), .B1(n24468), .B2(
        \xmem_data[33][4] ), .ZN(n10679) );
  AOI22_X1 U14790 ( .A1(n27500), .A2(\xmem_data[34][4] ), .B1(n27499), .B2(
        \xmem_data[35][4] ), .ZN(n10678) );
  AOI22_X1 U14791 ( .A1(n3384), .A2(\xmem_data[36][4] ), .B1(n27501), .B2(
        \xmem_data[37][4] ), .ZN(n10677) );
  AOI22_X1 U14792 ( .A1(n27502), .A2(\xmem_data[38][4] ), .B1(n3221), .B2(
        \xmem_data[39][4] ), .ZN(n10676) );
  NAND4_X1 U14793 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10695) );
  AOI22_X1 U14794 ( .A1(n23770), .A2(\xmem_data[40][4] ), .B1(n27507), .B2(
        \xmem_data[41][4] ), .ZN(n10683) );
  AOI22_X1 U14795 ( .A1(n25449), .A2(\xmem_data[42][4] ), .B1(n13444), .B2(
        \xmem_data[43][4] ), .ZN(n10682) );
  AOI22_X1 U14796 ( .A1(n3132), .A2(\xmem_data[44][4] ), .B1(n28510), .B2(
        \xmem_data[45][4] ), .ZN(n10681) );
  AOI22_X1 U14797 ( .A1(n27508), .A2(\xmem_data[46][4] ), .B1(n28415), .B2(
        \xmem_data[47][4] ), .ZN(n10680) );
  NAND4_X1 U14798 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10694) );
  AOI22_X1 U14799 ( .A1(n27514), .A2(\xmem_data[48][4] ), .B1(n27513), .B2(
        \xmem_data[49][4] ), .ZN(n10687) );
  AOI22_X1 U14800 ( .A1(n27515), .A2(\xmem_data[50][4] ), .B1(n30513), .B2(
        \xmem_data[51][4] ), .ZN(n10686) );
  AOI22_X1 U14801 ( .A1(n29605), .A2(\xmem_data[52][4] ), .B1(n27516), .B2(
        \xmem_data[53][4] ), .ZN(n10685) );
  AOI22_X1 U14802 ( .A1(n28096), .A2(\xmem_data[54][4] ), .B1(n27518), .B2(
        \xmem_data[55][4] ), .ZN(n10684) );
  NAND4_X1 U14803 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10693) );
  AOI22_X1 U14804 ( .A1(n31255), .A2(\xmem_data[56][4] ), .B1(n27523), .B2(
        \xmem_data[57][4] ), .ZN(n10691) );
  AOI22_X1 U14805 ( .A1(n27524), .A2(\xmem_data[58][4] ), .B1(n28291), .B2(
        \xmem_data[59][4] ), .ZN(n10690) );
  AOI22_X1 U14806 ( .A1(n20950), .A2(\xmem_data[60][4] ), .B1(n27525), .B2(
        \xmem_data[61][4] ), .ZN(n10689) );
  AOI22_X1 U14807 ( .A1(n29325), .A2(\xmem_data[62][4] ), .B1(n27526), .B2(
        \xmem_data[63][4] ), .ZN(n10688) );
  NAND4_X1 U14808 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10692) );
  OR4_X1 U14809 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10721) );
  AOI22_X1 U14810 ( .A1(n27568), .A2(\xmem_data[0][4] ), .B1(n27567), .B2(
        \xmem_data[1][4] ), .ZN(n10699) );
  AOI22_X1 U14811 ( .A1(n27564), .A2(\xmem_data[2][4] ), .B1(n27563), .B2(
        \xmem_data[3][4] ), .ZN(n10698) );
  AOI22_X1 U14812 ( .A1(n28718), .A2(\xmem_data[4][4] ), .B1(n3247), .B2(
        \xmem_data[5][4] ), .ZN(n10697) );
  AOI22_X1 U14813 ( .A1(n30592), .A2(\xmem_data[6][4] ), .B1(n3221), .B2(
        \xmem_data[7][4] ), .ZN(n10696) );
  AOI22_X1 U14814 ( .A1(n3342), .A2(\xmem_data[10][4] ), .B1(n27550), .B2(
        \xmem_data[11][4] ), .ZN(n10706) );
  AOI22_X1 U14815 ( .A1(n27551), .A2(\xmem_data[14][4] ), .B1(n3358), .B2(
        \xmem_data[15][4] ), .ZN(n10700) );
  INV_X1 U14816 ( .A(n10700), .ZN(n10704) );
  AND2_X1 U14817 ( .A1(n3375), .A2(\xmem_data[12][4] ), .ZN(n10703) );
  AOI22_X1 U14818 ( .A1(n31368), .A2(\xmem_data[8][4] ), .B1(n13469), .B2(
        \xmem_data[9][4] ), .ZN(n10701) );
  INV_X1 U14819 ( .A(n10701), .ZN(n10702) );
  NOR3_X1 U14820 ( .A1(n10704), .A2(n10703), .A3(n10702), .ZN(n10705) );
  NAND2_X1 U14821 ( .A1(n10706), .A2(n10705), .ZN(n10718) );
  AOI22_X1 U14822 ( .A1(n20716), .A2(\xmem_data[16][4] ), .B1(n27535), .B2(
        \xmem_data[17][4] ), .ZN(n10710) );
  AOI22_X1 U14823 ( .A1(n29023), .A2(\xmem_data[18][4] ), .B1(n27536), .B2(
        \xmem_data[19][4] ), .ZN(n10709) );
  AOI22_X1 U14824 ( .A1(n28752), .A2(\xmem_data[20][4] ), .B1(n20938), .B2(
        \xmem_data[21][4] ), .ZN(n10708) );
  AOI22_X1 U14825 ( .A1(n25573), .A2(\xmem_data[22][4] ), .B1(n24645), .B2(
        \xmem_data[23][4] ), .ZN(n10707) );
  NAND4_X1 U14826 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(
        n10716) );
  AOI22_X1 U14827 ( .A1(n20942), .A2(\xmem_data[24][4] ), .B1(n13452), .B2(
        \xmem_data[25][4] ), .ZN(n10714) );
  AOI22_X1 U14828 ( .A1(n28428), .A2(\xmem_data[26][4] ), .B1(n23778), .B2(
        \xmem_data[27][4] ), .ZN(n10713) );
  AOI22_X1 U14829 ( .A1(n29297), .A2(\xmem_data[28][4] ), .B1(n22685), .B2(
        \xmem_data[29][4] ), .ZN(n10712) );
  AOI22_X1 U14830 ( .A1(n27542), .A2(\xmem_data[30][4] ), .B1(n17003), .B2(
        \xmem_data[31][4] ), .ZN(n10711) );
  NAND4_X1 U14831 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10715) );
  OR3_X1 U14832 ( .A1(n10716), .A2(n10715), .A3(n3976), .ZN(n10717) );
  NOR2_X1 U14833 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  INV_X1 U14834 ( .A(n19410), .ZN(n27573) );
  AOI21_X1 U14835 ( .B1(n3786), .B2(n10719), .A(n27573), .ZN(n10720) );
  AOI21_X1 U14836 ( .B1(n10721), .B2(n27577), .A(n10720), .ZN(n10766) );
  AOI22_X1 U14837 ( .A1(n28036), .A2(\xmem_data[96][4] ), .B1(n27435), .B2(
        \xmem_data[97][4] ), .ZN(n10725) );
  AOI22_X1 U14838 ( .A1(n27436), .A2(\xmem_data[98][4] ), .B1(n31262), .B2(
        \xmem_data[99][4] ), .ZN(n10724) );
  AOI22_X1 U14839 ( .A1(n25443), .A2(\xmem_data[100][4] ), .B1(n27437), .B2(
        \xmem_data[101][4] ), .ZN(n10723) );
  AOI22_X1 U14840 ( .A1(n27439), .A2(\xmem_data[102][4] ), .B1(n3222), .B2(
        \xmem_data[103][4] ), .ZN(n10722) );
  NAND4_X1 U14841 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(
        n10741) );
  AOI22_X1 U14842 ( .A1(n27445), .A2(\xmem_data[104][4] ), .B1(n27444), .B2(
        \xmem_data[105][4] ), .ZN(n10729) );
  AOI22_X1 U14843 ( .A1(n22758), .A2(\xmem_data[106][4] ), .B1(n27903), .B2(
        \xmem_data[107][4] ), .ZN(n10728) );
  AOI22_X1 U14844 ( .A1(n3137), .A2(\xmem_data[108][4] ), .B1(n27446), .B2(
        \xmem_data[109][4] ), .ZN(n10727) );
  AOI22_X1 U14845 ( .A1(n27447), .A2(\xmem_data[110][4] ), .B1(n20546), .B2(
        \xmem_data[111][4] ), .ZN(n10726) );
  NAND4_X1 U14846 ( .A1(n10729), .A2(n10728), .A3(n10727), .A4(n10726), .ZN(
        n10740) );
  AOI22_X1 U14847 ( .A1(n27453), .A2(\xmem_data[112][4] ), .B1(n27452), .B2(
        \xmem_data[113][4] ), .ZN(n10733) );
  AOI22_X1 U14848 ( .A1(n28298), .A2(\xmem_data[114][4] ), .B1(n25458), .B2(
        \xmem_data[115][4] ), .ZN(n10732) );
  AOI22_X1 U14849 ( .A1(n27755), .A2(\xmem_data[116][4] ), .B1(n27454), .B2(
        \xmem_data[117][4] ), .ZN(n10731) );
  AOI22_X1 U14850 ( .A1(n13149), .A2(\xmem_data[118][4] ), .B1(n28427), .B2(
        \xmem_data[119][4] ), .ZN(n10730) );
  NAND4_X1 U14851 ( .A1(n10733), .A2(n10732), .A3(n10731), .A4(n10730), .ZN(
        n10739) );
  AOI22_X1 U14852 ( .A1(n29012), .A2(\xmem_data[120][4] ), .B1(n27460), .B2(
        \xmem_data[121][4] ), .ZN(n10737) );
  AOI22_X1 U14853 ( .A1(n27462), .A2(\xmem_data[122][4] ), .B1(n27461), .B2(
        \xmem_data[123][4] ), .ZN(n10736) );
  AOI22_X1 U14854 ( .A1(n20984), .A2(\xmem_data[124][4] ), .B1(n30599), .B2(
        \xmem_data[125][4] ), .ZN(n10735) );
  AOI22_X1 U14855 ( .A1(n20552), .A2(\xmem_data[126][4] ), .B1(n27463), .B2(
        \xmem_data[127][4] ), .ZN(n10734) );
  NAND4_X1 U14856 ( .A1(n10737), .A2(n10736), .A3(n10735), .A4(n10734), .ZN(
        n10738) );
  OR4_X1 U14857 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10764) );
  AOI22_X1 U14858 ( .A1(n27498), .A2(\xmem_data[64][4] ), .B1(n29125), .B2(
        \xmem_data[65][4] ), .ZN(n10746) );
  AOI22_X1 U14859 ( .A1(n27500), .A2(\xmem_data[66][4] ), .B1(n27499), .B2(
        \xmem_data[67][4] ), .ZN(n10745) );
  AOI22_X1 U14860 ( .A1(n21308), .A2(\xmem_data[68][4] ), .B1(n27501), .B2(
        \xmem_data[69][4] ), .ZN(n10744) );
  AND2_X1 U14861 ( .A1(n3218), .A2(\xmem_data[71][4] ), .ZN(n10742) );
  AOI21_X1 U14862 ( .B1(n27502), .B2(\xmem_data[70][4] ), .A(n10742), .ZN(
        n10743) );
  NAND4_X1 U14863 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10762) );
  AOI22_X1 U14864 ( .A1(n21050), .A2(\xmem_data[88][4] ), .B1(n27523), .B2(
        \xmem_data[89][4] ), .ZN(n10750) );
  AOI22_X1 U14865 ( .A1(n27524), .A2(\xmem_data[90][4] ), .B1(n24222), .B2(
        \xmem_data[91][4] ), .ZN(n10749) );
  AOI22_X1 U14866 ( .A1(n17004), .A2(\xmem_data[92][4] ), .B1(n27525), .B2(
        \xmem_data[93][4] ), .ZN(n10748) );
  AOI22_X1 U14867 ( .A1(n24685), .A2(\xmem_data[94][4] ), .B1(n27526), .B2(
        \xmem_data[95][4] ), .ZN(n10747) );
  NAND4_X1 U14868 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10761) );
  AOI22_X1 U14869 ( .A1(n27514), .A2(\xmem_data[80][4] ), .B1(n27513), .B2(
        \xmem_data[81][4] ), .ZN(n10754) );
  AOI22_X1 U14870 ( .A1(n27515), .A2(\xmem_data[82][4] ), .B1(n24160), .B2(
        \xmem_data[83][4] ), .ZN(n10753) );
  AOI22_X1 U14871 ( .A1(n27945), .A2(\xmem_data[84][4] ), .B1(n27516), .B2(
        \xmem_data[85][4] ), .ZN(n10752) );
  AOI22_X1 U14872 ( .A1(n23717), .A2(\xmem_data[86][4] ), .B1(n27518), .B2(
        \xmem_data[87][4] ), .ZN(n10751) );
  NAND4_X1 U14873 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10760) );
  AOI22_X1 U14874 ( .A1(n30964), .A2(\xmem_data[72][4] ), .B1(n27507), .B2(
        \xmem_data[73][4] ), .ZN(n10758) );
  AOI22_X1 U14875 ( .A1(n23741), .A2(\xmem_data[74][4] ), .B1(n13444), .B2(
        \xmem_data[75][4] ), .ZN(n10757) );
  AOI22_X1 U14876 ( .A1(n3134), .A2(\xmem_data[76][4] ), .B1(n25514), .B2(
        \xmem_data[77][4] ), .ZN(n10756) );
  AOI22_X1 U14877 ( .A1(n27508), .A2(\xmem_data[78][4] ), .B1(n3357), .B2(
        \xmem_data[79][4] ), .ZN(n10755) );
  NAND4_X1 U14878 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10759) );
  OR4_X1 U14879 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  AOI22_X1 U14880 ( .A1(n10764), .A2(n27496), .B1(n10763), .B2(n27494), .ZN(
        n10765) );
  NAND2_X1 U14881 ( .A1(n10766), .A2(n10765), .ZN(n31900) );
  XNOR2_X1 U14882 ( .A(n31900), .B(\fmem_data[20][5] ), .ZN(n31986) );
  XOR2_X1 U14883 ( .A(\fmem_data[20][5] ), .B(\fmem_data[20][4] ), .Z(n10767)
         );
  OAI22_X1 U14884 ( .A1(n33253), .A2(n35036), .B1(n31986), .B2(n35037), .ZN(
        n17750) );
  AOI22_X1 U14885 ( .A1(n29395), .A2(\xmem_data[64][7] ), .B1(n26884), .B2(
        \xmem_data[65][7] ), .ZN(n10771) );
  AOI22_X1 U14886 ( .A1(n29438), .A2(\xmem_data[66][7] ), .B1(n30666), .B2(
        \xmem_data[67][7] ), .ZN(n10770) );
  AOI22_X1 U14887 ( .A1(n3166), .A2(\xmem_data[68][7] ), .B1(n3191), .B2(
        \xmem_data[69][7] ), .ZN(n10769) );
  AOI22_X1 U14888 ( .A1(n23901), .A2(\xmem_data[70][7] ), .B1(n29439), .B2(
        \xmem_data[71][7] ), .ZN(n10768) );
  NAND4_X1 U14889 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10777) );
  NAND2_X1 U14890 ( .A1(n29433), .A2(\xmem_data[84][7] ), .ZN(n10775) );
  AOI22_X1 U14891 ( .A1(n29449), .A2(\xmem_data[82][7] ), .B1(n23754), .B2(
        \xmem_data[83][7] ), .ZN(n10774) );
  AOI22_X1 U14892 ( .A1(n29447), .A2(\xmem_data[80][7] ), .B1(n27723), .B2(
        \xmem_data[81][7] ), .ZN(n10773) );
  NAND2_X1 U14893 ( .A1(n30222), .A2(\xmem_data[85][7] ), .ZN(n10772) );
  NAND4_X1 U14894 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10776) );
  NOR2_X1 U14895 ( .A1(n10777), .A2(n10776), .ZN(n10788) );
  AOI22_X1 U14896 ( .A1(n30280), .A2(\xmem_data[88][7] ), .B1(n30217), .B2(
        \xmem_data[89][7] ), .ZN(n10781) );
  AOI22_X1 U14897 ( .A1(n29450), .A2(\xmem_data[90][7] ), .B1(n29350), .B2(
        \xmem_data[91][7] ), .ZN(n10780) );
  AOI22_X1 U14898 ( .A1(n29801), .A2(\xmem_data[92][7] ), .B1(n3368), .B2(
        \xmem_data[93][7] ), .ZN(n10779) );
  AOI22_X1 U14899 ( .A1(n7282), .A2(\xmem_data[94][7] ), .B1(n29451), .B2(
        \xmem_data[95][7] ), .ZN(n10778) );
  AOI22_X1 U14900 ( .A1(n30279), .A2(\xmem_data[86][7] ), .B1(n29431), .B2(
        \xmem_data[87][7] ), .ZN(n10786) );
  AOI22_X1 U14901 ( .A1(n29547), .A2(\xmem_data[72][7] ), .B1(n29640), .B2(
        \xmem_data[73][7] ), .ZN(n10785) );
  AOI22_X1 U14902 ( .A1(n29461), .A2(\xmem_data[74][7] ), .B1(n3151), .B2(
        \xmem_data[75][7] ), .ZN(n10784) );
  AOI22_X1 U14903 ( .A1(n29463), .A2(\xmem_data[76][7] ), .B1(n29462), .B2(
        \xmem_data[77][7] ), .ZN(n10783) );
  AOI22_X1 U14904 ( .A1(n29464), .A2(\xmem_data[78][7] ), .B1(n20826), .B2(
        \xmem_data[79][7] ), .ZN(n10782) );
  NAND4_X1 U14905 ( .A1(n10788), .A2(n10787), .A3(n10786), .A4(n3763), .ZN(
        n10812) );
  AOI22_X1 U14906 ( .A1(n29419), .A2(\xmem_data[112][7] ), .B1(n29418), .B2(
        \xmem_data[113][7] ), .ZN(n10793) );
  AOI22_X1 U14907 ( .A1(n29420), .A2(\xmem_data[114][7] ), .B1(n25725), .B2(
        \xmem_data[115][7] ), .ZN(n10792) );
  AOI22_X1 U14908 ( .A1(n30708), .A2(\xmem_data[116][7] ), .B1(n26510), .B2(
        \xmem_data[117][7] ), .ZN(n10791) );
  AND2_X1 U14909 ( .A1(n29422), .A2(\xmem_data[119][7] ), .ZN(n10789) );
  AOI21_X1 U14910 ( .B1(n29628), .B2(\xmem_data[118][7] ), .A(n10789), .ZN(
        n10790) );
  NAND4_X1 U14911 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10810) );
  AOI22_X1 U14912 ( .A1(n27754), .A2(\xmem_data[96][7] ), .B1(n29648), .B2(
        \xmem_data[97][7] ), .ZN(n10797) );
  AOI22_X1 U14913 ( .A1(n29397), .A2(\xmem_data[98][7] ), .B1(n23795), .B2(
        \xmem_data[99][7] ), .ZN(n10796) );
  AOI22_X1 U14914 ( .A1(n3165), .A2(\xmem_data[100][7] ), .B1(n3185), .B2(
        \xmem_data[101][7] ), .ZN(n10795) );
  AOI22_X1 U14915 ( .A1(n30684), .A2(\xmem_data[102][7] ), .B1(n29410), .B2(
        \xmem_data[103][7] ), .ZN(n10794) );
  NAND4_X1 U14916 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n10809) );
  AOI22_X1 U14917 ( .A1(n29590), .A2(\xmem_data[124][7] ), .B1(n28238), .B2(
        \xmem_data[125][7] ), .ZN(n10801) );
  AOI22_X1 U14918 ( .A1(n29402), .A2(\xmem_data[122][7] ), .B1(n29350), .B2(
        \xmem_data[123][7] ), .ZN(n10800) );
  AOI22_X1 U14919 ( .A1(n29400), .A2(\xmem_data[120][7] ), .B1(n29629), .B2(
        \xmem_data[121][7] ), .ZN(n10799) );
  AOI22_X1 U14920 ( .A1(n29404), .A2(\xmem_data[126][7] ), .B1(n29403), .B2(
        \xmem_data[127][7] ), .ZN(n10798) );
  NAND4_X1 U14921 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10808) );
  BUF_X1 U14922 ( .A(n10802), .Z(n30198) );
  AOI22_X1 U14923 ( .A1(n29815), .A2(\xmem_data[104][7] ), .B1(n30266), .B2(
        \xmem_data[105][7] ), .ZN(n10806) );
  AOI22_X1 U14924 ( .A1(n29380), .A2(\xmem_data[106][7] ), .B1(n29379), .B2(
        \xmem_data[107][7] ), .ZN(n10805) );
  AOI22_X1 U14925 ( .A1(n29382), .A2(\xmem_data[108][7] ), .B1(n29381), .B2(
        \xmem_data[109][7] ), .ZN(n10804) );
  AOI22_X1 U14926 ( .A1(n29384), .A2(\xmem_data[110][7] ), .B1(n29383), .B2(
        \xmem_data[111][7] ), .ZN(n10803) );
  NAND4_X1 U14927 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10807) );
  OR4_X1 U14928 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10811) );
  AOI22_X1 U14929 ( .A1(n10812), .A2(n29376), .B1(n29428), .B2(n10811), .ZN(
        n10856) );
  AOI22_X1 U14930 ( .A1(n30635), .A2(\xmem_data[32][7] ), .B1(n30634), .B2(
        \xmem_data[33][7] ), .ZN(n10816) );
  AOI22_X1 U14931 ( .A1(n29438), .A2(\xmem_data[34][7] ), .B1(n28752), .B2(
        \xmem_data[35][7] ), .ZN(n10815) );
  AOI22_X1 U14932 ( .A1(n3163), .A2(\xmem_data[36][7] ), .B1(n3187), .B2(
        \xmem_data[37][7] ), .ZN(n10814) );
  AOI22_X1 U14933 ( .A1(n30062), .A2(\xmem_data[38][7] ), .B1(n29439), .B2(
        \xmem_data[39][7] ), .ZN(n10813) );
  NAND4_X1 U14934 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n10832) );
  AOI22_X1 U14935 ( .A1(n27713), .A2(\xmem_data[40][7] ), .B1(n29721), .B2(
        \xmem_data[41][7] ), .ZN(n10820) );
  AOI22_X1 U14936 ( .A1(n29461), .A2(\xmem_data[42][7] ), .B1(n3151), .B2(
        \xmem_data[43][7] ), .ZN(n10819) );
  AOI22_X1 U14937 ( .A1(n29463), .A2(\xmem_data[44][7] ), .B1(n29462), .B2(
        \xmem_data[45][7] ), .ZN(n10818) );
  AOI22_X1 U14938 ( .A1(n29464), .A2(\xmem_data[46][7] ), .B1(n27852), .B2(
        \xmem_data[47][7] ), .ZN(n10817) );
  NAND4_X1 U14939 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        n10831) );
  AOI22_X1 U14940 ( .A1(n29447), .A2(\xmem_data[48][7] ), .B1(n27812), .B2(
        \xmem_data[49][7] ), .ZN(n10824) );
  AOI22_X1 U14941 ( .A1(n29449), .A2(\xmem_data[50][7] ), .B1(n28973), .B2(
        \xmem_data[51][7] ), .ZN(n10823) );
  AOI22_X1 U14942 ( .A1(n27741), .A2(\xmem_data[52][7] ), .B1(n28766), .B2(
        \xmem_data[53][7] ), .ZN(n10822) );
  AOI22_X1 U14943 ( .A1(n27740), .A2(\xmem_data[54][7] ), .B1(n29431), .B2(
        \xmem_data[55][7] ), .ZN(n10821) );
  NAND4_X1 U14944 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10830) );
  AOI22_X1 U14945 ( .A1(n30280), .A2(\xmem_data[56][7] ), .B1(n29761), .B2(
        \xmem_data[57][7] ), .ZN(n10828) );
  AOI22_X1 U14946 ( .A1(n29450), .A2(\xmem_data[58][7] ), .B1(n3134), .B2(
        \xmem_data[59][7] ), .ZN(n10827) );
  AOI22_X1 U14947 ( .A1(n29590), .A2(\xmem_data[60][7] ), .B1(n29646), .B2(
        \xmem_data[61][7] ), .ZN(n10826) );
  AOI22_X1 U14948 ( .A1(n29802), .A2(\xmem_data[62][7] ), .B1(n29451), .B2(
        \xmem_data[63][7] ), .ZN(n10825) );
  NAND4_X1 U14949 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  AOI22_X1 U14950 ( .A1(n27811), .A2(\xmem_data[0][7] ), .B1(n29592), .B2(
        \xmem_data[1][7] ), .ZN(n10836) );
  AOI22_X1 U14951 ( .A1(n29438), .A2(\xmem_data[2][7] ), .B1(n27755), .B2(
        \xmem_data[3][7] ), .ZN(n10835) );
  AOI22_X1 U14952 ( .A1(n3167), .A2(\xmem_data[4][7] ), .B1(n3182), .B2(
        \xmem_data[5][7] ), .ZN(n10834) );
  AOI22_X1 U14953 ( .A1(n28689), .A2(\xmem_data[6][7] ), .B1(n23777), .B2(
        \xmem_data[7][7] ), .ZN(n10833) );
  NAND4_X1 U14954 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10852) );
  AOI22_X1 U14955 ( .A1(n27713), .A2(\xmem_data[8][7] ), .B1(n29640), .B2(
        \xmem_data[9][7] ), .ZN(n10840) );
  AOI22_X1 U14956 ( .A1(n29461), .A2(\xmem_data[10][7] ), .B1(n3301), .B2(
        \xmem_data[11][7] ), .ZN(n10839) );
  AOI22_X1 U14957 ( .A1(n29463), .A2(\xmem_data[12][7] ), .B1(n29462), .B2(
        \xmem_data[13][7] ), .ZN(n10838) );
  AOI22_X1 U14958 ( .A1(n29489), .A2(\xmem_data[14][7] ), .B1(n20985), .B2(
        \xmem_data[15][7] ), .ZN(n10837) );
  NAND4_X1 U14959 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10851) );
  AOI22_X1 U14960 ( .A1(n28765), .A2(\xmem_data[16][7] ), .B1(n29497), .B2(
        \xmem_data[17][7] ), .ZN(n10844) );
  AOI22_X1 U14961 ( .A1(n29499), .A2(\xmem_data[18][7] ), .B1(n3383), .B2(
        \xmem_data[19][7] ), .ZN(n10843) );
  AOI22_X1 U14962 ( .A1(n30223), .A2(\xmem_data[20][7] ), .B1(n28206), .B2(
        \xmem_data[21][7] ), .ZN(n10842) );
  AOI22_X1 U14963 ( .A1(n29699), .A2(\xmem_data[22][7] ), .B1(n29494), .B2(
        \xmem_data[23][7] ), .ZN(n10841) );
  NAND4_X1 U14964 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        n10850) );
  AOI22_X1 U14965 ( .A1(n29647), .A2(\xmem_data[28][7] ), .B1(n29704), .B2(
        \xmem_data[29][7] ), .ZN(n10848) );
  AOI22_X1 U14966 ( .A1(n29501), .A2(\xmem_data[26][7] ), .B1(n3282), .B2(
        \xmem_data[27][7] ), .ZN(n10847) );
  AOI22_X1 U14967 ( .A1(n28787), .A2(\xmem_data[24][7] ), .B1(n3169), .B2(
        \xmem_data[25][7] ), .ZN(n10846) );
  AOI22_X1 U14968 ( .A1(n29500), .A2(\xmem_data[30][7] ), .B1(n30663), .B2(
        \xmem_data[31][7] ), .ZN(n10845) );
  NAND4_X1 U14969 ( .A1(n10848), .A2(n10847), .A3(n10846), .A4(n10845), .ZN(
        n10849) );
  OR4_X2 U14970 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10853) );
  AOI22_X1 U14971 ( .A1(n29471), .A2(n10854), .B1(n29511), .B2(n10853), .ZN(
        n10855) );
  NAND2_X1 U14972 ( .A1(n10856), .A2(n10855), .ZN(n35240) );
  XNOR2_X1 U14973 ( .A(n35240), .B(\fmem_data[3][3] ), .ZN(n30442) );
  AOI22_X1 U14974 ( .A1(n30766), .A2(\xmem_data[72][6] ), .B1(n30170), .B2(
        \xmem_data[73][6] ), .ZN(n10860) );
  AOI22_X1 U14975 ( .A1(n29461), .A2(\xmem_data[74][6] ), .B1(n3151), .B2(
        \xmem_data[75][6] ), .ZN(n10859) );
  AOI22_X1 U14976 ( .A1(n29463), .A2(\xmem_data[76][6] ), .B1(n29462), .B2(
        \xmem_data[77][6] ), .ZN(n10858) );
  AOI22_X1 U14977 ( .A1(n29464), .A2(\xmem_data[78][6] ), .B1(n29327), .B2(
        \xmem_data[79][6] ), .ZN(n10857) );
  NAND4_X1 U14978 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10865) );
  AND2_X1 U14979 ( .A1(n29697), .A2(\xmem_data[85][6] ), .ZN(n10862) );
  AOI21_X1 U14980 ( .B1(n27710), .B2(\xmem_data[84][6] ), .A(n10862), .ZN(
        n10863) );
  INV_X1 U14981 ( .A(n10863), .ZN(n10864) );
  NOR2_X1 U14982 ( .A1(n10865), .A2(n10864), .ZN(n10872) );
  INV_X1 U14983 ( .A(n10866), .ZN(n10870) );
  AOI22_X1 U14984 ( .A1(n29449), .A2(\xmem_data[82][6] ), .B1(n25443), .B2(
        \xmem_data[83][6] ), .ZN(n10868) );
  AOI22_X1 U14985 ( .A1(n29447), .A2(\xmem_data[80][6] ), .B1(n27812), .B2(
        \xmem_data[81][6] ), .ZN(n10867) );
  NAND2_X1 U14986 ( .A1(n10868), .A2(n10867), .ZN(n10869) );
  NOR2_X1 U14987 ( .A1(n10870), .A2(n10869), .ZN(n10871) );
  NAND2_X1 U14988 ( .A1(n10872), .A2(n10871), .ZN(n10883) );
  AOI22_X1 U14989 ( .A1(n3174), .A2(\xmem_data[64][6] ), .B1(n29739), .B2(
        \xmem_data[65][6] ), .ZN(n10876) );
  AOI22_X1 U14990 ( .A1(n29438), .A2(n20682), .B1(n3158), .B2(
        \xmem_data[67][6] ), .ZN(n10875) );
  AOI22_X1 U14991 ( .A1(n3164), .A2(\xmem_data[68][6] ), .B1(n3188), .B2(
        \xmem_data[69][6] ), .ZN(n10874) );
  AOI22_X1 U14992 ( .A1(n30075), .A2(\xmem_data[70][6] ), .B1(n29439), .B2(
        \xmem_data[71][6] ), .ZN(n10873) );
  AOI22_X1 U14993 ( .A1(n27771), .A2(\xmem_data[88][6] ), .B1(n30217), .B2(
        \xmem_data[89][6] ), .ZN(n10880) );
  AOI22_X1 U14994 ( .A1(n29450), .A2(\xmem_data[90][6] ), .B1(n3135), .B2(
        \xmem_data[91][6] ), .ZN(n10879) );
  AOI22_X1 U14995 ( .A1(n29602), .A2(\xmem_data[92][6] ), .B1(n29389), .B2(
        \xmem_data[93][6] ), .ZN(n10878) );
  AOI22_X1 U14996 ( .A1(n29500), .A2(\xmem_data[94][6] ), .B1(n29451), .B2(
        \xmem_data[95][6] ), .ZN(n10877) );
  NAND2_X1 U14997 ( .A1(n3775), .A2(n10881), .ZN(n10882) );
  OAI21_X1 U14998 ( .B1(n10883), .B2(n10882), .A(n29376), .ZN(n10942) );
  AOI22_X1 U14999 ( .A1(n29447), .A2(\xmem_data[48][6] ), .B1(n29418), .B2(
        \xmem_data[49][6] ), .ZN(n10887) );
  AOI22_X1 U15000 ( .A1(n29449), .A2(\xmem_data[50][6] ), .B1(n3153), .B2(
        \xmem_data[51][6] ), .ZN(n10886) );
  AOI22_X1 U15001 ( .A1(n29626), .A2(\xmem_data[52][6] ), .B1(n30775), .B2(
        \xmem_data[53][6] ), .ZN(n10885) );
  AOI22_X1 U15002 ( .A1(n28700), .A2(\xmem_data[54][6] ), .B1(n29431), .B2(
        \xmem_data[55][6] ), .ZN(n10884) );
  NAND4_X1 U15003 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10903) );
  AOI22_X1 U15004 ( .A1(n30280), .A2(\xmem_data[56][6] ), .B1(n29761), .B2(
        \xmem_data[57][6] ), .ZN(n10891) );
  AOI22_X1 U15005 ( .A1(n29450), .A2(\xmem_data[58][6] ), .B1(n3375), .B2(
        \xmem_data[59][6] ), .ZN(n10890) );
  AOI22_X1 U15006 ( .A1(n30191), .A2(\xmem_data[60][6] ), .B1(n28145), .B2(
        \xmem_data[61][6] ), .ZN(n10889) );
  AOI22_X1 U15007 ( .A1(n29500), .A2(\xmem_data[62][6] ), .B1(n29451), .B2(
        \xmem_data[63][6] ), .ZN(n10888) );
  NAND4_X1 U15008 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10902) );
  AOI22_X1 U15009 ( .A1(n30665), .A2(\xmem_data[32][6] ), .B1(n30249), .B2(
        \xmem_data[33][6] ), .ZN(n10895) );
  AOI22_X1 U15010 ( .A1(n29438), .A2(\xmem_data[34][6] ), .B1(n27755), .B2(
        \xmem_data[35][6] ), .ZN(n10894) );
  AOI22_X1 U15011 ( .A1(n3167), .A2(\xmem_data[36][6] ), .B1(n3182), .B2(
        \xmem_data[37][6] ), .ZN(n10893) );
  AOI22_X1 U15012 ( .A1(n30062), .A2(\xmem_data[38][6] ), .B1(n29439), .B2(
        \xmem_data[39][6] ), .ZN(n10892) );
  NAND4_X1 U15013 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10901) );
  AOI22_X1 U15014 ( .A1(n29547), .A2(\xmem_data[40][6] ), .B1(n29721), .B2(
        \xmem_data[41][6] ), .ZN(n10899) );
  AOI22_X1 U15015 ( .A1(n29461), .A2(\xmem_data[42][6] ), .B1(n3151), .B2(
        \xmem_data[43][6] ), .ZN(n10898) );
  AOI22_X1 U15016 ( .A1(n29463), .A2(\xmem_data[44][6] ), .B1(n29462), .B2(
        \xmem_data[45][6] ), .ZN(n10897) );
  AOI22_X1 U15017 ( .A1(n29464), .A2(\xmem_data[46][6] ), .B1(n28241), .B2(
        \xmem_data[47][6] ), .ZN(n10896) );
  NAND4_X1 U15018 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10900) );
  NAND2_X1 U15019 ( .A1(n10904), .A2(n29471), .ZN(n10941) );
  AOI22_X1 U15020 ( .A1(n3249), .A2(\xmem_data[28][6] ), .B1(n3369), .B2(
        \xmem_data[29][6] ), .ZN(n10908) );
  AOI22_X1 U15021 ( .A1(n29501), .A2(\xmem_data[26][6] ), .B1(n29350), .B2(
        \xmem_data[27][6] ), .ZN(n10907) );
  AOI22_X1 U15022 ( .A1(n29674), .A2(\xmem_data[24][6] ), .B1(n27833), .B2(
        \xmem_data[25][6] ), .ZN(n10906) );
  AOI22_X1 U15023 ( .A1(n29500), .A2(\xmem_data[30][6] ), .B1(n29591), .B2(
        \xmem_data[31][6] ), .ZN(n10905) );
  AOI22_X1 U15024 ( .A1(n28717), .A2(\xmem_data[16][6] ), .B1(n29497), .B2(
        \xmem_data[17][6] ), .ZN(n10912) );
  AOI22_X1 U15025 ( .A1(n29499), .A2(\xmem_data[18][6] ), .B1(n3149), .B2(
        \xmem_data[19][6] ), .ZN(n10911) );
  AOI22_X1 U15026 ( .A1(n29626), .A2(\xmem_data[20][6] ), .B1(n30707), .B2(
        \xmem_data[21][6] ), .ZN(n10910) );
  AOI22_X1 U15027 ( .A1(n29628), .A2(\xmem_data[22][6] ), .B1(n29494), .B2(
        \xmem_data[23][6] ), .ZN(n10909) );
  AOI22_X1 U15028 ( .A1(n30635), .A2(\xmem_data[0][6] ), .B1(n28778), .B2(
        \xmem_data[1][6] ), .ZN(n10916) );
  AOI22_X1 U15029 ( .A1(n29475), .A2(\xmem_data[2][6] ), .B1(n28231), .B2(
        \xmem_data[3][6] ), .ZN(n10915) );
  AOI22_X1 U15030 ( .A1(n3167), .A2(\xmem_data[4][6] ), .B1(n3186), .B2(
        \xmem_data[5][6] ), .ZN(n10914) );
  AOI22_X1 U15031 ( .A1(n30684), .A2(\xmem_data[6][6] ), .B1(n28232), .B2(
        \xmem_data[7][6] ), .ZN(n10913) );
  AOI22_X1 U15032 ( .A1(n30198), .A2(\xmem_data[8][6] ), .B1(n29721), .B2(
        \xmem_data[9][6] ), .ZN(n10920) );
  AOI22_X1 U15033 ( .A1(n29461), .A2(\xmem_data[10][6] ), .B1(n3151), .B2(
        \xmem_data[11][6] ), .ZN(n10919) );
  AOI22_X1 U15034 ( .A1(n29463), .A2(\xmem_data[12][6] ), .B1(n29723), .B2(
        \xmem_data[13][6] ), .ZN(n10918) );
  AOI22_X1 U15035 ( .A1(n29489), .A2(\xmem_data[14][6] ), .B1(n20826), .B2(
        \xmem_data[15][6] ), .ZN(n10917) );
  NAND2_X1 U15036 ( .A1(n10921), .A2(n29511), .ZN(n10940) );
  AOI22_X1 U15037 ( .A1(n29419), .A2(\xmem_data[112][6] ), .B1(n29418), .B2(
        \xmem_data[113][6] ), .ZN(n10925) );
  AOI22_X1 U15038 ( .A1(n29420), .A2(\xmem_data[114][6] ), .B1(n3449), .B2(
        \xmem_data[115][6] ), .ZN(n10924) );
  AOI22_X1 U15039 ( .A1(n28734), .A2(\xmem_data[116][6] ), .B1(n29753), .B2(
        \xmem_data[117][6] ), .ZN(n10923) );
  AOI22_X1 U15040 ( .A1(n30279), .A2(\xmem_data[118][6] ), .B1(n29422), .B2(
        \xmem_data[119][6] ), .ZN(n10922) );
  AOI22_X1 U15041 ( .A1(n29400), .A2(\xmem_data[120][6] ), .B1(n28208), .B2(
        \xmem_data[121][6] ), .ZN(n10929) );
  AOI22_X1 U15042 ( .A1(n29402), .A2(\xmem_data[122][6] ), .B1(n3134), .B2(
        \xmem_data[123][6] ), .ZN(n10928) );
  AOI22_X1 U15043 ( .A1(n29801), .A2(\xmem_data[124][6] ), .B1(n29704), .B2(
        \xmem_data[125][6] ), .ZN(n10927) );
  AOI22_X1 U15044 ( .A1(n29404), .A2(\xmem_data[126][6] ), .B1(n29403), .B2(
        \xmem_data[127][6] ), .ZN(n10926) );
  AOI22_X1 U15045 ( .A1(n30745), .A2(\xmem_data[96][6] ), .B1(n28110), .B2(
        \xmem_data[97][6] ), .ZN(n10933) );
  AOI22_X1 U15046 ( .A1(n29397), .A2(\xmem_data[98][6] ), .B1(n28091), .B2(
        \xmem_data[99][6] ), .ZN(n10932) );
  AOI22_X1 U15047 ( .A1(n3160), .A2(\xmem_data[100][6] ), .B1(n3190), .B2(
        \xmem_data[101][6] ), .ZN(n10931) );
  AOI22_X1 U15048 ( .A1(n30075), .A2(\xmem_data[102][6] ), .B1(n29410), .B2(
        \xmem_data[103][6] ), .ZN(n10930) );
  AOI22_X1 U15049 ( .A1(n30766), .A2(\xmem_data[104][6] ), .B1(n30685), .B2(
        \xmem_data[105][6] ), .ZN(n10937) );
  AOI22_X1 U15050 ( .A1(n29380), .A2(\xmem_data[106][6] ), .B1(n29379), .B2(
        \xmem_data[107][6] ), .ZN(n10936) );
  AOI22_X1 U15051 ( .A1(n29382), .A2(\xmem_data[108][6] ), .B1(n29381), .B2(
        \xmem_data[109][6] ), .ZN(n10935) );
  AOI22_X1 U15052 ( .A1(n29384), .A2(\xmem_data[110][6] ), .B1(n29383), .B2(
        \xmem_data[111][6] ), .ZN(n10934) );
  NAND2_X1 U15053 ( .A1(n10938), .A2(n29428), .ZN(n10939) );
  NAND4_X2 U15054 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n32188) );
  XNOR2_X1 U15055 ( .A(n32188), .B(\fmem_data[3][3] ), .ZN(n28403) );
  XOR2_X1 U15056 ( .A(\fmem_data[3][2] ), .B(\fmem_data[3][3] ), .Z(n10943) );
  BUF_X1 U15057 ( .A(n14936), .Z(n29279) );
  AOI22_X1 U15058 ( .A1(n27755), .A2(\xmem_data[8][5] ), .B1(n29279), .B2(
        \xmem_data[9][5] ), .ZN(n10947) );
  BUF_X1 U15059 ( .A(n14935), .Z(n29271) );
  BUF_X1 U15060 ( .A(n14882), .Z(n29281) );
  AOI22_X1 U15061 ( .A1(n29271), .A2(\xmem_data[7][5] ), .B1(n29055), .B2(
        \xmem_data[15][5] ), .ZN(n10946) );
  NAND2_X1 U15062 ( .A1(n10947), .A2(n10946), .ZN(n10952) );
  AOI22_X1 U15063 ( .A1(n24509), .A2(\xmem_data[10][5] ), .B1(n31270), .B2(
        \xmem_data[11][5] ), .ZN(n10948) );
  INV_X1 U15064 ( .A(n10948), .ZN(n10951) );
  AOI22_X1 U15065 ( .A1(n28050), .A2(\xmem_data[2][5] ), .B1(n27863), .B2(
        \xmem_data[3][5] ), .ZN(n10949) );
  INV_X1 U15066 ( .A(n10949), .ZN(n10950) );
  NOR3_X1 U15067 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n10955) );
  AOI22_X1 U15068 ( .A1(n29591), .A2(\xmem_data[4][5] ), .B1(n21015), .B2(
        \xmem_data[5][5] ), .ZN(n10954) );
  BUF_X1 U15069 ( .A(n13481), .Z(n29280) );
  AOI22_X1 U15070 ( .A1(n27855), .A2(\xmem_data[12][5] ), .B1(n29280), .B2(
        \xmem_data[13][5] ), .ZN(n10953) );
  NAND3_X1 U15071 ( .A1(n10955), .A2(n10954), .A3(n10953), .ZN(n10971) );
  BUF_X1 U15072 ( .A(n13468), .Z(n29286) );
  AOI22_X1 U15073 ( .A1(n3334), .A2(\xmem_data[24][5] ), .B1(n29286), .B2(
        \xmem_data[25][5] ), .ZN(n10959) );
  AOI22_X1 U15074 ( .A1(n24443), .A2(\xmem_data[26][5] ), .B1(n3220), .B2(
        \xmem_data[27][5] ), .ZN(n10958) );
  BUF_X1 U15075 ( .A(n14988), .Z(n29288) );
  AOI22_X1 U15076 ( .A1(n29288), .A2(\xmem_data[28][5] ), .B1(n28508), .B2(
        \xmem_data[29][5] ), .ZN(n10957) );
  BUF_X1 U15077 ( .A(n14926), .Z(n29289) );
  AOI22_X1 U15078 ( .A1(n29289), .A2(\xmem_data[30][5] ), .B1(n13444), .B2(
        \xmem_data[31][5] ), .ZN(n10956) );
  NAND4_X1 U15079 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10970) );
  BUF_X1 U15080 ( .A(n14974), .Z(n29297) );
  AOI22_X1 U15081 ( .A1(n29297), .A2(\xmem_data[16][5] ), .B1(n28062), .B2(
        \xmem_data[17][5] ), .ZN(n10963) );
  AOI22_X1 U15082 ( .A1(n24467), .A2(\xmem_data[18][5] ), .B1(n28468), .B2(
        \xmem_data[19][5] ), .ZN(n10962) );
  AOI22_X1 U15083 ( .A1(n29298), .A2(\xmem_data[20][5] ), .B1(n27567), .B2(
        \xmem_data[21][5] ), .ZN(n10961) );
  AOI22_X1 U15084 ( .A1(n25630), .A2(\xmem_data[22][5] ), .B1(n21309), .B2(
        \xmem_data[23][5] ), .ZN(n10960) );
  NAND4_X1 U15085 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10969) );
  BUF_X1 U15086 ( .A(n13436), .Z(n29272) );
  NAND2_X1 U15087 ( .A1(n29272), .A2(\xmem_data[6][5] ), .ZN(n10965) );
  NAND2_X1 U15088 ( .A1(n24190), .A2(\xmem_data[14][5] ), .ZN(n10964) );
  NAND2_X1 U15089 ( .A1(n10965), .A2(n10964), .ZN(n10967) );
  AND2_X1 U15090 ( .A1(n30295), .A2(\xmem_data[0][5] ), .ZN(n10966) );
  OR2_X1 U15091 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  OR4_X1 U15092 ( .A1(n10971), .A2(n10970), .A3(n10969), .A4(n10968), .ZN(
        n10976) );
  AOI21_X1 U15093 ( .B1(n4499), .B2(n10972), .A(n10973), .ZN(n11043) );
  AOI22_X1 U15094 ( .A1(load_xaddr_val[6]), .A2(n10973), .B1(n11381), .B2(
        n39040), .ZN(n10998) );
  NOR2_X1 U15095 ( .A1(n11043), .A2(n10998), .ZN(n25790) );
  INV_X1 U15096 ( .A(n25790), .ZN(n29341) );
  NOR2_X1 U15097 ( .A1(n29341), .A2(n39030), .ZN(n10974) );
  AND2_X1 U15098 ( .A1(n29306), .A2(n10974), .ZN(n10975) );
  AND2_X1 U15099 ( .A1(n11043), .A2(n10998), .ZN(n29269) );
  BUF_X1 U15100 ( .A(n14991), .Z(n29231) );
  AOI22_X1 U15101 ( .A1(n29231), .A2(\xmem_data[96][5] ), .B1(n28307), .B2(
        \xmem_data[97][5] ), .ZN(n10981) );
  AOI22_X1 U15102 ( .A1(n25670), .A2(\xmem_data[98][5] ), .B1(n24130), .B2(
        \xmem_data[99][5] ), .ZN(n10980) );
  BUF_X1 U15103 ( .A(n13435), .Z(n29232) );
  AOI22_X1 U15104 ( .A1(n30508), .A2(\xmem_data[100][5] ), .B1(n29232), .B2(
        \xmem_data[101][5] ), .ZN(n10979) );
  AOI22_X1 U15105 ( .A1(n25425), .A2(\xmem_data[102][5] ), .B1(n27912), .B2(
        \xmem_data[103][5] ), .ZN(n10978) );
  NAND4_X1 U15106 ( .A1(n10981), .A2(n10980), .A3(n10979), .A4(n10978), .ZN(
        n10997) );
  BUF_X1 U15107 ( .A(n29187), .Z(n29237) );
  AOI22_X1 U15108 ( .A1(n27818), .A2(\xmem_data[104][5] ), .B1(n23716), .B2(
        \xmem_data[105][5] ), .ZN(n10985) );
  AOI22_X1 U15109 ( .A1(n25573), .A2(\xmem_data[106][5] ), .B1(n31355), .B2(
        \xmem_data[107][5] ), .ZN(n10984) );
  BUF_X1 U15110 ( .A(n14971), .Z(n29239) );
  AOI22_X1 U15111 ( .A1(n29239), .A2(\xmem_data[108][5] ), .B1(n29238), .B2(
        \xmem_data[109][5] ), .ZN(n10983) );
  BUF_X1 U15112 ( .A(n14881), .Z(n29240) );
  AOI22_X1 U15113 ( .A1(n29240), .A2(\xmem_data[110][5] ), .B1(n27461), .B2(
        \xmem_data[111][5] ), .ZN(n10982) );
  NAND4_X1 U15114 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10996) );
  BUF_X1 U15115 ( .A(n14974), .Z(n29246) );
  BUF_X1 U15116 ( .A(n14883), .Z(n29245) );
  AOI22_X1 U15117 ( .A1(n29246), .A2(\xmem_data[112][5] ), .B1(n29245), .B2(
        \xmem_data[113][5] ), .ZN(n10989) );
  BUF_X1 U15118 ( .A(n14919), .Z(n29247) );
  AOI22_X1 U15119 ( .A1(n24572), .A2(\xmem_data[114][5] ), .B1(n29247), .B2(
        \xmem_data[115][5] ), .ZN(n10988) );
  BUF_X1 U15120 ( .A(n13457), .Z(n29248) );
  AOI22_X1 U15121 ( .A1(n20826), .A2(\xmem_data[116][5] ), .B1(n29248), .B2(
        \xmem_data[117][5] ), .ZN(n10987) );
  AOI22_X1 U15122 ( .A1(n25724), .A2(\xmem_data[118][5] ), .B1(n24573), .B2(
        \xmem_data[119][5] ), .ZN(n10986) );
  NAND4_X1 U15123 ( .A1(n10989), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n10995) );
  BUF_X1 U15124 ( .A(n13468), .Z(n29253) );
  AOI22_X1 U15125 ( .A1(n3351), .A2(\xmem_data[120][5] ), .B1(n29253), .B2(
        \xmem_data[121][5] ), .ZN(n10993) );
  BUF_X1 U15126 ( .A(n29064), .Z(n29254) );
  AOI22_X1 U15127 ( .A1(n29254), .A2(\xmem_data[122][5] ), .B1(n3222), .B2(
        \xmem_data[123][5] ), .ZN(n10992) );
  BUF_X1 U15128 ( .A(n14988), .Z(n29256) );
  BUF_X1 U15129 ( .A(n14989), .Z(n29255) );
  AOI22_X1 U15130 ( .A1(n29256), .A2(\xmem_data[124][5] ), .B1(n29255), .B2(
        \xmem_data[125][5] ), .ZN(n10991) );
  BUF_X1 U15131 ( .A(n14926), .Z(n29257) );
  AOI22_X1 U15132 ( .A1(n29257), .A2(\xmem_data[126][5] ), .B1(n20559), .B2(
        \xmem_data[127][5] ), .ZN(n10990) );
  NAND4_X1 U15133 ( .A1(n10993), .A2(n10992), .A3(n10991), .A4(n10990), .ZN(
        n10994) );
  OR4_X1 U15134 ( .A1(n10997), .A2(n10996), .A3(n10995), .A4(n10994), .ZN(
        n11022) );
  INV_X1 U15135 ( .A(n10998), .ZN(n11044) );
  NOR2_X1 U15136 ( .A1(n11043), .A2(n11044), .ZN(n29267) );
  BUF_X1 U15137 ( .A(n14928), .Z(n29306) );
  AOI22_X1 U15138 ( .A1(n27396), .A2(\xmem_data[64][5] ), .B1(n3231), .B2(
        \xmem_data[65][5] ), .ZN(n11003) );
  BUF_X1 U15139 ( .A(n10999), .Z(n29307) );
  AOI22_X1 U15140 ( .A1(n27910), .A2(\xmem_data[66][5] ), .B1(n29307), .B2(
        \xmem_data[67][5] ), .ZN(n11002) );
  BUF_X1 U15141 ( .A(n14997), .Z(n29308) );
  AOI22_X1 U15142 ( .A1(n29308), .A2(\xmem_data[68][5] ), .B1(n22675), .B2(
        \xmem_data[69][5] ), .ZN(n11001) );
  BUF_X1 U15143 ( .A(n13476), .Z(n29310) );
  BUF_X1 U15144 ( .A(n14898), .Z(n29309) );
  AOI22_X1 U15145 ( .A1(n29310), .A2(\xmem_data[70][5] ), .B1(n29309), .B2(
        \xmem_data[71][5] ), .ZN(n11000) );
  NAND4_X1 U15146 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11020) );
  BUF_X1 U15147 ( .A(n29187), .Z(n29315) );
  AOI22_X1 U15148 ( .A1(n27517), .A2(\xmem_data[72][5] ), .B1(n3213), .B2(
        \xmem_data[73][5] ), .ZN(n11007) );
  BUF_X1 U15149 ( .A(n13149), .Z(n29317) );
  BUF_X1 U15150 ( .A(n14970), .Z(n29316) );
  AOI22_X1 U15151 ( .A1(n29317), .A2(\xmem_data[74][5] ), .B1(n29316), .B2(
        \xmem_data[75][5] ), .ZN(n11006) );
  BUF_X1 U15152 ( .A(n14971), .Z(n29319) );
  AOI22_X1 U15153 ( .A1(n29319), .A2(\xmem_data[76][5] ), .B1(n29318), .B2(
        \xmem_data[77][5] ), .ZN(n11005) );
  AOI22_X1 U15154 ( .A1(n28061), .A2(\xmem_data[78][5] ), .B1(n20506), .B2(
        \xmem_data[79][5] ), .ZN(n11004) );
  NAND4_X1 U15155 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n11019) );
  BUF_X1 U15156 ( .A(n14974), .Z(n29324) );
  AOI22_X1 U15157 ( .A1(n29324), .A2(\xmem_data[80][5] ), .B1(n14975), .B2(
        \xmem_data[81][5] ), .ZN(n11012) );
  AOI22_X1 U15158 ( .A1(n29325), .A2(\xmem_data[82][5] ), .B1(n27463), .B2(
        \xmem_data[83][5] ), .ZN(n11011) );
  BUF_X1 U15159 ( .A(n13420), .Z(n29327) );
  BUF_X1 U15160 ( .A(n13487), .Z(n29326) );
  AOI22_X1 U15161 ( .A1(n29327), .A2(\xmem_data[84][5] ), .B1(n29326), .B2(
        \xmem_data[85][5] ), .ZN(n11010) );
  BUF_X1 U15162 ( .A(n28947), .Z(n29328) );
  AOI22_X1 U15163 ( .A1(n25630), .A2(\xmem_data[86][5] ), .B1(n29328), .B2(
        \xmem_data[87][5] ), .ZN(n11009) );
  NAND4_X1 U15164 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11018) );
  AOI22_X1 U15165 ( .A1(n3383), .A2(\xmem_data[88][5] ), .B1(n27437), .B2(
        \xmem_data[89][5] ), .ZN(n11016) );
  AOI22_X1 U15166 ( .A1(n28470), .A2(\xmem_data[90][5] ), .B1(n3219), .B2(
        \xmem_data[91][5] ), .ZN(n11015) );
  AOI22_X1 U15167 ( .A1(n24533), .A2(\xmem_data[92][5] ), .B1(n25562), .B2(
        \xmem_data[93][5] ), .ZN(n11014) );
  AOI22_X1 U15168 ( .A1(n28083), .A2(\xmem_data[94][5] ), .B1(n25415), .B2(
        \xmem_data[95][5] ), .ZN(n11013) );
  NAND4_X1 U15169 ( .A1(n11016), .A2(n11015), .A3(n11014), .A4(n11013), .ZN(
        n11017) );
  OR4_X1 U15170 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  AOI22_X1 U15171 ( .A1(n29269), .A2(n11022), .B1(n29267), .B2(n11021), .ZN(
        n11047) );
  AOI22_X1 U15172 ( .A1(n3134), .A2(\xmem_data[32][5] ), .B1(n3231), .B2(
        \xmem_data[33][5] ), .ZN(n11026) );
  AOI22_X1 U15173 ( .A1(n25422), .A2(\xmem_data[34][5] ), .B1(n29307), .B2(
        \xmem_data[35][5] ), .ZN(n11025) );
  AOI22_X1 U15174 ( .A1(n29308), .A2(\xmem_data[36][5] ), .B1(n22702), .B2(
        \xmem_data[37][5] ), .ZN(n11024) );
  AOI22_X1 U15175 ( .A1(n29310), .A2(\xmem_data[38][5] ), .B1(n29309), .B2(
        \xmem_data[39][5] ), .ZN(n11023) );
  NAND4_X1 U15176 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n11042) );
  AOI22_X1 U15177 ( .A1(n25519), .A2(\xmem_data[40][5] ), .B1(n25460), .B2(
        \xmem_data[41][5] ), .ZN(n11030) );
  AOI22_X1 U15178 ( .A1(n29317), .A2(\xmem_data[42][5] ), .B1(n29316), .B2(
        \xmem_data[43][5] ), .ZN(n11029) );
  AOI22_X1 U15179 ( .A1(n29319), .A2(\xmem_data[44][5] ), .B1(n29318), .B2(
        \xmem_data[45][5] ), .ZN(n11028) );
  AOI22_X1 U15180 ( .A1(n22683), .A2(\xmem_data[46][5] ), .B1(n24222), .B2(
        \xmem_data[47][5] ), .ZN(n11027) );
  NAND4_X1 U15181 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11041) );
  AOI22_X1 U15182 ( .A1(n29324), .A2(\xmem_data[48][5] ), .B1(n14975), .B2(
        \xmem_data[49][5] ), .ZN(n11034) );
  AOI22_X1 U15183 ( .A1(n29325), .A2(\xmem_data[50][5] ), .B1(n28500), .B2(
        \xmem_data[51][5] ), .ZN(n11033) );
  AOI22_X1 U15184 ( .A1(n29327), .A2(\xmem_data[52][5] ), .B1(n29326), .B2(
        \xmem_data[53][5] ), .ZN(n11032) );
  AOI22_X1 U15185 ( .A1(n27436), .A2(\xmem_data[54][5] ), .B1(n29328), .B2(
        \xmem_data[55][5] ), .ZN(n11031) );
  NAND4_X1 U15186 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11040) );
  AOI22_X1 U15187 ( .A1(n3383), .A2(\xmem_data[56][5] ), .B1(n24439), .B2(
        \xmem_data[57][5] ), .ZN(n11038) );
  AOI22_X1 U15188 ( .A1(n28318), .A2(\xmem_data[58][5] ), .B1(n3221), .B2(
        \xmem_data[59][5] ), .ZN(n11037) );
  AOI22_X1 U15189 ( .A1(n24533), .A2(\xmem_data[60][5] ), .B1(n20787), .B2(
        \xmem_data[61][5] ), .ZN(n11036) );
  AOI22_X1 U15190 ( .A1(n22666), .A2(\xmem_data[62][5] ), .B1(n17061), .B2(
        \xmem_data[63][5] ), .ZN(n11035) );
  NAND4_X1 U15191 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n11039) );
  OR4_X1 U15192 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11045) );
  AND2_X1 U15193 ( .A1(n11044), .A2(n11043), .ZN(n29343) );
  NAND2_X1 U15194 ( .A1(n11045), .A2(n29343), .ZN(n11046) );
  XOR2_X1 U15195 ( .A(\fmem_data[8][4] ), .B(\fmem_data[8][5] ), .Z(n11049) );
  AOI22_X1 U15196 ( .A1(n25451), .A2(\xmem_data[64][6] ), .B1(n23771), .B2(
        \xmem_data[65][6] ), .ZN(n11053) );
  AOI22_X1 U15197 ( .A1(n24638), .A2(n20682), .B1(n29307), .B2(
        \xmem_data[67][6] ), .ZN(n11052) );
  AOI22_X1 U15198 ( .A1(n29308), .A2(\xmem_data[68][6] ), .B1(n29232), .B2(
        \xmem_data[69][6] ), .ZN(n11051) );
  AOI22_X1 U15199 ( .A1(n29310), .A2(\xmem_data[70][6] ), .B1(n29309), .B2(
        \xmem_data[71][6] ), .ZN(n11050) );
  NAND4_X1 U15200 ( .A1(n11053), .A2(n11052), .A3(n11051), .A4(n11050), .ZN(
        n11069) );
  AOI22_X1 U15201 ( .A1(n30892), .A2(\xmem_data[72][6] ), .B1(n3213), .B2(
        \xmem_data[73][6] ), .ZN(n11057) );
  AOI22_X1 U15202 ( .A1(n29317), .A2(\xmem_data[74][6] ), .B1(n29316), .B2(
        \xmem_data[75][6] ), .ZN(n11056) );
  AOI22_X1 U15203 ( .A1(n29319), .A2(\xmem_data[76][6] ), .B1(n29318), .B2(
        \xmem_data[77][6] ), .ZN(n11055) );
  AOI22_X1 U15204 ( .A1(n27524), .A2(\xmem_data[78][6] ), .B1(n27856), .B2(
        \xmem_data[79][6] ), .ZN(n11054) );
  NAND4_X1 U15205 ( .A1(n11057), .A2(n11056), .A3(n11055), .A4(n11054), .ZN(
        n11068) );
  AOI22_X1 U15206 ( .A1(n29324), .A2(\xmem_data[80][6] ), .B1(n14975), .B2(
        \xmem_data[81][6] ), .ZN(n11061) );
  AOI22_X1 U15207 ( .A1(n29325), .A2(\xmem_data[82][6] ), .B1(n28292), .B2(
        \xmem_data[83][6] ), .ZN(n11060) );
  AOI22_X1 U15208 ( .A1(n29327), .A2(\xmem_data[84][6] ), .B1(n29326), .B2(
        \xmem_data[85][6] ), .ZN(n11059) );
  AOI22_X1 U15209 ( .A1(n3380), .A2(\xmem_data[86][6] ), .B1(n29328), .B2(
        \xmem_data[87][6] ), .ZN(n11058) );
  NAND4_X1 U15210 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n11067) );
  AOI22_X1 U15211 ( .A1(n3383), .A2(\xmem_data[88][6] ), .B1(n29253), .B2(
        \xmem_data[89][6] ), .ZN(n11065) );
  AOI22_X1 U15212 ( .A1(n28470), .A2(\xmem_data[90][6] ), .B1(n3219), .B2(
        \xmem_data[91][6] ), .ZN(n11064) );
  AOI22_X1 U15213 ( .A1(n29065), .A2(\xmem_data[92][6] ), .B1(n28476), .B2(
        \xmem_data[93][6] ), .ZN(n11063) );
  AOI22_X1 U15214 ( .A1(n29257), .A2(\xmem_data[94][6] ), .B1(n14890), .B2(
        \xmem_data[95][6] ), .ZN(n11062) );
  NAND4_X1 U15215 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11066) );
  OR4_X1 U15216 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11070) );
  NAND2_X1 U15217 ( .A1(n11070), .A2(n29267), .ZN(n11143) );
  AOI22_X1 U15218 ( .A1(n23754), .A2(\xmem_data[120][6] ), .B1(n29253), .B2(
        \xmem_data[121][6] ), .ZN(n11074) );
  AOI22_X1 U15219 ( .A1(n29254), .A2(\xmem_data[122][6] ), .B1(n3222), .B2(
        \xmem_data[123][6] ), .ZN(n11073) );
  AOI22_X1 U15220 ( .A1(n29256), .A2(\xmem_data[124][6] ), .B1(n29255), .B2(
        \xmem_data[125][6] ), .ZN(n11072) );
  AOI22_X1 U15221 ( .A1(n29257), .A2(\xmem_data[126][6] ), .B1(n29104), .B2(
        \xmem_data[127][6] ), .ZN(n11071) );
  NAND4_X1 U15222 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11090) );
  AOI22_X1 U15223 ( .A1(n29246), .A2(\xmem_data[112][6] ), .B1(n29245), .B2(
        \xmem_data[113][6] ), .ZN(n11078) );
  AOI22_X1 U15224 ( .A1(n20552), .A2(\xmem_data[114][6] ), .B1(n29247), .B2(
        \xmem_data[115][6] ), .ZN(n11077) );
  AOI22_X1 U15225 ( .A1(n24687), .A2(\xmem_data[116][6] ), .B1(n29248), .B2(
        \xmem_data[117][6] ), .ZN(n11076) );
  AOI22_X1 U15226 ( .A1(n3380), .A2(\xmem_data[118][6] ), .B1(n25561), .B2(
        \xmem_data[119][6] ), .ZN(n11075) );
  NAND4_X1 U15227 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11089) );
  AOI22_X1 U15228 ( .A1(n25422), .A2(\xmem_data[98][6] ), .B1(n22739), .B2(
        \xmem_data[99][6] ), .ZN(n11081) );
  AOI22_X1 U15229 ( .A1(n23762), .A2(\xmem_data[100][6] ), .B1(n29232), .B2(
        \xmem_data[101][6] ), .ZN(n11080) );
  AOI22_X1 U15230 ( .A1(n17041), .A2(\xmem_data[102][6] ), .B1(n20798), .B2(
        \xmem_data[103][6] ), .ZN(n11079) );
  NAND4_X1 U15231 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11088) );
  AOI22_X1 U15232 ( .A1(n27945), .A2(\xmem_data[104][6] ), .B1(n31269), .B2(
        \xmem_data[105][6] ), .ZN(n11086) );
  AOI22_X1 U15233 ( .A1(n21007), .A2(\xmem_data[106][6] ), .B1(n31355), .B2(
        \xmem_data[107][6] ), .ZN(n11085) );
  AOI22_X1 U15234 ( .A1(n29239), .A2(\xmem_data[108][6] ), .B1(n29238), .B2(
        \xmem_data[109][6] ), .ZN(n11084) );
  AOI22_X1 U15235 ( .A1(n29240), .A2(\xmem_data[110][6] ), .B1(n30495), .B2(
        \xmem_data[111][6] ), .ZN(n11083) );
  NAND4_X1 U15236 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11087) );
  OR4_X1 U15237 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11091) );
  NAND2_X1 U15238 ( .A1(n11091), .A2(n29269), .ZN(n11142) );
  AOI22_X1 U15239 ( .A1(n29297), .A2(\xmem_data[16][6] ), .B1(n20507), .B2(
        \xmem_data[17][6] ), .ZN(n11097) );
  AOI22_X1 U15240 ( .A1(n24467), .A2(\xmem_data[18][6] ), .B1(n29247), .B2(
        \xmem_data[19][6] ), .ZN(n11096) );
  AND2_X1 U15241 ( .A1(n27957), .A2(\xmem_data[21][6] ), .ZN(n11092) );
  AOI21_X1 U15242 ( .B1(n29298), .B2(\xmem_data[20][6] ), .A(n11092), .ZN(
        n11095) );
  AND2_X1 U15243 ( .A1(n25441), .A2(\xmem_data[22][6] ), .ZN(n11093) );
  AOI21_X1 U15244 ( .B1(n3203), .B2(\xmem_data[23][6] ), .A(n11093), .ZN(
        n11094) );
  AOI22_X1 U15245 ( .A1(n3158), .A2(\xmem_data[8][6] ), .B1(n29279), .B2(
        \xmem_data[9][6] ), .ZN(n11101) );
  AOI22_X1 U15246 ( .A1(n30949), .A2(\xmem_data[10][6] ), .B1(n29048), .B2(
        \xmem_data[11][6] ), .ZN(n11100) );
  AOI22_X1 U15247 ( .A1(n30893), .A2(\xmem_data[12][6] ), .B1(n29280), .B2(
        \xmem_data[13][6] ), .ZN(n11099) );
  AOI22_X1 U15248 ( .A1(n29100), .A2(\xmem_data[14][6] ), .B1(n21009), .B2(
        \xmem_data[15][6] ), .ZN(n11098) );
  NAND4_X1 U15249 ( .A1(n11101), .A2(n11100), .A3(n11099), .A4(n11098), .ZN(
        n11102) );
  NOR2_X1 U15250 ( .A1(n11102), .A2(n3734), .ZN(n11114) );
  AOI22_X1 U15251 ( .A1(n3334), .A2(\xmem_data[24][6] ), .B1(n29286), .B2(
        \xmem_data[25][6] ), .ZN(n11106) );
  AOI22_X1 U15252 ( .A1(n30503), .A2(\xmem_data[26][6] ), .B1(n3220), .B2(
        \xmem_data[27][6] ), .ZN(n11105) );
  AOI22_X1 U15253 ( .A1(n29288), .A2(\xmem_data[28][6] ), .B1(n31367), .B2(
        \xmem_data[29][6] ), .ZN(n11104) );
  AOI22_X1 U15254 ( .A1(n29289), .A2(\xmem_data[30][6] ), .B1(n25415), .B2(
        \xmem_data[31][6] ), .ZN(n11103) );
  AND4_X1 U15255 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11113) );
  AOI22_X1 U15256 ( .A1(n29272), .A2(\xmem_data[6][6] ), .B1(n29271), .B2(
        \xmem_data[7][6] ), .ZN(n11109) );
  AOI22_X1 U15257 ( .A1(n25422), .A2(\xmem_data[2][6] ), .B1(n3358), .B2(
        \xmem_data[3][6] ), .ZN(n11108) );
  NAND2_X1 U15258 ( .A1(n27396), .A2(\xmem_data[0][6] ), .ZN(n11107) );
  NAND3_X1 U15259 ( .A1(n11109), .A2(n11108), .A3(n11107), .ZN(n11112) );
  AOI22_X1 U15260 ( .A1(n31353), .A2(\xmem_data[4][6] ), .B1(n24212), .B2(
        \xmem_data[5][6] ), .ZN(n11110) );
  INV_X1 U15261 ( .A(n11110), .ZN(n11111) );
  NAND4_X1 U15262 ( .A1(n3543), .A2(n11114), .A3(n11113), .A4(n3939), .ZN(
        n11140) );
  AOI22_X1 U15263 ( .A1(n30592), .A2(\xmem_data[58][6] ), .B1(n3222), .B2(
        \xmem_data[59][6] ), .ZN(n11115) );
  INV_X1 U15264 ( .A(n11115), .ZN(n11123) );
  AOI22_X1 U15265 ( .A1(n29325), .A2(\xmem_data[50][6] ), .B1(n22751), .B2(
        \xmem_data[51][6] ), .ZN(n11117) );
  AOI22_X1 U15266 ( .A1(n28367), .A2(\xmem_data[60][6] ), .B1(n20723), .B2(
        \xmem_data[61][6] ), .ZN(n11116) );
  NAND2_X1 U15267 ( .A1(n11117), .A2(n11116), .ZN(n11122) );
  AOI22_X1 U15268 ( .A1(n24534), .A2(\xmem_data[62][6] ), .B1(n28372), .B2(
        \xmem_data[63][6] ), .ZN(n11120) );
  AOI22_X1 U15269 ( .A1(n29324), .A2(\xmem_data[48][6] ), .B1(n14975), .B2(
        \xmem_data[49][6] ), .ZN(n11119) );
  AOI22_X1 U15270 ( .A1(n3384), .A2(\xmem_data[56][6] ), .B1(n27437), .B2(
        \xmem_data[57][6] ), .ZN(n11118) );
  NOR3_X1 U15271 ( .A1(n11123), .A2(n11122), .A3(n11121), .ZN(n11138) );
  AOI22_X1 U15272 ( .A1(n20962), .A2(\xmem_data[32][6] ), .B1(n25450), .B2(
        \xmem_data[33][6] ), .ZN(n11127) );
  AOI22_X1 U15273 ( .A1(n25422), .A2(\xmem_data[34][6] ), .B1(n29307), .B2(
        \xmem_data[35][6] ), .ZN(n11126) );
  AOI22_X1 U15274 ( .A1(n29308), .A2(\xmem_data[36][6] ), .B1(n23761), .B2(
        \xmem_data[37][6] ), .ZN(n11125) );
  AOI22_X1 U15275 ( .A1(n29310), .A2(\xmem_data[38][6] ), .B1(n29309), .B2(
        \xmem_data[39][6] ), .ZN(n11124) );
  NAND4_X1 U15276 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11131) );
  AND2_X1 U15277 ( .A1(n27959), .A2(\xmem_data[54][6] ), .ZN(n11128) );
  AOI21_X1 U15278 ( .B1(n29328), .B2(\xmem_data[55][6] ), .A(n11128), .ZN(
        n11129) );
  INV_X1 U15279 ( .A(n11129), .ZN(n11130) );
  NOR2_X1 U15280 ( .A1(n11131), .A2(n11130), .ZN(n11137) );
  AOI22_X1 U15281 ( .A1(n28752), .A2(\xmem_data[40][6] ), .B1(n3213), .B2(
        \xmem_data[41][6] ), .ZN(n11135) );
  AOI22_X1 U15282 ( .A1(n29317), .A2(\xmem_data[42][6] ), .B1(n29316), .B2(
        \xmem_data[43][6] ), .ZN(n11134) );
  AOI22_X1 U15283 ( .A1(n29319), .A2(\xmem_data[44][6] ), .B1(n29318), .B2(
        \xmem_data[45][6] ), .ZN(n11133) );
  AOI22_X1 U15284 ( .A1(n30557), .A2(\xmem_data[46][6] ), .B1(n30955), .B2(
        \xmem_data[47][6] ), .ZN(n11132) );
  AOI22_X1 U15285 ( .A1(n29327), .A2(\xmem_data[52][6] ), .B1(n29326), .B2(
        \xmem_data[53][6] ), .ZN(n11136) );
  NAND4_X1 U15286 ( .A1(n11138), .A2(n11137), .A3(n3752), .A4(n11136), .ZN(
        n11139) );
  AOI22_X1 U15287 ( .A1(n11140), .A2(n25790), .B1(n11139), .B2(n29343), .ZN(
        n11141) );
  AOI22_X1 U15288 ( .A1(n27852), .A2(\xmem_data[96][3] ), .B1(n27435), .B2(
        \xmem_data[97][3] ), .ZN(n11147) );
  AOI22_X1 U15289 ( .A1(n27436), .A2(\xmem_data[98][3] ), .B1(n27499), .B2(
        \xmem_data[99][3] ), .ZN(n11146) );
  AOI22_X1 U15290 ( .A1(n21308), .A2(\xmem_data[100][3] ), .B1(n27437), .B2(
        \xmem_data[101][3] ), .ZN(n11145) );
  AOI22_X1 U15291 ( .A1(n27439), .A2(\xmem_data[102][3] ), .B1(n3221), .B2(
        \xmem_data[103][3] ), .ZN(n11144) );
  NAND4_X1 U15292 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11163) );
  AOI22_X1 U15293 ( .A1(n27445), .A2(\xmem_data[104][3] ), .B1(n27444), .B2(
        \xmem_data[105][3] ), .ZN(n11151) );
  AOI22_X1 U15294 ( .A1(n23741), .A2(\xmem_data[106][3] ), .B1(n30882), .B2(
        \xmem_data[107][3] ), .ZN(n11150) );
  AOI22_X1 U15295 ( .A1(n3129), .A2(\xmem_data[108][3] ), .B1(n27446), .B2(
        \xmem_data[109][3] ), .ZN(n11149) );
  AOI22_X1 U15296 ( .A1(n27447), .A2(\xmem_data[110][3] ), .B1(n20982), .B2(
        \xmem_data[111][3] ), .ZN(n11148) );
  NAND4_X1 U15297 ( .A1(n11151), .A2(n11150), .A3(n11149), .A4(n11148), .ZN(
        n11162) );
  AOI22_X1 U15298 ( .A1(n27453), .A2(\xmem_data[112][3] ), .B1(n27452), .B2(
        \xmem_data[113][3] ), .ZN(n11155) );
  AOI22_X1 U15299 ( .A1(n31268), .A2(\xmem_data[114][3] ), .B1(n20717), .B2(
        \xmem_data[115][3] ), .ZN(n11154) );
  AOI22_X1 U15300 ( .A1(n17018), .A2(\xmem_data[116][3] ), .B1(n27454), .B2(
        \xmem_data[117][3] ), .ZN(n11153) );
  AOI22_X1 U15301 ( .A1(n29010), .A2(\xmem_data[118][3] ), .B1(n21006), .B2(
        \xmem_data[119][3] ), .ZN(n11152) );
  NAND4_X1 U15302 ( .A1(n11155), .A2(n11154), .A3(n11153), .A4(n11152), .ZN(
        n11161) );
  AOI22_X1 U15303 ( .A1(n23722), .A2(\xmem_data[120][3] ), .B1(n27460), .B2(
        \xmem_data[121][3] ), .ZN(n11159) );
  AOI22_X1 U15304 ( .A1(n27462), .A2(\xmem_data[122][3] ), .B1(n27461), .B2(
        \xmem_data[123][3] ), .ZN(n11158) );
  AOI22_X1 U15305 ( .A1(n30269), .A2(\xmem_data[124][3] ), .B1(n28062), .B2(
        \xmem_data[125][3] ), .ZN(n11157) );
  AOI22_X1 U15306 ( .A1(n3172), .A2(\xmem_data[126][3] ), .B1(n27463), .B2(
        \xmem_data[127][3] ), .ZN(n11156) );
  NAND4_X1 U15307 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11160) );
  OR4_X1 U15308 ( .A1(n11163), .A2(n11162), .A3(n11161), .A4(n11160), .ZN(
        n11186) );
  AOI22_X1 U15309 ( .A1(n30754), .A2(\xmem_data[64][3] ), .B1(n27435), .B2(
        \xmem_data[65][3] ), .ZN(n11168) );
  AOI22_X1 U15310 ( .A1(n27436), .A2(\xmem_data[66][3] ), .B1(n20489), .B2(
        \xmem_data[67][3] ), .ZN(n11167) );
  AOI22_X1 U15311 ( .A1(n3350), .A2(\xmem_data[68][3] ), .B1(n27437), .B2(
        \xmem_data[69][3] ), .ZN(n11166) );
  AND2_X1 U15312 ( .A1(n3222), .A2(\xmem_data[71][3] ), .ZN(n11164) );
  AOI21_X1 U15313 ( .B1(n27439), .B2(\xmem_data[70][3] ), .A(n11164), .ZN(
        n11165) );
  NAND4_X1 U15314 ( .A1(n11168), .A2(n11167), .A3(n11166), .A4(n11165), .ZN(
        n11184) );
  AOI22_X1 U15315 ( .A1(n27445), .A2(\xmem_data[72][3] ), .B1(n27444), .B2(
        \xmem_data[73][3] ), .ZN(n11172) );
  AOI22_X1 U15316 ( .A1(n21069), .A2(\xmem_data[74][3] ), .B1(n25415), .B2(
        \xmem_data[75][3] ), .ZN(n11171) );
  AOI22_X1 U15317 ( .A1(n28084), .A2(\xmem_data[76][3] ), .B1(n27446), .B2(
        \xmem_data[77][3] ), .ZN(n11170) );
  AOI22_X1 U15318 ( .A1(n27447), .A2(\xmem_data[78][3] ), .B1(n28415), .B2(
        \xmem_data[79][3] ), .ZN(n11169) );
  NAND4_X1 U15319 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11183) );
  AOI22_X1 U15320 ( .A1(n27453), .A2(\xmem_data[80][3] ), .B1(n27452), .B2(
        \xmem_data[81][3] ), .ZN(n11176) );
  AOI22_X1 U15321 ( .A1(n31268), .A2(\xmem_data[82][3] ), .B1(n24597), .B2(
        \xmem_data[83][3] ), .ZN(n11175) );
  AOI22_X1 U15322 ( .A1(n27755), .A2(\xmem_data[84][3] ), .B1(n27454), .B2(
        \xmem_data[85][3] ), .ZN(n11174) );
  AOI22_X1 U15323 ( .A1(n22676), .A2(\xmem_data[86][3] ), .B1(n28427), .B2(
        \xmem_data[87][3] ), .ZN(n11173) );
  NAND4_X1 U15324 ( .A1(n11176), .A2(n11175), .A3(n11174), .A4(n11173), .ZN(
        n11182) );
  AOI22_X1 U15325 ( .A1(n17044), .A2(\xmem_data[88][3] ), .B1(n27460), .B2(
        \xmem_data[89][3] ), .ZN(n11180) );
  AOI22_X1 U15326 ( .A1(n27462), .A2(\xmem_data[90][3] ), .B1(n27461), .B2(
        \xmem_data[91][3] ), .ZN(n11179) );
  AOI22_X1 U15327 ( .A1(n25636), .A2(\xmem_data[92][3] ), .B1(n28062), .B2(
        \xmem_data[93][3] ), .ZN(n11178) );
  AOI22_X1 U15328 ( .A1(n20818), .A2(\xmem_data[94][3] ), .B1(n27463), .B2(
        \xmem_data[95][3] ), .ZN(n11177) );
  NAND4_X1 U15329 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11181) );
  OR4_X1 U15330 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n11185) );
  AOI22_X1 U15331 ( .A1(n27496), .A2(n11186), .B1(n27494), .B2(n11185), .ZN(
        n11237) );
  AOI22_X1 U15332 ( .A1(n27502), .A2(\xmem_data[6][3] ), .B1(n3220), .B2(
        \xmem_data[7][3] ), .ZN(n11197) );
  AOI22_X1 U15333 ( .A1(n24710), .A2(\xmem_data[24][3] ), .B1(n13452), .B2(
        \xmem_data[25][3] ), .ZN(n11190) );
  AOI22_X1 U15334 ( .A1(n27524), .A2(\xmem_data[26][3] ), .B1(n25716), .B2(
        \xmem_data[27][3] ), .ZN(n11189) );
  AOI22_X1 U15335 ( .A1(n29297), .A2(\xmem_data[28][3] ), .B1(n29245), .B2(
        \xmem_data[29][3] ), .ZN(n11188) );
  AOI22_X1 U15336 ( .A1(n27542), .A2(\xmem_data[30][3] ), .B1(n29086), .B2(
        \xmem_data[31][3] ), .ZN(n11187) );
  NAND4_X1 U15337 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11193) );
  AOI22_X1 U15338 ( .A1(n3413), .A2(\xmem_data[4][3] ), .B1(n25360), .B2(
        \xmem_data[5][3] ), .ZN(n11191) );
  AOI22_X1 U15339 ( .A1(n27564), .A2(\xmem_data[2][3] ), .B1(n27563), .B2(
        \xmem_data[3][3] ), .ZN(n11195) );
  AOI22_X1 U15340 ( .A1(n27568), .A2(\xmem_data[0][3] ), .B1(n27567), .B2(
        \xmem_data[1][3] ), .ZN(n11194) );
  NAND4_X1 U15341 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(
        n11212) );
  AOI22_X1 U15342 ( .A1(n25612), .A2(\xmem_data[8][3] ), .B1(n29095), .B2(
        \xmem_data[9][3] ), .ZN(n11198) );
  AOI22_X1 U15343 ( .A1(n27551), .A2(\xmem_data[14][3] ), .B1(n3358), .B2(
        \xmem_data[15][3] ), .ZN(n11200) );
  NAND2_X1 U15344 ( .A1(n25451), .A2(\xmem_data[12][3] ), .ZN(n11199) );
  NAND2_X1 U15345 ( .A1(n11200), .A2(n11199), .ZN(n11203) );
  AOI22_X1 U15346 ( .A1(n25617), .A2(\xmem_data[10][3] ), .B1(n27550), .B2(
        \xmem_data[11][3] ), .ZN(n11201) );
  INV_X1 U15347 ( .A(n11201), .ZN(n11202) );
  OR3_X1 U15348 ( .A1(n11204), .A2(n11203), .A3(n11202), .ZN(n11210) );
  AOI22_X1 U15349 ( .A1(n28309), .A2(\xmem_data[16][3] ), .B1(n27535), .B2(
        \xmem_data[17][3] ), .ZN(n11208) );
  AOI22_X1 U15350 ( .A1(n25710), .A2(\xmem_data[18][3] ), .B1(n27536), .B2(
        \xmem_data[19][3] ), .ZN(n11207) );
  AOI22_X1 U15351 ( .A1(n28053), .A2(\xmem_data[20][3] ), .B1(n25383), .B2(
        \xmem_data[21][3] ), .ZN(n11206) );
  AOI22_X1 U15352 ( .A1(n25434), .A2(\xmem_data[22][3] ), .B1(n28427), .B2(
        \xmem_data[23][3] ), .ZN(n11205) );
  NAND4_X1 U15353 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11209) );
  OR2_X1 U15354 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  NOR2_X1 U15355 ( .A1(n11212), .A2(n11211), .ZN(n11213) );
  AOI22_X1 U15356 ( .A1(n27498), .A2(\xmem_data[32][3] ), .B1(n28035), .B2(
        \xmem_data[33][3] ), .ZN(n11217) );
  AOI22_X1 U15357 ( .A1(n27500), .A2(\xmem_data[34][3] ), .B1(n27499), .B2(
        \xmem_data[35][3] ), .ZN(n11216) );
  AOI22_X1 U15358 ( .A1(n25725), .A2(\xmem_data[36][3] ), .B1(n27501), .B2(
        \xmem_data[37][3] ), .ZN(n11215) );
  AOI22_X1 U15359 ( .A1(n27502), .A2(\xmem_data[38][3] ), .B1(n3221), .B2(
        \xmem_data[39][3] ), .ZN(n11214) );
  NAND4_X1 U15360 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11233) );
  AOI22_X1 U15361 ( .A1(n22708), .A2(\xmem_data[40][3] ), .B1(n27507), .B2(
        \xmem_data[41][3] ), .ZN(n11221) );
  AOI22_X1 U15362 ( .A1(n20725), .A2(\xmem_data[42][3] ), .B1(n13444), .B2(
        \xmem_data[43][3] ), .ZN(n11220) );
  AOI22_X1 U15363 ( .A1(n3128), .A2(\xmem_data[44][3] ), .B1(n31252), .B2(
        \xmem_data[45][3] ), .ZN(n11219) );
  AOI22_X1 U15364 ( .A1(n27508), .A2(\xmem_data[46][3] ), .B1(n24590), .B2(
        \xmem_data[47][3] ), .ZN(n11218) );
  NAND4_X1 U15365 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11232) );
  AOI22_X1 U15366 ( .A1(n27514), .A2(\xmem_data[48][3] ), .B1(n27513), .B2(
        \xmem_data[49][3] ), .ZN(n11225) );
  AOI22_X1 U15367 ( .A1(n27515), .A2(\xmem_data[50][3] ), .B1(n14999), .B2(
        \xmem_data[51][3] ), .ZN(n11224) );
  AOI22_X1 U15368 ( .A1(n30303), .A2(\xmem_data[52][3] ), .B1(n27516), .B2(
        \xmem_data[53][3] ), .ZN(n11223) );
  AOI22_X1 U15369 ( .A1(n24214), .A2(\xmem_data[54][3] ), .B1(n27518), .B2(
        \xmem_data[55][3] ), .ZN(n11222) );
  NAND4_X1 U15370 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11231) );
  AOI22_X1 U15371 ( .A1(n28687), .A2(\xmem_data[56][3] ), .B1(n27523), .B2(
        \xmem_data[57][3] ), .ZN(n11229) );
  AOI22_X1 U15372 ( .A1(n27524), .A2(\xmem_data[58][3] ), .B1(n30955), .B2(
        \xmem_data[59][3] ), .ZN(n11228) );
  AOI22_X1 U15373 ( .A1(n24522), .A2(\xmem_data[60][3] ), .B1(n27525), .B2(
        \xmem_data[61][3] ), .ZN(n11227) );
  AOI22_X1 U15374 ( .A1(n27847), .A2(\xmem_data[62][3] ), .B1(n27526), .B2(
        \xmem_data[63][3] ), .ZN(n11226) );
  NAND4_X1 U15375 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11230) );
  OR4_X1 U15376 ( .A1(n11233), .A2(n11232), .A3(n11231), .A4(n11230), .ZN(
        n11235) );
  NOR2_X1 U15377 ( .A1(n27573), .A2(n39018), .ZN(n11234) );
  AOI21_X1 U15378 ( .B1(n11235), .B2(n27577), .A(n3897), .ZN(n11236) );
  XNOR2_X1 U15379 ( .A(n31899), .B(\fmem_data[20][7] ), .ZN(n30459) );
  XOR2_X1 U15380 ( .A(\fmem_data[20][6] ), .B(\fmem_data[20][7] ), .Z(n11238)
         );
  XNOR2_X1 U15381 ( .A(n31900), .B(\fmem_data[20][7] ), .ZN(n31643) );
  XOR2_X1 U15382 ( .A(\fmem_data[0][2] ), .B(\fmem_data[0][3] ), .Z(n11239) );
  AOI22_X1 U15383 ( .A1(n20939), .A2(\xmem_data[32][7] ), .B1(n20938), .B2(
        \xmem_data[33][7] ), .ZN(n11243) );
  AOI22_X1 U15384 ( .A1(n20542), .A2(\xmem_data[34][7] ), .B1(n20940), .B2(
        \xmem_data[35][7] ), .ZN(n11242) );
  AOI22_X1 U15385 ( .A1(n20942), .A2(\xmem_data[36][7] ), .B1(n20941), .B2(
        \xmem_data[37][7] ), .ZN(n11241) );
  AOI22_X1 U15386 ( .A1(n28385), .A2(\xmem_data[38][7] ), .B1(n20943), .B2(
        \xmem_data[39][7] ), .ZN(n11240) );
  NAND4_X1 U15387 ( .A1(n11243), .A2(n11242), .A3(n11241), .A4(n11240), .ZN(
        n11249) );
  AOI22_X1 U15388 ( .A1(n20962), .A2(\xmem_data[56][7] ), .B1(n29306), .B2(
        \xmem_data[57][7] ), .ZN(n11247) );
  AOI22_X1 U15389 ( .A1(n20961), .A2(\xmem_data[58][7] ), .B1(n3357), .B2(
        \xmem_data[59][7] ), .ZN(n11246) );
  AOI22_X1 U15390 ( .A1(n17064), .A2(\xmem_data[60][7] ), .B1(n20958), .B2(
        \xmem_data[61][7] ), .ZN(n11245) );
  AOI22_X1 U15391 ( .A1(n20959), .A2(\xmem_data[62][7] ), .B1(n25671), .B2(
        \xmem_data[63][7] ), .ZN(n11244) );
  NAND4_X1 U15392 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11248) );
  NOR2_X1 U15393 ( .A1(n11249), .A2(n11248), .ZN(n11263) );
  NAND2_X1 U15394 ( .A1(n20952), .A2(\xmem_data[44][7] ), .ZN(n11251) );
  NAND2_X1 U15395 ( .A1(n20951), .A2(\xmem_data[45][7] ), .ZN(n11250) );
  NAND2_X1 U15396 ( .A1(n11251), .A2(n11250), .ZN(n11259) );
  AOI22_X1 U15397 ( .A1(n24606), .A2(\xmem_data[42][7] ), .B1(n29017), .B2(
        \xmem_data[43][7] ), .ZN(n11254) );
  AOI22_X1 U15398 ( .A1(n30864), .A2(\xmem_data[48][7] ), .B1(n24172), .B2(
        \xmem_data[49][7] ), .ZN(n11253) );
  AOI22_X1 U15399 ( .A1(n20950), .A2(\xmem_data[40][7] ), .B1(n20949), .B2(
        \xmem_data[41][7] ), .ZN(n11252) );
  AOI22_X1 U15400 ( .A1(n20969), .A2(\xmem_data[54][7] ), .B1(n28342), .B2(
        \xmem_data[55][7] ), .ZN(n11256) );
  AOI22_X1 U15401 ( .A1(n25731), .A2(\xmem_data[52][7] ), .B1(n30963), .B2(
        \xmem_data[53][7] ), .ZN(n11255) );
  NAND2_X1 U15402 ( .A1(n11256), .A2(n11255), .ZN(n11257) );
  NOR3_X1 U15403 ( .A1(n11259), .A2(n11258), .A3(n11257), .ZN(n11262) );
  AOI22_X1 U15404 ( .A1(n28082), .A2(\xmem_data[50][7] ), .B1(n3220), .B2(
        \xmem_data[51][7] ), .ZN(n11261) );
  AOI22_X1 U15405 ( .A1(n20953), .A2(\xmem_data[46][7] ), .B1(n27563), .B2(
        \xmem_data[47][7] ), .ZN(n11260) );
  NAND4_X1 U15406 ( .A1(n11263), .A2(n11262), .A3(n11261), .A4(n11260), .ZN(
        n11289) );
  AOI22_X1 U15407 ( .A1(n21005), .A2(\xmem_data[0][7] ), .B1(n29162), .B2(
        \xmem_data[1][7] ), .ZN(n11267) );
  AOI22_X1 U15408 ( .A1(n21007), .A2(\xmem_data[2][7] ), .B1(n21006), .B2(
        \xmem_data[3][7] ), .ZN(n11266) );
  AOI22_X1 U15409 ( .A1(n21008), .A2(\xmem_data[4][7] ), .B1(n29318), .B2(
        \xmem_data[5][7] ), .ZN(n11265) );
  AOI22_X1 U15410 ( .A1(n21010), .A2(\xmem_data[6][7] ), .B1(n25581), .B2(
        \xmem_data[7][7] ), .ZN(n11264) );
  NAND4_X1 U15411 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(
        n11268) );
  OR2_X1 U15412 ( .A1(n11268), .A2(n3969), .ZN(n11287) );
  AOI22_X1 U15413 ( .A1(n3433), .A2(\xmem_data[16][7] ), .B1(n25687), .B2(
        \xmem_data[17][7] ), .ZN(n11272) );
  AOI22_X1 U15414 ( .A1(n20991), .A2(\xmem_data[18][7] ), .B1(n3220), .B2(
        \xmem_data[19][7] ), .ZN(n11271) );
  AOI22_X1 U15415 ( .A1(n29789), .A2(\xmem_data[20][7] ), .B1(n20992), .B2(
        \xmem_data[21][7] ), .ZN(n11270) );
  AOI22_X1 U15416 ( .A1(n20994), .A2(\xmem_data[22][7] ), .B1(n20993), .B2(
        \xmem_data[23][7] ), .ZN(n11269) );
  NAND4_X1 U15417 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11286) );
  AOI22_X1 U15418 ( .A1(n28152), .A2(\xmem_data[28][7] ), .B1(n21015), .B2(
        \xmem_data[29][7] ), .ZN(n11279) );
  AOI22_X1 U15419 ( .A1(n25567), .A2(\xmem_data[30][7] ), .B1(n29271), .B2(
        \xmem_data[31][7] ), .ZN(n11273) );
  INV_X1 U15420 ( .A(n11273), .ZN(n11277) );
  AOI22_X1 U15421 ( .A1(n23813), .A2(\xmem_data[26][7] ), .B1(n20982), .B2(
        \xmem_data[27][7] ), .ZN(n11275) );
  NAND2_X1 U15422 ( .A1(n25377), .A2(\xmem_data[24][7] ), .ZN(n11274) );
  NAND2_X1 U15423 ( .A1(n11275), .A2(n11274), .ZN(n11276) );
  NOR2_X1 U15424 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  NAND2_X1 U15425 ( .A1(n11279), .A2(n11278), .ZN(n11285) );
  AOI22_X1 U15426 ( .A1(n20984), .A2(\xmem_data[8][7] ), .B1(n20983), .B2(
        \xmem_data[9][7] ), .ZN(n11283) );
  AOI22_X1 U15427 ( .A1(n24685), .A2(\xmem_data[10][7] ), .B1(n22751), .B2(
        \xmem_data[11][7] ), .ZN(n11282) );
  AOI22_X1 U15428 ( .A1(n20985), .A2(\xmem_data[12][7] ), .B1(n10456), .B2(
        \xmem_data[13][7] ), .ZN(n11281) );
  AOI22_X1 U15429 ( .A1(n20986), .A2(\xmem_data[14][7] ), .B1(n24470), .B2(
        \xmem_data[15][7] ), .ZN(n11280) );
  NAND4_X1 U15430 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n11284) );
  OR4_X1 U15431 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11288) );
  AOI22_X1 U15432 ( .A1(n20311), .A2(n11289), .B1(n11288), .B2(n20980), .ZN(
        n11333) );
  AOI22_X1 U15433 ( .A1(n21048), .A2(\xmem_data[96][7] ), .B1(n3208), .B2(
        \xmem_data[97][7] ), .ZN(n11293) );
  AOI22_X1 U15434 ( .A1(n23764), .A2(\xmem_data[98][7] ), .B1(n28427), .B2(
        \xmem_data[99][7] ), .ZN(n11292) );
  AOI22_X1 U15435 ( .A1(n21050), .A2(\xmem_data[100][7] ), .B1(n21049), .B2(
        \xmem_data[101][7] ), .ZN(n11291) );
  AOI22_X1 U15436 ( .A1(n28460), .A2(\xmem_data[102][7] ), .B1(n25679), .B2(
        \xmem_data[103][7] ), .ZN(n11290) );
  NAND4_X1 U15437 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n11309) );
  AOI22_X1 U15438 ( .A1(n21056), .A2(\xmem_data[104][7] ), .B1(n27975), .B2(
        \xmem_data[105][7] ), .ZN(n11297) );
  AOI22_X1 U15439 ( .A1(n21058), .A2(\xmem_data[106][7] ), .B1(n21057), .B2(
        \xmem_data[107][7] ), .ZN(n11296) );
  AOI22_X1 U15440 ( .A1(n21060), .A2(\xmem_data[108][7] ), .B1(n21059), .B2(
        \xmem_data[109][7] ), .ZN(n11295) );
  AOI22_X1 U15441 ( .A1(n21061), .A2(\xmem_data[110][7] ), .B1(n31346), .B2(
        \xmem_data[111][7] ), .ZN(n11294) );
  NAND4_X1 U15442 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11308) );
  AOI22_X1 U15443 ( .A1(n25624), .A2(\xmem_data[112][7] ), .B1(n25485), .B2(
        \xmem_data[113][7] ), .ZN(n11301) );
  AOI22_X1 U15444 ( .A1(n21066), .A2(\xmem_data[114][7] ), .B1(n3219), .B2(
        \xmem_data[115][7] ), .ZN(n11300) );
  AOI22_X1 U15445 ( .A1(n21067), .A2(\xmem_data[116][7] ), .B1(n20723), .B2(
        \xmem_data[117][7] ), .ZN(n11299) );
  AOI22_X1 U15446 ( .A1(n21069), .A2(\xmem_data[118][7] ), .B1(n21068), .B2(
        \xmem_data[119][7] ), .ZN(n11298) );
  NAND4_X1 U15447 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11307) );
  AOI22_X1 U15448 ( .A1(n21074), .A2(\xmem_data[120][7] ), .B1(n27547), .B2(
        \xmem_data[121][7] ), .ZN(n11305) );
  AOI22_X1 U15449 ( .A1(n27551), .A2(\xmem_data[122][7] ), .B1(n27943), .B2(
        \xmem_data[123][7] ), .ZN(n11304) );
  AOI22_X1 U15450 ( .A1(n29403), .A2(\xmem_data[124][7] ), .B1(n21075), .B2(
        \xmem_data[125][7] ), .ZN(n11303) );
  AOI22_X1 U15451 ( .A1(n30891), .A2(\xmem_data[126][7] ), .B1(n21076), .B2(
        \xmem_data[127][7] ), .ZN(n11302) );
  NAND4_X1 U15452 ( .A1(n11305), .A2(n11304), .A3(n11303), .A4(n11302), .ZN(
        n11306) );
  OR4_X1 U15453 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11331) );
  AOI22_X1 U15454 ( .A1(n20939), .A2(\xmem_data[64][7] ), .B1(n20938), .B2(
        \xmem_data[65][7] ), .ZN(n11313) );
  AOI22_X1 U15455 ( .A1(n20585), .A2(\xmem_data[66][7] ), .B1(n20940), .B2(
        \xmem_data[67][7] ), .ZN(n11312) );
  AOI22_X1 U15456 ( .A1(n20942), .A2(\xmem_data[68][7] ), .B1(n20941), .B2(
        \xmem_data[69][7] ), .ZN(n11311) );
  AOI22_X1 U15457 ( .A1(n24647), .A2(\xmem_data[70][7] ), .B1(n20943), .B2(
        \xmem_data[71][7] ), .ZN(n11310) );
  NAND4_X1 U15458 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11329) );
  AOI22_X1 U15459 ( .A1(n20950), .A2(\xmem_data[72][7] ), .B1(n20949), .B2(
        \xmem_data[73][7] ), .ZN(n11317) );
  AOI22_X1 U15460 ( .A1(n27542), .A2(\xmem_data[74][7] ), .B1(n23781), .B2(
        \xmem_data[75][7] ), .ZN(n11316) );
  AOI22_X1 U15461 ( .A1(n20952), .A2(\xmem_data[76][7] ), .B1(n20951), .B2(
        \xmem_data[77][7] ), .ZN(n11315) );
  AOI22_X1 U15462 ( .A1(n20953), .A2(\xmem_data[78][7] ), .B1(n21309), .B2(
        \xmem_data[79][7] ), .ZN(n11314) );
  NAND4_X1 U15463 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11328) );
  AOI22_X1 U15464 ( .A1(n25443), .A2(\xmem_data[80][7] ), .B1(n30863), .B2(
        \xmem_data[81][7] ), .ZN(n11321) );
  AOI22_X1 U15465 ( .A1(n20518), .A2(\xmem_data[82][7] ), .B1(n3221), .B2(
        \xmem_data[83][7] ), .ZN(n11320) );
  AOI22_X1 U15466 ( .A1(n25448), .A2(\xmem_data[84][7] ), .B1(n23739), .B2(
        \xmem_data[85][7] ), .ZN(n11319) );
  AOI22_X1 U15467 ( .A1(n20969), .A2(\xmem_data[86][7] ), .B1(n30882), .B2(
        \xmem_data[87][7] ), .ZN(n11318) );
  NAND4_X1 U15468 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11327) );
  AOI22_X1 U15469 ( .A1(n20962), .A2(\xmem_data[88][7] ), .B1(n28007), .B2(
        \xmem_data[89][7] ), .ZN(n11325) );
  AOI22_X1 U15470 ( .A1(n20961), .A2(\xmem_data[90][7] ), .B1(n30884), .B2(
        \xmem_data[91][7] ), .ZN(n11324) );
  AOI22_X1 U15471 ( .A1(n17013), .A2(\xmem_data[92][7] ), .B1(n20958), .B2(
        \xmem_data[93][7] ), .ZN(n11323) );
  AOI22_X1 U15472 ( .A1(n20959), .A2(\xmem_data[94][7] ), .B1(n21076), .B2(
        \xmem_data[95][7] ), .ZN(n11322) );
  NAND4_X1 U15473 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  OR4_X1 U15474 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11330) );
  AOI22_X1 U15475 ( .A1(n21088), .A2(n11331), .B1(n21086), .B2(n11330), .ZN(
        n11332) );
  XNOR2_X1 U15476 ( .A(n35401), .B(\fmem_data[0][3] ), .ZN(n30414) );
  AOI21_X1 U15477 ( .B1(n34537), .B2(n34535), .A(n30414), .ZN(n11334) );
  INV_X1 U15478 ( .A(n11334), .ZN(n34875) );
  FA_X1 U15479 ( .A(n11336), .B(n11335), .CI(n3906), .CO(n35173), .S(n12722)
         );
  OAI21_X1 U15480 ( .B1(n12721), .B2(n12720), .A(n12722), .ZN(n11338) );
  NAND2_X1 U15481 ( .A1(n12721), .A2(n12720), .ZN(n11337) );
  NAND2_X1 U15482 ( .A1(n11338), .A2(n11337), .ZN(n35154) );
  XNOR2_X1 U15483 ( .A(n35155), .B(n35154), .ZN(n12716) );
  FA_X1 U15484 ( .A(n11341), .B(n11340), .CI(n11339), .CO(n35096), .S(n12719)
         );
  BUF_X1 U15485 ( .A(n11436), .Z(n29590) );
  BUF_X2 U15486 ( .A(n11437), .Z(n29589) );
  AOI22_X1 U15487 ( .A1(n29481), .A2(\xmem_data[96][3] ), .B1(n30190), .B2(
        \xmem_data[97][3] ), .ZN(n11348) );
  NOR2_X1 U15488 ( .A1(n11344), .A2(n3377), .ZN(n11438) );
  BUF_X1 U15489 ( .A(n14997), .Z(n29591) );
  AOI22_X1 U15490 ( .A1(n3239), .A2(\xmem_data[98][3] ), .B1(n29591), .B2(
        \xmem_data[99][3] ), .ZN(n11347) );
  AOI22_X1 U15491 ( .A1(n29604), .A2(\xmem_data[100][3] ), .B1(n29648), .B2(
        \xmem_data[101][3] ), .ZN(n11346) );
  NAND3_X1 U15492 ( .A1(n11343), .A2(n11342), .A3(n6173), .ZN(n11370) );
  NOR2_X1 U15493 ( .A1(n11344), .A2(n11370), .ZN(n15833) );
  BUF_X1 U15494 ( .A(n15833), .Z(n29593) );
  AOI22_X1 U15495 ( .A1(n29593), .A2(\xmem_data[102][3] ), .B1(n25607), .B2(
        \xmem_data[103][3] ), .ZN(n11345) );
  AOI22_X1 U15496 ( .A1(n3166), .A2(\xmem_data[104][3] ), .B1(n3182), .B2(
        \xmem_data[105][3] ), .ZN(n11355) );
  AOI22_X1 U15497 ( .A1(n29610), .A2(\xmem_data[106][3] ), .B1(n29012), .B2(
        \xmem_data[107][3] ), .ZN(n11354) );
  AOI22_X1 U15498 ( .A1(n30198), .A2(\xmem_data[108][3] ), .B1(n30644), .B2(
        \xmem_data[109][3] ), .ZN(n11353) );
  NAND2_X1 U15499 ( .A1(n11350), .A2(n11349), .ZN(n11351) );
  NOR2_X1 U15500 ( .A1(n11370), .A2(n11351), .ZN(n15844) );
  BUF_X1 U15501 ( .A(n15844), .Z(n29574) );
  BUF_X1 U15502 ( .A(n14974), .Z(n29573) );
  AOI22_X1 U15503 ( .A1(n29574), .A2(\xmem_data[110][3] ), .B1(n29573), .B2(
        \xmem_data[111][3] ), .ZN(n11352) );
  BUF_X1 U15504 ( .A(n14988), .Z(n29565) );
  AOI22_X1 U15505 ( .A1(n29699), .A2(\xmem_data[122][3] ), .B1(n29565), .B2(
        \xmem_data[123][3] ), .ZN(n11379) );
  AOI22_X1 U15506 ( .A1(n30291), .A2(\xmem_data[120][3] ), .B1(n29831), .B2(
        \xmem_data[121][3] ), .ZN(n11356) );
  INV_X1 U15507 ( .A(n11356), .ZN(n11377) );
  BUF_X1 U15508 ( .A(n11484), .Z(n29566) );
  BUF_X1 U15509 ( .A(n11780), .Z(n29556) );
  AOI22_X1 U15510 ( .A1(n29566), .A2(\xmem_data[124][3] ), .B1(n27833), .B2(
        \xmem_data[125][3] ), .ZN(n11375) );
  NOR2_X1 U15511 ( .A1(n11358), .A2(n11363), .ZN(n11475) );
  BUF_X1 U15512 ( .A(n11475), .Z(n29580) );
  NOR2_X1 U15513 ( .A1(n11359), .A2(n11363), .ZN(n11453) );
  AOI22_X1 U15514 ( .A1(n29580), .A2(\xmem_data[112][3] ), .B1(n29615), .B2(
        \xmem_data[113][3] ), .ZN(n11367) );
  NOR2_X1 U15515 ( .A1(n11360), .A2(n11363), .ZN(n11476) );
  BUF_X1 U15516 ( .A(n11476), .Z(n29581) );
  AOI22_X1 U15517 ( .A1(n29581), .A2(\xmem_data[114][3] ), .B1(n20770), .B2(
        \xmem_data[115][3] ), .ZN(n11366) );
  NOR2_X1 U15518 ( .A1(n11361), .A2(n11363), .ZN(n11454) );
  NOR2_X1 U15519 ( .A1(n3246), .A2(n11363), .ZN(n11455) );
  BUF_X2 U15520 ( .A(n11455), .Z(n29582) );
  AOI22_X1 U15521 ( .A1(n29583), .A2(\xmem_data[116][3] ), .B1(n29582), .B2(
        \xmem_data[117][3] ), .ZN(n11365) );
  NOR2_X1 U15522 ( .A1(n11370), .A2(n11363), .ZN(n11456) );
  AOI22_X1 U15523 ( .A1(n29584), .A2(\xmem_data[118][3] ), .B1(n25443), .B2(
        \xmem_data[119][3] ), .ZN(n11364) );
  NAND4_X1 U15524 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11373) );
  NAND2_X1 U15525 ( .A1(n11368), .A2(n11350), .ZN(n11369) );
  NOR2_X1 U15526 ( .A1(n11370), .A2(n11369), .ZN(n11561) );
  AOI22_X1 U15527 ( .A1(n29568), .A2(\xmem_data[126][3] ), .B1(n3345), .B2(
        \xmem_data[127][3] ), .ZN(n11371) );
  INV_X1 U15528 ( .A(n11371), .ZN(n11372) );
  NOR2_X1 U15529 ( .A1(n11373), .A2(n11372), .ZN(n11374) );
  NAND2_X1 U15530 ( .A1(n11375), .A2(n11374), .ZN(n11376) );
  NOR2_X1 U15531 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  NAND4_X1 U15532 ( .A1(n3849), .A2(n3539), .A3(n11379), .A4(n11378), .ZN(
        n11384) );
  INV_X1 U15533 ( .A(n11380), .ZN(n37192) );
  NOR2_X1 U15534 ( .A1(n37192), .A2(n11381), .ZN(n11383) );
  XOR2_X1 U15535 ( .A(n11383), .B(load_xaddr_val[6]), .Z(n11434) );
  AND2_X1 U15536 ( .A1(n11467), .A2(n11434), .ZN(n29598) );
  NAND2_X1 U15537 ( .A1(n11384), .A2(n29598), .ZN(n11474) );
  AOI22_X1 U15538 ( .A1(n29446), .A2(\xmem_data[64][3] ), .B1(n3369), .B2(
        \xmem_data[65][3] ), .ZN(n11388) );
  AOI22_X1 U15539 ( .A1(n3239), .A2(\xmem_data[66][3] ), .B1(n29591), .B2(
        \xmem_data[67][3] ), .ZN(n11387) );
  AOI22_X1 U15540 ( .A1(n27754), .A2(\xmem_data[68][3] ), .B1(n30301), .B2(
        \xmem_data[69][3] ), .ZN(n11386) );
  AOI22_X1 U15541 ( .A1(n29593), .A2(\xmem_data[70][3] ), .B1(n17018), .B2(
        \xmem_data[71][3] ), .ZN(n11385) );
  NAND4_X1 U15542 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(
        n11394) );
  AOI22_X1 U15543 ( .A1(n3163), .A2(\xmem_data[72][3] ), .B1(n3190), .B2(
        \xmem_data[73][3] ), .ZN(n11392) );
  AOI22_X1 U15544 ( .A1(n30062), .A2(\xmem_data[74][3] ), .B1(n28687), .B2(
        \xmem_data[75][3] ), .ZN(n11391) );
  AOI22_X1 U15545 ( .A1(n29815), .A2(\xmem_data[76][3] ), .B1(n30644), .B2(
        \xmem_data[77][3] ), .ZN(n11390) );
  AOI22_X1 U15546 ( .A1(n29574), .A2(\xmem_data[78][3] ), .B1(n29573), .B2(
        \xmem_data[79][3] ), .ZN(n11389) );
  NAND4_X1 U15547 ( .A1(n11392), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(
        n11393) );
  OR2_X1 U15548 ( .A1(n11394), .A2(n11393), .ZN(n11410) );
  AOI22_X1 U15549 ( .A1(n27740), .A2(\xmem_data[90][3] ), .B1(n29565), .B2(
        \xmem_data[91][3] ), .ZN(n11408) );
  BUF_X1 U15550 ( .A(n11484), .Z(n29630) );
  BUF_X1 U15551 ( .A(n11780), .Z(n29629) );
  AOI22_X1 U15552 ( .A1(n29630), .A2(\xmem_data[92][3] ), .B1(n3197), .B2(
        \xmem_data[93][3] ), .ZN(n11395) );
  INV_X1 U15553 ( .A(n11395), .ZN(n11406) );
  AOI22_X1 U15554 ( .A1(n30223), .A2(\xmem_data[88][3] ), .B1(n27832), .B2(
        \xmem_data[89][3] ), .ZN(n11404) );
  BUF_X1 U15555 ( .A(n11475), .Z(n29616) );
  AOI22_X1 U15556 ( .A1(n29616), .A2(\xmem_data[80][3] ), .B1(n29655), .B2(
        \xmem_data[81][3] ), .ZN(n11399) );
  AOI22_X1 U15557 ( .A1(n29617), .A2(\xmem_data[82][3] ), .B1(n30901), .B2(
        \xmem_data[83][3] ), .ZN(n11398) );
  AOI22_X1 U15558 ( .A1(n29583), .A2(\xmem_data[84][3] ), .B1(n29582), .B2(
        \xmem_data[85][3] ), .ZN(n11397) );
  AOI22_X1 U15559 ( .A1(n29584), .A2(\xmem_data[86][3] ), .B1(n28164), .B2(
        \xmem_data[87][3] ), .ZN(n11396) );
  NAND4_X1 U15560 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11402) );
  AOI22_X1 U15561 ( .A1(n29568), .A2(\xmem_data[94][3] ), .B1(n3345), .B2(
        \xmem_data[95][3] ), .ZN(n11400) );
  INV_X1 U15562 ( .A(n11400), .ZN(n11401) );
  NOR2_X1 U15563 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U15564 ( .A1(n11404), .A2(n11403), .ZN(n11405) );
  NOR2_X1 U15565 ( .A1(n11406), .A2(n11405), .ZN(n11407) );
  NAND2_X1 U15566 ( .A1(n11408), .A2(n11407), .ZN(n11409) );
  INV_X1 U15567 ( .A(n11434), .ZN(n11468) );
  NOR2_X1 U15568 ( .A1(n11467), .A2(n11468), .ZN(n29600) );
  OAI21_X1 U15569 ( .B1(n11410), .B2(n11409), .A(n29600), .ZN(n11473) );
  BUF_X1 U15570 ( .A(n11436), .Z(n29647) );
  AOI22_X1 U15571 ( .A1(n29602), .A2(\xmem_data[0][3] ), .B1(n27761), .B2(
        \xmem_data[1][3] ), .ZN(n11414) );
  AOI22_X1 U15572 ( .A1(n3239), .A2(\xmem_data[2][3] ), .B1(n28152), .B2(
        \xmem_data[3][3] ), .ZN(n11413) );
  AOI22_X1 U15573 ( .A1(n28779), .A2(\xmem_data[4][3] ), .B1(n29768), .B2(
        \xmem_data[5][3] ), .ZN(n11412) );
  AOI22_X1 U15574 ( .A1(n15833), .A2(\xmem_data[6][3] ), .B1(n29605), .B2(
        \xmem_data[7][3] ), .ZN(n11411) );
  NAND4_X1 U15575 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11425) );
  AOI22_X1 U15576 ( .A1(n29580), .A2(\xmem_data[16][3] ), .B1(n29579), .B2(
        \xmem_data[17][3] ), .ZN(n11418) );
  BUF_X1 U15577 ( .A(n13420), .Z(n29657) );
  AOI22_X1 U15578 ( .A1(n29581), .A2(\xmem_data[18][3] ), .B1(n29657), .B2(
        \xmem_data[19][3] ), .ZN(n11417) );
  BUF_X1 U15579 ( .A(n11454), .Z(n29660) );
  AOI22_X1 U15580 ( .A1(n29660), .A2(\xmem_data[20][3] ), .B1(n29659), .B2(
        \xmem_data[21][3] ), .ZN(n11416) );
  BUF_X1 U15581 ( .A(n11456), .Z(n29662) );
  BUF_X1 U15582 ( .A(n28973), .Z(n29661) );
  AOI22_X1 U15583 ( .A1(n29662), .A2(\xmem_data[22][3] ), .B1(n29661), .B2(
        \xmem_data[23][3] ), .ZN(n11415) );
  NAND4_X1 U15584 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11421) );
  AOI22_X1 U15585 ( .A1(n11561), .A2(\xmem_data[30][3] ), .B1(n3146), .B2(
        \xmem_data[31][3] ), .ZN(n11419) );
  INV_X1 U15586 ( .A(n11419), .ZN(n11420) );
  NOR2_X1 U15587 ( .A1(n11421), .A2(n11420), .ZN(n11423) );
  AOI22_X1 U15588 ( .A1(n30217), .A2(\xmem_data[29][3] ), .B1(n29566), .B2(
        \xmem_data[28][3] ), .ZN(n11422) );
  NAND2_X1 U15589 ( .A1(n11423), .A2(n11422), .ZN(n11424) );
  NOR2_X1 U15590 ( .A1(n11425), .A2(n11424), .ZN(n11433) );
  AOI22_X1 U15591 ( .A1(n3164), .A2(\xmem_data[8][3] ), .B1(n3191), .B2(
        \xmem_data[9][3] ), .ZN(n11430) );
  BUF_X1 U15592 ( .A(n14971), .Z(n29639) );
  AOI22_X1 U15593 ( .A1(n27031), .A2(\xmem_data[10][3] ), .B1(n29639), .B2(
        \xmem_data[11][3] ), .ZN(n11429) );
  AOI22_X1 U15594 ( .A1(n29488), .A2(\xmem_data[12][3] ), .B1(n30266), .B2(
        \xmem_data[13][3] ), .ZN(n11428) );
  AOI22_X1 U15595 ( .A1(n15844), .A2(\xmem_data[14][3] ), .B1(n29324), .B2(
        \xmem_data[15][3] ), .ZN(n11427) );
  AOI22_X1 U15596 ( .A1(n30279), .A2(\xmem_data[26][3] ), .B1(n28218), .B2(
        \xmem_data[27][3] ), .ZN(n11432) );
  AOI22_X1 U15597 ( .A1(n29626), .A2(\xmem_data[24][3] ), .B1(n30106), .B2(
        \xmem_data[25][3] ), .ZN(n11431) );
  NAND4_X1 U15598 ( .A1(n11433), .A2(n3799), .A3(n11432), .A4(n11431), .ZN(
        n11435) );
  NOR2_X1 U15599 ( .A1(n11467), .A2(n11434), .ZN(n29681) );
  NAND2_X1 U15600 ( .A1(n11435), .A2(n29681), .ZN(n11472) );
  BUF_X1 U15601 ( .A(n11436), .Z(n29602) );
  AOI22_X1 U15602 ( .A1(n30633), .A2(\xmem_data[32][3] ), .B1(n28665), .B2(
        \xmem_data[33][3] ), .ZN(n11443) );
  BUF_X1 U15603 ( .A(n11438), .Z(n29603) );
  AOI22_X1 U15604 ( .A1(n29603), .A2(\xmem_data[34][3] ), .B1(n24157), .B2(
        \xmem_data[35][3] ), .ZN(n11442) );
  BUF_X1 U15605 ( .A(n11439), .Z(n29604) );
  AOI22_X1 U15606 ( .A1(n30250), .A2(\xmem_data[36][3] ), .B1(n26884), .B2(
        \xmem_data[37][3] ), .ZN(n11441) );
  BUF_X2 U15607 ( .A(n15833), .Z(n29649) );
  BUF_X1 U15608 ( .A(n29187), .Z(n29605) );
  AOI22_X1 U15609 ( .A1(n29649), .A2(\xmem_data[38][3] ), .B1(n27818), .B2(
        \xmem_data[39][3] ), .ZN(n11440) );
  NAND4_X1 U15610 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11450) );
  AOI22_X1 U15611 ( .A1(n3166), .A2(\xmem_data[40][3] ), .B1(n3190), .B2(
        \xmem_data[41][3] ), .ZN(n11448) );
  AOI22_X1 U15612 ( .A1(n30764), .A2(\xmem_data[42][3] ), .B1(n23722), .B2(
        \xmem_data[43][3] ), .ZN(n11447) );
  AOI22_X1 U15613 ( .A1(n28680), .A2(\xmem_data[44][3] ), .B1(n30170), .B2(
        \xmem_data[45][3] ), .ZN(n11446) );
  AOI22_X1 U15614 ( .A1(n29641), .A2(\xmem_data[46][3] ), .B1(n3300), .B2(
        \xmem_data[47][3] ), .ZN(n11445) );
  NAND4_X1 U15615 ( .A1(n11448), .A2(n11447), .A3(n11446), .A4(n11445), .ZN(
        n11449) );
  OR2_X1 U15616 ( .A1(n11450), .A2(n11449), .ZN(n11470) );
  BUF_X1 U15617 ( .A(n14988), .Z(n29627) );
  AOI22_X1 U15618 ( .A1(n29790), .A2(\xmem_data[58][3] ), .B1(n29627), .B2(
        \xmem_data[59][3] ), .ZN(n11466) );
  AOI22_X1 U15619 ( .A1(n29630), .A2(\xmem_data[60][3] ), .B1(n29556), .B2(
        \xmem_data[61][3] ), .ZN(n11465) );
  AOI22_X1 U15620 ( .A1(n28734), .A2(\xmem_data[56][3] ), .B1(n29697), .B2(
        \xmem_data[57][3] ), .ZN(n11464) );
  AOI22_X1 U15621 ( .A1(n29667), .A2(\xmem_data[62][3] ), .B1(n3374), .B2(
        \xmem_data[63][3] ), .ZN(n11452) );
  INV_X1 U15622 ( .A(n11452), .ZN(n11462) );
  BUF_X1 U15623 ( .A(n11453), .Z(n29615) );
  AOI22_X1 U15624 ( .A1(n29616), .A2(\xmem_data[48][3] ), .B1(n29615), .B2(
        \xmem_data[49][3] ), .ZN(n11460) );
  AOI22_X1 U15625 ( .A1(n29617), .A2(\xmem_data[50][3] ), .B1(n20567), .B2(
        \xmem_data[51][3] ), .ZN(n11459) );
  BUF_X1 U15626 ( .A(n11454), .Z(n29619) );
  BUF_X1 U15627 ( .A(n11455), .Z(n29618) );
  AOI22_X1 U15628 ( .A1(n29619), .A2(\xmem_data[52][3] ), .B1(n29618), .B2(
        \xmem_data[53][3] ), .ZN(n11458) );
  BUF_X1 U15629 ( .A(n11456), .Z(n29621) );
  BUF_X1 U15630 ( .A(n28973), .Z(n29620) );
  AOI22_X1 U15631 ( .A1(n29621), .A2(\xmem_data[54][3] ), .B1(n3142), .B2(
        \xmem_data[55][3] ), .ZN(n11457) );
  NAND4_X1 U15632 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11461) );
  NOR2_X1 U15633 ( .A1(n11462), .A2(n11461), .ZN(n11463) );
  NAND4_X1 U15634 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11469) );
  AND2_X1 U15635 ( .A1(n11468), .A2(n11467), .ZN(n29683) );
  OAI21_X1 U15636 ( .B1(n11470), .B2(n11469), .A(n29683), .ZN(n11471) );
  NAND4_X2 U15637 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n32440) );
  XNOR2_X1 U15638 ( .A(n32440), .B(\fmem_data[7][7] ), .ZN(n31939) );
  AOI22_X1 U15639 ( .A1(n28207), .A2(\xmem_data[90][2] ), .B1(n29565), .B2(
        \xmem_data[91][2] ), .ZN(n11488) );
  BUF_X1 U15640 ( .A(n11475), .Z(n29656) );
  AOI22_X1 U15641 ( .A1(n29656), .A2(\xmem_data[80][2] ), .B1(n29579), .B2(
        \xmem_data[81][2] ), .ZN(n11480) );
  BUF_X1 U15642 ( .A(n11476), .Z(n29658) );
  AOI22_X1 U15643 ( .A1(n29658), .A2(\xmem_data[82][2] ), .B1(n23753), .B2(
        \xmem_data[83][2] ), .ZN(n11479) );
  AOI22_X1 U15644 ( .A1(n29583), .A2(\xmem_data[84][2] ), .B1(n29582), .B2(
        \xmem_data[85][2] ), .ZN(n11478) );
  AOI22_X1 U15645 ( .A1(n29584), .A2(\xmem_data[86][2] ), .B1(n23754), .B2(
        \xmem_data[87][2] ), .ZN(n11477) );
  NAND4_X1 U15646 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(
        n11483) );
  AOI22_X1 U15647 ( .A1(n29568), .A2(\xmem_data[94][2] ), .B1(n3345), .B2(
        \xmem_data[95][2] ), .ZN(n11481) );
  INV_X1 U15648 ( .A(n11481), .ZN(n11482) );
  NOR2_X1 U15649 ( .A1(n11483), .A2(n11482), .ZN(n11487) );
  AOI22_X1 U15650 ( .A1(n28146), .A2(\xmem_data[64][2] ), .B1(n28665), .B2(
        \xmem_data[65][2] ), .ZN(n11486) );
  BUF_X1 U15651 ( .A(n11484), .Z(n29674) );
  AOI22_X1 U15652 ( .A1(n29674), .A2(\xmem_data[92][2] ), .B1(n27833), .B2(
        \xmem_data[93][2] ), .ZN(n11485) );
  NAND4_X1 U15653 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11506) );
  AOI22_X1 U15654 ( .A1(n30070), .A2(\xmem_data[74][2] ), .B1(n30617), .B2(
        \xmem_data[75][2] ), .ZN(n11504) );
  NAND2_X1 U15655 ( .A1(n29433), .A2(\xmem_data[88][2] ), .ZN(n11503) );
  AOI22_X1 U15656 ( .A1(n28680), .A2(\xmem_data[76][2] ), .B1(n29487), .B2(
        \xmem_data[77][2] ), .ZN(n11490) );
  INV_X1 U15657 ( .A(n11490), .ZN(n11493) );
  AOI22_X1 U15658 ( .A1(n29395), .A2(\xmem_data[68][2] ), .B1(n30237), .B2(
        \xmem_data[69][2] ), .ZN(n11491) );
  INV_X1 U15659 ( .A(n11491), .ZN(n11492) );
  NOR2_X1 U15660 ( .A1(n11493), .A2(n11492), .ZN(n11502) );
  AOI22_X1 U15661 ( .A1(n3166), .A2(\xmem_data[72][2] ), .B1(n3182), .B2(
        \xmem_data[73][2] ), .ZN(n11494) );
  INV_X1 U15662 ( .A(n11494), .ZN(n11500) );
  AOI22_X1 U15663 ( .A1(n29593), .A2(\xmem_data[70][2] ), .B1(n3466), .B2(
        \xmem_data[71][2] ), .ZN(n11498) );
  NAND2_X1 U15664 ( .A1(n28206), .A2(\xmem_data[89][2] ), .ZN(n11497) );
  AOI22_X1 U15665 ( .A1(n29574), .A2(\xmem_data[78][2] ), .B1(n29573), .B2(
        \xmem_data[79][2] ), .ZN(n11496) );
  AOI22_X1 U15666 ( .A1(n3239), .A2(\xmem_data[66][2] ), .B1(n29591), .B2(
        \xmem_data[67][2] ), .ZN(n11495) );
  NAND4_X1 U15667 ( .A1(n11498), .A2(n11497), .A3(n11496), .A4(n11495), .ZN(
        n11499) );
  NOR2_X1 U15668 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  NAND4_X1 U15669 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  OAI21_X1 U15670 ( .B1(n11506), .B2(n11505), .A(n29600), .ZN(n11584) );
  AOI22_X1 U15671 ( .A1(n28146), .A2(\xmem_data[32][2] ), .B1(n3368), .B2(
        \xmem_data[33][2] ), .ZN(n11510) );
  AOI22_X1 U15672 ( .A1(n29603), .A2(\xmem_data[34][2] ), .B1(n28743), .B2(
        \xmem_data[35][2] ), .ZN(n11509) );
  AOI22_X1 U15673 ( .A1(n30302), .A2(\xmem_data[36][2] ), .B1(n28684), .B2(
        \xmem_data[37][2] ), .ZN(n11508) );
  AOI22_X1 U15674 ( .A1(n29649), .A2(\xmem_data[38][2] ), .B1(n28053), .B2(
        \xmem_data[39][2] ), .ZN(n11507) );
  AOI22_X1 U15675 ( .A1(n26812), .A2(\xmem_data[42][2] ), .B1(n29639), .B2(
        \xmem_data[43][2] ), .ZN(n11514) );
  AOI22_X1 U15676 ( .A1(n3163), .A2(\xmem_data[40][2] ), .B1(n3188), .B2(
        \xmem_data[41][2] ), .ZN(n11513) );
  AOI22_X1 U15677 ( .A1(n30076), .A2(\xmem_data[44][2] ), .B1(n30266), .B2(
        \xmem_data[45][2] ), .ZN(n11512) );
  AOI22_X1 U15678 ( .A1(n29641), .A2(\xmem_data[46][2] ), .B1(n3328), .B2(
        \xmem_data[47][2] ), .ZN(n11511) );
  AOI22_X1 U15679 ( .A1(n29566), .A2(\xmem_data[60][2] ), .B1(n29629), .B2(
        \xmem_data[61][2] ), .ZN(n11515) );
  INV_X1 U15680 ( .A(n11515), .ZN(n11523) );
  AOI22_X1 U15681 ( .A1(n29580), .A2(\xmem_data[48][2] ), .B1(n29579), .B2(
        \xmem_data[49][2] ), .ZN(n11519) );
  AOI22_X1 U15682 ( .A1(n29581), .A2(\xmem_data[50][2] ), .B1(n31345), .B2(
        \xmem_data[51][2] ), .ZN(n11518) );
  AOI22_X1 U15683 ( .A1(n29619), .A2(\xmem_data[52][2] ), .B1(n29618), .B2(
        \xmem_data[53][2] ), .ZN(n11517) );
  AOI22_X1 U15684 ( .A1(n29621), .A2(\xmem_data[54][2] ), .B1(n3142), .B2(
        \xmem_data[55][2] ), .ZN(n11516) );
  NAND4_X1 U15685 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11522) );
  AOI22_X1 U15686 ( .A1(n29667), .A2(\xmem_data[62][2] ), .B1(n3126), .B2(
        \xmem_data[63][2] ), .ZN(n11520) );
  INV_X1 U15687 ( .A(n11520), .ZN(n11521) );
  NOR3_X1 U15688 ( .A1(n11523), .A2(n11522), .A3(n11521), .ZN(n11529) );
  AOI22_X1 U15689 ( .A1(n29788), .A2(\xmem_data[56][2] ), .B1(n29831), .B2(
        \xmem_data[57][2] ), .ZN(n11524) );
  INV_X1 U15690 ( .A(n11524), .ZN(n11527) );
  AOI22_X1 U15691 ( .A1(n28138), .A2(\xmem_data[58][2] ), .B1(n29627), .B2(
        \xmem_data[59][2] ), .ZN(n11525) );
  INV_X1 U15692 ( .A(n11525), .ZN(n11526) );
  NOR2_X1 U15693 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  NAND4_X1 U15694 ( .A1(n11530), .A2(n3814), .A3(n11529), .A4(n11528), .ZN(
        n11531) );
  NAND2_X1 U15695 ( .A1(n11531), .A2(n29683), .ZN(n11583) );
  NAND2_X1 U15696 ( .A1(n27710), .A2(\xmem_data[120][2] ), .ZN(n11533) );
  NAND2_X1 U15697 ( .A1(n29672), .A2(\xmem_data[121][2] ), .ZN(n11532) );
  NAND2_X1 U15698 ( .A1(n11533), .A2(n11532), .ZN(n11544) );
  AOI22_X1 U15699 ( .A1(n29674), .A2(\xmem_data[124][2] ), .B1(n30696), .B2(
        \xmem_data[125][2] ), .ZN(n11542) );
  AOI22_X1 U15700 ( .A1(n29656), .A2(\xmem_data[112][2] ), .B1(n29655), .B2(
        \xmem_data[113][2] ), .ZN(n11537) );
  AOI22_X1 U15701 ( .A1(n29658), .A2(\xmem_data[114][2] ), .B1(n20826), .B2(
        \xmem_data[115][2] ), .ZN(n11536) );
  AOI22_X1 U15702 ( .A1(n29583), .A2(\xmem_data[116][2] ), .B1(n29582), .B2(
        \xmem_data[117][2] ), .ZN(n11535) );
  AOI22_X1 U15703 ( .A1(n29584), .A2(\xmem_data[118][2] ), .B1(n28677), .B2(
        \xmem_data[119][2] ), .ZN(n11534) );
  NAND4_X1 U15704 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11540) );
  AOI22_X1 U15705 ( .A1(n29568), .A2(\xmem_data[126][2] ), .B1(n3345), .B2(
        \xmem_data[127][2] ), .ZN(n11538) );
  INV_X1 U15706 ( .A(n11538), .ZN(n11539) );
  NOR2_X1 U15707 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  NAND2_X1 U15708 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  NOR2_X1 U15709 ( .A1(n11544), .A2(n11543), .ZN(n11555) );
  AOI22_X1 U15710 ( .A1(n26812), .A2(\xmem_data[106][2] ), .B1(n20942), .B2(
        \xmem_data[107][2] ), .ZN(n11548) );
  AOI22_X1 U15711 ( .A1(n3166), .A2(\xmem_data[104][2] ), .B1(n3186), .B2(
        \xmem_data[105][2] ), .ZN(n11547) );
  AOI22_X1 U15712 ( .A1(n27713), .A2(\xmem_data[108][2] ), .B1(n30170), .B2(
        \xmem_data[109][2] ), .ZN(n11546) );
  AOI22_X1 U15713 ( .A1(n29574), .A2(\xmem_data[110][2] ), .B1(n29573), .B2(
        \xmem_data[111][2] ), .ZN(n11545) );
  AOI22_X1 U15714 ( .A1(n27740), .A2(\xmem_data[122][2] ), .B1(n29565), .B2(
        \xmem_data[123][2] ), .ZN(n11554) );
  AOI22_X1 U15715 ( .A1(n30743), .A2(\xmem_data[96][2] ), .B1(n3369), .B2(
        \xmem_data[97][2] ), .ZN(n11552) );
  AOI22_X1 U15716 ( .A1(n3239), .A2(\xmem_data[98][2] ), .B1(n29591), .B2(
        \xmem_data[99][2] ), .ZN(n11551) );
  AOI22_X1 U15717 ( .A1(n27754), .A2(\xmem_data[100][2] ), .B1(n27753), .B2(
        \xmem_data[101][2] ), .ZN(n11550) );
  AOI22_X1 U15718 ( .A1(n29593), .A2(\xmem_data[102][2] ), .B1(n21005), .B2(
        \xmem_data[103][2] ), .ZN(n11549) );
  AND4_X1 U15719 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11553) );
  NAND4_X1 U15720 ( .A1(n11555), .A2(n3815), .A3(n11554), .A4(n11553), .ZN(
        n11556) );
  NAND2_X1 U15721 ( .A1(n11556), .A2(n29598), .ZN(n11582) );
  AOI22_X1 U15722 ( .A1(n30633), .A2(\xmem_data[0][2] ), .B1(n29589), .B2(
        \xmem_data[1][2] ), .ZN(n11560) );
  AOI22_X1 U15723 ( .A1(n3239), .A2(\xmem_data[2][2] ), .B1(n28743), .B2(
        \xmem_data[3][2] ), .ZN(n11559) );
  AOI22_X1 U15724 ( .A1(n28751), .A2(\xmem_data[4][2] ), .B1(n29739), .B2(
        \xmem_data[5][2] ), .ZN(n11558) );
  AOI22_X1 U15725 ( .A1(n29649), .A2(\xmem_data[6][2] ), .B1(n25461), .B2(
        \xmem_data[7][2] ), .ZN(n11557) );
  NAND4_X1 U15726 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11572) );
  AOI22_X1 U15727 ( .A1(n29626), .A2(\xmem_data[24][2] ), .B1(n29697), .B2(
        \xmem_data[25][2] ), .ZN(n11570) );
  AOI22_X1 U15728 ( .A1(n11561), .A2(\xmem_data[30][2] ), .B1(n3131), .B2(
        \xmem_data[31][2] ), .ZN(n11562) );
  INV_X1 U15729 ( .A(n11562), .ZN(n11568) );
  AOI22_X1 U15730 ( .A1(n29616), .A2(\xmem_data[16][2] ), .B1(n29655), .B2(
        \xmem_data[17][2] ), .ZN(n11566) );
  AOI22_X1 U15731 ( .A1(n29617), .A2(\xmem_data[18][2] ), .B1(n29657), .B2(
        \xmem_data[19][2] ), .ZN(n11565) );
  AOI22_X1 U15732 ( .A1(n29660), .A2(\xmem_data[20][2] ), .B1(n29659), .B2(
        \xmem_data[21][2] ), .ZN(n11564) );
  AOI22_X1 U15733 ( .A1(n29662), .A2(\xmem_data[22][2] ), .B1(n29661), .B2(
        \xmem_data[23][2] ), .ZN(n11563) );
  NAND4_X1 U15734 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11567) );
  NOR2_X1 U15735 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  NAND2_X1 U15736 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  NOR2_X1 U15737 ( .A1(n11572), .A2(n11571), .ZN(n11579) );
  AOI22_X1 U15738 ( .A1(n3167), .A2(\xmem_data[8][2] ), .B1(n3187), .B2(
        \xmem_data[9][2] ), .ZN(n11576) );
  AOI22_X1 U15739 ( .A1(n28755), .A2(\xmem_data[10][2] ), .B1(n24115), .B2(
        \xmem_data[11][2] ), .ZN(n11575) );
  AOI22_X1 U15740 ( .A1(n30766), .A2(\xmem_data[12][2] ), .B1(n30170), .B2(
        \xmem_data[13][2] ), .ZN(n11574) );
  AOI22_X1 U15741 ( .A1(n29641), .A2(\xmem_data[14][2] ), .B1(n29246), .B2(
        \xmem_data[15][2] ), .ZN(n11573) );
  AOI22_X1 U15742 ( .A1(n29630), .A2(\xmem_data[28][2] ), .B1(n28208), .B2(
        \xmem_data[29][2] ), .ZN(n11578) );
  AOI22_X1 U15743 ( .A1(n29628), .A2(\xmem_data[26][2] ), .B1(n30278), .B2(
        \xmem_data[27][2] ), .ZN(n11577) );
  NAND4_X1 U15744 ( .A1(n11579), .A2(n3810), .A3(n11578), .A4(n11577), .ZN(
        n11580) );
  NAND2_X1 U15745 ( .A1(n11580), .A2(n29681), .ZN(n11581) );
  XNOR2_X1 U15746 ( .A(n33459), .B(\fmem_data[7][7] ), .ZN(n29684) );
  XOR2_X1 U15747 ( .A(\fmem_data[7][6] ), .B(\fmem_data[7][7] ), .Z(n11585) );
  OAI22_X1 U15748 ( .A1(n31939), .A2(n35619), .B1(n29684), .B2(n35618), .ZN(
        n20291) );
  AOI22_X1 U15749 ( .A1(n29849), .A2(\xmem_data[32][2] ), .B1(n29848), .B2(
        \xmem_data[33][2] ), .ZN(n11589) );
  AOI22_X1 U15750 ( .A1(n29851), .A2(\xmem_data[34][2] ), .B1(n29850), .B2(
        \xmem_data[35][2] ), .ZN(n11588) );
  AOI22_X1 U15751 ( .A1(n29853), .A2(\xmem_data[36][2] ), .B1(n29852), .B2(
        \xmem_data[37][2] ), .ZN(n11587) );
  AOI22_X1 U15752 ( .A1(n29855), .A2(\xmem_data[38][2] ), .B1(n29854), .B2(
        \xmem_data[39][2] ), .ZN(n11586) );
  NAND4_X1 U15753 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11605) );
  AOI22_X1 U15754 ( .A1(n29860), .A2(\xmem_data[40][2] ), .B1(n29976), .B2(
        \xmem_data[41][2] ), .ZN(n11593) );
  AOI22_X1 U15755 ( .A1(n29978), .A2(\xmem_data[42][2] ), .B1(n3194), .B2(
        \xmem_data[43][2] ), .ZN(n11592) );
  AOI22_X1 U15756 ( .A1(n29980), .A2(\xmem_data[44][2] ), .B1(n29979), .B2(
        \xmem_data[45][2] ), .ZN(n11591) );
  AOI22_X1 U15757 ( .A1(n29982), .A2(\xmem_data[46][2] ), .B1(n29981), .B2(
        \xmem_data[47][2] ), .ZN(n11590) );
  NAND4_X1 U15758 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11604) );
  AOI22_X1 U15759 ( .A1(n29866), .A2(\xmem_data[48][2] ), .B1(n29865), .B2(
        \xmem_data[49][2] ), .ZN(n11597) );
  AOI22_X1 U15760 ( .A1(n29868), .A2(\xmem_data[50][2] ), .B1(n29916), .B2(
        \xmem_data[51][2] ), .ZN(n11596) );
  AOI22_X1 U15761 ( .A1(n29870), .A2(\xmem_data[52][2] ), .B1(n29869), .B2(
        \xmem_data[53][2] ), .ZN(n11595) );
  AOI22_X1 U15762 ( .A1(n29871), .A2(\xmem_data[54][2] ), .B1(n29952), .B2(
        \xmem_data[55][2] ), .ZN(n11594) );
  NAND4_X1 U15763 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11603) );
  AOI22_X1 U15764 ( .A1(n29877), .A2(\xmem_data[56][2] ), .B1(n29876), .B2(
        \xmem_data[57][2] ), .ZN(n11601) );
  AOI22_X1 U15765 ( .A1(n29879), .A2(\xmem_data[58][2] ), .B1(n29878), .B2(
        \xmem_data[59][2] ), .ZN(n11600) );
  AOI22_X1 U15766 ( .A1(n29881), .A2(\xmem_data[60][2] ), .B1(n29880), .B2(
        \xmem_data[61][2] ), .ZN(n11599) );
  AOI22_X1 U15767 ( .A1(n29883), .A2(\xmem_data[62][2] ), .B1(n29882), .B2(
        \xmem_data[63][2] ), .ZN(n11598) );
  NAND4_X1 U15768 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11602) );
  INV_X1 U15769 ( .A(n29937), .ZN(n11669) );
  AOI22_X1 U15770 ( .A1(n29988), .A2(\xmem_data[112][2] ), .B1(n29987), .B2(
        \xmem_data[113][2] ), .ZN(n11609) );
  AOI22_X1 U15771 ( .A1(n29990), .A2(\xmem_data[114][2] ), .B1(n29989), .B2(
        \xmem_data[115][2] ), .ZN(n11608) );
  AOI22_X1 U15772 ( .A1(n29992), .A2(\xmem_data[116][2] ), .B1(n29991), .B2(
        \xmem_data[117][2] ), .ZN(n11607) );
  AOI22_X1 U15773 ( .A1(n29994), .A2(\xmem_data[118][2] ), .B1(n29920), .B2(
        \xmem_data[119][2] ), .ZN(n11606) );
  AOI22_X1 U15774 ( .A1(n3243), .A2(\xmem_data[120][2] ), .B1(n3242), .B2(
        \xmem_data[121][2] ), .ZN(n11613) );
  AOI22_X1 U15775 ( .A1(n3235), .A2(\xmem_data[122][2] ), .B1(n3238), .B2(
        \xmem_data[123][2] ), .ZN(n11612) );
  AOI22_X1 U15776 ( .A1(n3236), .A2(\xmem_data[124][2] ), .B1(n3225), .B2(
        \xmem_data[125][2] ), .ZN(n11611) );
  AOI22_X1 U15777 ( .A1(n3237), .A2(\xmem_data[126][2] ), .B1(n3234), .B2(
        \xmem_data[127][2] ), .ZN(n11610) );
  NAND4_X1 U15778 ( .A1(n11613), .A2(n11612), .A3(n11611), .A4(n11610), .ZN(
        n11619) );
  AOI22_X1 U15779 ( .A1(n29966), .A2(\xmem_data[96][2] ), .B1(n29965), .B2(
        \xmem_data[97][2] ), .ZN(n11617) );
  AOI22_X1 U15780 ( .A1(n29968), .A2(\xmem_data[98][2] ), .B1(n29967), .B2(
        \xmem_data[99][2] ), .ZN(n11616) );
  AOI22_X1 U15781 ( .A1(n29969), .A2(\xmem_data[100][2] ), .B1(n29896), .B2(
        \xmem_data[101][2] ), .ZN(n11615) );
  AOI22_X1 U15782 ( .A1(n29971), .A2(\xmem_data[102][2] ), .B1(n29970), .B2(
        \xmem_data[103][2] ), .ZN(n11614) );
  NAND4_X1 U15783 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11618) );
  AOI22_X1 U15784 ( .A1(n29977), .A2(\xmem_data[104][2] ), .B1(n29976), .B2(
        \xmem_data[105][2] ), .ZN(n11623) );
  AOI22_X1 U15785 ( .A1(n29905), .A2(\xmem_data[106][2] ), .B1(n3196), .B2(
        \xmem_data[107][2] ), .ZN(n11622) );
  AOI22_X1 U15786 ( .A1(n29907), .A2(\xmem_data[108][2] ), .B1(n29906), .B2(
        \xmem_data[109][2] ), .ZN(n11621) );
  AOI22_X1 U15787 ( .A1(n29909), .A2(\xmem_data[110][2] ), .B1(n29908), .B2(
        \xmem_data[111][2] ), .ZN(n11620) );
  NAND3_X1 U15788 ( .A1(n3537), .A2(n11624), .A3(n3905), .ZN(n11625) );
  NAND2_X1 U15789 ( .A1(n11625), .A2(n30007), .ZN(n11668) );
  AOI22_X1 U15790 ( .A1(n29988), .A2(\xmem_data[80][2] ), .B1(n29987), .B2(
        \xmem_data[81][2] ), .ZN(n11629) );
  AOI22_X1 U15791 ( .A1(n29990), .A2(\xmem_data[82][2] ), .B1(n29989), .B2(
        \xmem_data[83][2] ), .ZN(n11628) );
  AOI22_X1 U15792 ( .A1(n29992), .A2(\xmem_data[84][2] ), .B1(n29991), .B2(
        \xmem_data[85][2] ), .ZN(n11627) );
  AOI22_X1 U15793 ( .A1(n29994), .A2(\xmem_data[86][2] ), .B1(n29952), .B2(
        \xmem_data[87][2] ), .ZN(n11626) );
  AOI22_X1 U15794 ( .A1(n29966), .A2(\xmem_data[64][2] ), .B1(n29965), .B2(
        \xmem_data[65][2] ), .ZN(n11633) );
  AOI22_X1 U15795 ( .A1(n29968), .A2(\xmem_data[66][2] ), .B1(n29967), .B2(
        \xmem_data[67][2] ), .ZN(n11632) );
  AOI22_X1 U15796 ( .A1(n29969), .A2(\xmem_data[68][2] ), .B1(n29896), .B2(
        \xmem_data[69][2] ), .ZN(n11631) );
  AOI22_X1 U15797 ( .A1(n29971), .A2(\xmem_data[70][2] ), .B1(n29970), .B2(
        \xmem_data[71][2] ), .ZN(n11630) );
  AOI22_X1 U15798 ( .A1(n3243), .A2(\xmem_data[88][2] ), .B1(n3242), .B2(
        \xmem_data[89][2] ), .ZN(n11637) );
  AOI22_X1 U15799 ( .A1(n3235), .A2(\xmem_data[90][2] ), .B1(n3238), .B2(
        \xmem_data[91][2] ), .ZN(n11636) );
  AOI22_X1 U15800 ( .A1(n3236), .A2(\xmem_data[92][2] ), .B1(n3225), .B2(
        \xmem_data[93][2] ), .ZN(n11635) );
  AOI22_X1 U15801 ( .A1(n3237), .A2(\xmem_data[94][2] ), .B1(n3234), .B2(
        \xmem_data[95][2] ), .ZN(n11634) );
  AOI22_X1 U15802 ( .A1(n29977), .A2(\xmem_data[72][2] ), .B1(n29976), .B2(
        \xmem_data[73][2] ), .ZN(n11641) );
  AOI22_X1 U15803 ( .A1(n29978), .A2(\xmem_data[74][2] ), .B1(n3194), .B2(
        \xmem_data[75][2] ), .ZN(n11640) );
  AOI22_X1 U15804 ( .A1(n29980), .A2(\xmem_data[76][2] ), .B1(n29906), .B2(
        \xmem_data[77][2] ), .ZN(n11639) );
  AOI22_X1 U15805 ( .A1(n29982), .A2(\xmem_data[78][2] ), .B1(n29908), .B2(
        \xmem_data[79][2] ), .ZN(n11638) );
  NAND4_X1 U15806 ( .A1(n3843), .A2(n3538), .A3(n3475), .A4(n3472), .ZN(n11666) );
  NAND2_X1 U15807 ( .A1(n3195), .A2(\xmem_data[11][2] ), .ZN(n11643) );
  NAND2_X1 U15808 ( .A1(n29905), .A2(\xmem_data[10][2] ), .ZN(n11642) );
  NAND2_X1 U15809 ( .A1(n11643), .A2(n11642), .ZN(n11649) );
  AOI22_X1 U15810 ( .A1(\xmem_data[6][2] ), .A2(n29899), .B1(n29895), .B2(
        \xmem_data[2][2] ), .ZN(n11647) );
  AOI22_X1 U15811 ( .A1(\xmem_data[5][2] ), .A2(n29896), .B1(n29892), .B2(
        \xmem_data[1][2] ), .ZN(n11646) );
  AOI22_X1 U15812 ( .A1(\xmem_data[0][2] ), .A2(n29893), .B1(n29894), .B2(
        \xmem_data[3][2] ), .ZN(n11645) );
  AOI22_X1 U15813 ( .A1(\xmem_data[7][2] ), .A2(n29898), .B1(n29897), .B2(
        \xmem_data[4][2] ), .ZN(n11644) );
  NAND4_X1 U15814 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11648) );
  NOR2_X1 U15815 ( .A1(n11649), .A2(n11648), .ZN(n11664) );
  AOI22_X1 U15816 ( .A1(n29915), .A2(\xmem_data[16][2] ), .B1(n29914), .B2(
        \xmem_data[17][2] ), .ZN(n11653) );
  AOI22_X1 U15817 ( .A1(n29917), .A2(\xmem_data[18][2] ), .B1(n29916), .B2(
        \xmem_data[19][2] ), .ZN(n11652) );
  AOI22_X1 U15818 ( .A1(n29919), .A2(\xmem_data[20][2] ), .B1(n29918), .B2(
        \xmem_data[21][2] ), .ZN(n11651) );
  AOI22_X1 U15819 ( .A1(n29921), .A2(\xmem_data[22][2] ), .B1(n29952), .B2(
        \xmem_data[23][2] ), .ZN(n11650) );
  AOI22_X1 U15820 ( .A1(n3243), .A2(\xmem_data[24][2] ), .B1(n3242), .B2(
        \xmem_data[25][2] ), .ZN(n11657) );
  AOI22_X1 U15821 ( .A1(n3235), .A2(\xmem_data[26][2] ), .B1(n3238), .B2(
        \xmem_data[27][2] ), .ZN(n11656) );
  AOI22_X1 U15822 ( .A1(n3236), .A2(\xmem_data[28][2] ), .B1(n3225), .B2(
        \xmem_data[29][2] ), .ZN(n11655) );
  AOI22_X1 U15823 ( .A1(n3237), .A2(\xmem_data[30][2] ), .B1(n3234), .B2(
        \xmem_data[31][2] ), .ZN(n11654) );
  NAND4_X1 U15824 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11662) );
  AOI22_X1 U15825 ( .A1(n29982), .A2(\xmem_data[14][2] ), .B1(n29981), .B2(
        \xmem_data[15][2] ), .ZN(n11660) );
  AOI22_X1 U15826 ( .A1(n29980), .A2(\xmem_data[12][2] ), .B1(n29979), .B2(
        \xmem_data[13][2] ), .ZN(n11659) );
  AOI22_X1 U15827 ( .A1(n29904), .A2(\xmem_data[8][2] ), .B1(n29942), .B2(
        \xmem_data[9][2] ), .ZN(n11658) );
  NAND3_X1 U15828 ( .A1(n11660), .A2(n11659), .A3(n11658), .ZN(n11661) );
  NOR2_X1 U15829 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  NAND3_X1 U15830 ( .A1(n11664), .A2(n3803), .A3(n11663), .ZN(n11665) );
  AOI22_X1 U15831 ( .A1(n11666), .A2(n30009), .B1(n11665), .B2(n29935), .ZN(
        n11667) );
  XOR2_X1 U15832 ( .A(\fmem_data[1][6] ), .B(\fmem_data[1][7] ), .Z(n11670) );
  AOI22_X1 U15833 ( .A1(n29849), .A2(\xmem_data[32][3] ), .B1(n29848), .B2(
        \xmem_data[33][3] ), .ZN(n11674) );
  AOI22_X1 U15834 ( .A1(n29851), .A2(\xmem_data[34][3] ), .B1(n29850), .B2(
        \xmem_data[35][3] ), .ZN(n11673) );
  AOI22_X1 U15835 ( .A1(n29853), .A2(\xmem_data[36][3] ), .B1(n29852), .B2(
        \xmem_data[37][3] ), .ZN(n11672) );
  AOI22_X1 U15836 ( .A1(n29855), .A2(\xmem_data[38][3] ), .B1(n29854), .B2(
        \xmem_data[39][3] ), .ZN(n11671) );
  NAND4_X1 U15837 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11690) );
  AOI22_X1 U15838 ( .A1(n29860), .A2(\xmem_data[40][3] ), .B1(n29942), .B2(
        \xmem_data[41][3] ), .ZN(n11678) );
  AOI22_X1 U15839 ( .A1(n29978), .A2(\xmem_data[42][3] ), .B1(n3194), .B2(
        \xmem_data[43][3] ), .ZN(n11677) );
  AOI22_X1 U15840 ( .A1(n29980), .A2(\xmem_data[44][3] ), .B1(n29979), .B2(
        \xmem_data[45][3] ), .ZN(n11676) );
  AOI22_X1 U15841 ( .A1(n29982), .A2(\xmem_data[46][3] ), .B1(n29981), .B2(
        \xmem_data[47][3] ), .ZN(n11675) );
  NAND4_X1 U15842 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11689) );
  AOI22_X1 U15843 ( .A1(n29866), .A2(\xmem_data[48][3] ), .B1(n29865), .B2(
        \xmem_data[49][3] ), .ZN(n11682) );
  AOI22_X1 U15844 ( .A1(n29868), .A2(\xmem_data[50][3] ), .B1(n29867), .B2(
        \xmem_data[51][3] ), .ZN(n11681) );
  AOI22_X1 U15845 ( .A1(n29870), .A2(\xmem_data[52][3] ), .B1(n29869), .B2(
        \xmem_data[53][3] ), .ZN(n11680) );
  AOI22_X1 U15846 ( .A1(n29871), .A2(\xmem_data[54][3] ), .B1(n29920), .B2(
        \xmem_data[55][3] ), .ZN(n11679) );
  NAND4_X1 U15847 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(
        n11688) );
  AOI22_X1 U15848 ( .A1(n29877), .A2(\xmem_data[56][3] ), .B1(n29876), .B2(
        \xmem_data[57][3] ), .ZN(n11686) );
  AOI22_X1 U15849 ( .A1(n29879), .A2(\xmem_data[58][3] ), .B1(n29878), .B2(
        \xmem_data[59][3] ), .ZN(n11685) );
  AOI22_X1 U15850 ( .A1(n29881), .A2(\xmem_data[60][3] ), .B1(n29880), .B2(
        \xmem_data[61][3] ), .ZN(n11684) );
  AOI22_X1 U15851 ( .A1(n29883), .A2(\xmem_data[62][3] ), .B1(n29882), .B2(
        \xmem_data[63][3] ), .ZN(n11683) );
  NAND4_X1 U15852 ( .A1(n11686), .A2(n11685), .A3(n11684), .A4(n11683), .ZN(
        n11687) );
  OR4_X1 U15853 ( .A1(n11690), .A2(n11689), .A3(n11688), .A4(n11687), .ZN(
        n11710) );
  AOI22_X1 U15854 ( .A1(n29904), .A2(\xmem_data[8][3] ), .B1(n29976), .B2(
        \xmem_data[9][3] ), .ZN(n11694) );
  AOI22_X1 U15855 ( .A1(n29978), .A2(\xmem_data[10][3] ), .B1(n3194), .B2(
        \xmem_data[11][3] ), .ZN(n11693) );
  AOI22_X1 U15856 ( .A1(n29980), .A2(\xmem_data[12][3] ), .B1(n29944), .B2(
        \xmem_data[13][3] ), .ZN(n11692) );
  AOI22_X1 U15857 ( .A1(n29982), .A2(\xmem_data[14][3] ), .B1(n29946), .B2(
        \xmem_data[15][3] ), .ZN(n11691) );
  AOI22_X1 U15858 ( .A1(n29915), .A2(\xmem_data[16][3] ), .B1(n29914), .B2(
        \xmem_data[17][3] ), .ZN(n11698) );
  AOI22_X1 U15859 ( .A1(n29917), .A2(\xmem_data[18][3] ), .B1(n29916), .B2(
        \xmem_data[19][3] ), .ZN(n11697) );
  AOI22_X1 U15860 ( .A1(n29919), .A2(\xmem_data[20][3] ), .B1(n29918), .B2(
        \xmem_data[21][3] ), .ZN(n11696) );
  AOI22_X1 U15861 ( .A1(n29921), .A2(\xmem_data[22][3] ), .B1(n29920), .B2(
        \xmem_data[23][3] ), .ZN(n11695) );
  AOI22_X1 U15862 ( .A1(n29893), .A2(\xmem_data[0][3] ), .B1(n29892), .B2(
        \xmem_data[1][3] ), .ZN(n11704) );
  AOI22_X1 U15863 ( .A1(n29895), .A2(\xmem_data[2][3] ), .B1(n29894), .B2(
        \xmem_data[3][3] ), .ZN(n11703) );
  AOI22_X1 U15864 ( .A1(n29897), .A2(\xmem_data[4][3] ), .B1(n11699), .B2(
        \xmem_data[5][3] ), .ZN(n11702) );
  AOI22_X1 U15865 ( .A1(n29899), .A2(\xmem_data[6][3] ), .B1(n11700), .B2(
        \xmem_data[7][3] ), .ZN(n11701) );
  AOI22_X1 U15866 ( .A1(n3243), .A2(\xmem_data[24][3] ), .B1(n3242), .B2(
        \xmem_data[25][3] ), .ZN(n11708) );
  AOI22_X1 U15867 ( .A1(n3235), .A2(\xmem_data[26][3] ), .B1(n3238), .B2(
        \xmem_data[27][3] ), .ZN(n11707) );
  AOI22_X1 U15868 ( .A1(n3236), .A2(\xmem_data[28][3] ), .B1(n3225), .B2(
        \xmem_data[29][3] ), .ZN(n11706) );
  AOI22_X1 U15869 ( .A1(n3237), .A2(\xmem_data[30][3] ), .B1(n3234), .B2(
        \xmem_data[31][3] ), .ZN(n11705) );
  AOI22_X1 U15870 ( .A1(n11710), .A2(n29937), .B1(n29935), .B2(n11709), .ZN(
        n11754) );
  AOI22_X1 U15871 ( .A1(n29966), .A2(\xmem_data[96][3] ), .B1(n29965), .B2(
        \xmem_data[97][3] ), .ZN(n11714) );
  AOI22_X1 U15872 ( .A1(n29968), .A2(\xmem_data[98][3] ), .B1(n29967), .B2(
        \xmem_data[99][3] ), .ZN(n11713) );
  AOI22_X1 U15873 ( .A1(n29969), .A2(\xmem_data[100][3] ), .B1(n29896), .B2(
        \xmem_data[101][3] ), .ZN(n11712) );
  AOI22_X1 U15874 ( .A1(n29971), .A2(\xmem_data[102][3] ), .B1(n29970), .B2(
        \xmem_data[103][3] ), .ZN(n11711) );
  AND4_X1 U15875 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11730) );
  AOI22_X1 U15876 ( .A1(n29982), .A2(\xmem_data[110][3] ), .B1(n29946), .B2(
        \xmem_data[111][3] ), .ZN(n11718) );
  AOI22_X1 U15877 ( .A1(n29978), .A2(\xmem_data[106][3] ), .B1(n3196), .B2(
        \xmem_data[107][3] ), .ZN(n11717) );
  AOI22_X1 U15878 ( .A1(n29980), .A2(\xmem_data[108][3] ), .B1(n29944), .B2(
        \xmem_data[109][3] ), .ZN(n11716) );
  AOI22_X1 U15879 ( .A1(n29977), .A2(\xmem_data[104][3] ), .B1(n29942), .B2(
        \xmem_data[105][3] ), .ZN(n11715) );
  AND4_X1 U15880 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n11729) );
  AOI22_X1 U15881 ( .A1(n29988), .A2(\xmem_data[112][3] ), .B1(n29987), .B2(
        \xmem_data[113][3] ), .ZN(n11722) );
  AOI22_X1 U15882 ( .A1(n29990), .A2(\xmem_data[114][3] ), .B1(n29989), .B2(
        \xmem_data[115][3] ), .ZN(n11721) );
  AOI22_X1 U15883 ( .A1(n29992), .A2(\xmem_data[116][3] ), .B1(n29991), .B2(
        \xmem_data[117][3] ), .ZN(n11720) );
  AOI22_X1 U15884 ( .A1(n29994), .A2(\xmem_data[118][3] ), .B1(n29993), .B2(
        \xmem_data[119][3] ), .ZN(n11719) );
  AND4_X1 U15885 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11728) );
  AOI22_X1 U15886 ( .A1(n3243), .A2(\xmem_data[120][3] ), .B1(n3242), .B2(
        \xmem_data[121][3] ), .ZN(n11726) );
  AOI22_X1 U15887 ( .A1(n3235), .A2(\xmem_data[122][3] ), .B1(n3238), .B2(
        \xmem_data[123][3] ), .ZN(n11725) );
  AOI22_X1 U15888 ( .A1(n3236), .A2(\xmem_data[124][3] ), .B1(n3225), .B2(
        \xmem_data[125][3] ), .ZN(n11724) );
  AOI22_X1 U15889 ( .A1(n3237), .A2(\xmem_data[126][3] ), .B1(n3234), .B2(
        \xmem_data[127][3] ), .ZN(n11723) );
  AND4_X1 U15890 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11727) );
  NAND4_X1 U15891 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11752) );
  AOI22_X1 U15892 ( .A1(n29966), .A2(\xmem_data[64][3] ), .B1(n29965), .B2(
        \xmem_data[65][3] ), .ZN(n11734) );
  AOI22_X1 U15893 ( .A1(n29968), .A2(\xmem_data[66][3] ), .B1(n29967), .B2(
        \xmem_data[67][3] ), .ZN(n11733) );
  AOI22_X1 U15894 ( .A1(n29969), .A2(\xmem_data[68][3] ), .B1(n29896), .B2(
        \xmem_data[69][3] ), .ZN(n11732) );
  AOI22_X1 U15895 ( .A1(n29971), .A2(\xmem_data[70][3] ), .B1(n29970), .B2(
        \xmem_data[71][3] ), .ZN(n11731) );
  AND4_X1 U15896 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11750) );
  AOI22_X1 U15897 ( .A1(n29977), .A2(\xmem_data[72][3] ), .B1(n29976), .B2(
        \xmem_data[73][3] ), .ZN(n11738) );
  AOI22_X1 U15898 ( .A1(n29905), .A2(\xmem_data[74][3] ), .B1(n3196), .B2(
        \xmem_data[75][3] ), .ZN(n11737) );
  AOI22_X1 U15899 ( .A1(n29980), .A2(\xmem_data[76][3] ), .B1(n29944), .B2(
        \xmem_data[77][3] ), .ZN(n11736) );
  AOI22_X1 U15900 ( .A1(n29982), .A2(\xmem_data[78][3] ), .B1(n29946), .B2(
        \xmem_data[79][3] ), .ZN(n11735) );
  AND4_X1 U15901 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11749) );
  AOI22_X1 U15902 ( .A1(n29988), .A2(\xmem_data[80][3] ), .B1(n29987), .B2(
        \xmem_data[81][3] ), .ZN(n11742) );
  AOI22_X1 U15903 ( .A1(n29990), .A2(\xmem_data[82][3] ), .B1(n29989), .B2(
        \xmem_data[83][3] ), .ZN(n11741) );
  AOI22_X1 U15904 ( .A1(n29992), .A2(\xmem_data[84][3] ), .B1(n29991), .B2(
        \xmem_data[85][3] ), .ZN(n11740) );
  AOI22_X1 U15905 ( .A1(n29994), .A2(\xmem_data[86][3] ), .B1(n29920), .B2(
        \xmem_data[87][3] ), .ZN(n11739) );
  AND4_X1 U15906 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11748) );
  AOI22_X1 U15907 ( .A1(n3243), .A2(\xmem_data[88][3] ), .B1(n3242), .B2(
        \xmem_data[89][3] ), .ZN(n11746) );
  AOI22_X1 U15908 ( .A1(n3235), .A2(\xmem_data[90][3] ), .B1(n3238), .B2(
        \xmem_data[91][3] ), .ZN(n11745) );
  AOI22_X1 U15909 ( .A1(n3236), .A2(\xmem_data[92][3] ), .B1(n3225), .B2(
        \xmem_data[93][3] ), .ZN(n11744) );
  AOI22_X1 U15910 ( .A1(n3237), .A2(\xmem_data[94][3] ), .B1(n3234), .B2(
        \xmem_data[95][3] ), .ZN(n11743) );
  AND4_X1 U15911 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11747) );
  NAND4_X1 U15912 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  AOI22_X1 U15913 ( .A1(n30007), .A2(n11752), .B1(n30009), .B2(n11751), .ZN(
        n11753) );
  AOI22_X1 U15914 ( .A1(n30766), .A2(\xmem_data[96][3] ), .B1(n30765), .B2(
        \xmem_data[97][3] ), .ZN(n11758) );
  AOI22_X1 U15915 ( .A1(n27804), .A2(\xmem_data[98][3] ), .B1(n24522), .B2(
        \xmem_data[99][3] ), .ZN(n11757) );
  AOI22_X1 U15916 ( .A1(n28725), .A2(\xmem_data[100][3] ), .B1(n27805), .B2(
        \xmem_data[101][3] ), .ZN(n11756) );
  AOI22_X1 U15917 ( .A1(n27806), .A2(\xmem_data[102][3] ), .B1(n29383), .B2(
        \xmem_data[103][3] ), .ZN(n11755) );
  AND4_X1 U15918 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11774) );
  AOI22_X1 U15919 ( .A1(n7451), .A2(\xmem_data[104][3] ), .B1(n27812), .B2(
        \xmem_data[105][3] ), .ZN(n11762) );
  AOI22_X1 U15920 ( .A1(n27814), .A2(\xmem_data[106][3] ), .B1(n27813), .B2(
        \xmem_data[107][3] ), .ZN(n11761) );
  AOI22_X1 U15921 ( .A1(n29788), .A2(\xmem_data[108][3] ), .B1(n29831), .B2(
        \xmem_data[109][3] ), .ZN(n11760) );
  AOI22_X1 U15922 ( .A1(n29790), .A2(\xmem_data[110][3] ), .B1(n27831), .B2(
        \xmem_data[111][3] ), .ZN(n11759) );
  AND4_X1 U15923 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11773) );
  AOI22_X1 U15924 ( .A1(n27834), .A2(\xmem_data[112][3] ), .B1(n29629), .B2(
        \xmem_data[113][3] ), .ZN(n11766) );
  AOI22_X1 U15925 ( .A1(n3223), .A2(\xmem_data[114][3] ), .B1(n3140), .B2(
        \xmem_data[115][3] ), .ZN(n11765) );
  AOI22_X1 U15926 ( .A1(n29446), .A2(\xmem_data[116][3] ), .B1(n28665), .B2(
        \xmem_data[117][3] ), .ZN(n11764) );
  AOI22_X1 U15927 ( .A1(n29500), .A2(\xmem_data[118][3] ), .B1(n27763), .B2(
        \xmem_data[119][3] ), .ZN(n11763) );
  AND4_X1 U15928 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11772) );
  AOI22_X1 U15929 ( .A1(n30665), .A2(\xmem_data[120][3] ), .B1(n27728), .B2(
        \xmem_data[121][3] ), .ZN(n11770) );
  AOI22_X1 U15930 ( .A1(n27819), .A2(\xmem_data[122][3] ), .B1(n29237), .B2(
        \xmem_data[123][3] ), .ZN(n11769) );
  AOI22_X1 U15931 ( .A1(n3167), .A2(\xmem_data[124][3] ), .B1(n3185), .B2(
        \xmem_data[125][3] ), .ZN(n11768) );
  AOI22_X1 U15932 ( .A1(n30075), .A2(\xmem_data[126][3] ), .B1(n27825), .B2(
        \xmem_data[127][3] ), .ZN(n11767) );
  AND4_X1 U15933 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11771) );
  NAND4_X1 U15934 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11798) );
  AOI22_X1 U15935 ( .A1(n7451), .A2(\xmem_data[72][3] ), .B1(n27812), .B2(
        \xmem_data[73][3] ), .ZN(n11779) );
  AOI22_X1 U15936 ( .A1(n27814), .A2(\xmem_data[74][3] ), .B1(n27813), .B2(
        \xmem_data[75][3] ), .ZN(n11778) );
  AOI22_X1 U15937 ( .A1(n29433), .A2(\xmem_data[76][3] ), .B1(n29672), .B2(
        \xmem_data[77][3] ), .ZN(n11777) );
  AND2_X1 U15938 ( .A1(n27831), .A2(\xmem_data[79][3] ), .ZN(n11775) );
  AOI21_X1 U15939 ( .B1(n28207), .B2(\xmem_data[78][3] ), .A(n11775), .ZN(
        n11776) );
  NAND4_X1 U15940 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11796) );
  AOI22_X1 U15941 ( .A1(n27834), .A2(\xmem_data[80][3] ), .B1(n28667), .B2(
        \xmem_data[81][3] ), .ZN(n11784) );
  AOI22_X1 U15942 ( .A1(n3223), .A2(\xmem_data[82][3] ), .B1(n3131), .B2(
        \xmem_data[83][3] ), .ZN(n11783) );
  AOI22_X1 U15943 ( .A1(n30633), .A2(\xmem_data[84][3] ), .B1(n29589), .B2(
        \xmem_data[85][3] ), .ZN(n11782) );
  AOI22_X1 U15944 ( .A1(n29500), .A2(\xmem_data[86][3] ), .B1(n30083), .B2(
        \xmem_data[87][3] ), .ZN(n11781) );
  NAND4_X1 U15945 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11795) );
  AOI22_X1 U15946 ( .A1(n30745), .A2(\xmem_data[88][3] ), .B1(n29739), .B2(
        \xmem_data[89][3] ), .ZN(n11788) );
  AOI22_X1 U15947 ( .A1(n27819), .A2(\xmem_data[90][3] ), .B1(n27455), .B2(
        \xmem_data[91][3] ), .ZN(n11787) );
  AOI22_X1 U15948 ( .A1(n3163), .A2(\xmem_data[92][3] ), .B1(n3187), .B2(
        \xmem_data[93][3] ), .ZN(n11786) );
  AOI22_X1 U15949 ( .A1(n30310), .A2(\xmem_data[94][3] ), .B1(n25400), .B2(
        \xmem_data[95][3] ), .ZN(n11785) );
  NAND4_X1 U15950 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11794) );
  AOI22_X1 U15951 ( .A1(n29488), .A2(\xmem_data[64][3] ), .B1(n30644), .B2(
        \xmem_data[65][3] ), .ZN(n11792) );
  AOI22_X1 U15952 ( .A1(n27804), .A2(\xmem_data[66][3] ), .B1(n20950), .B2(
        \xmem_data[67][3] ), .ZN(n11791) );
  AOI22_X1 U15953 ( .A1(n29382), .A2(\xmem_data[68][3] ), .B1(n27805), .B2(
        \xmem_data[69][3] ), .ZN(n11790) );
  AOI22_X1 U15954 ( .A1(n27806), .A2(\xmem_data[70][3] ), .B1(n27717), .B2(
        \xmem_data[71][3] ), .ZN(n11789) );
  NAND4_X1 U15955 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  AOI22_X1 U15956 ( .A1(n11798), .A2(n27801), .B1(n27839), .B2(n11797), .ZN(
        n27329) );
  AOI22_X1 U15957 ( .A1(n29722), .A2(\xmem_data[0][3] ), .B1(n30170), .B2(
        \xmem_data[1][3] ), .ZN(n11803) );
  AOI22_X1 U15958 ( .A1(n28681), .A2(\xmem_data[6][3] ), .B1(n29327), .B2(
        \xmem_data[7][3] ), .ZN(n11801) );
  AOI22_X1 U15959 ( .A1(n29463), .A2(\xmem_data[4][3] ), .B1(n29723), .B2(
        \xmem_data[5][3] ), .ZN(n11800) );
  AOI22_X1 U15960 ( .A1(n27804), .A2(\xmem_data[2][3] ), .B1(n28701), .B2(
        \xmem_data[3][3] ), .ZN(n11799) );
  AND3_X1 U15961 ( .A1(n11801), .A2(n11800), .A3(n11799), .ZN(n11802) );
  NAND2_X1 U15962 ( .A1(n11803), .A2(n11802), .ZN(n11819) );
  AOI22_X1 U15963 ( .A1(n28765), .A2(\xmem_data[8][3] ), .B1(n27743), .B2(
        \xmem_data[9][3] ), .ZN(n11807) );
  AOI22_X1 U15964 ( .A1(n27742), .A2(\xmem_data[10][3] ), .B1(n3144), .B2(
        \xmem_data[11][3] ), .ZN(n11806) );
  AOI22_X1 U15965 ( .A1(n28136), .A2(\xmem_data[12][3] ), .B1(n30100), .B2(
        \xmem_data[13][3] ), .ZN(n11805) );
  AOI22_X1 U15966 ( .A1(n29628), .A2(\xmem_data[14][3] ), .B1(n28218), .B2(
        \xmem_data[15][3] ), .ZN(n11804) );
  NAND4_X1 U15967 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11818) );
  AOI22_X1 U15968 ( .A1(n27811), .A2(\xmem_data[24][3] ), .B1(n28684), .B2(
        \xmem_data[25][3] ), .ZN(n11811) );
  AOI22_X1 U15969 ( .A1(n27756), .A2(\xmem_data[26][3] ), .B1(n28154), .B2(
        \xmem_data[27][3] ), .ZN(n11810) );
  AOI22_X1 U15970 ( .A1(n3165), .A2(\xmem_data[28][3] ), .B1(n11426), .B2(
        \xmem_data[29][3] ), .ZN(n11809) );
  AOI22_X1 U15971 ( .A1(n30764), .A2(\xmem_data[30][3] ), .B1(n27825), .B2(
        \xmem_data[31][3] ), .ZN(n11808) );
  NAND4_X1 U15972 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11817) );
  AOI22_X1 U15973 ( .A1(n30743), .A2(\xmem_data[20][3] ), .B1(n29482), .B2(
        \xmem_data[21][3] ), .ZN(n11815) );
  AOI22_X1 U15974 ( .A1(n3223), .A2(\xmem_data[18][3] ), .B1(n3131), .B2(
        \xmem_data[19][3] ), .ZN(n11814) );
  AOI22_X1 U15975 ( .A1(n27771), .A2(\xmem_data[16][3] ), .B1(n29556), .B2(
        \xmem_data[17][3] ), .ZN(n11813) );
  AOI22_X1 U15976 ( .A1(n29709), .A2(\xmem_data[22][3] ), .B1(n30083), .B2(
        \xmem_data[23][3] ), .ZN(n11812) );
  NAND4_X1 U15977 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11816) );
  OR4_X1 U15978 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11841) );
  AOI22_X1 U15979 ( .A1(n29786), .A2(\xmem_data[40][3] ), .B1(n27723), .B2(
        \xmem_data[41][3] ), .ZN(n11823) );
  AOI22_X1 U15980 ( .A1(n27742), .A2(\xmem_data[42][3] ), .B1(n3149), .B2(
        \xmem_data[43][3] ), .ZN(n11822) );
  AOI22_X1 U15981 ( .A1(n29421), .A2(\xmem_data[44][3] ), .B1(n29432), .B2(
        \xmem_data[45][3] ), .ZN(n11821) );
  AOI22_X1 U15982 ( .A1(n29628), .A2(\xmem_data[46][3] ), .B1(n27708), .B2(
        \xmem_data[47][3] ), .ZN(n11820) );
  NAND4_X1 U15983 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11839) );
  AOI22_X1 U15984 ( .A1(n27701), .A2(\xmem_data[48][3] ), .B1(n29761), .B2(
        \xmem_data[49][3] ), .ZN(n11827) );
  AOI22_X1 U15985 ( .A1(n27702), .A2(\xmem_data[50][3] ), .B1(n3132), .B2(
        \xmem_data[51][3] ), .ZN(n11826) );
  AOI22_X1 U15986 ( .A1(n29705), .A2(\xmem_data[52][3] ), .B1(n3369), .B2(
        \xmem_data[53][3] ), .ZN(n11825) );
  AOI22_X1 U15987 ( .A1(n26879), .A2(\xmem_data[54][3] ), .B1(n30083), .B2(
        \xmem_data[55][3] ), .ZN(n11824) );
  NAND4_X1 U15988 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11838) );
  AOI22_X1 U15989 ( .A1(n30635), .A2(\xmem_data[56][3] ), .B1(n27728), .B2(
        \xmem_data[57][3] ), .ZN(n11831) );
  AOI22_X1 U15990 ( .A1(n27729), .A2(\xmem_data[58][3] ), .B1(n21048), .B2(
        \xmem_data[59][3] ), .ZN(n11830) );
  AOI22_X1 U15991 ( .A1(n3167), .A2(\xmem_data[60][3] ), .B1(n3186), .B2(
        \xmem_data[61][3] ), .ZN(n11829) );
  AOI22_X1 U15992 ( .A1(n29716), .A2(\xmem_data[62][3] ), .B1(n29639), .B2(
        \xmem_data[63][3] ), .ZN(n11828) );
  NAND4_X1 U15993 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11837) );
  AOI22_X1 U15994 ( .A1(n30063), .A2(\xmem_data[32][3] ), .B1(n30765), .B2(
        \xmem_data[33][3] ), .ZN(n11835) );
  AOI22_X1 U15995 ( .A1(n27714), .A2(\xmem_data[34][3] ), .B1(n23780), .B2(
        \xmem_data[35][3] ), .ZN(n11834) );
  AOI22_X1 U15996 ( .A1(n27716), .A2(\xmem_data[36][3] ), .B1(n27715), .B2(
        \xmem_data[37][3] ), .ZN(n11833) );
  AOI22_X1 U15997 ( .A1(n27718), .A2(\xmem_data[38][3] ), .B1(n27717), .B2(
        \xmem_data[39][3] ), .ZN(n11832) );
  NAND4_X1 U15998 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11836) );
  AOI22_X1 U15999 ( .A1(n11841), .A2(n27778), .B1(n11840), .B2(n27737), .ZN(
        n27328) );
  NAND2_X1 U16000 ( .A1(n3258), .A2(n27328), .ZN(n11842) );
  XNOR2_X1 U16001 ( .A(n11842), .B(\fmem_data[27][7] ), .ZN(n31937) );
  AOI22_X1 U16002 ( .A1(n30743), .A2(\xmem_data[84][2] ), .B1(n3369), .B2(
        \xmem_data[85][2] ), .ZN(n11843) );
  INV_X1 U16003 ( .A(n11843), .ZN(n11858) );
  AOI22_X1 U16004 ( .A1(n3162), .A2(\xmem_data[92][2] ), .B1(n3185), .B2(
        \xmem_data[93][2] ), .ZN(n11856) );
  NAND2_X1 U16005 ( .A1(n27812), .A2(\xmem_data[73][2] ), .ZN(n11845) );
  NAND2_X1 U16006 ( .A1(n7451), .A2(\xmem_data[72][2] ), .ZN(n11844) );
  NAND2_X1 U16007 ( .A1(n11845), .A2(n11844), .ZN(n11854) );
  AOI22_X1 U16008 ( .A1(n26879), .A2(\xmem_data[86][2] ), .B1(n27763), .B2(
        \xmem_data[87][2] ), .ZN(n11849) );
  AOI22_X1 U16009 ( .A1(n11846), .A2(\xmem_data[90][2] ), .B1(n28336), .B2(
        \xmem_data[91][2] ), .ZN(n11848) );
  AOI22_X1 U16010 ( .A1(n26878), .A2(\xmem_data[82][2] ), .B1(n3140), .B2(
        \xmem_data[83][2] ), .ZN(n11847) );
  NAND3_X1 U16011 ( .A1(n11849), .A2(n11848), .A3(n11847), .ZN(n11853) );
  AOI22_X1 U16012 ( .A1(n11850), .A2(\xmem_data[74][2] ), .B1(n27813), .B2(
        \xmem_data[75][2] ), .ZN(n11851) );
  INV_X1 U16013 ( .A(n11851), .ZN(n11852) );
  NOR3_X1 U16014 ( .A1(n11854), .A2(n11853), .A3(n11852), .ZN(n11855) );
  NAND2_X1 U16015 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  NOR2_X1 U16016 ( .A1(n11858), .A2(n11857), .ZN(n11866) );
  AOI22_X1 U16017 ( .A1(n27834), .A2(\xmem_data[80][2] ), .B1(n3198), .B2(
        \xmem_data[81][2] ), .ZN(n11865) );
  AOI22_X1 U16018 ( .A1(n30684), .A2(\xmem_data[94][2] ), .B1(n28754), .B2(
        \xmem_data[95][2] ), .ZN(n11859) );
  INV_X1 U16019 ( .A(n11859), .ZN(n11862) );
  AOI22_X1 U16020 ( .A1(n29769), .A2(\xmem_data[88][2] ), .B1(n29592), .B2(
        \xmem_data[89][2] ), .ZN(n11860) );
  INV_X1 U16021 ( .A(n11860), .ZN(n11861) );
  NOR2_X1 U16022 ( .A1(n11862), .A2(n11861), .ZN(n11864) );
  AOI22_X1 U16023 ( .A1(n28207), .A2(\xmem_data[78][2] ), .B1(n27831), .B2(
        \xmem_data[79][2] ), .ZN(n11863) );
  NAND4_X1 U16024 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11874) );
  AND2_X1 U16025 ( .A1(n29432), .A2(\xmem_data[77][2] ), .ZN(n11867) );
  AOI21_X1 U16026 ( .B1(n28136), .B2(\xmem_data[76][2] ), .A(n11867), .ZN(
        n11872) );
  AOI22_X1 U16027 ( .A1(n27713), .A2(\xmem_data[64][2] ), .B1(n29487), .B2(
        \xmem_data[65][2] ), .ZN(n11871) );
  AOI22_X1 U16028 ( .A1(n27804), .A2(\xmem_data[66][2] ), .B1(n20732), .B2(
        \xmem_data[67][2] ), .ZN(n11870) );
  AOI22_X1 U16029 ( .A1(n29382), .A2(\xmem_data[68][2] ), .B1(n27805), .B2(
        \xmem_data[69][2] ), .ZN(n11869) );
  AOI22_X1 U16030 ( .A1(n27806), .A2(\xmem_data[70][2] ), .B1(n29657), .B2(
        \xmem_data[71][2] ), .ZN(n11868) );
  NAND2_X1 U16031 ( .A1(n11872), .A2(n3750), .ZN(n11873) );
  OAI21_X1 U16032 ( .B1(n11874), .B2(n11873), .A(n27839), .ZN(n11954) );
  AOI22_X1 U16033 ( .A1(n30076), .A2(\xmem_data[0][2] ), .B1(n30644), .B2(
        \xmem_data[1][2] ), .ZN(n11878) );
  AOI22_X1 U16034 ( .A1(n7446), .A2(\xmem_data[2][2] ), .B1(n29379), .B2(
        \xmem_data[3][2] ), .ZN(n11877) );
  AOI22_X1 U16035 ( .A1(n29777), .A2(\xmem_data[4][2] ), .B1(n29462), .B2(
        \xmem_data[5][2] ), .ZN(n11876) );
  AOI22_X1 U16036 ( .A1(n29464), .A2(\xmem_data[6][2] ), .B1(n23753), .B2(
        \xmem_data[7][2] ), .ZN(n11875) );
  AOI22_X1 U16037 ( .A1(n29705), .A2(\xmem_data[20][2] ), .B1(n29589), .B2(
        \xmem_data[21][2] ), .ZN(n11879) );
  INV_X1 U16038 ( .A(n11879), .ZN(n11885) );
  NAND2_X1 U16039 ( .A1(n29626), .A2(\xmem_data[12][2] ), .ZN(n11883) );
  AOI22_X1 U16040 ( .A1(n27742), .A2(\xmem_data[10][2] ), .B1(n28245), .B2(
        \xmem_data[11][2] ), .ZN(n11882) );
  AOI22_X1 U16041 ( .A1(n28765), .A2(\xmem_data[8][2] ), .B1(n27743), .B2(
        \xmem_data[9][2] ), .ZN(n11881) );
  NAND2_X1 U16042 ( .A1(n29831), .A2(\xmem_data[13][2] ), .ZN(n11880) );
  NAND4_X1 U16043 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11884) );
  NOR2_X1 U16044 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  NAND2_X1 U16045 ( .A1(n3804), .A2(n11886), .ZN(n11900) );
  AOI22_X1 U16046 ( .A1(n3165), .A2(\xmem_data[28][2] ), .B1(n3187), .B2(
        \xmem_data[29][2] ), .ZN(n11895) );
  AOI22_X1 U16047 ( .A1(n29476), .A2(\xmem_data[30][2] ), .B1(n27825), .B2(
        \xmem_data[31][2] ), .ZN(n11894) );
  AOI22_X1 U16048 ( .A1(n30250), .A2(\xmem_data[24][2] ), .B1(n30193), .B2(
        \xmem_data[25][2] ), .ZN(n11893) );
  AOI22_X1 U16049 ( .A1(n29709), .A2(\xmem_data[22][2] ), .B1(n27763), .B2(
        \xmem_data[23][2] ), .ZN(n11887) );
  INV_X1 U16050 ( .A(n11887), .ZN(n11891) );
  AOI22_X1 U16051 ( .A1(n3223), .A2(\xmem_data[18][2] ), .B1(n3140), .B2(
        \xmem_data[19][2] ), .ZN(n11889) );
  AOI22_X1 U16052 ( .A1(n27756), .A2(\xmem_data[26][2] ), .B1(n30303), .B2(
        \xmem_data[27][2] ), .ZN(n11888) );
  NAND2_X1 U16053 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  NOR2_X1 U16054 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  AOI22_X1 U16055 ( .A1(n29423), .A2(\xmem_data[14][2] ), .B1(n30278), .B2(
        \xmem_data[15][2] ), .ZN(n11897) );
  AOI22_X1 U16056 ( .A1(n27771), .A2(\xmem_data[16][2] ), .B1(n30293), .B2(
        \xmem_data[17][2] ), .ZN(n11896) );
  OAI21_X1 U16057 ( .B1(n11900), .B2(n11899), .A(n27778), .ZN(n11953) );
  AOI22_X1 U16058 ( .A1(n3162), .A2(\xmem_data[124][2] ), .B1(n3185), .B2(
        \xmem_data[125][2] ), .ZN(n11901) );
  INV_X1 U16059 ( .A(n11901), .ZN(n11907) );
  AOI22_X1 U16060 ( .A1(n28751), .A2(\xmem_data[120][2] ), .B1(n29768), .B2(
        \xmem_data[121][2] ), .ZN(n11903) );
  AOI22_X1 U16061 ( .A1(n27819), .A2(\xmem_data[122][2] ), .B1(n24213), .B2(
        \xmem_data[123][2] ), .ZN(n11902) );
  NAND2_X1 U16062 ( .A1(n11903), .A2(n11902), .ZN(n11906) );
  NAND2_X1 U16063 ( .A1(n30310), .A2(\xmem_data[126][2] ), .ZN(n11904) );
  NAND2_X1 U16064 ( .A1(n11904), .A2(n3980), .ZN(n11905) );
  NOR3_X1 U16065 ( .A1(n11907), .A2(n11906), .A3(n11905), .ZN(n11920) );
  AOI22_X1 U16066 ( .A1(n29801), .A2(\xmem_data[116][2] ), .B1(n29347), .B2(
        \xmem_data[117][2] ), .ZN(n11908) );
  INV_X1 U16067 ( .A(n11908), .ZN(n11912) );
  AOI22_X1 U16068 ( .A1(n29500), .A2(\xmem_data[118][2] ), .B1(n27763), .B2(
        \xmem_data[119][2] ), .ZN(n11910) );
  AOI22_X1 U16069 ( .A1(n3223), .A2(\xmem_data[114][2] ), .B1(n3140), .B2(
        \xmem_data[115][2] ), .ZN(n11909) );
  NAND2_X1 U16070 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  NOR2_X1 U16071 ( .A1(n11912), .A2(n11911), .ZN(n11919) );
  AOI22_X1 U16072 ( .A1(n28173), .A2(\xmem_data[96][2] ), .B1(n30685), .B2(
        \xmem_data[97][2] ), .ZN(n11916) );
  AOI22_X1 U16073 ( .A1(n27804), .A2(\xmem_data[98][2] ), .B1(n29573), .B2(
        \xmem_data[99][2] ), .ZN(n11915) );
  AOI22_X1 U16074 ( .A1(n28725), .A2(\xmem_data[100][2] ), .B1(n27805), .B2(
        \xmem_data[101][2] ), .ZN(n11914) );
  AOI22_X1 U16075 ( .A1(n27806), .A2(\xmem_data[102][2] ), .B1(n27717), .B2(
        \xmem_data[103][2] ), .ZN(n11913) );
  AOI22_X1 U16076 ( .A1(n27834), .A2(\xmem_data[112][2] ), .B1(n29708), .B2(
        \xmem_data[113][2] ), .ZN(n11917) );
  NAND4_X1 U16077 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11926) );
  AOI22_X1 U16078 ( .A1(n7451), .A2(\xmem_data[104][2] ), .B1(n27812), .B2(
        \xmem_data[105][2] ), .ZN(n11924) );
  AOI22_X1 U16079 ( .A1(n27814), .A2(\xmem_data[106][2] ), .B1(n27813), .B2(
        \xmem_data[107][2] ), .ZN(n11923) );
  AOI22_X1 U16080 ( .A1(n30291), .A2(\xmem_data[108][2] ), .B1(n27832), .B2(
        \xmem_data[109][2] ), .ZN(n11922) );
  AOI22_X1 U16081 ( .A1(n30215), .A2(\xmem_data[110][2] ), .B1(n27831), .B2(
        \xmem_data[111][2] ), .ZN(n11921) );
  NAND4_X1 U16082 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11925) );
  OAI21_X1 U16083 ( .B1(n11926), .B2(n11925), .A(n27801), .ZN(n11952) );
  NAND2_X1 U16084 ( .A1(n23901), .A2(\xmem_data[62][2] ), .ZN(n11928) );
  NAND2_X1 U16085 ( .A1(n29047), .A2(\xmem_data[63][2] ), .ZN(n11927) );
  NAND2_X1 U16086 ( .A1(n11928), .A2(n11927), .ZN(n11933) );
  AOI22_X1 U16087 ( .A1(n3163), .A2(\xmem_data[60][2] ), .B1(n3182), .B2(
        \xmem_data[61][2] ), .ZN(n11931) );
  AOI22_X1 U16088 ( .A1(n27729), .A2(\xmem_data[58][2] ), .B1(n24545), .B2(
        \xmem_data[59][2] ), .ZN(n11930) );
  AOI22_X1 U16089 ( .A1(n28751), .A2(\xmem_data[56][2] ), .B1(n29592), .B2(
        \xmem_data[57][2] ), .ZN(n11929) );
  NAND3_X1 U16090 ( .A1(n11931), .A2(n11930), .A3(n11929), .ZN(n11932) );
  NOR2_X1 U16091 ( .A1(n11933), .A2(n11932), .ZN(n11944) );
  AOI22_X1 U16092 ( .A1(n30198), .A2(\xmem_data[32][2] ), .B1(n29640), .B2(
        \xmem_data[33][2] ), .ZN(n11937) );
  AOI22_X1 U16093 ( .A1(n27714), .A2(\xmem_data[34][2] ), .B1(n30600), .B2(
        \xmem_data[35][2] ), .ZN(n11936) );
  AOI22_X1 U16094 ( .A1(n27716), .A2(\xmem_data[36][2] ), .B1(n27715), .B2(
        \xmem_data[37][2] ), .ZN(n11935) );
  AOI22_X1 U16095 ( .A1(n27718), .A2(\xmem_data[38][2] ), .B1(n27717), .B2(
        \xmem_data[39][2] ), .ZN(n11934) );
  AOI22_X1 U16096 ( .A1(n27701), .A2(\xmem_data[48][2] ), .B1(n30776), .B2(
        \xmem_data[49][2] ), .ZN(n11943) );
  AOI22_X1 U16097 ( .A1(n26879), .A2(\xmem_data[54][2] ), .B1(n27763), .B2(
        \xmem_data[55][2] ), .ZN(n11939) );
  AOI22_X1 U16098 ( .A1(n27702), .A2(\xmem_data[50][2] ), .B1(n3140), .B2(
        \xmem_data[51][2] ), .ZN(n11938) );
  NAND2_X1 U16099 ( .A1(n11939), .A2(n11938), .ZN(n11941) );
  NOR3_X1 U16100 ( .A1(n11941), .A2(n3861), .A3(n11940), .ZN(n11942) );
  NAND4_X1 U16101 ( .A1(n11944), .A2(n3792), .A3(n11943), .A4(n11942), .ZN(
        n11950) );
  AOI22_X1 U16102 ( .A1(n29419), .A2(\xmem_data[40][2] ), .B1(n27723), .B2(
        \xmem_data[41][2] ), .ZN(n11948) );
  AOI22_X1 U16103 ( .A1(n27814), .A2(\xmem_data[42][2] ), .B1(n3149), .B2(
        \xmem_data[43][2] ), .ZN(n11947) );
  AOI22_X1 U16104 ( .A1(n27710), .A2(\xmem_data[44][2] ), .B1(n30775), .B2(
        \xmem_data[45][2] ), .ZN(n11946) );
  AOI22_X1 U16105 ( .A1(n29790), .A2(\xmem_data[46][2] ), .B1(n27708), .B2(
        \xmem_data[47][2] ), .ZN(n11945) );
  NAND4_X1 U16106 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11949) );
  OAI21_X1 U16107 ( .B1(n11950), .B2(n11949), .A(n27737), .ZN(n11951) );
  XNOR2_X1 U16108 ( .A(n3260), .B(\fmem_data[27][7] ), .ZN(n30831) );
  XOR2_X1 U16109 ( .A(\fmem_data[27][6] ), .B(\fmem_data[27][7] ), .Z(n11955)
         );
  OAI22_X1 U16110 ( .A1(n31937), .A2(n35642), .B1(n30831), .B2(n35641), .ZN(
        n20289) );
  AOI22_X1 U16111 ( .A1(n27710), .A2(\xmem_data[48][5] ), .B1(n28766), .B2(
        \xmem_data[49][5] ), .ZN(n11958) );
  AOI22_X1 U16112 ( .A1(n28139), .A2(\xmem_data[52][5] ), .B1(n30776), .B2(
        \xmem_data[53][5] ), .ZN(n11957) );
  AOI22_X1 U16113 ( .A1(n28140), .A2(\xmem_data[54][5] ), .B1(n27905), .B2(
        \xmem_data[55][5] ), .ZN(n11956) );
  NAND4_X1 U16114 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11975) );
  AOI22_X1 U16115 ( .A1(n30764), .A2(\xmem_data[34][5] ), .B1(n28147), .B2(
        \xmem_data[35][5] ), .ZN(n11963) );
  AOI22_X1 U16116 ( .A1(n3162), .A2(\xmem_data[32][5] ), .B1(n3187), .B2(
        \xmem_data[33][5] ), .ZN(n11962) );
  AOI22_X1 U16117 ( .A1(n30766), .A2(\xmem_data[36][5] ), .B1(n30765), .B2(
        \xmem_data[37][5] ), .ZN(n11961) );
  AOI22_X1 U16118 ( .A1(n28151), .A2(\xmem_data[38][5] ), .B1(n24522), .B2(
        \xmem_data[39][5] ), .ZN(n11960) );
  NAND4_X1 U16119 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11974) );
  AOI22_X1 U16120 ( .A1(n27703), .A2(\xmem_data[56][5] ), .B1(n28738), .B2(
        \xmem_data[57][5] ), .ZN(n11967) );
  AOI22_X1 U16121 ( .A1(n28153), .A2(\xmem_data[58][5] ), .B1(n28152), .B2(
        \xmem_data[59][5] ), .ZN(n11966) );
  AOI22_X1 U16122 ( .A1(n29395), .A2(\xmem_data[60][5] ), .B1(n26884), .B2(
        \xmem_data[61][5] ), .ZN(n11965) );
  AOI22_X1 U16123 ( .A1(n28155), .A2(\xmem_data[62][5] ), .B1(n28154), .B2(
        \xmem_data[63][5] ), .ZN(n11964) );
  NAND4_X1 U16124 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11973) );
  AOI22_X1 U16125 ( .A1(n28160), .A2(\xmem_data[40][5] ), .B1(n28159), .B2(
        \xmem_data[41][5] ), .ZN(n11971) );
  AOI22_X1 U16126 ( .A1(n28161), .A2(\xmem_data[42][5] ), .B1(n31308), .B2(
        \xmem_data[43][5] ), .ZN(n11970) );
  AOI22_X1 U16127 ( .A1(n28163), .A2(\xmem_data[44][5] ), .B1(n28162), .B2(
        \xmem_data[45][5] ), .ZN(n11969) );
  AOI22_X1 U16128 ( .A1(n28165), .A2(\xmem_data[46][5] ), .B1(n28164), .B2(
        \xmem_data[47][5] ), .ZN(n11968) );
  NAND4_X1 U16129 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11972) );
  OR4_X1 U16130 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n11999) );
  AOI22_X1 U16131 ( .A1(n29647), .A2(\xmem_data[24][5] ), .B1(n30662), .B2(
        \xmem_data[25][5] ), .ZN(n11986) );
  AOI22_X1 U16132 ( .A1(n27754), .A2(\xmem_data[28][5] ), .B1(n29768), .B2(
        \xmem_data[29][5] ), .ZN(n11985) );
  AOI22_X1 U16133 ( .A1(n28191), .A2(\xmem_data[8][5] ), .B1(n28190), .B2(
        \xmem_data[9][5] ), .ZN(n11979) );
  AOI22_X1 U16134 ( .A1(n28193), .A2(\xmem_data[10][5] ), .B1(n28192), .B2(
        \xmem_data[11][5] ), .ZN(n11978) );
  AOI22_X1 U16135 ( .A1(n28195), .A2(\xmem_data[12][5] ), .B1(n28194), .B2(
        \xmem_data[13][5] ), .ZN(n11977) );
  AOI22_X1 U16136 ( .A1(n28196), .A2(\xmem_data[14][5] ), .B1(n28245), .B2(
        \xmem_data[15][5] ), .ZN(n11976) );
  NAND4_X1 U16137 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11983) );
  AOI22_X1 U16138 ( .A1(n3240), .A2(\xmem_data[30][5] ), .B1(n30746), .B2(
        \xmem_data[31][5] ), .ZN(n11981) );
  AOI22_X1 U16139 ( .A1(n3241), .A2(\xmem_data[26][5] ), .B1(n28152), .B2(
        \xmem_data[27][5] ), .ZN(n11980) );
  NAND3_X1 U16140 ( .A1(n11986), .A2(n11985), .A3(n11984), .ZN(n11997) );
  AOI22_X1 U16141 ( .A1(n29421), .A2(\xmem_data[16][5] ), .B1(n29753), .B2(
        \xmem_data[17][5] ), .ZN(n11990) );
  AOI22_X1 U16142 ( .A1(n28700), .A2(\xmem_data[18][5] ), .B1(n30292), .B2(
        \xmem_data[19][5] ), .ZN(n11989) );
  AOI22_X1 U16143 ( .A1(n28209), .A2(\xmem_data[20][5] ), .B1(n30776), .B2(
        \xmem_data[21][5] ), .ZN(n11988) );
  AOI22_X1 U16144 ( .A1(n28210), .A2(\xmem_data[22][5] ), .B1(n30698), .B2(
        \xmem_data[23][5] ), .ZN(n11987) );
  NAND4_X1 U16145 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11996) );
  AOI22_X1 U16146 ( .A1(n3164), .A2(\xmem_data[0][5] ), .B1(n3187), .B2(
        \xmem_data[1][5] ), .ZN(n11994) );
  AOI22_X1 U16147 ( .A1(n29610), .A2(\xmem_data[2][5] ), .B1(n28147), .B2(
        \xmem_data[3][5] ), .ZN(n11993) );
  AOI22_X1 U16148 ( .A1(n28680), .A2(\xmem_data[4][5] ), .B1(n30765), .B2(
        \xmem_data[5][5] ), .ZN(n11992) );
  AOI22_X1 U16149 ( .A1(n3233), .A2(\xmem_data[6][5] ), .B1(n28202), .B2(
        \xmem_data[7][5] ), .ZN(n11991) );
  NAND4_X1 U16150 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  AOI22_X1 U16151 ( .A1(n11999), .A2(n28177), .B1(n28215), .B2(n11998), .ZN(
        n12044) );
  AOI22_X1 U16152 ( .A1(n3166), .A2(\xmem_data[64][5] ), .B1(n3184), .B2(
        \xmem_data[65][5] ), .ZN(n12003) );
  AOI22_X1 U16153 ( .A1(n30070), .A2(\xmem_data[66][5] ), .B1(n28147), .B2(
        \xmem_data[67][5] ), .ZN(n12002) );
  AOI22_X1 U16154 ( .A1(n30717), .A2(\xmem_data[68][5] ), .B1(n30685), .B2(
        \xmem_data[69][5] ), .ZN(n12001) );
  AOI22_X1 U16155 ( .A1(n28151), .A2(\xmem_data[70][5] ), .B1(n28226), .B2(
        \xmem_data[71][5] ), .ZN(n12000) );
  NAND4_X1 U16156 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12019) );
  AOI22_X1 U16157 ( .A1(n28160), .A2(\xmem_data[72][5] ), .B1(n28159), .B2(
        \xmem_data[73][5] ), .ZN(n12007) );
  AOI22_X1 U16158 ( .A1(n28161), .A2(\xmem_data[74][5] ), .B1(n30674), .B2(
        \xmem_data[75][5] ), .ZN(n12006) );
  AOI22_X1 U16159 ( .A1(n28163), .A2(\xmem_data[76][5] ), .B1(n28162), .B2(
        \xmem_data[77][5] ), .ZN(n12005) );
  AOI22_X1 U16160 ( .A1(n28165), .A2(\xmem_data[78][5] ), .B1(n28164), .B2(
        \xmem_data[79][5] ), .ZN(n12004) );
  NAND4_X1 U16161 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12018) );
  AOI22_X1 U16162 ( .A1(n30215), .A2(\xmem_data[82][5] ), .B1(n28137), .B2(
        \xmem_data[83][5] ), .ZN(n12011) );
  AOI22_X1 U16163 ( .A1(n28136), .A2(\xmem_data[80][5] ), .B1(n26616), .B2(
        \xmem_data[81][5] ), .ZN(n12010) );
  AOI22_X1 U16164 ( .A1(n28139), .A2(\xmem_data[84][5] ), .B1(n29708), .B2(
        \xmem_data[85][5] ), .ZN(n12009) );
  AOI22_X1 U16165 ( .A1(n28140), .A2(\xmem_data[86][5] ), .B1(n29350), .B2(
        \xmem_data[87][5] ), .ZN(n12008) );
  NAND4_X1 U16166 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12017) );
  AOI22_X1 U16167 ( .A1(n30248), .A2(\xmem_data[88][5] ), .B1(n30662), .B2(
        \xmem_data[89][5] ), .ZN(n12015) );
  AOI22_X1 U16168 ( .A1(n28153), .A2(\xmem_data[90][5] ), .B1(n28152), .B2(
        \xmem_data[91][5] ), .ZN(n12014) );
  AOI22_X1 U16169 ( .A1(n29395), .A2(\xmem_data[92][5] ), .B1(n27728), .B2(
        \xmem_data[93][5] ), .ZN(n12013) );
  AOI22_X1 U16170 ( .A1(n28155), .A2(\xmem_data[94][5] ), .B1(n28154), .B2(
        \xmem_data[95][5] ), .ZN(n12012) );
  NAND4_X1 U16171 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  OR4_X1 U16172 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  AOI22_X1 U16173 ( .A1(n3167), .A2(\xmem_data[96][5] ), .B1(n3191), .B2(
        \xmem_data[97][5] ), .ZN(n12024) );
  AOI22_X1 U16174 ( .A1(n23901), .A2(\xmem_data[98][5] ), .B1(n28232), .B2(
        \xmem_data[99][5] ), .ZN(n12023) );
  AOI22_X1 U16175 ( .A1(n30766), .A2(\xmem_data[100][5] ), .B1(n29721), .B2(
        \xmem_data[101][5] ), .ZN(n12022) );
  AOI22_X1 U16176 ( .A1(n3233), .A2(\xmem_data[102][5] ), .B1(n28226), .B2(
        \xmem_data[103][5] ), .ZN(n12021) );
  NAND4_X1 U16177 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12040) );
  AOI22_X1 U16178 ( .A1(n28240), .A2(\xmem_data[104][5] ), .B1(n28239), .B2(
        \xmem_data[105][5] ), .ZN(n12028) );
  AOI22_X1 U16179 ( .A1(n28242), .A2(\xmem_data[106][5] ), .B1(n28241), .B2(
        \xmem_data[107][5] ), .ZN(n12027) );
  AOI22_X1 U16180 ( .A1(n28244), .A2(\xmem_data[108][5] ), .B1(n28243), .B2(
        \xmem_data[109][5] ), .ZN(n12026) );
  AOI22_X1 U16181 ( .A1(n28246), .A2(\xmem_data[110][5] ), .B1(n28245), .B2(
        \xmem_data[111][5] ), .ZN(n12025) );
  NAND4_X1 U16182 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12039) );
  AOI22_X1 U16183 ( .A1(n29628), .A2(\xmem_data[114][5] ), .B1(n28218), .B2(
        \xmem_data[115][5] ), .ZN(n12032) );
  AOI22_X1 U16184 ( .A1(n29433), .A2(\xmem_data[112][5] ), .B1(n29432), .B2(
        \xmem_data[113][5] ), .ZN(n12031) );
  AOI22_X1 U16185 ( .A1(n28219), .A2(\xmem_data[116][5] ), .B1(n29761), .B2(
        \xmem_data[117][5] ), .ZN(n12030) );
  AOI22_X1 U16186 ( .A1(n28220), .A2(\xmem_data[118][5] ), .B1(n30698), .B2(
        \xmem_data[119][5] ), .ZN(n12029) );
  NAND4_X1 U16187 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12038) );
  AOI22_X1 U16188 ( .A1(n30743), .A2(\xmem_data[120][5] ), .B1(n3368), .B2(
        \xmem_data[121][5] ), .ZN(n12036) );
  AOI22_X1 U16189 ( .A1(n3241), .A2(\xmem_data[122][5] ), .B1(n28233), .B2(
        \xmem_data[123][5] ), .ZN(n12035) );
  AOI22_X1 U16190 ( .A1(n28751), .A2(\xmem_data[124][5] ), .B1(n30634), .B2(
        \xmem_data[125][5] ), .ZN(n12034) );
  AOI22_X1 U16191 ( .A1(n3240), .A2(\xmem_data[126][5] ), .B1(n28231), .B2(
        \xmem_data[127][5] ), .ZN(n12033) );
  NAND4_X1 U16192 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12037) );
  OR4_X1 U16193 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12041) );
  NAND2_X1 U16194 ( .A1(n12041), .A2(n28133), .ZN(n12042) );
  XNOR2_X1 U16195 ( .A(n31386), .B(\fmem_data[31][5] ), .ZN(n31971) );
  AOI22_X1 U16196 ( .A1(n28700), .A2(\xmem_data[114][4] ), .B1(n28218), .B2(
        \xmem_data[115][4] ), .ZN(n12048) );
  AOI22_X1 U16197 ( .A1(n28219), .A2(\xmem_data[116][4] ), .B1(n3170), .B2(
        \xmem_data[117][4] ), .ZN(n12047) );
  AOI22_X1 U16198 ( .A1(n28734), .A2(\xmem_data[112][4] ), .B1(n30775), .B2(
        \xmem_data[113][4] ), .ZN(n12046) );
  AOI22_X1 U16199 ( .A1(n28220), .A2(\xmem_data[118][4] ), .B1(n16973), .B2(
        \xmem_data[119][4] ), .ZN(n12045) );
  AOI22_X1 U16200 ( .A1(n3163), .A2(\xmem_data[96][4] ), .B1(n3183), .B2(
        \xmem_data[97][4] ), .ZN(n12052) );
  AOI22_X1 U16201 ( .A1(n30310), .A2(\xmem_data[98][4] ), .B1(n28232), .B2(
        \xmem_data[99][4] ), .ZN(n12051) );
  AOI22_X1 U16202 ( .A1(n29722), .A2(\xmem_data[100][4] ), .B1(n30266), .B2(
        \xmem_data[101][4] ), .ZN(n12050) );
  AOI22_X1 U16203 ( .A1(n3233), .A2(\xmem_data[102][4] ), .B1(n28226), .B2(
        \xmem_data[103][4] ), .ZN(n12049) );
  AOI22_X1 U16204 ( .A1(n28240), .A2(\xmem_data[104][4] ), .B1(n28239), .B2(
        \xmem_data[105][4] ), .ZN(n12056) );
  AOI22_X1 U16205 ( .A1(n28242), .A2(\xmem_data[106][4] ), .B1(n28241), .B2(
        \xmem_data[107][4] ), .ZN(n12055) );
  AOI22_X1 U16206 ( .A1(n28244), .A2(\xmem_data[108][4] ), .B1(n28243), .B2(
        \xmem_data[109][4] ), .ZN(n12054) );
  AOI22_X1 U16207 ( .A1(n28246), .A2(\xmem_data[110][4] ), .B1(n28245), .B2(
        \xmem_data[111][4] ), .ZN(n12053) );
  AOI22_X1 U16208 ( .A1(n29481), .A2(\xmem_data[120][4] ), .B1(n28738), .B2(
        \xmem_data[121][4] ), .ZN(n12060) );
  AOI22_X1 U16209 ( .A1(n3241), .A2(\xmem_data[122][4] ), .B1(n28233), .B2(
        \xmem_data[123][4] ), .ZN(n12059) );
  AOI22_X1 U16210 ( .A1(n29604), .A2(\xmem_data[124][4] ), .B1(n30249), .B2(
        \xmem_data[125][4] ), .ZN(n12058) );
  AOI22_X1 U16211 ( .A1(n3240), .A2(\xmem_data[126][4] ), .B1(n28231), .B2(
        \xmem_data[127][4] ), .ZN(n12057) );
  AOI22_X1 U16212 ( .A1(n3165), .A2(\xmem_data[64][4] ), .B1(n3187), .B2(
        \xmem_data[65][4] ), .ZN(n12064) );
  AOI22_X1 U16213 ( .A1(n30715), .A2(\xmem_data[66][4] ), .B1(n28147), .B2(
        \xmem_data[67][4] ), .ZN(n12063) );
  AOI22_X1 U16214 ( .A1(n30063), .A2(\xmem_data[68][4] ), .B1(n30644), .B2(
        \xmem_data[69][4] ), .ZN(n12062) );
  AOI22_X1 U16215 ( .A1(n28151), .A2(\xmem_data[70][4] ), .B1(n3271), .B2(
        \xmem_data[71][4] ), .ZN(n12061) );
  NAND4_X1 U16216 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12081) );
  AOI22_X1 U16217 ( .A1(n28160), .A2(\xmem_data[72][4] ), .B1(n28159), .B2(
        \xmem_data[73][4] ), .ZN(n12068) );
  AOI22_X1 U16218 ( .A1(n28161), .A2(\xmem_data[74][4] ), .B1(n29657), .B2(
        \xmem_data[75][4] ), .ZN(n12067) );
  AOI22_X1 U16219 ( .A1(n28163), .A2(\xmem_data[76][4] ), .B1(n28162), .B2(
        \xmem_data[77][4] ), .ZN(n12066) );
  AOI22_X1 U16220 ( .A1(n28165), .A2(\xmem_data[78][4] ), .B1(n28164), .B2(
        \xmem_data[79][4] ), .ZN(n12065) );
  NAND4_X1 U16221 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12080) );
  AOI22_X1 U16222 ( .A1(n28139), .A2(\xmem_data[84][4] ), .B1(n28208), .B2(
        \xmem_data[85][4] ), .ZN(n12073) );
  AOI22_X1 U16223 ( .A1(n28136), .A2(\xmem_data[80][4] ), .B1(n28206), .B2(
        \xmem_data[81][4] ), .ZN(n12072) );
  AND2_X1 U16224 ( .A1(n28137), .A2(\xmem_data[83][4] ), .ZN(n12069) );
  AOI21_X1 U16225 ( .B1(n30215), .B2(\xmem_data[82][4] ), .A(n12069), .ZN(
        n12071) );
  AOI22_X1 U16226 ( .A1(n28140), .A2(\xmem_data[86][4] ), .B1(n29231), .B2(
        \xmem_data[87][4] ), .ZN(n12070) );
  NAND4_X1 U16227 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12079) );
  AOI22_X1 U16228 ( .A1(n30248), .A2(\xmem_data[88][4] ), .B1(n3368), .B2(
        \xmem_data[89][4] ), .ZN(n12077) );
  AOI22_X1 U16229 ( .A1(n28153), .A2(\xmem_data[90][4] ), .B1(n28152), .B2(
        \xmem_data[91][4] ), .ZN(n12076) );
  AOI22_X1 U16230 ( .A1(n3173), .A2(\xmem_data[92][4] ), .B1(n28778), .B2(
        \xmem_data[93][4] ), .ZN(n12075) );
  AOI22_X1 U16231 ( .A1(n28155), .A2(\xmem_data[94][4] ), .B1(n28154), .B2(
        \xmem_data[95][4] ), .ZN(n12074) );
  NAND4_X1 U16232 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12078) );
  AOI22_X1 U16233 ( .A1(n12083), .A2(n28133), .B1(n12082), .B2(n28258), .ZN(
        n12127) );
  AOI22_X1 U16234 ( .A1(n3166), .A2(\xmem_data[32][4] ), .B1(n3185), .B2(
        \xmem_data[33][4] ), .ZN(n12087) );
  AOI22_X1 U16235 ( .A1(n30715), .A2(\xmem_data[34][4] ), .B1(n28147), .B2(
        \xmem_data[35][4] ), .ZN(n12086) );
  AOI22_X1 U16236 ( .A1(n29547), .A2(\xmem_data[36][4] ), .B1(n30170), .B2(
        \xmem_data[37][4] ), .ZN(n12085) );
  AOI22_X1 U16237 ( .A1(n28151), .A2(\xmem_data[38][4] ), .B1(n29297), .B2(
        \xmem_data[39][4] ), .ZN(n12084) );
  NAND4_X1 U16238 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12103) );
  AOI22_X1 U16239 ( .A1(n28160), .A2(\xmem_data[40][4] ), .B1(n28159), .B2(
        \xmem_data[41][4] ), .ZN(n12091) );
  AOI22_X1 U16240 ( .A1(n28161), .A2(\xmem_data[42][4] ), .B1(n29298), .B2(
        \xmem_data[43][4] ), .ZN(n12090) );
  AOI22_X1 U16241 ( .A1(n28163), .A2(\xmem_data[44][4] ), .B1(n28162), .B2(
        \xmem_data[45][4] ), .ZN(n12089) );
  AOI22_X1 U16242 ( .A1(n28165), .A2(\xmem_data[46][4] ), .B1(n28164), .B2(
        \xmem_data[47][4] ), .ZN(n12088) );
  NAND4_X1 U16243 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12102) );
  AOI22_X1 U16244 ( .A1(n29423), .A2(\xmem_data[50][4] ), .B1(n28137), .B2(
        \xmem_data[51][4] ), .ZN(n12095) );
  AOI22_X1 U16245 ( .A1(n29788), .A2(\xmem_data[48][4] ), .B1(n28206), .B2(
        \xmem_data[49][4] ), .ZN(n12094) );
  AOI22_X1 U16246 ( .A1(n28139), .A2(\xmem_data[52][4] ), .B1(n30696), .B2(
        \xmem_data[53][4] ), .ZN(n12093) );
  AOI22_X1 U16247 ( .A1(n28140), .A2(\xmem_data[54][4] ), .B1(n25417), .B2(
        \xmem_data[55][4] ), .ZN(n12092) );
  NAND4_X1 U16248 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(
        n12101) );
  AOI22_X1 U16249 ( .A1(n29801), .A2(\xmem_data[56][4] ), .B1(n30662), .B2(
        \xmem_data[57][4] ), .ZN(n12099) );
  AOI22_X1 U16250 ( .A1(n28153), .A2(\xmem_data[58][4] ), .B1(n28152), .B2(
        \xmem_data[59][4] ), .ZN(n12098) );
  AOI22_X1 U16251 ( .A1(n29714), .A2(\xmem_data[60][4] ), .B1(n27728), .B2(
        \xmem_data[61][4] ), .ZN(n12097) );
  AOI22_X1 U16252 ( .A1(n28155), .A2(\xmem_data[62][4] ), .B1(n28154), .B2(
        \xmem_data[63][4] ), .ZN(n12096) );
  NAND4_X1 U16253 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n12100) );
  OR4_X2 U16254 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(
        n12125) );
  AOI22_X1 U16255 ( .A1(n28136), .A2(\xmem_data[16][4] ), .B1(n28766), .B2(
        \xmem_data[17][4] ), .ZN(n12107) );
  AOI22_X1 U16256 ( .A1(n29699), .A2(\xmem_data[18][4] ), .B1(n29832), .B2(
        \xmem_data[19][4] ), .ZN(n12106) );
  AOI22_X1 U16257 ( .A1(n28209), .A2(\xmem_data[20][4] ), .B1(n28786), .B2(
        \xmem_data[21][4] ), .ZN(n12105) );
  AOI22_X1 U16258 ( .A1(n28210), .A2(\xmem_data[22][4] ), .B1(n3375), .B2(
        \xmem_data[23][4] ), .ZN(n12104) );
  NAND4_X1 U16259 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12123) );
  AOI22_X1 U16260 ( .A1(n3165), .A2(\xmem_data[0][4] ), .B1(n3182), .B2(
        \xmem_data[1][4] ), .ZN(n12111) );
  AOI22_X1 U16261 ( .A1(n29810), .A2(\xmem_data[2][4] ), .B1(n29639), .B2(
        \xmem_data[3][4] ), .ZN(n12110) );
  AOI22_X1 U16262 ( .A1(n29722), .A2(\xmem_data[4][4] ), .B1(n30685), .B2(
        \xmem_data[5][4] ), .ZN(n12109) );
  AOI22_X1 U16263 ( .A1(n3233), .A2(\xmem_data[6][4] ), .B1(n28202), .B2(
        \xmem_data[7][4] ), .ZN(n12108) );
  NAND4_X1 U16264 ( .A1(n12111), .A2(n12110), .A3(n12109), .A4(n12108), .ZN(
        n12122) );
  AOI22_X1 U16265 ( .A1(n29481), .A2(\xmem_data[24][4] ), .B1(n3369), .B2(
        \xmem_data[25][4] ), .ZN(n12115) );
  AOI22_X1 U16266 ( .A1(n3241), .A2(\xmem_data[26][4] ), .B1(n20545), .B2(
        \xmem_data[27][4] ), .ZN(n12114) );
  AOI22_X1 U16267 ( .A1(n29714), .A2(\xmem_data[28][4] ), .B1(n30249), .B2(
        \xmem_data[29][4] ), .ZN(n12113) );
  AOI22_X1 U16268 ( .A1(n3240), .A2(\xmem_data[30][4] ), .B1(n28516), .B2(
        \xmem_data[31][4] ), .ZN(n12112) );
  NAND4_X1 U16269 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12121) );
  AOI22_X1 U16270 ( .A1(n28191), .A2(\xmem_data[8][4] ), .B1(n28190), .B2(
        \xmem_data[9][4] ), .ZN(n12119) );
  AOI22_X1 U16271 ( .A1(n28193), .A2(\xmem_data[10][4] ), .B1(n28192), .B2(
        \xmem_data[11][4] ), .ZN(n12118) );
  AOI22_X1 U16272 ( .A1(n28195), .A2(\xmem_data[12][4] ), .B1(n28194), .B2(
        \xmem_data[13][4] ), .ZN(n12117) );
  AOI22_X1 U16273 ( .A1(n28196), .A2(\xmem_data[14][4] ), .B1(n28718), .B2(
        \xmem_data[15][4] ), .ZN(n12116) );
  NAND4_X1 U16274 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12120) );
  NAND2_X1 U16275 ( .A1(n12127), .A2(n12126), .ZN(n32110) );
  XNOR2_X1 U16276 ( .A(n32110), .B(\fmem_data[31][5] ), .ZN(n28938) );
  XOR2_X1 U16277 ( .A(\fmem_data[31][4] ), .B(\fmem_data[31][5] ), .Z(n12128)
         );
  OAI22_X1 U16278 ( .A1(n31971), .A2(n34944), .B1(n28938), .B2(n34945), .ZN(
        n34226) );
  AOI22_X1 U16279 ( .A1(n29446), .A2(\xmem_data[100][7] ), .B1(n30190), .B2(
        \xmem_data[101][7] ), .ZN(n12135) );
  AOI22_X1 U16280 ( .A1(n28740), .A2(\xmem_data[96][7] ), .B1(n30293), .B2(
        \xmem_data[97][7] ), .ZN(n12134) );
  AOI22_X1 U16281 ( .A1(n3244), .A2(\xmem_data[98][7] ), .B1(n3126), .B2(
        \xmem_data[99][7] ), .ZN(n12129) );
  AOI22_X1 U16282 ( .A1(n28744), .A2(\xmem_data[102][7] ), .B1(n28743), .B2(
        \xmem_data[103][7] ), .ZN(n12130) );
  NAND3_X1 U16283 ( .A1(n12135), .A2(n12134), .A3(n12133), .ZN(n12141) );
  AOI22_X1 U16284 ( .A1(n28685), .A2(\xmem_data[104][7] ), .B1(n27753), .B2(
        \xmem_data[105][7] ), .ZN(n12139) );
  AOI22_X1 U16285 ( .A1(n28753), .A2(\xmem_data[106][7] ), .B1(n28053), .B2(
        \xmem_data[107][7] ), .ZN(n12138) );
  AOI22_X1 U16286 ( .A1(n3164), .A2(\xmem_data[108][7] ), .B1(n3183), .B2(
        \xmem_data[109][7] ), .ZN(n12137) );
  AOI22_X1 U16287 ( .A1(n28689), .A2(\xmem_data[110][7] ), .B1(n28781), .B2(
        \xmem_data[111][7] ), .ZN(n12136) );
  NAND4_X1 U16288 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  OR2_X1 U16289 ( .A1(n12141), .A2(n12140), .ZN(n12157) );
  AOI22_X1 U16290 ( .A1(n29815), .A2(\xmem_data[112][7] ), .B1(n30716), .B2(
        \xmem_data[113][7] ), .ZN(n12145) );
  AOI22_X1 U16291 ( .A1(n28720), .A2(\xmem_data[114][7] ), .B1(n3151), .B2(
        \xmem_data[115][7] ), .ZN(n12144) );
  AOI22_X1 U16292 ( .A1(n28725), .A2(\xmem_data[116][7] ), .B1(n28724), .B2(
        \xmem_data[117][7] ), .ZN(n12143) );
  AOI22_X1 U16293 ( .A1(n28727), .A2(\xmem_data[118][7] ), .B1(n29327), .B2(
        \xmem_data[119][7] ), .ZN(n12142) );
  AOI22_X1 U16294 ( .A1(n28765), .A2(\xmem_data[120][7] ), .B1(n3124), .B2(
        \xmem_data[121][7] ), .ZN(n12146) );
  INV_X1 U16295 ( .A(n12146), .ZN(n12147) );
  AOI21_X1 U16296 ( .B1(n30215), .B2(\xmem_data[126][7] ), .A(n12147), .ZN(
        n12155) );
  AOI22_X1 U16297 ( .A1(n28719), .A2(\xmem_data[122][7] ), .B1(n28718), .B2(
        \xmem_data[123][7] ), .ZN(n12148) );
  INV_X1 U16298 ( .A(n12148), .ZN(n12152) );
  NAND2_X1 U16299 ( .A1(n30106), .A2(\xmem_data[125][7] ), .ZN(n12150) );
  NAND2_X1 U16300 ( .A1(n28733), .A2(\xmem_data[127][7] ), .ZN(n12149) );
  NAND2_X1 U16301 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND3_X1 U16302 ( .A1(n3822), .A2(n12155), .A3(n12154), .ZN(n12156) );
  OAI21_X1 U16303 ( .B1(n12157), .B2(n12156), .A(n28762), .ZN(n12230) );
  AOI22_X1 U16304 ( .A1(n29436), .A2(\xmem_data[8][7] ), .B1(n30084), .B2(
        \xmem_data[9][7] ), .ZN(n12161) );
  AOI22_X1 U16305 ( .A1(n28686), .A2(\xmem_data[10][7] ), .B1(n3466), .B2(
        \xmem_data[11][7] ), .ZN(n12160) );
  AOI22_X1 U16306 ( .A1(n3166), .A2(\xmem_data[12][7] ), .B1(n3185), .B2(
        \xmem_data[13][7] ), .ZN(n12159) );
  AOI22_X1 U16307 ( .A1(n29810), .A2(\xmem_data[14][7] ), .B1(n28687), .B2(
        \xmem_data[15][7] ), .ZN(n12158) );
  AOI22_X1 U16308 ( .A1(n28787), .A2(\xmem_data[0][7] ), .B1(n30696), .B2(
        \xmem_data[1][7] ), .ZN(n12165) );
  AOI22_X1 U16309 ( .A1(n3244), .A2(\xmem_data[2][7] ), .B1(n30698), .B2(
        \xmem_data[3][7] ), .ZN(n12164) );
  AOI22_X1 U16310 ( .A1(n29446), .A2(\xmem_data[4][7] ), .B1(n28665), .B2(
        \xmem_data[5][7] ), .ZN(n12163) );
  AOI22_X1 U16311 ( .A1(n28788), .A2(\xmem_data[6][7] ), .B1(n20799), .B2(
        \xmem_data[7][7] ), .ZN(n12162) );
  AOI22_X1 U16312 ( .A1(n30198), .A2(\xmem_data[16][7] ), .B1(n30644), .B2(
        \xmem_data[17][7] ), .ZN(n12169) );
  AOI22_X1 U16313 ( .A1(n28702), .A2(\xmem_data[18][7] ), .B1(n29379), .B2(
        \xmem_data[19][7] ), .ZN(n12168) );
  AOI22_X1 U16314 ( .A1(n27716), .A2(\xmem_data[20][7] ), .B1(n28724), .B2(
        \xmem_data[21][7] ), .ZN(n12167) );
  AOI22_X1 U16315 ( .A1(n29489), .A2(\xmem_data[22][7] ), .B1(n28772), .B2(
        \xmem_data[23][7] ), .ZN(n12166) );
  AOI22_X1 U16316 ( .A1(n30291), .A2(\xmem_data[28][7] ), .B1(n29432), .B2(
        \xmem_data[29][7] ), .ZN(n12170) );
  INV_X1 U16317 ( .A(n12170), .ZN(n12176) );
  AOI22_X1 U16318 ( .A1(n30279), .A2(\xmem_data[30][7] ), .B1(n28218), .B2(
        \xmem_data[31][7] ), .ZN(n12171) );
  INV_X1 U16319 ( .A(n12171), .ZN(n12175) );
  AOI22_X1 U16320 ( .A1(n29786), .A2(\xmem_data[24][7] ), .B1(n27743), .B2(
        \xmem_data[25][7] ), .ZN(n12173) );
  AOI22_X1 U16321 ( .A1(n3227), .A2(\xmem_data[26][7] ), .B1(n3142), .B2(
        \xmem_data[27][7] ), .ZN(n12172) );
  NAND2_X1 U16322 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NOR3_X1 U16323 ( .A1(n12176), .A2(n12175), .A3(n12174), .ZN(n12177) );
  NAND4_X1 U16324 ( .A1(n3850), .A2(n3540), .A3(n3474), .A4(n12177), .ZN(
        n12178) );
  NAND2_X1 U16325 ( .A1(n12178), .A2(n28794), .ZN(n12229) );
  AOI22_X1 U16326 ( .A1(n28207), .A2(\xmem_data[94][7] ), .B1(n28218), .B2(
        \xmem_data[95][7] ), .ZN(n12181) );
  AOI22_X1 U16327 ( .A1(n3163), .A2(\xmem_data[76][7] ), .B1(n3189), .B2(
        \xmem_data[77][7] ), .ZN(n12180) );
  AOI22_X1 U16328 ( .A1(n28686), .A2(\xmem_data[74][7] ), .B1(n27945), .B2(
        \xmem_data[75][7] ), .ZN(n12179) );
  AOI22_X1 U16329 ( .A1(n29363), .A2(\xmem_data[80][7] ), .B1(n30716), .B2(
        \xmem_data[81][7] ), .ZN(n12185) );
  AOI22_X1 U16330 ( .A1(n28702), .A2(\xmem_data[82][7] ), .B1(n28701), .B2(
        \xmem_data[83][7] ), .ZN(n12184) );
  AOI22_X1 U16331 ( .A1(n28725), .A2(\xmem_data[84][7] ), .B1(n28696), .B2(
        \xmem_data[85][7] ), .ZN(n12183) );
  AOI22_X1 U16332 ( .A1(n28681), .A2(\xmem_data[86][7] ), .B1(n25407), .B2(
        \xmem_data[87][7] ), .ZN(n12182) );
  NAND4_X1 U16333 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  OR2_X1 U16334 ( .A1(n12187), .A2(n12186), .ZN(n12202) );
  AOI22_X1 U16335 ( .A1(n29788), .A2(\xmem_data[92][7] ), .B1(n30182), .B2(
        \xmem_data[93][7] ), .ZN(n12188) );
  INV_X1 U16336 ( .A(n12188), .ZN(n12196) );
  AOI22_X1 U16337 ( .A1(n3173), .A2(\xmem_data[72][7] ), .B1(n30090), .B2(
        \xmem_data[73][7] ), .ZN(n12189) );
  INV_X1 U16338 ( .A(n12189), .ZN(n12195) );
  AOI22_X1 U16339 ( .A1(n28670), .A2(\xmem_data[66][7] ), .B1(n27905), .B2(
        \xmem_data[67][7] ), .ZN(n12193) );
  AOI22_X1 U16340 ( .A1(n29419), .A2(\xmem_data[88][7] ), .B1(n29418), .B2(
        \xmem_data[89][7] ), .ZN(n12192) );
  AOI22_X1 U16341 ( .A1(n3227), .A2(\xmem_data[90][7] ), .B1(n28677), .B2(
        \xmem_data[91][7] ), .ZN(n12191) );
  AOI22_X1 U16342 ( .A1(n28744), .A2(\xmem_data[70][7] ), .B1(n28671), .B2(
        \xmem_data[71][7] ), .ZN(n12190) );
  NAND4_X1 U16343 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12194) );
  NOR3_X1 U16344 ( .A1(n12196), .A2(n12195), .A3(n12194), .ZN(n12200) );
  AOI22_X1 U16345 ( .A1(n30633), .A2(\xmem_data[68][7] ), .B1(n28738), .B2(
        \xmem_data[69][7] ), .ZN(n12199) );
  AOI22_X1 U16346 ( .A1(n30280), .A2(\xmem_data[64][7] ), .B1(n30696), .B2(
        \xmem_data[65][7] ), .ZN(n12198) );
  AOI22_X1 U16347 ( .A1(n29716), .A2(\xmem_data[78][7] ), .B1(n28754), .B2(
        \xmem_data[79][7] ), .ZN(n12197) );
  NAND4_X1 U16348 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  OAI21_X1 U16349 ( .B1(n12202), .B2(n12201), .A(n28662), .ZN(n12228) );
  AOI22_X1 U16350 ( .A1(n29790), .A2(\xmem_data[62][7] ), .B1(n30292), .B2(
        \xmem_data[63][7] ), .ZN(n12209) );
  AOI22_X1 U16351 ( .A1(n28734), .A2(\xmem_data[60][7] ), .B1(n29831), .B2(
        \xmem_data[61][7] ), .ZN(n12208) );
  AOI22_X1 U16352 ( .A1(n29447), .A2(\xmem_data[56][7] ), .B1(n3124), .B2(
        \xmem_data[57][7] ), .ZN(n12203) );
  INV_X1 U16353 ( .A(n12203), .ZN(n12206) );
  AOI22_X1 U16354 ( .A1(n3227), .A2(\xmem_data[58][7] ), .B1(n28677), .B2(
        \xmem_data[59][7] ), .ZN(n12204) );
  INV_X1 U16355 ( .A(n12204), .ZN(n12205) );
  NOR2_X1 U16356 ( .A1(n12206), .A2(n12205), .ZN(n12207) );
  AOI22_X1 U16357 ( .A1(n29395), .A2(\xmem_data[40][7] ), .B1(n26884), .B2(
        \xmem_data[41][7] ), .ZN(n12213) );
  AOI22_X1 U16358 ( .A1(n28686), .A2(\xmem_data[42][7] ), .B1(n28091), .B2(
        \xmem_data[43][7] ), .ZN(n12212) );
  AOI22_X1 U16359 ( .A1(n3162), .A2(\xmem_data[44][7] ), .B1(n3186), .B2(
        \xmem_data[45][7] ), .ZN(n12211) );
  AOI22_X1 U16360 ( .A1(n30715), .A2(\xmem_data[46][7] ), .B1(n28754), .B2(
        \xmem_data[47][7] ), .ZN(n12210) );
  NAND4_X1 U16361 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12219) );
  AOI22_X1 U16362 ( .A1(n30766), .A2(\xmem_data[48][7] ), .B1(n29487), .B2(
        \xmem_data[49][7] ), .ZN(n12217) );
  AOI22_X1 U16363 ( .A1(n28702), .A2(\xmem_data[50][7] ), .B1(n28701), .B2(
        \xmem_data[51][7] ), .ZN(n12216) );
  AOI22_X1 U16364 ( .A1(n28725), .A2(\xmem_data[52][7] ), .B1(n28696), .B2(
        \xmem_data[53][7] ), .ZN(n12215) );
  AOI22_X1 U16365 ( .A1(n28681), .A2(\xmem_data[54][7] ), .B1(n28772), .B2(
        \xmem_data[55][7] ), .ZN(n12214) );
  NAND4_X1 U16366 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12218) );
  OR3_X1 U16367 ( .A1(n12220), .A2(n12219), .A3(n12218), .ZN(n12226) );
  AOI22_X1 U16368 ( .A1(n28787), .A2(\xmem_data[32][7] ), .B1(n30293), .B2(
        \xmem_data[33][7] ), .ZN(n12224) );
  AOI22_X1 U16369 ( .A1(n28670), .A2(\xmem_data[34][7] ), .B1(n3146), .B2(
        \xmem_data[35][7] ), .ZN(n12223) );
  AOI22_X1 U16370 ( .A1(n30633), .A2(\xmem_data[36][7] ), .B1(n29482), .B2(
        \xmem_data[37][7] ), .ZN(n12222) );
  AOI22_X1 U16371 ( .A1(n28788), .A2(\xmem_data[38][7] ), .B1(n28671), .B2(
        \xmem_data[39][7] ), .ZN(n12221) );
  NAND4_X1 U16372 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12225) );
  OAI21_X1 U16373 ( .B1(n12226), .B2(n12225), .A(n28713), .ZN(n12227) );
  XNOR2_X1 U16374 ( .A(n35238), .B(\fmem_data[11][3] ), .ZN(n30353) );
  AOI22_X1 U16375 ( .A1(n29769), .A2(\xmem_data[40][6] ), .B1(n26884), .B2(
        \xmem_data[41][6] ), .ZN(n12234) );
  AOI22_X1 U16376 ( .A1(n28686), .A2(\xmem_data[42][6] ), .B1(n23795), .B2(
        \xmem_data[43][6] ), .ZN(n12233) );
  AOI22_X1 U16377 ( .A1(n3162), .A2(\xmem_data[44][6] ), .B1(n3180), .B2(
        \xmem_data[45][6] ), .ZN(n12232) );
  AOI22_X1 U16378 ( .A1(n26812), .A2(\xmem_data[46][6] ), .B1(n28687), .B2(
        \xmem_data[47][6] ), .ZN(n12231) );
  AOI22_X1 U16379 ( .A1(n29433), .A2(\xmem_data[60][6] ), .B1(n30775), .B2(
        \xmem_data[61][6] ), .ZN(n12235) );
  INV_X1 U16380 ( .A(n12235), .ZN(n12242) );
  AOI22_X1 U16381 ( .A1(n28670), .A2(\xmem_data[34][6] ), .B1(n3132), .B2(
        \xmem_data[35][6] ), .ZN(n12239) );
  AOI22_X1 U16382 ( .A1(n29419), .A2(\xmem_data[56][6] ), .B1(n27743), .B2(
        \xmem_data[57][6] ), .ZN(n12238) );
  AOI22_X1 U16383 ( .A1(n3227), .A2(\xmem_data[58][6] ), .B1(n28677), .B2(
        \xmem_data[59][6] ), .ZN(n12237) );
  AOI22_X1 U16384 ( .A1(n28744), .A2(\xmem_data[38][6] ), .B1(n28671), .B2(
        \xmem_data[39][6] ), .ZN(n12236) );
  NAND2_X1 U16385 ( .A1(n3776), .A2(n12240), .ZN(n12241) );
  NOR2_X1 U16386 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  NAND2_X1 U16387 ( .A1(n3777), .A2(n12243), .ZN(n12251) );
  AOI22_X1 U16388 ( .A1(n30766), .A2(\xmem_data[48][6] ), .B1(n30765), .B2(
        \xmem_data[49][6] ), .ZN(n12247) );
  AOI22_X1 U16389 ( .A1(n28702), .A2(\xmem_data[50][6] ), .B1(n28701), .B2(
        \xmem_data[51][6] ), .ZN(n12246) );
  AOI22_X1 U16390 ( .A1(n28725), .A2(\xmem_data[52][6] ), .B1(n28696), .B2(
        \xmem_data[53][6] ), .ZN(n12245) );
  AOI22_X1 U16391 ( .A1(n28681), .A2(\xmem_data[54][6] ), .B1(n25628), .B2(
        \xmem_data[55][6] ), .ZN(n12244) );
  AOI22_X1 U16392 ( .A1(n29628), .A2(\xmem_data[62][6] ), .B1(n29832), .B2(
        \xmem_data[63][6] ), .ZN(n12249) );
  AOI22_X1 U16393 ( .A1(n27834), .A2(\xmem_data[32][6] ), .B1(n29708), .B2(
        \xmem_data[33][6] ), .ZN(n12248) );
  OAI21_X1 U16394 ( .B1(n12251), .B2(n12250), .A(n28713), .ZN(n12341) );
  AOI22_X1 U16395 ( .A1(n29628), .A2(\xmem_data[94][6] ), .B1(n29565), .B2(
        \xmem_data[95][6] ), .ZN(n12258) );
  AOI22_X1 U16396 ( .A1(n29433), .A2(\xmem_data[92][6] ), .B1(n30182), .B2(
        \xmem_data[93][6] ), .ZN(n12257) );
  AOI22_X1 U16397 ( .A1(n8088), .A2(\xmem_data[88][6] ), .B1(n3124), .B2(
        \xmem_data[89][6] ), .ZN(n12252) );
  INV_X1 U16398 ( .A(n12252), .ZN(n12255) );
  AOI22_X1 U16399 ( .A1(n3227), .A2(\xmem_data[90][6] ), .B1(n28677), .B2(
        \xmem_data[91][6] ), .ZN(n12253) );
  INV_X1 U16400 ( .A(n12253), .ZN(n12254) );
  NOR2_X1 U16401 ( .A1(n12255), .A2(n12254), .ZN(n12256) );
  AOI22_X1 U16402 ( .A1(n28685), .A2(\xmem_data[72][6] ), .B1(n30193), .B2(
        \xmem_data[73][6] ), .ZN(n12262) );
  AOI22_X1 U16403 ( .A1(n28686), .A2(\xmem_data[74][6] ), .B1(n25461), .B2(
        \xmem_data[75][6] ), .ZN(n12261) );
  AOI22_X1 U16404 ( .A1(n3163), .A2(\xmem_data[76][6] ), .B1(n3184), .B2(
        \xmem_data[77][6] ), .ZN(n12260) );
  AOI22_X1 U16405 ( .A1(n27031), .A2(\xmem_data[78][6] ), .B1(n28687), .B2(
        \xmem_data[79][6] ), .ZN(n12259) );
  NAND4_X1 U16406 ( .A1(n12259), .A2(n12261), .A3(n12260), .A4(n12262), .ZN(
        n12268) );
  AOI22_X1 U16407 ( .A1(n30766), .A2(\xmem_data[80][6] ), .B1(n29640), .B2(
        \xmem_data[81][6] ), .ZN(n12266) );
  AOI22_X1 U16408 ( .A1(n28702), .A2(\xmem_data[82][6] ), .B1(n28701), .B2(
        \xmem_data[83][6] ), .ZN(n12265) );
  AOI22_X1 U16409 ( .A1(n28725), .A2(\xmem_data[84][6] ), .B1(n28696), .B2(
        \xmem_data[85][6] ), .ZN(n12264) );
  AOI22_X1 U16410 ( .A1(n28681), .A2(\xmem_data[86][6] ), .B1(n20567), .B2(
        \xmem_data[87][6] ), .ZN(n12263) );
  NAND4_X1 U16411 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12267) );
  OR3_X1 U16412 ( .A1(n12269), .A2(n12268), .A3(n12267), .ZN(n12275) );
  AOI22_X1 U16413 ( .A1(n27701), .A2(\xmem_data[64][6] ), .B1(n29629), .B2(
        \xmem_data[65][6] ), .ZN(n12273) );
  AOI22_X1 U16414 ( .A1(n28670), .A2(n20682), .B1(n3282), .B2(
        \xmem_data[67][6] ), .ZN(n12272) );
  AOI22_X1 U16415 ( .A1(n3249), .A2(\xmem_data[68][6] ), .B1(n28238), .B2(
        \xmem_data[69][6] ), .ZN(n12271) );
  AOI22_X1 U16416 ( .A1(n28744), .A2(\xmem_data[70][6] ), .B1(n28671), .B2(
        \xmem_data[71][6] ), .ZN(n12270) );
  NAND4_X1 U16417 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  OAI21_X1 U16418 ( .B1(n12275), .B2(n12274), .A(n28662), .ZN(n12340) );
  AND2_X1 U16419 ( .A1(n28754), .A2(\xmem_data[111][6] ), .ZN(n12276) );
  AOI21_X1 U16420 ( .B1(n29716), .B2(\xmem_data[110][6] ), .A(n12276), .ZN(
        n12279) );
  AOI22_X1 U16421 ( .A1(n28753), .A2(\xmem_data[106][6] ), .B1(n29237), .B2(
        \xmem_data[107][6] ), .ZN(n12278) );
  AOI22_X1 U16422 ( .A1(n30076), .A2(\xmem_data[112][6] ), .B1(n30765), .B2(
        \xmem_data[113][6] ), .ZN(n12283) );
  AOI22_X1 U16423 ( .A1(n28720), .A2(\xmem_data[114][6] ), .B1(n25401), .B2(
        \xmem_data[115][6] ), .ZN(n12282) );
  AOI22_X1 U16424 ( .A1(n28725), .A2(\xmem_data[116][6] ), .B1(n28724), .B2(
        \xmem_data[117][6] ), .ZN(n12281) );
  AOI22_X1 U16425 ( .A1(n28727), .A2(\xmem_data[118][6] ), .B1(n14982), .B2(
        \xmem_data[119][6] ), .ZN(n12280) );
  NAND4_X1 U16426 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12284) );
  OR2_X1 U16427 ( .A1(n12285), .A2(n12284), .ZN(n12302) );
  AND2_X1 U16428 ( .A1(n28733), .A2(\xmem_data[127][6] ), .ZN(n12286) );
  AOI21_X1 U16429 ( .B1(n3392), .B2(\xmem_data[126][6] ), .A(n12286), .ZN(
        n12300) );
  NAND2_X1 U16430 ( .A1(n28734), .A2(\xmem_data[124][6] ), .ZN(n12288) );
  NAND2_X1 U16431 ( .A1(n30106), .A2(\xmem_data[125][6] ), .ZN(n12287) );
  NAND2_X1 U16432 ( .A1(n12288), .A2(n12287), .ZN(n12296) );
  AOI22_X1 U16433 ( .A1(n3163), .A2(\xmem_data[108][6] ), .B1(n3185), .B2(
        \xmem_data[109][6] ), .ZN(n12289) );
  INV_X1 U16434 ( .A(n12289), .ZN(n12295) );
  AOI22_X1 U16435 ( .A1(n3244), .A2(\xmem_data[98][6] ), .B1(n3126), .B2(
        \xmem_data[99][6] ), .ZN(n12293) );
  AOI22_X1 U16436 ( .A1(n29829), .A2(\xmem_data[120][6] ), .B1(n3124), .B2(
        \xmem_data[121][6] ), .ZN(n12292) );
  AOI22_X1 U16437 ( .A1(n28719), .A2(\xmem_data[122][6] ), .B1(n28718), .B2(
        \xmem_data[123][6] ), .ZN(n12291) );
  AOI22_X1 U16438 ( .A1(n28744), .A2(\xmem_data[102][6] ), .B1(n28743), .B2(
        \xmem_data[103][6] ), .ZN(n12290) );
  NAND4_X1 U16439 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  NOR3_X1 U16440 ( .A1(n12296), .A2(n12295), .A3(n12294), .ZN(n12299) );
  AOI22_X1 U16441 ( .A1(n30191), .A2(\xmem_data[100][6] ), .B1(n29589), .B2(
        \xmem_data[101][6] ), .ZN(n12298) );
  AOI22_X1 U16442 ( .A1(n28740), .A2(\xmem_data[96][6] ), .B1(n28667), .B2(
        \xmem_data[97][6] ), .ZN(n12297) );
  NAND4_X1 U16443 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  OAI21_X1 U16444 ( .B1(n12302), .B2(n12301), .A(n28762), .ZN(n12339) );
  AOI22_X1 U16445 ( .A1(n27716), .A2(\xmem_data[20][6] ), .B1(n29381), .B2(
        \xmem_data[21][6] ), .ZN(n12306) );
  AOI22_X1 U16446 ( .A1(n28765), .A2(\xmem_data[24][6] ), .B1(n27743), .B2(
        \xmem_data[25][6] ), .ZN(n12305) );
  AOI22_X1 U16447 ( .A1(n28702), .A2(\xmem_data[18][6] ), .B1(n3301), .B2(
        \xmem_data[19][6] ), .ZN(n12304) );
  NAND2_X1 U16448 ( .A1(n29721), .A2(\xmem_data[17][6] ), .ZN(n12303) );
  NAND4_X1 U16449 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12309) );
  AOI22_X1 U16450 ( .A1(n28787), .A2(\xmem_data[0][6] ), .B1(n29761), .B2(
        \xmem_data[1][6] ), .ZN(n12307) );
  INV_X1 U16451 ( .A(n12307), .ZN(n12308) );
  NOR2_X1 U16452 ( .A1(n12309), .A2(n12308), .ZN(n12336) );
  AOI22_X1 U16453 ( .A1(n26812), .A2(\xmem_data[14][6] ), .B1(n28781), .B2(
        \xmem_data[15][6] ), .ZN(n12311) );
  AOI22_X1 U16454 ( .A1(n3165), .A2(\xmem_data[12][6] ), .B1(n3191), .B2(
        \xmem_data[13][6] ), .ZN(n12310) );
  NAND2_X1 U16455 ( .A1(n12311), .A2(n12310), .ZN(n12314) );
  AOI22_X1 U16456 ( .A1(n29590), .A2(\xmem_data[4][6] ), .B1(n30730), .B2(
        \xmem_data[5][6] ), .ZN(n12312) );
  INV_X1 U16457 ( .A(n12312), .ZN(n12313) );
  NOR2_X1 U16458 ( .A1(n12314), .A2(n12313), .ZN(n12335) );
  AND2_X1 U16459 ( .A1(n29423), .A2(\xmem_data[30][6] ), .ZN(n12320) );
  AND2_X1 U16460 ( .A1(n29565), .A2(\xmem_data[31][6] ), .ZN(n12315) );
  AOI21_X1 U16461 ( .B1(n29753), .B2(\xmem_data[29][6] ), .A(n12315), .ZN(
        n12318) );
  AOI22_X1 U16462 ( .A1(n3227), .A2(\xmem_data[26][6] ), .B1(n3153), .B2(
        \xmem_data[27][6] ), .ZN(n12317) );
  NAND2_X1 U16463 ( .A1(n28173), .A2(\xmem_data[16][6] ), .ZN(n12316) );
  NOR2_X1 U16464 ( .A1(n12320), .A2(n12319), .ZN(n12334) );
  AOI22_X1 U16465 ( .A1(n30250), .A2(\xmem_data[8][6] ), .B1(n27753), .B2(
        \xmem_data[9][6] ), .ZN(n12321) );
  INV_X1 U16466 ( .A(n12321), .ZN(n12332) );
  AOI22_X1 U16467 ( .A1(n29489), .A2(\xmem_data[22][6] ), .B1(n28772), .B2(
        \xmem_data[23][6] ), .ZN(n12329) );
  AOI22_X1 U16468 ( .A1(n28780), .A2(\xmem_data[10][6] ), .B1(n27517), .B2(
        \xmem_data[11][6] ), .ZN(n12322) );
  INV_X1 U16469 ( .A(n12322), .ZN(n12327) );
  AND2_X1 U16470 ( .A1(n3244), .A2(\xmem_data[2][6] ), .ZN(n12326) );
  NAND2_X1 U16471 ( .A1(n28788), .A2(\xmem_data[6][6] ), .ZN(n12324) );
  AOI22_X1 U16472 ( .A1(\xmem_data[7][6] ), .A2(n30744), .B1(n3129), .B2(
        \xmem_data[3][6] ), .ZN(n12323) );
  NAND2_X1 U16473 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  NOR3_X1 U16474 ( .A1(n12327), .A2(n12326), .A3(n12325), .ZN(n12328) );
  NAND2_X1 U16475 ( .A1(n12329), .A2(n12328), .ZN(n12330) );
  NOR3_X1 U16476 ( .A1(n12332), .A2(n12331), .A3(n12330), .ZN(n12333) );
  NAND4_X1 U16477 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12337) );
  NAND2_X1 U16478 ( .A1(n12337), .A2(n28794), .ZN(n12338) );
  XNOR2_X1 U16479 ( .A(n35112), .B(\fmem_data[11][3] ), .ZN(n26152) );
  XOR2_X1 U16480 ( .A(\fmem_data[11][2] ), .B(\fmem_data[11][3] ), .Z(n12342)
         );
  OAI22_X1 U16481 ( .A1(n30353), .A2(n34533), .B1(n26152), .B2(n34429), .ZN(
        n34225) );
  XNOR2_X1 U16482 ( .A(n32225), .B(\fmem_data[9][3] ), .ZN(n26252) );
  XOR2_X1 U16483 ( .A(\fmem_data[9][2] ), .B(\fmem_data[9][3] ), .Z(n12343) );
  AOI22_X1 U16484 ( .A1(n27903), .A2(\xmem_data[96][6] ), .B1(n3375), .B2(
        \xmem_data[97][6] ), .ZN(n12347) );
  AOI22_X1 U16485 ( .A1(n25450), .A2(\xmem_data[98][6] ), .B1(n28972), .B2(
        \xmem_data[99][6] ), .ZN(n12346) );
  AOI22_X1 U16486 ( .A1(n3358), .A2(\xmem_data[100][6] ), .B1(n28346), .B2(
        \xmem_data[101][6] ), .ZN(n12345) );
  AOI22_X1 U16487 ( .A1(n22675), .A2(\xmem_data[102][6] ), .B1(n30891), .B2(
        \xmem_data[103][6] ), .ZN(n12344) );
  NAND4_X1 U16488 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12365) );
  AOI22_X1 U16489 ( .A1(n29009), .A2(\xmem_data[104][6] ), .B1(n29008), .B2(
        \xmem_data[105][6] ), .ZN(n12351) );
  AOI22_X1 U16490 ( .A1(n3212), .A2(\xmem_data[106][6] ), .B1(n29010), .B2(
        \xmem_data[107][6] ), .ZN(n12350) );
  AOI22_X1 U16491 ( .A1(n21006), .A2(\xmem_data[108][6] ), .B1(n29012), .B2(
        \xmem_data[109][6] ), .ZN(n12349) );
  AOI22_X1 U16492 ( .A1(n23776), .A2(\xmem_data[110][6] ), .B1(n28428), .B2(
        \xmem_data[111][6] ), .ZN(n12348) );
  NAND4_X1 U16493 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12364) );
  AOI22_X1 U16494 ( .A1(n20816), .A2(\xmem_data[112][6] ), .B1(n28955), .B2(
        \xmem_data[113][6] ), .ZN(n12356) );
  AOI22_X1 U16495 ( .A1(n20553), .A2(\xmem_data[114][6] ), .B1(n24467), .B2(
        \xmem_data[115][6] ), .ZN(n12355) );
  AND2_X1 U16496 ( .A1(n29017), .A2(\xmem_data[116][6] ), .ZN(n12352) );
  AOI21_X1 U16497 ( .B1(n30674), .B2(\xmem_data[117][6] ), .A(n12352), .ZN(
        n12354) );
  AOI22_X1 U16498 ( .A1(n20579), .A2(\xmem_data[118][6] ), .B1(n25686), .B2(
        \xmem_data[119][6] ), .ZN(n12353) );
  NAND4_X1 U16499 ( .A1(n12356), .A2(n12355), .A3(n12354), .A4(n12353), .ZN(
        n12363) );
  AOI22_X1 U16500 ( .A1(n28947), .A2(\xmem_data[120][6] ), .B1(n21308), .B2(
        \xmem_data[121][6] ), .ZN(n12361) );
  AND2_X1 U16501 ( .A1(n30589), .A2(\xmem_data[122][6] ), .ZN(n12357) );
  AOI21_X1 U16502 ( .B1(n30906), .B2(\xmem_data[123][6] ), .A(n12357), .ZN(
        n12360) );
  AOI22_X1 U16503 ( .A1(n3218), .A2(\xmem_data[124][6] ), .B1(n29026), .B2(
        \xmem_data[125][6] ), .ZN(n12359) );
  AOI22_X1 U16504 ( .A1(n29028), .A2(\xmem_data[126][6] ), .B1(n29027), .B2(
        \xmem_data[127][6] ), .ZN(n12358) );
  NAND4_X1 U16505 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  OR4_X1 U16506 ( .A1(n12365), .A2(n12364), .A3(n12363), .A4(n12362), .ZN(
        n12389) );
  AOI22_X1 U16507 ( .A1(n29055), .A2(\xmem_data[80][6] ), .B1(n29054), .B2(
        \xmem_data[81][6] ), .ZN(n12370) );
  AOI22_X1 U16508 ( .A1(n27525), .A2(\xmem_data[82][6] ), .B1(n3179), .B2(
        \xmem_data[83][6] ), .ZN(n12369) );
  AND2_X1 U16509 ( .A1(n27526), .A2(\xmem_data[84][6] ), .ZN(n12366) );
  AOI21_X1 U16510 ( .B1(n20985), .B2(\xmem_data[85][6] ), .A(n12366), .ZN(
        n12368) );
  AOI22_X1 U16511 ( .A1(n24468), .A2(\xmem_data[86][6] ), .B1(n29057), .B2(
        \xmem_data[87][6] ), .ZN(n12367) );
  NAND4_X1 U16512 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12387) );
  AND2_X1 U16513 ( .A1(n29253), .A2(\xmem_data[90][6] ), .ZN(n12371) );
  AOI21_X1 U16514 ( .B1(n24631), .B2(\xmem_data[91][6] ), .A(n12371), .ZN(
        n12375) );
  AOI22_X1 U16515 ( .A1(n12471), .A2(\xmem_data[88][6] ), .B1(n3228), .B2(
        \xmem_data[89][6] ), .ZN(n12374) );
  AOI22_X1 U16516 ( .A1(n3218), .A2(\xmem_data[92][6] ), .B1(n29065), .B2(
        \xmem_data[93][6] ), .ZN(n12373) );
  AOI22_X1 U16517 ( .A1(n23739), .A2(\xmem_data[94][6] ), .B1(n29257), .B2(
        \xmem_data[95][6] ), .ZN(n12372) );
  NAND4_X1 U16518 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12386) );
  AOI22_X1 U16519 ( .A1(n20559), .A2(\xmem_data[64][6] ), .B1(n29350), .B2(
        \xmem_data[65][6] ), .ZN(n12379) );
  AOI22_X1 U16520 ( .A1(n25492), .A2(n20682), .B1(n28972), .B2(
        \xmem_data[67][6] ), .ZN(n12378) );
  AOI22_X1 U16521 ( .A1(n13475), .A2(\xmem_data[68][6] ), .B1(n20716), .B2(
        \xmem_data[69][6] ), .ZN(n12377) );
  AOI22_X1 U16522 ( .A1(n25605), .A2(\xmem_data[70][6] ), .B1(n29023), .B2(
        \xmem_data[71][6] ), .ZN(n12376) );
  NAND4_X1 U16523 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12376), .ZN(
        n12385) );
  AOI22_X1 U16524 ( .A1(n29046), .A2(\xmem_data[72][6] ), .B1(n20776), .B2(
        \xmem_data[73][6] ), .ZN(n12383) );
  AOI22_X1 U16525 ( .A1(n29188), .A2(\xmem_data[74][6] ), .B1(n24593), .B2(
        \xmem_data[75][6] ), .ZN(n12382) );
  AOI22_X1 U16526 ( .A1(n29048), .A2(\xmem_data[76][6] ), .B1(n29047), .B2(
        \xmem_data[77][6] ), .ZN(n12381) );
  AOI22_X1 U16527 ( .A1(n29049), .A2(\xmem_data[78][6] ), .B1(n28428), .B2(
        \xmem_data[79][6] ), .ZN(n12380) );
  NAND4_X1 U16528 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12384) );
  AOI22_X1 U16529 ( .A1(n12389), .A2(n28968), .B1(n12388), .B2(n29041), .ZN(
        n12437) );
  AOI22_X1 U16530 ( .A1(n25486), .A2(\xmem_data[0][6] ), .B1(n28344), .B2(
        \xmem_data[1][6] ), .ZN(n12393) );
  AOI22_X1 U16531 ( .A1(n29045), .A2(\xmem_data[2][6] ), .B1(n27447), .B2(
        \xmem_data[3][6] ), .ZN(n12392) );
  AOI22_X1 U16532 ( .A1(n22739), .A2(\xmem_data[4][6] ), .B1(n30744), .B2(
        \xmem_data[5][6] ), .ZN(n12391) );
  AOI22_X1 U16533 ( .A1(n22675), .A2(\xmem_data[6][6] ), .B1(n30891), .B2(
        \xmem_data[7][6] ), .ZN(n12390) );
  NAND4_X1 U16534 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        n12411) );
  AOI22_X1 U16535 ( .A1(n22703), .A2(\xmem_data[8][6] ), .B1(n29807), .B2(
        \xmem_data[9][6] ), .ZN(n12397) );
  AOI22_X1 U16536 ( .A1(n28993), .A2(\xmem_data[10][6] ), .B1(n29317), .B2(
        \xmem_data[11][6] ), .ZN(n12396) );
  AOI22_X1 U16537 ( .A1(n20940), .A2(\xmem_data[12][6] ), .B1(n28994), .B2(
        \xmem_data[13][6] ), .ZN(n12395) );
  AOI22_X1 U16538 ( .A1(n28380), .A2(\xmem_data[14][6] ), .B1(n28061), .B2(
        \xmem_data[15][6] ), .ZN(n12394) );
  NAND4_X1 U16539 ( .A1(n12397), .A2(n12396), .A3(n12395), .A4(n12394), .ZN(
        n12410) );
  AOI22_X1 U16540 ( .A1(n25581), .A2(\xmem_data[16][6] ), .B1(n28202), .B2(
        \xmem_data[17][6] ), .ZN(n12402) );
  AOI22_X1 U16541 ( .A1(n28983), .A2(\xmem_data[18][6] ), .B1(n22684), .B2(
        \xmem_data[19][6] ), .ZN(n12401) );
  AND2_X1 U16542 ( .A1(n28979), .A2(\xmem_data[20][6] ), .ZN(n12398) );
  AOI21_X1 U16543 ( .B1(n20826), .B2(\xmem_data[21][6] ), .A(n12398), .ZN(
        n12400) );
  AOI22_X1 U16544 ( .A1(n20951), .A2(\xmem_data[22][6] ), .B1(n21061), .B2(
        \xmem_data[23][6] ), .ZN(n12399) );
  NAND4_X1 U16545 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12409) );
  AOI22_X1 U16546 ( .A1(n21309), .A2(\xmem_data[24][6] ), .B1(n25443), .B2(
        \xmem_data[25][6] ), .ZN(n12407) );
  AND2_X1 U16547 ( .A1(n24172), .A2(\xmem_data[26][6] ), .ZN(n12403) );
  AOI21_X1 U16548 ( .B1(n20991), .B2(\xmem_data[27][6] ), .A(n12403), .ZN(
        n12406) );
  AOI22_X1 U16549 ( .A1(n3217), .A2(\xmem_data[28][6] ), .B1(n23740), .B2(
        \xmem_data[29][6] ), .ZN(n12405) );
  AOI22_X1 U16550 ( .A1(n29095), .A2(\xmem_data[30][6] ), .B1(n24438), .B2(
        \xmem_data[31][6] ), .ZN(n12404) );
  NAND4_X1 U16551 ( .A1(n12407), .A2(n12406), .A3(n12405), .A4(n12404), .ZN(
        n12408) );
  OR4_X1 U16552 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12435) );
  AOI22_X1 U16553 ( .A1(n24555), .A2(\xmem_data[38][6] ), .B1(n16986), .B2(
        \xmem_data[39][6] ), .ZN(n12415) );
  AOI22_X1 U16554 ( .A1(n21068), .A2(\xmem_data[32][6] ), .B1(n28952), .B2(
        \xmem_data[33][6] ), .ZN(n12414) );
  AOI22_X1 U16555 ( .A1(n31252), .A2(\xmem_data[34][6] ), .B1(n20961), .B2(
        \xmem_data[35][6] ), .ZN(n12413) );
  AOI22_X1 U16556 ( .A1(n30884), .A2(\xmem_data[36][6] ), .B1(n30886), .B2(
        \xmem_data[37][6] ), .ZN(n12412) );
  NAND4_X1 U16557 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12433) );
  AOI22_X1 U16558 ( .A1(n29046), .A2(\xmem_data[40][6] ), .B1(n27517), .B2(
        \xmem_data[41][6] ), .ZN(n12419) );
  AOI22_X1 U16559 ( .A1(n24457), .A2(\xmem_data[42][6] ), .B1(n20800), .B2(
        \xmem_data[43][6] ), .ZN(n12418) );
  AOI22_X1 U16560 ( .A1(n29048), .A2(\xmem_data[44][6] ), .B1(n29047), .B2(
        \xmem_data[45][6] ), .ZN(n12417) );
  AOI22_X1 U16561 ( .A1(n29049), .A2(\xmem_data[46][6] ), .B1(n28385), .B2(
        \xmem_data[47][6] ), .ZN(n12416) );
  NAND4_X1 U16562 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        n12432) );
  AND2_X1 U16563 ( .A1(n28501), .A2(\xmem_data[58][6] ), .ZN(n12420) );
  AOI21_X1 U16564 ( .B1(n24631), .B2(\xmem_data[59][6] ), .A(n12420), .ZN(
        n12424) );
  AOI22_X1 U16565 ( .A1(n21309), .A2(\xmem_data[56][6] ), .B1(n3384), .B2(
        \xmem_data[57][6] ), .ZN(n12423) );
  AOI22_X1 U16566 ( .A1(n3218), .A2(\xmem_data[60][6] ), .B1(n29065), .B2(
        \xmem_data[61][6] ), .ZN(n12422) );
  AOI22_X1 U16567 ( .A1(n23739), .A2(\xmem_data[62][6] ), .B1(n29174), .B2(
        \xmem_data[63][6] ), .ZN(n12421) );
  NAND4_X1 U16568 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12431) );
  AOI22_X1 U16569 ( .A1(n29055), .A2(\xmem_data[48][6] ), .B1(n29054), .B2(
        \xmem_data[49][6] ), .ZN(n12429) );
  AOI22_X1 U16570 ( .A1(n24223), .A2(\xmem_data[50][6] ), .B1(n29325), .B2(
        \xmem_data[51][6] ), .ZN(n12428) );
  AND2_X1 U16571 ( .A1(n29017), .A2(\xmem_data[52][6] ), .ZN(n12425) );
  AOI21_X1 U16572 ( .B1(n20770), .B2(\xmem_data[53][6] ), .A(n12425), .ZN(
        n12427) );
  AOI22_X1 U16573 ( .A1(n24624), .A2(\xmem_data[54][6] ), .B1(n29057), .B2(
        \xmem_data[55][6] ), .ZN(n12426) );
  NAND4_X1 U16574 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12430) );
  OR4_X1 U16575 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12434) );
  AOI22_X1 U16576 ( .A1(n12435), .A2(n29002), .B1(n12434), .B2(n29078), .ZN(
        n12436) );
  NAND2_X1 U16577 ( .A1(n12437), .A2(n12436), .ZN(n35021) );
  XNOR2_X1 U16578 ( .A(n35021), .B(\fmem_data[9][3] ), .ZN(n33043) );
  OAI22_X1 U16579 ( .A1(n26252), .A2(n33875), .B1(n33043), .B2(n33873), .ZN(
        n33934) );
  AOI22_X1 U16580 ( .A1(n27550), .A2(\xmem_data[32][2] ), .B1(n28952), .B2(
        \xmem_data[33][2] ), .ZN(n12441) );
  AOI22_X1 U16581 ( .A1(n28007), .A2(\xmem_data[34][2] ), .B1(n28050), .B2(
        \xmem_data[35][2] ), .ZN(n12440) );
  AOI22_X1 U16582 ( .A1(n30854), .A2(\xmem_data[36][2] ), .B1(n30744), .B2(
        \xmem_data[37][2] ), .ZN(n12439) );
  AOI22_X1 U16583 ( .A1(n27513), .A2(\xmem_data[38][2] ), .B1(n28298), .B2(
        \xmem_data[39][2] ), .ZN(n12438) );
  NAND4_X1 U16584 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n12438), .ZN(
        n12457) );
  AOI22_X1 U16585 ( .A1(n29046), .A2(\xmem_data[40][2] ), .B1(n3466), .B2(
        \xmem_data[41][2] ), .ZN(n12445) );
  AOI22_X1 U16586 ( .A1(n3208), .A2(\xmem_data[42][2] ), .B1(n24593), .B2(
        \xmem_data[43][2] ), .ZN(n12444) );
  AOI22_X1 U16587 ( .A1(n29048), .A2(\xmem_data[44][2] ), .B1(n29047), .B2(
        \xmem_data[45][2] ), .ZN(n12443) );
  AOI22_X1 U16588 ( .A1(n29049), .A2(\xmem_data[46][2] ), .B1(n28061), .B2(
        \xmem_data[47][2] ), .ZN(n12442) );
  NAND4_X1 U16589 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12456) );
  AOI22_X1 U16590 ( .A1(n29055), .A2(\xmem_data[48][2] ), .B1(n29054), .B2(
        \xmem_data[49][2] ), .ZN(n12449) );
  AOI22_X1 U16591 ( .A1(n27365), .A2(\xmem_data[50][2] ), .B1(n30497), .B2(
        \xmem_data[51][2] ), .ZN(n12448) );
  AOI22_X1 U16592 ( .A1(n27526), .A2(\xmem_data[52][2] ), .B1(n20826), .B2(
        \xmem_data[53][2] ), .ZN(n12447) );
  AOI22_X1 U16593 ( .A1(n25528), .A2(\xmem_data[54][2] ), .B1(n29057), .B2(
        \xmem_data[55][2] ), .ZN(n12446) );
  NAND4_X1 U16594 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12455) );
  AOI22_X1 U16595 ( .A1(n25629), .A2(\xmem_data[56][2] ), .B1(n29661), .B2(
        \xmem_data[57][2] ), .ZN(n12453) );
  AOI22_X1 U16596 ( .A1(n25687), .A2(\xmem_data[58][2] ), .B1(n29254), .B2(
        \xmem_data[59][2] ), .ZN(n12452) );
  AOI22_X1 U16597 ( .A1(n3220), .A2(\xmem_data[60][2] ), .B1(n29065), .B2(
        \xmem_data[61][2] ), .ZN(n12451) );
  AOI22_X1 U16598 ( .A1(n23739), .A2(\xmem_data[62][2] ), .B1(n28083), .B2(
        \xmem_data[63][2] ), .ZN(n12450) );
  NAND4_X1 U16599 ( .A1(n12453), .A2(n12452), .A3(n12451), .A4(n12450), .ZN(
        n12454) );
  OR4_X1 U16600 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12458) );
  NAND2_X1 U16601 ( .A1(n12458), .A2(n29078), .ZN(n12528) );
  AOI22_X1 U16602 ( .A1(n25616), .A2(\xmem_data[0][2] ), .B1(n3375), .B2(
        \xmem_data[1][2] ), .ZN(n12462) );
  AOI22_X1 U16603 ( .A1(n29045), .A2(\xmem_data[2][2] ), .B1(n25422), .B2(
        \xmem_data[3][2] ), .ZN(n12461) );
  AOI22_X1 U16604 ( .A1(n27863), .A2(\xmem_data[4][2] ), .B1(n25424), .B2(
        \xmem_data[5][2] ), .ZN(n12460) );
  AOI22_X1 U16605 ( .A1(n24212), .A2(\xmem_data[6][2] ), .B1(n20541), .B2(
        \xmem_data[7][2] ), .ZN(n12459) );
  NAND4_X1 U16606 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12479) );
  AOI22_X1 U16607 ( .A1(n22703), .A2(\xmem_data[8][2] ), .B1(n20718), .B2(
        \xmem_data[9][2] ), .ZN(n12466) );
  AOI22_X1 U16608 ( .A1(n28993), .A2(\xmem_data[10][2] ), .B1(n24509), .B2(
        \xmem_data[11][2] ), .ZN(n12465) );
  AOI22_X1 U16609 ( .A1(n25715), .A2(\xmem_data[12][2] ), .B1(n28994), .B2(
        \xmem_data[13][2] ), .ZN(n12464) );
  AOI22_X1 U16610 ( .A1(n29238), .A2(\xmem_data[14][2] ), .B1(n20731), .B2(
        \xmem_data[15][2] ), .ZN(n12463) );
  NAND4_X1 U16611 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12478) );
  AOI22_X1 U16612 ( .A1(n28429), .A2(\xmem_data[16][2] ), .B1(n24522), .B2(
        \xmem_data[17][2] ), .ZN(n12470) );
  AOI22_X1 U16613 ( .A1(n28983), .A2(\xmem_data[18][2] ), .B1(n25582), .B2(
        \xmem_data[19][2] ), .ZN(n12469) );
  AOI22_X1 U16614 ( .A1(n28979), .A2(\xmem_data[20][2] ), .B1(n30901), .B2(
        \xmem_data[21][2] ), .ZN(n12468) );
  AOI22_X1 U16615 ( .A1(n27435), .A2(\xmem_data[22][2] ), .B1(n29057), .B2(
        \xmem_data[23][2] ), .ZN(n12467) );
  NAND4_X1 U16616 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12477) );
  AOI22_X1 U16617 ( .A1(n12471), .A2(\xmem_data[24][2] ), .B1(n3305), .B2(
        \xmem_data[25][2] ), .ZN(n12475) );
  AOI22_X1 U16618 ( .A1(n27437), .A2(\xmem_data[26][2] ), .B1(n23734), .B2(
        \xmem_data[27][2] ), .ZN(n12474) );
  AOI22_X1 U16619 ( .A1(n3218), .A2(\xmem_data[28][2] ), .B1(n28367), .B2(
        \xmem_data[29][2] ), .ZN(n12473) );
  AOI22_X1 U16620 ( .A1(n28319), .A2(\xmem_data[30][2] ), .B1(n25416), .B2(
        \xmem_data[31][2] ), .ZN(n12472) );
  NAND4_X1 U16621 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12476) );
  OR4_X1 U16622 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  NAND2_X1 U16623 ( .A1(n12480), .A2(n29002), .ZN(n12527) );
  AOI22_X1 U16624 ( .A1(n28342), .A2(\xmem_data[96][2] ), .B1(n3129), .B2(
        \xmem_data[97][2] ), .ZN(n12484) );
  AOI22_X1 U16625 ( .A1(n24657), .A2(\xmem_data[98][2] ), .B1(n28972), .B2(
        \xmem_data[99][2] ), .ZN(n12483) );
  AOI22_X1 U16626 ( .A1(n27943), .A2(\xmem_data[100][2] ), .B1(n30608), .B2(
        \xmem_data[101][2] ), .ZN(n12482) );
  AOI22_X1 U16627 ( .A1(n17012), .A2(\xmem_data[102][2] ), .B1(n27537), .B2(
        \xmem_data[103][2] ), .ZN(n12481) );
  NAND4_X1 U16628 ( .A1(n12484), .A2(n12483), .A3(n12482), .A4(n12481), .ZN(
        n12500) );
  AOI22_X1 U16629 ( .A1(n29009), .A2(\xmem_data[104][2] ), .B1(n29008), .B2(
        \xmem_data[105][2] ), .ZN(n12488) );
  AOI22_X1 U16630 ( .A1(n3213), .A2(\xmem_data[106][2] ), .B1(n29010), .B2(
        \xmem_data[107][2] ), .ZN(n12487) );
  AOI22_X1 U16631 ( .A1(n27918), .A2(\xmem_data[108][2] ), .B1(n29012), .B2(
        \xmem_data[109][2] ), .ZN(n12486) );
  AOI22_X1 U16632 ( .A1(n30616), .A2(\xmem_data[110][2] ), .B1(n3177), .B2(
        \xmem_data[111][2] ), .ZN(n12485) );
  NAND4_X1 U16633 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(
        n12499) );
  AOI22_X1 U16634 ( .A1(n27856), .A2(\xmem_data[112][2] ), .B1(n28955), .B2(
        \xmem_data[113][2] ), .ZN(n12492) );
  AOI22_X1 U16635 ( .A1(n20553), .A2(\xmem_data[114][2] ), .B1(n29151), .B2(
        \xmem_data[115][2] ), .ZN(n12491) );
  AOI22_X1 U16636 ( .A1(n29017), .A2(\xmem_data[116][2] ), .B1(n25628), .B2(
        \xmem_data[117][2] ), .ZN(n12490) );
  AOI22_X1 U16637 ( .A1(n27435), .A2(\xmem_data[118][2] ), .B1(n25441), .B2(
        \xmem_data[119][2] ), .ZN(n12489) );
  NAND4_X1 U16638 ( .A1(n12492), .A2(n12491), .A3(n12490), .A4(n12489), .ZN(
        n12498) );
  AOI22_X1 U16639 ( .A1(n23731), .A2(\xmem_data[122][2] ), .B1(n25413), .B2(
        \xmem_data[123][2] ), .ZN(n12496) );
  AOI22_X1 U16640 ( .A1(n21309), .A2(\xmem_data[120][2] ), .B1(n21308), .B2(
        \xmem_data[121][2] ), .ZN(n12495) );
  AOI22_X1 U16641 ( .A1(n3219), .A2(\xmem_data[124][2] ), .B1(n29026), .B2(
        \xmem_data[125][2] ), .ZN(n12494) );
  AOI22_X1 U16642 ( .A1(n29028), .A2(\xmem_data[126][2] ), .B1(n29027), .B2(
        \xmem_data[127][2] ), .ZN(n12493) );
  NAND4_X1 U16643 ( .A1(n12496), .A2(n12495), .A3(n12494), .A4(n12493), .ZN(
        n12497) );
  OR4_X1 U16644 ( .A1(n12500), .A2(n12499), .A3(n12498), .A4(n12497), .ZN(
        n12501) );
  NAND2_X1 U16645 ( .A1(n12501), .A2(n28968), .ZN(n12526) );
  AOI22_X1 U16646 ( .A1(n28075), .A2(\xmem_data[88][2] ), .B1(n21308), .B2(
        \xmem_data[89][2] ), .ZN(n12506) );
  AND2_X1 U16647 ( .A1(n25360), .A2(\xmem_data[90][2] ), .ZN(n12502) );
  AOI21_X1 U16648 ( .B1(n30592), .B2(\xmem_data[91][2] ), .A(n12502), .ZN(
        n12505) );
  AOI22_X1 U16649 ( .A1(n3221), .A2(\xmem_data[92][2] ), .B1(n29026), .B2(
        \xmem_data[93][2] ), .ZN(n12504) );
  AOI22_X1 U16650 ( .A1(n29028), .A2(\xmem_data[94][2] ), .B1(n29027), .B2(
        \xmem_data[95][2] ), .ZN(n12503) );
  NAND4_X1 U16651 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12523) );
  AOI22_X1 U16652 ( .A1(n25581), .A2(\xmem_data[80][2] ), .B1(n28955), .B2(
        \xmem_data[81][2] ), .ZN(n12511) );
  AOI22_X1 U16653 ( .A1(n24622), .A2(\xmem_data[82][2] ), .B1(n20782), .B2(
        \xmem_data[83][2] ), .ZN(n12510) );
  AND2_X1 U16654 ( .A1(n29017), .A2(\xmem_data[84][2] ), .ZN(n12507) );
  AOI21_X1 U16655 ( .B1(n29657), .B2(\xmem_data[85][2] ), .A(n12507), .ZN(
        n12509) );
  AOI22_X1 U16656 ( .A1(n24468), .A2(\xmem_data[86][2] ), .B1(n20827), .B2(
        \xmem_data[87][2] ), .ZN(n12508) );
  NAND4_X1 U16657 ( .A1(n12511), .A2(n12510), .A3(n12509), .A4(n12508), .ZN(
        n12522) );
  AOI22_X1 U16658 ( .A1(n25616), .A2(\xmem_data[64][2] ), .B1(n3374), .B2(
        \xmem_data[65][2] ), .ZN(n12515) );
  AOI22_X1 U16659 ( .A1(n29045), .A2(\xmem_data[66][2] ), .B1(n27447), .B2(
        \xmem_data[67][2] ), .ZN(n12514) );
  AOI22_X1 U16660 ( .A1(n28481), .A2(\xmem_data[68][2] ), .B1(n29308), .B2(
        \xmem_data[69][2] ), .ZN(n12513) );
  AOI22_X1 U16661 ( .A1(n22675), .A2(\xmem_data[70][2] ), .B1(n20495), .B2(
        \xmem_data[71][2] ), .ZN(n12512) );
  NAND4_X1 U16662 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12521) );
  AOI22_X1 U16663 ( .A1(n29009), .A2(\xmem_data[72][2] ), .B1(n29008), .B2(
        \xmem_data[73][2] ), .ZN(n12519) );
  AOI22_X1 U16664 ( .A1(n3212), .A2(\xmem_data[74][2] ), .B1(n29010), .B2(
        \xmem_data[75][2] ), .ZN(n12518) );
  AOI22_X1 U16665 ( .A1(n17043), .A2(\xmem_data[76][2] ), .B1(n29012), .B2(
        \xmem_data[77][2] ), .ZN(n12517) );
  AOI22_X1 U16666 ( .A1(n29238), .A2(\xmem_data[78][2] ), .B1(n3204), .B2(
        \xmem_data[79][2] ), .ZN(n12516) );
  NAND4_X1 U16667 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12520) );
  OR4_X1 U16668 ( .A1(n12523), .A2(n12522), .A3(n12521), .A4(n12520), .ZN(
        n12524) );
  NAND2_X1 U16669 ( .A1(n12524), .A2(n29041), .ZN(n12525) );
  XNOR2_X1 U16670 ( .A(n33743), .B(\fmem_data[9][7] ), .ZN(n34241) );
  AOI22_X1 U16671 ( .A1(n22669), .A2(\xmem_data[0][1] ), .B1(n28952), .B2(
        \xmem_data[1][1] ), .ZN(n12532) );
  AOI22_X1 U16672 ( .A1(n25514), .A2(\xmem_data[2][1] ), .B1(n25422), .B2(
        \xmem_data[3][1] ), .ZN(n12531) );
  AOI22_X1 U16673 ( .A1(n22739), .A2(\xmem_data[4][1] ), .B1(n30943), .B2(
        \xmem_data[5][1] ), .ZN(n12530) );
  AOI22_X1 U16674 ( .A1(n13168), .A2(\xmem_data[6][1] ), .B1(n29023), .B2(
        \xmem_data[7][1] ), .ZN(n12529) );
  NAND4_X1 U16675 ( .A1(n12532), .A2(n12531), .A3(n12530), .A4(n12529), .ZN(
        n12548) );
  AOI22_X1 U16676 ( .A1(n28517), .A2(\xmem_data[8][1] ), .B1(n29008), .B2(
        \xmem_data[9][1] ), .ZN(n12536) );
  AOI22_X1 U16677 ( .A1(n28993), .A2(\xmem_data[10][1] ), .B1(n20585), .B2(
        \xmem_data[11][1] ), .ZN(n12535) );
  AOI22_X1 U16678 ( .A1(n24219), .A2(\xmem_data[12][1] ), .B1(n28994), .B2(
        \xmem_data[13][1] ), .ZN(n12534) );
  AOI22_X1 U16679 ( .A1(n29238), .A2(\xmem_data[14][1] ), .B1(n24190), .B2(
        \xmem_data[15][1] ), .ZN(n12533) );
  NAND4_X1 U16680 ( .A1(n12536), .A2(n12535), .A3(n12534), .A4(n12533), .ZN(
        n12547) );
  AOI22_X1 U16681 ( .A1(n25679), .A2(\xmem_data[16][1] ), .B1(n28461), .B2(
        \xmem_data[17][1] ), .ZN(n12540) );
  AOI22_X1 U16682 ( .A1(n28983), .A2(\xmem_data[18][1] ), .B1(n22684), .B2(
        \xmem_data[19][1] ), .ZN(n12539) );
  AOI22_X1 U16683 ( .A1(n28979), .A2(\xmem_data[20][1] ), .B1(n17051), .B2(
        \xmem_data[21][1] ), .ZN(n12538) );
  AOI22_X1 U16684 ( .A1(n20769), .A2(\xmem_data[22][1] ), .B1(n25686), .B2(
        \xmem_data[23][1] ), .ZN(n12537) );
  NAND4_X1 U16685 ( .A1(n12540), .A2(n12539), .A3(n12538), .A4(n12537), .ZN(
        n12546) );
  AOI22_X1 U16686 ( .A1(n28974), .A2(\xmem_data[24][1] ), .B1(n21308), .B2(
        \xmem_data[25][1] ), .ZN(n12544) );
  AOI22_X1 U16687 ( .A1(n31347), .A2(\xmem_data[26][1] ), .B1(n29064), .B2(
        \xmem_data[27][1] ), .ZN(n12543) );
  AOI22_X1 U16688 ( .A1(n3222), .A2(\xmem_data[28][1] ), .B1(n25612), .B2(
        \xmem_data[29][1] ), .ZN(n12542) );
  AOI22_X1 U16689 ( .A1(n28356), .A2(\xmem_data[30][1] ), .B1(n25617), .B2(
        \xmem_data[31][1] ), .ZN(n12541) );
  NAND4_X1 U16690 ( .A1(n12544), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n12545) );
  OR4_X1 U16691 ( .A1(n12548), .A2(n12547), .A3(n12546), .A4(n12545), .ZN(
        n12549) );
  NAND2_X1 U16692 ( .A1(n12549), .A2(n29002), .ZN(n12617) );
  AOI22_X1 U16693 ( .A1(n23811), .A2(\xmem_data[32][1] ), .B1(n28952), .B2(
        \xmem_data[33][1] ), .ZN(n12553) );
  AOI22_X1 U16694 ( .A1(n29045), .A2(\xmem_data[34][1] ), .B1(n27447), .B2(
        \xmem_data[35][1] ), .ZN(n12552) );
  AOI22_X1 U16695 ( .A1(n20588), .A2(\xmem_data[36][1] ), .B1(n25424), .B2(
        \xmem_data[37][1] ), .ZN(n12551) );
  AOI22_X1 U16696 ( .A1(n24212), .A2(\xmem_data[38][1] ), .B1(n25425), .B2(
        \xmem_data[39][1] ), .ZN(n12550) );
  NAND4_X1 U16697 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12569) );
  AOI22_X1 U16698 ( .A1(n29046), .A2(\xmem_data[40][1] ), .B1(n31328), .B2(
        \xmem_data[41][1] ), .ZN(n12557) );
  AOI22_X1 U16699 ( .A1(n3212), .A2(\xmem_data[42][1] ), .B1(n20585), .B2(
        \xmem_data[43][1] ), .ZN(n12556) );
  AOI22_X1 U16700 ( .A1(n29048), .A2(\xmem_data[44][1] ), .B1(n29047), .B2(
        \xmem_data[45][1] ), .ZN(n12555) );
  AOI22_X1 U16701 ( .A1(n29049), .A2(\xmem_data[46][1] ), .B1(n30899), .B2(
        \xmem_data[47][1] ), .ZN(n12554) );
  NAND4_X1 U16702 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12568) );
  AOI22_X1 U16703 ( .A1(n29055), .A2(\xmem_data[48][1] ), .B1(n29054), .B2(
        \xmem_data[49][1] ), .ZN(n12561) );
  AOI22_X1 U16704 ( .A1(n27975), .A2(\xmem_data[50][1] ), .B1(n27542), .B2(
        \xmem_data[51][1] ), .ZN(n12560) );
  AOI22_X1 U16705 ( .A1(n11008), .A2(\xmem_data[52][1] ), .B1(n27852), .B2(
        \xmem_data[53][1] ), .ZN(n12559) );
  AOI22_X1 U16706 ( .A1(n24122), .A2(\xmem_data[54][1] ), .B1(n29057), .B2(
        \xmem_data[55][1] ), .ZN(n12558) );
  NAND4_X1 U16707 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12567) );
  AOI22_X1 U16708 ( .A1(n27958), .A2(\xmem_data[56][1] ), .B1(n21308), .B2(
        \xmem_data[57][1] ), .ZN(n12565) );
  AOI22_X1 U16709 ( .A1(n27437), .A2(\xmem_data[58][1] ), .B1(n29064), .B2(
        \xmem_data[59][1] ), .ZN(n12564) );
  AOI22_X1 U16710 ( .A1(n3219), .A2(\xmem_data[60][1] ), .B1(n29065), .B2(
        \xmem_data[61][1] ), .ZN(n12563) );
  AOI22_X1 U16711 ( .A1(n23739), .A2(\xmem_data[62][1] ), .B1(n27938), .B2(
        \xmem_data[63][1] ), .ZN(n12562) );
  NAND4_X1 U16712 ( .A1(n12565), .A2(n12564), .A3(n12563), .A4(n12562), .ZN(
        n12566) );
  OR4_X1 U16713 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12570) );
  NAND2_X1 U16714 ( .A1(n12570), .A2(n29078), .ZN(n12616) );
  AOI22_X1 U16715 ( .A1(n27903), .A2(\xmem_data[96][1] ), .B1(n3344), .B2(
        \xmem_data[97][1] ), .ZN(n12574) );
  AOI22_X1 U16716 ( .A1(n25514), .A2(\xmem_data[98][1] ), .B1(n28972), .B2(
        \xmem_data[99][1] ), .ZN(n12573) );
  AOI22_X1 U16717 ( .A1(n27943), .A2(\xmem_data[100][1] ), .B1(n20587), .B2(
        \xmem_data[101][1] ), .ZN(n12572) );
  AOI22_X1 U16718 ( .A1(n22702), .A2(\xmem_data[102][1] ), .B1(n30891), .B2(
        \xmem_data[103][1] ), .ZN(n12571) );
  NAND4_X1 U16719 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12590) );
  AOI22_X1 U16720 ( .A1(n29009), .A2(\xmem_data[104][1] ), .B1(n29008), .B2(
        \xmem_data[105][1] ), .ZN(n12578) );
  AOI22_X1 U16721 ( .A1(n3212), .A2(\xmem_data[106][1] ), .B1(n29010), .B2(
        \xmem_data[107][1] ), .ZN(n12577) );
  AOI22_X1 U16722 ( .A1(n23796), .A2(\xmem_data[108][1] ), .B1(n29012), .B2(
        \xmem_data[109][1] ), .ZN(n12576) );
  AOI22_X1 U16723 ( .A1(n29238), .A2(\xmem_data[110][1] ), .B1(n3177), .B2(
        \xmem_data[111][1] ), .ZN(n12575) );
  NAND4_X1 U16724 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12589) );
  AOI22_X1 U16725 ( .A1(n20506), .A2(\xmem_data[112][1] ), .B1(n28955), .B2(
        \xmem_data[113][1] ), .ZN(n12582) );
  AOI22_X1 U16726 ( .A1(n23723), .A2(\xmem_data[114][1] ), .B1(n27542), .B2(
        \xmem_data[115][1] ), .ZN(n12581) );
  AOI22_X1 U16727 ( .A1(n29017), .A2(\xmem_data[116][1] ), .B1(n25584), .B2(
        \xmem_data[117][1] ), .ZN(n12580) );
  AOI22_X1 U16728 ( .A1(n25388), .A2(\xmem_data[118][1] ), .B1(n20953), .B2(
        \xmem_data[119][1] ), .ZN(n12579) );
  NAND4_X1 U16729 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12588) );
  AOI22_X1 U16730 ( .A1(n28947), .A2(\xmem_data[120][1] ), .B1(n21308), .B2(
        \xmem_data[121][1] ), .ZN(n12586) );
  AOI22_X1 U16731 ( .A1(n22753), .A2(\xmem_data[122][1] ), .B1(n29064), .B2(
        \xmem_data[123][1] ), .ZN(n12585) );
  AOI22_X1 U16732 ( .A1(n3221), .A2(\xmem_data[124][1] ), .B1(n29026), .B2(
        \xmem_data[125][1] ), .ZN(n12584) );
  AOI22_X1 U16733 ( .A1(n29028), .A2(\xmem_data[126][1] ), .B1(n29027), .B2(
        \xmem_data[127][1] ), .ZN(n12583) );
  NAND4_X1 U16734 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12587) );
  OR4_X1 U16735 ( .A1(n12590), .A2(n12589), .A3(n12588), .A4(n12587), .ZN(
        n12591) );
  NAND2_X1 U16736 ( .A1(n12591), .A2(n28968), .ZN(n12615) );
  AOI22_X1 U16737 ( .A1(n25716), .A2(\xmem_data[80][1] ), .B1(n28955), .B2(
        \xmem_data[81][1] ), .ZN(n12596) );
  AOI22_X1 U16738 ( .A1(n25583), .A2(\xmem_data[82][1] ), .B1(n24166), .B2(
        \xmem_data[83][1] ), .ZN(n12595) );
  AND2_X1 U16739 ( .A1(n29017), .A2(\xmem_data[84][1] ), .ZN(n12592) );
  AOI21_X1 U16740 ( .B1(n28192), .B2(\xmem_data[85][1] ), .A(n12592), .ZN(
        n12594) );
  AOI22_X1 U16741 ( .A1(n29248), .A2(\xmem_data[86][1] ), .B1(n20827), .B2(
        \xmem_data[87][1] ), .ZN(n12593) );
  NAND4_X1 U16742 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12612) );
  AOI22_X1 U16743 ( .A1(n29009), .A2(\xmem_data[72][1] ), .B1(n29008), .B2(
        \xmem_data[73][1] ), .ZN(n12600) );
  AOI22_X1 U16744 ( .A1(n3212), .A2(\xmem_data[74][1] ), .B1(n29010), .B2(
        \xmem_data[75][1] ), .ZN(n12599) );
  AOI22_X1 U16745 ( .A1(n25520), .A2(\xmem_data[76][1] ), .B1(n29012), .B2(
        \xmem_data[77][1] ), .ZN(n12598) );
  AOI22_X1 U16746 ( .A1(n28380), .A2(\xmem_data[78][1] ), .B1(n25717), .B2(
        \xmem_data[79][1] ), .ZN(n12597) );
  NAND4_X1 U16747 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12611) );
  AOI22_X1 U16748 ( .A1(n24573), .A2(\xmem_data[88][1] ), .B1(n3386), .B2(
        \xmem_data[89][1] ), .ZN(n12604) );
  AOI22_X1 U16749 ( .A1(n22753), .A2(\xmem_data[90][1] ), .B1(n29064), .B2(
        \xmem_data[91][1] ), .ZN(n12603) );
  AOI22_X1 U16750 ( .A1(n3220), .A2(\xmem_data[92][1] ), .B1(n29026), .B2(
        \xmem_data[93][1] ), .ZN(n12602) );
  AOI22_X1 U16751 ( .A1(n29028), .A2(\xmem_data[94][1] ), .B1(n29027), .B2(
        \xmem_data[95][1] ), .ZN(n12601) );
  NAND4_X1 U16752 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12610) );
  AOI22_X1 U16753 ( .A1(n30550), .A2(\xmem_data[64][1] ), .B1(n3374), .B2(
        \xmem_data[65][1] ), .ZN(n12608) );
  AOI22_X1 U16754 ( .A1(n29045), .A2(\xmem_data[66][1] ), .B1(n28972), .B2(
        \xmem_data[67][1] ), .ZN(n12607) );
  AOI22_X1 U16755 ( .A1(n24590), .A2(\xmem_data[68][1] ), .B1(n17064), .B2(
        \xmem_data[69][1] ), .ZN(n12606) );
  AOI22_X1 U16756 ( .A1(n28345), .A2(\xmem_data[70][1] ), .B1(n20495), .B2(
        \xmem_data[71][1] ), .ZN(n12605) );
  NAND4_X1 U16757 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        n12609) );
  OR4_X1 U16758 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        n12613) );
  NAND2_X1 U16759 ( .A1(n12613), .A2(n29041), .ZN(n12614) );
  XNOR2_X1 U16760 ( .A(n33451), .B(\fmem_data[9][7] ), .ZN(n26254) );
  OAI22_X1 U16761 ( .A1(n35726), .A2(n34241), .B1(n26254), .B2(n35725), .ZN(
        n33933) );
  AOI22_X1 U16762 ( .A1(n22701), .A2(\xmem_data[32][3] ), .B1(n29451), .B2(
        \xmem_data[33][3] ), .ZN(n12621) );
  AOI22_X1 U16763 ( .A1(n22702), .A2(\xmem_data[34][3] ), .B1(n13436), .B2(
        \xmem_data[35][3] ), .ZN(n12620) );
  AOI22_X1 U16764 ( .A1(n22703), .A2(\xmem_data[36][3] ), .B1(n28091), .B2(
        \xmem_data[37][3] ), .ZN(n12619) );
  AOI22_X1 U16765 ( .A1(n20586), .A2(\xmem_data[38][3] ), .B1(n27919), .B2(
        \xmem_data[39][3] ), .ZN(n12618) );
  NAND4_X1 U16766 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12637) );
  AOI22_X1 U16767 ( .A1(n22718), .A2(\xmem_data[40][3] ), .B1(n22717), .B2(
        \xmem_data[41][3] ), .ZN(n12625) );
  AOI22_X1 U16768 ( .A1(n28097), .A2(\xmem_data[42][3] ), .B1(n25632), .B2(
        \xmem_data[43][3] ), .ZN(n12624) );
  AOI22_X1 U16769 ( .A1(n27461), .A2(\xmem_data[44][3] ), .B1(n3329), .B2(
        \xmem_data[45][3] ), .ZN(n12623) );
  AOI22_X1 U16770 ( .A1(n27365), .A2(\xmem_data[46][3] ), .B1(n22719), .B2(
        \xmem_data[47][3] ), .ZN(n12622) );
  NAND4_X1 U16771 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12636) );
  AOI22_X1 U16772 ( .A1(n27526), .A2(\xmem_data[48][3] ), .B1(n17051), .B2(
        \xmem_data[49][3] ), .ZN(n12629) );
  AOI22_X1 U16773 ( .A1(n22727), .A2(\xmem_data[50][3] ), .B1(n25724), .B2(
        \xmem_data[51][3] ), .ZN(n12628) );
  AOI22_X1 U16774 ( .A1(n22729), .A2(\xmem_data[52][3] ), .B1(n22728), .B2(
        \xmem_data[53][3] ), .ZN(n12627) );
  AOI22_X1 U16775 ( .A1(n28501), .A2(\xmem_data[54][3] ), .B1(n29254), .B2(
        \xmem_data[55][3] ), .ZN(n12626) );
  NAND4_X1 U16776 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12635) );
  AOI22_X1 U16777 ( .A1(n3218), .A2(\xmem_data[56][3] ), .B1(n22708), .B2(
        \xmem_data[57][3] ), .ZN(n12633) );
  AOI22_X1 U16778 ( .A1(n22710), .A2(\xmem_data[58][3] ), .B1(n22709), .B2(
        \xmem_data[59][3] ), .ZN(n12632) );
  AOI22_X1 U16779 ( .A1(n22711), .A2(\xmem_data[60][3] ), .B1(n20808), .B2(
        \xmem_data[61][3] ), .ZN(n12631) );
  AOI22_X1 U16780 ( .A1(n28045), .A2(\xmem_data[62][3] ), .B1(n22712), .B2(
        \xmem_data[63][3] ), .ZN(n12630) );
  NAND4_X1 U16781 ( .A1(n12633), .A2(n12632), .A3(n12631), .A4(n12630), .ZN(
        n12634) );
  OR4_X1 U16782 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        n12666) );
  AND2_X1 U16783 ( .A1(n22751), .A2(\xmem_data[16][3] ), .ZN(n12638) );
  AOI21_X1 U16784 ( .B1(n29657), .B2(\xmem_data[17][3] ), .A(n12638), .ZN(
        n12642) );
  AOI22_X1 U16785 ( .A1(n24122), .A2(\xmem_data[18][3] ), .B1(n25630), .B2(
        \xmem_data[19][3] ), .ZN(n12641) );
  AOI22_X1 U16786 ( .A1(n22752), .A2(\xmem_data[20][3] ), .B1(n3228), .B2(
        \xmem_data[21][3] ), .ZN(n12640) );
  AOI22_X1 U16787 ( .A1(n22753), .A2(\xmem_data[22][3] ), .B1(n29064), .B2(
        \xmem_data[23][3] ), .ZN(n12639) );
  NAND4_X1 U16788 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12648) );
  AOI22_X1 U16789 ( .A1(n25520), .A2(\xmem_data[8][3] ), .B1(n30872), .B2(
        \xmem_data[9][3] ), .ZN(n12646) );
  AOI22_X1 U16790 ( .A1(n29238), .A2(\xmem_data[10][3] ), .B1(n3177), .B2(
        \xmem_data[11][3] ), .ZN(n12645) );
  AOI22_X1 U16791 ( .A1(n27856), .A2(\xmem_data[12][3] ), .B1(n3328), .B2(
        \xmem_data[13][3] ), .ZN(n12644) );
  AOI22_X1 U16792 ( .A1(n28983), .A2(\xmem_data[14][3] ), .B1(n25582), .B2(
        \xmem_data[15][3] ), .ZN(n12643) );
  NAND4_X1 U16793 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12647) );
  OR2_X1 U16794 ( .A1(n12648), .A2(n12647), .ZN(n12663) );
  AOI22_X1 U16795 ( .A1(n3221), .A2(\xmem_data[24][3] ), .B1(n27445), .B2(
        \xmem_data[25][3] ), .ZN(n12655) );
  AOI22_X1 U16796 ( .A1(n22759), .A2(\xmem_data[28][3] ), .B1(n3280), .B2(
        \xmem_data[29][3] ), .ZN(n12649) );
  INV_X1 U16797 ( .A(n12649), .ZN(n12653) );
  AOI22_X1 U16798 ( .A1(n13469), .A2(\xmem_data[26][3] ), .B1(n22758), .B2(
        \xmem_data[27][3] ), .ZN(n12651) );
  NAND2_X1 U16799 ( .A1(n23813), .A2(\xmem_data[31][3] ), .ZN(n12650) );
  NAND2_X1 U16800 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  NOR2_X1 U16801 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  NAND2_X1 U16802 ( .A1(n12655), .A2(n12654), .ZN(n12661) );
  AOI22_X1 U16803 ( .A1(n22739), .A2(\xmem_data[0][3] ), .B1(n22738), .B2(
        \xmem_data[1][3] ), .ZN(n12659) );
  AOI22_X1 U16804 ( .A1(n22740), .A2(\xmem_data[2][3] ), .B1(n20495), .B2(
        \xmem_data[3][3] ), .ZN(n12658) );
  AOI22_X1 U16805 ( .A1(n22741), .A2(\xmem_data[4][3] ), .B1(n3119), .B2(
        \xmem_data[5][3] ), .ZN(n12657) );
  AOI22_X1 U16806 ( .A1(n22742), .A2(\xmem_data[6][3] ), .B1(n25573), .B2(
        \xmem_data[7][3] ), .ZN(n12656) );
  NAND4_X1 U16807 ( .A1(n12659), .A2(n12658), .A3(n12657), .A4(n12656), .ZN(
        n12660) );
  OR2_X1 U16808 ( .A1(n12661), .A2(n12660), .ZN(n12662) );
  NOR2_X1 U16809 ( .A1(n12663), .A2(n12662), .ZN(n12664) );
  NOR2_X1 U16810 ( .A1(n12664), .A2(n22022), .ZN(n12665) );
  AOI21_X1 U16811 ( .B1(n12666), .B2(n22735), .A(n12665), .ZN(n12714) );
  AOI22_X1 U16812 ( .A1(n20546), .A2(\xmem_data[64][3] ), .B1(n27944), .B2(
        \xmem_data[65][3] ), .ZN(n12670) );
  AOI22_X1 U16813 ( .A1(n22675), .A2(\xmem_data[66][3] ), .B1(n16986), .B2(
        \xmem_data[67][3] ), .ZN(n12669) );
  AOI22_X1 U16814 ( .A1(n22674), .A2(\xmem_data[68][3] ), .B1(n29437), .B2(
        \xmem_data[69][3] ), .ZN(n12668) );
  AOI22_X1 U16815 ( .A1(n22677), .A2(\xmem_data[70][3] ), .B1(n22676), .B2(
        \xmem_data[71][3] ), .ZN(n12667) );
  NAND4_X1 U16816 ( .A1(n12670), .A2(n12669), .A3(n12668), .A4(n12667), .ZN(
        n12687) );
  AOI22_X1 U16817 ( .A1(n28058), .A2(\xmem_data[72][3] ), .B1(n22682), .B2(
        \xmem_data[73][3] ), .ZN(n12674) );
  AOI22_X1 U16818 ( .A1(n24510), .A2(\xmem_data[74][3] ), .B1(n22683), .B2(
        \xmem_data[75][3] ), .ZN(n12673) );
  AOI22_X1 U16819 ( .A1(n23778), .A2(\xmem_data[76][3] ), .B1(n3337), .B2(
        \xmem_data[77][3] ), .ZN(n12672) );
  AOI22_X1 U16820 ( .A1(n22685), .A2(\xmem_data[78][3] ), .B1(n22684), .B2(
        \xmem_data[79][3] ), .ZN(n12671) );
  NAND4_X1 U16821 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12686) );
  AOI22_X1 U16822 ( .A1(n20733), .A2(\xmem_data[80][3] ), .B1(n20985), .B2(
        \xmem_data[81][3] ), .ZN(n12679) );
  AOI22_X1 U16823 ( .A1(n31261), .A2(\xmem_data[82][3] ), .B1(n27959), .B2(
        \xmem_data[83][3] ), .ZN(n12678) );
  AOI22_X1 U16824 ( .A1(n20709), .A2(\xmem_data[84][3] ), .B1(n3386), .B2(
        \xmem_data[85][3] ), .ZN(n12677) );
  AND2_X1 U16825 ( .A1(n30589), .A2(\xmem_data[86][3] ), .ZN(n12675) );
  AOI21_X1 U16826 ( .B1(n24631), .B2(\xmem_data[87][3] ), .A(n12675), .ZN(
        n12676) );
  NAND4_X1 U16827 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n12676), .ZN(
        n12685) );
  AOI22_X1 U16828 ( .A1(n3222), .A2(\xmem_data[88][3] ), .B1(n28367), .B2(
        \xmem_data[89][3] ), .ZN(n12683) );
  AOI22_X1 U16829 ( .A1(n22667), .A2(\xmem_data[90][3] ), .B1(n22666), .B2(
        \xmem_data[91][3] ), .ZN(n12682) );
  AOI22_X1 U16830 ( .A1(n22669), .A2(\xmem_data[92][3] ), .B1(n22668), .B2(
        \xmem_data[93][3] ), .ZN(n12681) );
  AOI22_X1 U16831 ( .A1(n25514), .A2(\xmem_data[94][3] ), .B1(n28374), .B2(
        \xmem_data[95][3] ), .ZN(n12680) );
  NAND4_X1 U16832 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12684) );
  OR4_X1 U16833 ( .A1(n12687), .A2(n12686), .A3(n12685), .A4(n12684), .ZN(
        n12689) );
  NOR2_X1 U16834 ( .A1(n22022), .A2(n39013), .ZN(n12688) );
  AOI21_X1 U16835 ( .B1(n12689), .B2(n22663), .A(n3883), .ZN(n12713) );
  AOI22_X1 U16836 ( .A1(n28415), .A2(\xmem_data[96][3] ), .B1(n27763), .B2(
        \xmem_data[97][3] ), .ZN(n12693) );
  AOI22_X1 U16837 ( .A1(n22675), .A2(\xmem_data[98][3] ), .B1(n29310), .B2(
        \xmem_data[99][3] ), .ZN(n12692) );
  AOI22_X1 U16838 ( .A1(n22674), .A2(\xmem_data[100][3] ), .B1(n29237), .B2(
        \xmem_data[101][3] ), .ZN(n12691) );
  AOI22_X1 U16839 ( .A1(n22677), .A2(\xmem_data[102][3] ), .B1(n22676), .B2(
        \xmem_data[103][3] ), .ZN(n12690) );
  NAND4_X1 U16840 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12710) );
  AOI22_X1 U16841 ( .A1(n20940), .A2(\xmem_data[104][3] ), .B1(n22682), .B2(
        \xmem_data[105][3] ), .ZN(n12697) );
  AOI22_X1 U16842 ( .A1(n29318), .A2(\xmem_data[106][3] ), .B1(n22683), .B2(
        \xmem_data[107][3] ), .ZN(n12696) );
  AOI22_X1 U16843 ( .A1(n25716), .A2(\xmem_data[108][3] ), .B1(n29297), .B2(
        \xmem_data[109][3] ), .ZN(n12695) );
  AOI22_X1 U16844 ( .A1(n22685), .A2(\xmem_data[110][3] ), .B1(n22684), .B2(
        \xmem_data[111][3] ), .ZN(n12694) );
  NAND4_X1 U16845 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12709) );
  AOI22_X1 U16846 ( .A1(n17049), .A2(\xmem_data[112][3] ), .B1(n20985), .B2(
        \xmem_data[113][3] ), .ZN(n12702) );
  AOI22_X1 U16847 ( .A1(n24686), .A2(\xmem_data[114][3] ), .B1(n3380), .B2(
        \xmem_data[115][3] ), .ZN(n12701) );
  AOI22_X1 U16848 ( .A1(n28037), .A2(\xmem_data[116][3] ), .B1(n3334), .B2(
        \xmem_data[117][3] ), .ZN(n12700) );
  AND2_X1 U16849 ( .A1(n28501), .A2(\xmem_data[118][3] ), .ZN(n12698) );
  AOI21_X1 U16850 ( .B1(n27439), .B2(\xmem_data[119][3] ), .A(n12698), .ZN(
        n12699) );
  NAND4_X1 U16851 ( .A1(n12702), .A2(n12701), .A3(n12700), .A4(n12699), .ZN(
        n12708) );
  AOI22_X1 U16852 ( .A1(n3220), .A2(\xmem_data[120][3] ), .B1(n27831), .B2(
        \xmem_data[121][3] ), .ZN(n12706) );
  AOI22_X1 U16853 ( .A1(n22667), .A2(\xmem_data[122][3] ), .B1(n22666), .B2(
        \xmem_data[123][3] ), .ZN(n12705) );
  AOI22_X1 U16854 ( .A1(n22669), .A2(\xmem_data[124][3] ), .B1(n22668), .B2(
        \xmem_data[125][3] ), .ZN(n12704) );
  AOI22_X1 U16855 ( .A1(n28007), .A2(\xmem_data[126][3] ), .B1(n28374), .B2(
        \xmem_data[127][3] ), .ZN(n12703) );
  NAND4_X1 U16856 ( .A1(n12706), .A2(n12705), .A3(n12704), .A4(n12703), .ZN(
        n12707) );
  OR4_X1 U16857 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  NAND2_X1 U16858 ( .A1(n12711), .A2(n22698), .ZN(n12712) );
  XOR2_X1 U16859 ( .A(\fmem_data[5][4] ), .B(\fmem_data[5][5] ), .Z(n12715) );
  XNOR2_X1 U16860 ( .A(n31233), .B(\fmem_data[5][5] ), .ZN(n30434) );
  OAI22_X1 U16861 ( .A1(n22778), .A2(n33857), .B1(n30434), .B2(n33859), .ZN(
        n33932) );
  XNOR2_X1 U16862 ( .A(n12716), .B(n35153), .ZN(n35210) );
  FA_X1 U16863 ( .A(n12719), .B(n12718), .CI(n12717), .CO(n35153), .S(n23594)
         );
  XNOR2_X1 U16864 ( .A(n12721), .B(n12720), .ZN(n12723) );
  XNOR2_X1 U16865 ( .A(n12723), .B(n12722), .ZN(n23593) );
  XNOR2_X1 U16866 ( .A(n12725), .B(n12724), .ZN(n12726) );
  XNOR2_X1 U16867 ( .A(n12727), .B(n12726), .ZN(n23592) );
  AOI22_X1 U16868 ( .A1(n30956), .A2(\xmem_data[8][5] ), .B1(n3372), .B2(
        \xmem_data[9][5] ), .ZN(n12732) );
  AOI22_X1 U16869 ( .A1(n30686), .A2(\xmem_data[10][5] ), .B1(n3200), .B2(
        \xmem_data[11][5] ), .ZN(n12731) );
  AOI22_X1 U16870 ( .A1(n20818), .A2(\xmem_data[12][5] ), .B1(n17049), .B2(
        \xmem_data[13][5] ), .ZN(n12730) );
  AND2_X1 U16871 ( .A1(n17050), .A2(\xmem_data[15][5] ), .ZN(n12728) );
  AOI21_X1 U16872 ( .B1(n17051), .B2(\xmem_data[14][5] ), .A(n12728), .ZN(
        n12729) );
  AND4_X1 U16873 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12744) );
  AOI22_X1 U16874 ( .A1(n20725), .A2(\xmem_data[24][5] ), .B1(n17061), .B2(
        \xmem_data[25][5] ), .ZN(n12736) );
  AOI22_X1 U16875 ( .A1(n17063), .A2(\xmem_data[26][5] ), .B1(n17062), .B2(
        \xmem_data[27][5] ), .ZN(n12735) );
  AOI22_X1 U16876 ( .A1(n25422), .A2(\xmem_data[28][5] ), .B1(n29180), .B2(
        \xmem_data[29][5] ), .ZN(n12734) );
  AOI22_X1 U16877 ( .A1(n17064), .A2(\xmem_data[30][5] ), .B1(n22740), .B2(
        \xmem_data[31][5] ), .ZN(n12733) );
  NAND4_X1 U16878 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12742) );
  AND2_X1 U16879 ( .A1(n17056), .A2(\xmem_data[16][5] ), .ZN(n12737) );
  AOI21_X1 U16880 ( .B1(n29118), .B2(\xmem_data[17][5] ), .A(n12737), .ZN(
        n12740) );
  AOI22_X1 U16881 ( .A1(n17033), .A2(\xmem_data[22][5] ), .B1(n23739), .B2(
        \xmem_data[23][5] ), .ZN(n12739) );
  AOI22_X1 U16882 ( .A1(n3333), .A2(\xmem_data[18][5] ), .B1(n16979), .B2(
        \xmem_data[19][5] ), .ZN(n12738) );
  NAND3_X1 U16883 ( .A1(n12740), .A2(n12739), .A3(n12738), .ZN(n12741) );
  NOR2_X1 U16884 ( .A1(n12742), .A2(n12741), .ZN(n12743) );
  AOI22_X1 U16885 ( .A1(n17041), .A2(\xmem_data[0][5] ), .B1(n14999), .B2(
        \xmem_data[1][5] ), .ZN(n12748) );
  AOI22_X1 U16886 ( .A1(n20939), .A2(\xmem_data[2][5] ), .B1(n17019), .B2(
        \xmem_data[3][5] ), .ZN(n12747) );
  AOI22_X1 U16887 ( .A1(n27919), .A2(\xmem_data[4][5] ), .B1(n17043), .B2(
        \xmem_data[5][5] ), .ZN(n12746) );
  AOI22_X1 U16888 ( .A1(n17044), .A2(\xmem_data[6][5] ), .B1(n24116), .B2(
        \xmem_data[7][5] ), .ZN(n12745) );
  NAND4_X1 U16889 ( .A1(n12748), .A2(n12747), .A3(n12746), .A4(n12745), .ZN(
        n12751) );
  AOI22_X1 U16890 ( .A1(n21066), .A2(\xmem_data[20][5] ), .B1(n3221), .B2(
        \xmem_data[21][5] ), .ZN(n12749) );
  INV_X1 U16891 ( .A(n12749), .ZN(n12750) );
  AOI22_X1 U16892 ( .A1(n16986), .A2(\xmem_data[96][5] ), .B1(n21076), .B2(
        \xmem_data[97][5] ), .ZN(n12755) );
  AOI22_X1 U16893 ( .A1(n16988), .A2(\xmem_data[98][5] ), .B1(n17019), .B2(
        \xmem_data[99][5] ), .ZN(n12754) );
  AOI22_X1 U16894 ( .A1(n20585), .A2(\xmem_data[100][5] ), .B1(n16989), .B2(
        \xmem_data[101][5] ), .ZN(n12753) );
  AOI22_X1 U16895 ( .A1(n16990), .A2(\xmem_data[102][5] ), .B1(n31254), .B2(
        \xmem_data[103][5] ), .ZN(n12752) );
  AOI22_X1 U16896 ( .A1(n30849), .A2(\xmem_data[104][5] ), .B1(n30598), .B2(
        \xmem_data[105][5] ), .ZN(n12759) );
  AOI22_X1 U16897 ( .A1(n3270), .A2(\xmem_data[106][5] ), .B1(n3201), .B2(
        \xmem_data[107][5] ), .ZN(n12758) );
  AOI22_X1 U16898 ( .A1(n31316), .A2(\xmem_data[108][5] ), .B1(n27463), .B2(
        \xmem_data[109][5] ), .ZN(n12757) );
  AOI22_X1 U16899 ( .A1(n13420), .A2(\xmem_data[110][5] ), .B1(n17050), .B2(
        \xmem_data[111][5] ), .ZN(n12756) );
  AOI22_X1 U16900 ( .A1(n27564), .A2(\xmem_data[112][5] ), .B1(n30908), .B2(
        \xmem_data[113][5] ), .ZN(n12763) );
  AOI22_X1 U16901 ( .A1(n16980), .A2(\xmem_data[114][5] ), .B1(n16979), .B2(
        \xmem_data[115][5] ), .ZN(n12762) );
  AOI22_X1 U16902 ( .A1(n21066), .A2(\xmem_data[116][5] ), .B1(n3218), .B2(
        \xmem_data[117][5] ), .ZN(n12761) );
  AOI22_X1 U16903 ( .A1(n17033), .A2(\xmem_data[118][5] ), .B1(n27507), .B2(
        \xmem_data[119][5] ), .ZN(n12760) );
  AOI22_X1 U16904 ( .A1(n24534), .A2(\xmem_data[120][5] ), .B1(n17061), .B2(
        \xmem_data[121][5] ), .ZN(n12767) );
  AOI22_X1 U16905 ( .A1(n16973), .A2(\xmem_data[122][5] ), .B1(n16972), .B2(
        \xmem_data[123][5] ), .ZN(n12766) );
  AOI22_X1 U16906 ( .A1(n16974), .A2(\xmem_data[124][5] ), .B1(n29180), .B2(
        \xmem_data[125][5] ), .ZN(n12765) );
  AOI22_X1 U16907 ( .A1(n25708), .A2(\xmem_data[126][5] ), .B1(n24448), .B2(
        \xmem_data[127][5] ), .ZN(n12764) );
  AOI22_X1 U16908 ( .A1(n31268), .A2(\xmem_data[64][5] ), .B1(n23715), .B2(
        \xmem_data[65][5] ), .ZN(n12771) );
  AOI22_X1 U16909 ( .A1(n30543), .A2(\xmem_data[66][5] ), .B1(n17019), .B2(
        \xmem_data[67][5] ), .ZN(n12770) );
  AOI22_X1 U16910 ( .A1(n17020), .A2(\xmem_data[68][5] ), .B1(n24219), .B2(
        \xmem_data[69][5] ), .ZN(n12769) );
  AOI22_X1 U16911 ( .A1(n17021), .A2(\xmem_data[70][5] ), .B1(n29238), .B2(
        \xmem_data[71][5] ), .ZN(n12768) );
  AOI22_X1 U16912 ( .A1(n25717), .A2(\xmem_data[72][5] ), .B1(n17001), .B2(
        \xmem_data[73][5] ), .ZN(n12775) );
  AOI22_X1 U16913 ( .A1(n17004), .A2(\xmem_data[74][5] ), .B1(n3200), .B2(
        \xmem_data[75][5] ), .ZN(n12774) );
  AOI22_X1 U16914 ( .A1(n20818), .A2(\xmem_data[76][5] ), .B1(n17003), .B2(
        \xmem_data[77][5] ), .ZN(n12773) );
  AOI22_X1 U16915 ( .A1(n13420), .A2(\xmem_data[78][5] ), .B1(n16999), .B2(
        \xmem_data[79][5] ), .ZN(n12772) );
  AOI22_X1 U16916 ( .A1(n17030), .A2(\xmem_data[80][5] ), .B1(n22752), .B2(
        \xmem_data[81][5] ), .ZN(n12779) );
  AOI22_X1 U16917 ( .A1(n3388), .A2(\xmem_data[82][5] ), .B1(n17031), .B2(
        \xmem_data[83][5] ), .ZN(n12778) );
  AOI22_X1 U16918 ( .A1(n29064), .A2(\xmem_data[84][5] ), .B1(n3218), .B2(
        \xmem_data[85][5] ), .ZN(n12777) );
  AOI22_X1 U16919 ( .A1(n17033), .A2(\xmem_data[86][5] ), .B1(n28356), .B2(
        \xmem_data[87][5] ), .ZN(n12776) );
  AOI22_X1 U16920 ( .A1(n17010), .A2(\xmem_data[88][5] ), .B1(n24564), .B2(
        \xmem_data[89][5] ), .ZN(n12783) );
  AOI22_X1 U16921 ( .A1(n28952), .A2(\xmem_data[90][5] ), .B1(n17011), .B2(
        \xmem_data[91][5] ), .ZN(n12782) );
  AOI22_X1 U16922 ( .A1(n23813), .A2(\xmem_data[92][5] ), .B1(n13475), .B2(
        \xmem_data[93][5] ), .ZN(n12781) );
  AOI22_X1 U16923 ( .A1(n17013), .A2(\xmem_data[94][5] ), .B1(n17012), .B2(
        \xmem_data[95][5] ), .ZN(n12780) );
  AOI22_X1 U16924 ( .A1(n16997), .A2(n12785), .B1(n16966), .B2(n12784), .ZN(
        n12808) );
  AOI22_X1 U16925 ( .A1(n27537), .A2(\xmem_data[32][5] ), .B1(n30613), .B2(
        \xmem_data[33][5] ), .ZN(n12789) );
  AOI22_X1 U16926 ( .A1(n30892), .A2(\xmem_data[34][5] ), .B1(n16987), .B2(
        \xmem_data[35][5] ), .ZN(n12788) );
  AOI22_X1 U16927 ( .A1(n17020), .A2(\xmem_data[36][5] ), .B1(n27918), .B2(
        \xmem_data[37][5] ), .ZN(n12787) );
  AOI22_X1 U16928 ( .A1(n17021), .A2(\xmem_data[38][5] ), .B1(n29238), .B2(
        \xmem_data[39][5] ), .ZN(n12786) );
  NAND4_X1 U16929 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12805) );
  AOI22_X1 U16930 ( .A1(n3326), .A2(\xmem_data[40][5] ), .B1(n17001), .B2(
        \xmem_data[41][5] ), .ZN(n12793) );
  AOI22_X1 U16931 ( .A1(n17004), .A2(\xmem_data[42][5] ), .B1(n3201), .B2(
        \xmem_data[43][5] ), .ZN(n12792) );
  AOI22_X1 U16932 ( .A1(n24606), .A2(\xmem_data[44][5] ), .B1(n17003), .B2(
        \xmem_data[45][5] ), .ZN(n12791) );
  AOI22_X1 U16933 ( .A1(n30901), .A2(\xmem_data[46][5] ), .B1(n16999), .B2(
        \xmem_data[47][5] ), .ZN(n12790) );
  NAND4_X1 U16934 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12804) );
  AOI22_X1 U16935 ( .A1(n17030), .A2(\xmem_data[48][5] ), .B1(n30571), .B2(
        \xmem_data[49][5] ), .ZN(n12797) );
  AOI22_X1 U16936 ( .A1(n3388), .A2(\xmem_data[50][5] ), .B1(n17031), .B2(
        \xmem_data[51][5] ), .ZN(n12796) );
  AOI22_X1 U16937 ( .A1(n28470), .A2(\xmem_data[52][5] ), .B1(n3219), .B2(
        \xmem_data[53][5] ), .ZN(n12795) );
  AOI22_X1 U16938 ( .A1(n17033), .A2(\xmem_data[54][5] ), .B1(n28476), .B2(
        \xmem_data[55][5] ), .ZN(n12794) );
  NAND4_X1 U16939 ( .A1(n12797), .A2(n12796), .A3(n12795), .A4(n12794), .ZN(
        n12803) );
  AOI22_X1 U16940 ( .A1(n17010), .A2(\xmem_data[56][5] ), .B1(n20993), .B2(
        \xmem_data[57][5] ), .ZN(n12801) );
  AOI22_X1 U16941 ( .A1(n3280), .A2(\xmem_data[58][5] ), .B1(n17011), .B2(
        \xmem_data[59][5] ), .ZN(n12800) );
  AOI22_X1 U16942 ( .A1(n27910), .A2(\xmem_data[60][5] ), .B1(n3357), .B2(
        \xmem_data[61][5] ), .ZN(n12799) );
  AOI22_X1 U16943 ( .A1(n17013), .A2(\xmem_data[62][5] ), .B1(n17012), .B2(
        \xmem_data[63][5] ), .ZN(n12798) );
  NAND4_X1 U16944 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12802) );
  OR4_X1 U16945 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12806) );
  NAND2_X1 U16946 ( .A1(n12806), .A2(n17038), .ZN(n12807) );
  OAI22_X1 U16947 ( .A1(n30158), .A2(n35018), .B1(n12809), .B2(n35019), .ZN(
        n26028) );
  XNOR2_X1 U16948 ( .A(n35336), .B(\fmem_data[2][3] ), .ZN(n32015) );
  XOR2_X1 U16949 ( .A(\fmem_data[0][6] ), .B(\fmem_data[0][7] ), .Z(n12811) );
  AOI22_X1 U16950 ( .A1(n3414), .A2(\xmem_data[80][3] ), .B1(n22753), .B2(
        \xmem_data[81][3] ), .ZN(n12816) );
  AND2_X1 U16951 ( .A1(n3221), .A2(\xmem_data[83][3] ), .ZN(n12812) );
  AOI21_X1 U16952 ( .B1(n21066), .B2(\xmem_data[82][3] ), .A(n12812), .ZN(
        n12815) );
  AOI22_X1 U16953 ( .A1(n21067), .A2(\xmem_data[84][3] ), .B1(n25562), .B2(
        \xmem_data[85][3] ), .ZN(n12814) );
  AOI22_X1 U16954 ( .A1(n21069), .A2(\xmem_data[86][3] ), .B1(n21068), .B2(
        \xmem_data[87][3] ), .ZN(n12813) );
  NAND4_X1 U16955 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12832) );
  AOI22_X1 U16956 ( .A1(n21056), .A2(\xmem_data[72][3] ), .B1(n28098), .B2(
        \xmem_data[73][3] ), .ZN(n12820) );
  AOI22_X1 U16957 ( .A1(n21058), .A2(\xmem_data[74][3] ), .B1(n21057), .B2(
        \xmem_data[75][3] ), .ZN(n12819) );
  AOI22_X1 U16958 ( .A1(n21060), .A2(\xmem_data[76][3] ), .B1(n21059), .B2(
        \xmem_data[77][3] ), .ZN(n12818) );
  AOI22_X1 U16959 ( .A1(n21061), .A2(\xmem_data[78][3] ), .B1(n28037), .B2(
        \xmem_data[79][3] ), .ZN(n12817) );
  NAND4_X1 U16960 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        n12831) );
  AOI22_X1 U16961 ( .A1(n21074), .A2(\xmem_data[88][3] ), .B1(n3231), .B2(
        \xmem_data[89][3] ), .ZN(n12824) );
  AOI22_X1 U16962 ( .A1(n25422), .A2(\xmem_data[90][3] ), .B1(n28415), .B2(
        \xmem_data[91][3] ), .ZN(n12823) );
  AOI22_X1 U16963 ( .A1(n20716), .A2(\xmem_data[92][3] ), .B1(n21075), .B2(
        \xmem_data[93][3] ), .ZN(n12822) );
  AOI22_X1 U16964 ( .A1(n30614), .A2(\xmem_data[94][3] ), .B1(n21076), .B2(
        \xmem_data[95][3] ), .ZN(n12821) );
  NAND4_X1 U16965 ( .A1(n12824), .A2(n12823), .A3(n12822), .A4(n12821), .ZN(
        n12830) );
  AOI22_X1 U16966 ( .A1(n21048), .A2(\xmem_data[64][3] ), .B1(n20938), .B2(
        \xmem_data[65][3] ), .ZN(n12828) );
  AOI22_X1 U16967 ( .A1(n24509), .A2(\xmem_data[66][3] ), .B1(n24219), .B2(
        \xmem_data[67][3] ), .ZN(n12827) );
  AOI22_X1 U16968 ( .A1(n21050), .A2(\xmem_data[68][3] ), .B1(n21049), .B2(
        \xmem_data[69][3] ), .ZN(n12826) );
  AOI22_X1 U16969 ( .A1(n28428), .A2(\xmem_data[70][3] ), .B1(n21051), .B2(
        \xmem_data[71][3] ), .ZN(n12825) );
  NAND4_X1 U16970 ( .A1(n12828), .A2(n12827), .A3(n12826), .A4(n12825), .ZN(
        n12829) );
  OR4_X1 U16971 ( .A1(n12832), .A2(n12831), .A3(n12830), .A4(n12829), .ZN(
        n12833) );
  NAND2_X1 U16972 ( .A1(n12833), .A2(n21086), .ZN(n12836) );
  NOR2_X1 U16973 ( .A1(n20386), .A2(n39027), .ZN(n12834) );
  NAND2_X1 U16974 ( .A1(n25492), .A2(n12834), .ZN(n12835) );
  NAND2_X1 U16975 ( .A1(n12836), .A2(n12835), .ZN(n12913) );
  AOI22_X1 U16976 ( .A1(n20950), .A2(\xmem_data[40][3] ), .B1(n20949), .B2(
        \xmem_data[41][3] ), .ZN(n12841) );
  AOI22_X1 U16977 ( .A1(n28293), .A2(\xmem_data[42][3] ), .B1(n17049), .B2(
        \xmem_data[43][3] ), .ZN(n12840) );
  AOI22_X1 U16978 ( .A1(n20952), .A2(\xmem_data[44][3] ), .B1(n20951), .B2(
        \xmem_data[45][3] ), .ZN(n12839) );
  AND2_X1 U16979 ( .A1(n20953), .A2(\xmem_data[46][3] ), .ZN(n12837) );
  AOI21_X1 U16980 ( .B1(n20489), .B2(\xmem_data[47][3] ), .A(n12837), .ZN(
        n12838) );
  NAND4_X1 U16981 ( .A1(n12841), .A2(n12840), .A3(n12839), .A4(n12838), .ZN(
        n12860) );
  AOI22_X1 U16982 ( .A1(n30503), .A2(\xmem_data[50][3] ), .B1(n3222), .B2(
        \xmem_data[51][3] ), .ZN(n12848) );
  AOI22_X1 U16983 ( .A1(n20969), .A2(\xmem_data[54][3] ), .B1(n23811), .B2(
        \xmem_data[55][3] ), .ZN(n12842) );
  INV_X1 U16984 ( .A(n12842), .ZN(n12846) );
  AOI22_X1 U16985 ( .A1(n29288), .A2(\xmem_data[52][3] ), .B1(n14925), .B2(
        \xmem_data[53][3] ), .ZN(n12844) );
  AOI22_X1 U16986 ( .A1(n3335), .A2(\xmem_data[48][3] ), .B1(n14875), .B2(
        \xmem_data[49][3] ), .ZN(n12843) );
  NAND2_X1 U16987 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NOR2_X1 U16988 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  NAND2_X1 U16989 ( .A1(n12848), .A2(n12847), .ZN(n12859) );
  AOI22_X1 U16990 ( .A1(n20962), .A2(\xmem_data[56][3] ), .B1(n3231), .B2(
        \xmem_data[57][3] ), .ZN(n12852) );
  AOI22_X1 U16991 ( .A1(n20961), .A2(\xmem_data[58][3] ), .B1(n27943), .B2(
        \xmem_data[59][3] ), .ZN(n12851) );
  AOI22_X1 U16992 ( .A1(n25457), .A2(\xmem_data[60][3] ), .B1(n20958), .B2(
        \xmem_data[61][3] ), .ZN(n12850) );
  AOI22_X1 U16993 ( .A1(n20959), .A2(\xmem_data[62][3] ), .B1(n29271), .B2(
        \xmem_data[63][3] ), .ZN(n12849) );
  NAND4_X1 U16994 ( .A1(n12852), .A2(n12851), .A3(n12850), .A4(n12849), .ZN(
        n12858) );
  AOI22_X1 U16995 ( .A1(n20939), .A2(\xmem_data[32][3] ), .B1(n20938), .B2(
        \xmem_data[33][3] ), .ZN(n12856) );
  AOI22_X1 U16996 ( .A1(n20800), .A2(\xmem_data[34][3] ), .B1(n20940), .B2(
        \xmem_data[35][3] ), .ZN(n12855) );
  AOI22_X1 U16997 ( .A1(n20942), .A2(\xmem_data[36][3] ), .B1(n20941), .B2(
        \xmem_data[37][3] ), .ZN(n12854) );
  AOI22_X1 U16998 ( .A1(n28385), .A2(\xmem_data[38][3] ), .B1(n20943), .B2(
        \xmem_data[39][3] ), .ZN(n12853) );
  NAND4_X1 U16999 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  AND2_X1 U17000 ( .A1(n12861), .A2(n20311), .ZN(n12912) );
  AOI22_X1 U17001 ( .A1(n21048), .A2(\xmem_data[96][3] ), .B1(n3213), .B2(
        \xmem_data[97][3] ), .ZN(n12865) );
  AOI22_X1 U17002 ( .A1(n24509), .A2(\xmem_data[98][3] ), .B1(n31329), .B2(
        \xmem_data[99][3] ), .ZN(n12864) );
  AOI22_X1 U17003 ( .A1(n21050), .A2(\xmem_data[100][3] ), .B1(n21049), .B2(
        \xmem_data[101][3] ), .ZN(n12863) );
  AOI22_X1 U17004 ( .A1(n28061), .A2(\xmem_data[102][3] ), .B1(n25581), .B2(
        \xmem_data[103][3] ), .ZN(n12862) );
  NAND4_X1 U17005 ( .A1(n12865), .A2(n12864), .A3(n12863), .A4(n12862), .ZN(
        n12881) );
  AOI22_X1 U17006 ( .A1(n21056), .A2(\xmem_data[104][3] ), .B1(n28098), .B2(
        \xmem_data[105][3] ), .ZN(n12869) );
  AOI22_X1 U17007 ( .A1(n21058), .A2(\xmem_data[106][3] ), .B1(n21057), .B2(
        \xmem_data[107][3] ), .ZN(n12868) );
  AOI22_X1 U17008 ( .A1(n21060), .A2(\xmem_data[108][3] ), .B1(n21059), .B2(
        \xmem_data[109][3] ), .ZN(n12867) );
  AOI22_X1 U17009 ( .A1(n21061), .A2(\xmem_data[110][3] ), .B1(n31309), .B2(
        \xmem_data[111][3] ), .ZN(n12866) );
  NAND4_X1 U17010 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12880) );
  AOI22_X1 U17011 ( .A1(n25624), .A2(\xmem_data[112][3] ), .B1(n31347), .B2(
        \xmem_data[113][3] ), .ZN(n12873) );
  AOI22_X1 U17012 ( .A1(n21066), .A2(\xmem_data[114][3] ), .B1(n3220), .B2(
        \xmem_data[115][3] ), .ZN(n12872) );
  AOI22_X1 U17013 ( .A1(n21067), .A2(\xmem_data[116][3] ), .B1(n30534), .B2(
        \xmem_data[117][3] ), .ZN(n12871) );
  AOI22_X1 U17014 ( .A1(n21069), .A2(\xmem_data[118][3] ), .B1(n21068), .B2(
        \xmem_data[119][3] ), .ZN(n12870) );
  NAND4_X1 U17015 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n12870), .ZN(
        n12879) );
  AOI22_X1 U17016 ( .A1(n21074), .A2(\xmem_data[120][3] ), .B1(n24553), .B2(
        \xmem_data[121][3] ), .ZN(n12877) );
  AOI22_X1 U17017 ( .A1(n28374), .A2(\xmem_data[122][3] ), .B1(n20546), .B2(
        \xmem_data[123][3] ), .ZN(n12876) );
  AOI22_X1 U17018 ( .A1(n17064), .A2(\xmem_data[124][3] ), .B1(n21075), .B2(
        \xmem_data[125][3] ), .ZN(n12875) );
  AOI22_X1 U17019 ( .A1(n13436), .A2(\xmem_data[126][3] ), .B1(n21076), .B2(
        \xmem_data[127][3] ), .ZN(n12874) );
  NAND4_X1 U17020 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        n12878) );
  OR4_X1 U17021 ( .A1(n12881), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12882) );
  AND2_X1 U17022 ( .A1(n12882), .A2(n21088), .ZN(n12911) );
  AOI22_X1 U17023 ( .A1(n3149), .A2(\xmem_data[16][3] ), .B1(n23731), .B2(
        \xmem_data[17][3] ), .ZN(n12887) );
  AND2_X1 U17024 ( .A1(n3222), .A2(\xmem_data[19][3] ), .ZN(n12883) );
  AOI21_X1 U17025 ( .B1(n20991), .B2(\xmem_data[18][3] ), .A(n12883), .ZN(
        n12886) );
  AOI22_X1 U17026 ( .A1(n27831), .A2(\xmem_data[20][3] ), .B1(n20992), .B2(
        \xmem_data[21][3] ), .ZN(n12885) );
  AOI22_X1 U17027 ( .A1(n20994), .A2(\xmem_data[22][3] ), .B1(n20993), .B2(
        \xmem_data[23][3] ), .ZN(n12884) );
  NAND4_X1 U17028 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12896) );
  AOI22_X1 U17029 ( .A1(n29451), .A2(\xmem_data[28][3] ), .B1(n21015), .B2(
        \xmem_data[29][3] ), .ZN(n12894) );
  AOI22_X1 U17030 ( .A1(n29272), .A2(\xmem_data[30][3] ), .B1(n22703), .B2(
        \xmem_data[31][3] ), .ZN(n12888) );
  INV_X1 U17031 ( .A(n12888), .ZN(n12892) );
  AOI22_X1 U17032 ( .A1(n23813), .A2(\xmem_data[26][3] ), .B1(n20982), .B2(
        \xmem_data[27][3] ), .ZN(n12890) );
  NAND2_X1 U17033 ( .A1(n27396), .A2(\xmem_data[24][3] ), .ZN(n12889) );
  NAND2_X1 U17034 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  NOR2_X1 U17035 ( .A1(n12892), .A2(n12891), .ZN(n12893) );
  NAND2_X1 U17036 ( .A1(n12894), .A2(n12893), .ZN(n12895) );
  OR2_X1 U17037 ( .A1(n12896), .A2(n12895), .ZN(n12908) );
  AOI22_X1 U17038 ( .A1(n21005), .A2(\xmem_data[0][3] ), .B1(n25460), .B2(
        \xmem_data[1][3] ), .ZN(n12900) );
  AOI22_X1 U17039 ( .A1(n21007), .A2(\xmem_data[2][3] ), .B1(n21006), .B2(
        \xmem_data[3][3] ), .ZN(n12899) );
  AOI22_X1 U17040 ( .A1(n21008), .A2(\xmem_data[4][3] ), .B1(n29318), .B2(
        \xmem_data[5][3] ), .ZN(n12898) );
  AOI22_X1 U17041 ( .A1(n21010), .A2(\xmem_data[6][3] ), .B1(n30598), .B2(
        \xmem_data[7][3] ), .ZN(n12897) );
  NAND4_X1 U17042 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12906) );
  AOI22_X1 U17043 ( .A1(n20984), .A2(\xmem_data[8][3] ), .B1(n20983), .B2(
        \xmem_data[9][3] ), .ZN(n12904) );
  AOI22_X1 U17044 ( .A1(n28293), .A2(\xmem_data[10][3] ), .B1(n20488), .B2(
        \xmem_data[11][3] ), .ZN(n12903) );
  AOI22_X1 U17045 ( .A1(n20985), .A2(\xmem_data[12][3] ), .B1(n24524), .B2(
        \xmem_data[13][3] ), .ZN(n12902) );
  AOI22_X1 U17046 ( .A1(n20986), .A2(\xmem_data[14][3] ), .B1(n25357), .B2(
        \xmem_data[15][3] ), .ZN(n12901) );
  NAND4_X1 U17047 ( .A1(n12904), .A2(n12903), .A3(n12902), .A4(n12901), .ZN(
        n12905) );
  OR2_X1 U17048 ( .A1(n12906), .A2(n12905), .ZN(n12907) );
  NOR2_X1 U17049 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  NOR2_X1 U17050 ( .A1(n12909), .A2(n20386), .ZN(n12910) );
  OR4_X2 U17051 ( .A1(n12913), .A2(n12912), .A3(n12911), .A4(n12910), .ZN(
        n32064) );
  XNOR2_X1 U17052 ( .A(n32064), .B(\fmem_data[0][7] ), .ZN(n30448) );
  OAI22_X1 U17053 ( .A1(n35493), .A2(n30448), .B1(n31641), .B2(n35494), .ZN(
        n26027) );
  AOI22_X1 U17054 ( .A1(n23730), .A2(\xmem_data[112][5] ), .B1(n24468), .B2(
        \xmem_data[113][5] ), .ZN(n12918) );
  AOI22_X1 U17055 ( .A1(n21061), .A2(\xmem_data[114][5] ), .B1(n28947), .B2(
        \xmem_data[115][5] ), .ZN(n12917) );
  AOI22_X1 U17056 ( .A1(n23732), .A2(\xmem_data[116][5] ), .B1(n23731), .B2(
        \xmem_data[117][5] ), .ZN(n12916) );
  AND2_X1 U17057 ( .A1(n3222), .A2(\xmem_data[119][5] ), .ZN(n12914) );
  AOI21_X1 U17058 ( .B1(n23734), .B2(\xmem_data[118][5] ), .A(n12914), .ZN(
        n12915) );
  NAND4_X1 U17059 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12935) );
  AOI22_X1 U17060 ( .A1(n23722), .A2(\xmem_data[104][5] ), .B1(n24460), .B2(
        \xmem_data[105][5] ), .ZN(n12922) );
  AOI22_X1 U17061 ( .A1(n24511), .A2(\xmem_data[106][5] ), .B1(n31361), .B2(
        \xmem_data[107][5] ), .ZN(n12921) );
  AOI22_X1 U17062 ( .A1(n23724), .A2(\xmem_data[108][5] ), .B1(n23723), .B2(
        \xmem_data[109][5] ), .ZN(n12920) );
  AOI22_X1 U17063 ( .A1(n20782), .A2(\xmem_data[110][5] ), .B1(n23725), .B2(
        \xmem_data[111][5] ), .ZN(n12919) );
  NAND4_X1 U17064 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12933) );
  AOI22_X1 U17065 ( .A1(n23740), .A2(\xmem_data[120][5] ), .B1(n23739), .B2(
        \xmem_data[121][5] ), .ZN(n12926) );
  AOI22_X1 U17066 ( .A1(n23741), .A2(\xmem_data[122][5] ), .B1(n27994), .B2(
        \xmem_data[123][5] ), .ZN(n12925) );
  AOI22_X1 U17067 ( .A1(n23742), .A2(\xmem_data[124][5] ), .B1(n25492), .B2(
        \xmem_data[125][5] ), .ZN(n12924) );
  AOI22_X1 U17068 ( .A1(n27447), .A2(\xmem_data[126][5] ), .B1(n13475), .B2(
        \xmem_data[127][5] ), .ZN(n12923) );
  NAND4_X1 U17069 ( .A1(n12926), .A2(n12925), .A3(n12924), .A4(n12923), .ZN(
        n12932) );
  AOI22_X1 U17070 ( .A1(n30744), .A2(\xmem_data[96][5] ), .B1(n24212), .B2(
        \xmem_data[97][5] ), .ZN(n12930) );
  AOI22_X1 U17071 ( .A1(n30614), .A2(\xmem_data[98][5] ), .B1(n23715), .B2(
        \xmem_data[99][5] ), .ZN(n12929) );
  AOI22_X1 U17072 ( .A1(n29008), .A2(\xmem_data[100][5] ), .B1(n23716), .B2(
        \xmem_data[101][5] ), .ZN(n12928) );
  AOI22_X1 U17073 ( .A1(n23717), .A2(\xmem_data[102][5] ), .B1(n25677), .B2(
        \xmem_data[103][5] ), .ZN(n12927) );
  NAND4_X1 U17074 ( .A1(n12930), .A2(n12929), .A3(n12928), .A4(n12927), .ZN(
        n12931) );
  OR3_X1 U17075 ( .A1(n12933), .A2(n12932), .A3(n12931), .ZN(n12934) );
  OAI21_X1 U17076 ( .B1(n12935), .B2(n12934), .A(n23751), .ZN(n12959) );
  AOI22_X1 U17077 ( .A1(n23753), .A2(\xmem_data[80][5] ), .B1(n20707), .B2(
        \xmem_data[81][5] ), .ZN(n12940) );
  AOI22_X1 U17078 ( .A1(n25441), .A2(\xmem_data[82][5] ), .B1(n28317), .B2(
        \xmem_data[83][5] ), .ZN(n12939) );
  AOI22_X1 U17079 ( .A1(n23754), .A2(\xmem_data[84][5] ), .B1(n27437), .B2(
        \xmem_data[85][5] ), .ZN(n12938) );
  AND2_X1 U17080 ( .A1(n3218), .A2(\xmem_data[87][5] ), .ZN(n12936) );
  AOI21_X1 U17081 ( .B1(n23756), .B2(\xmem_data[86][5] ), .A(n12936), .ZN(
        n12937) );
  NAND4_X1 U17082 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12957) );
  AOI22_X1 U17083 ( .A1(n23777), .A2(\xmem_data[72][5] ), .B1(n23776), .B2(
        \xmem_data[73][5] ), .ZN(n12944) );
  AOI22_X1 U17084 ( .A1(n3205), .A2(\xmem_data[74][5] ), .B1(n23778), .B2(
        \xmem_data[75][5] ), .ZN(n12943) );
  AOI22_X1 U17085 ( .A1(n23780), .A2(\xmem_data[76][5] ), .B1(n23779), .B2(
        \xmem_data[77][5] ), .ZN(n12942) );
  AOI22_X1 U17086 ( .A1(n20734), .A2(\xmem_data[78][5] ), .B1(n23781), .B2(
        \xmem_data[79][5] ), .ZN(n12941) );
  NAND4_X1 U17087 ( .A1(n12944), .A2(n12943), .A3(n12942), .A4(n12941), .ZN(
        n12955) );
  AOI22_X1 U17088 ( .A1(n23770), .A2(\xmem_data[88][5] ), .B1(n23769), .B2(
        \xmem_data[89][5] ), .ZN(n12948) );
  AOI22_X1 U17089 ( .A1(n23812), .A2(\xmem_data[90][5] ), .B1(n25486), .B2(
        \xmem_data[91][5] ), .ZN(n12947) );
  AOI22_X1 U17090 ( .A1(n3280), .A2(\xmem_data[92][5] ), .B1(n3231), .B2(
        \xmem_data[93][5] ), .ZN(n12946) );
  AOI22_X1 U17091 ( .A1(n27447), .A2(\xmem_data[94][5] ), .B1(n3357), .B2(
        \xmem_data[95][5] ), .ZN(n12945) );
  NAND4_X1 U17092 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12954) );
  AOI22_X1 U17093 ( .A1(n23762), .A2(\xmem_data[64][5] ), .B1(n23761), .B2(
        \xmem_data[65][5] ), .ZN(n12952) );
  AOI22_X1 U17094 ( .A1(n23763), .A2(\xmem_data[66][5] ), .B1(n22703), .B2(
        \xmem_data[67][5] ), .ZN(n12951) );
  AOI22_X1 U17095 ( .A1(n29315), .A2(\xmem_data[68][5] ), .B1(n15000), .B2(
        \xmem_data[69][5] ), .ZN(n12950) );
  AOI22_X1 U17096 ( .A1(n23764), .A2(\xmem_data[70][5] ), .B1(n14970), .B2(
        \xmem_data[71][5] ), .ZN(n12949) );
  NAND4_X1 U17097 ( .A1(n12952), .A2(n12951), .A3(n12950), .A4(n12949), .ZN(
        n12953) );
  NAND2_X1 U17098 ( .A1(n12959), .A2(n12958), .ZN(n13014) );
  AOI22_X1 U17099 ( .A1(n23762), .A2(\xmem_data[32][5] ), .B1(n23761), .B2(
        \xmem_data[33][5] ), .ZN(n12963) );
  AOI22_X1 U17100 ( .A1(n23763), .A2(\xmem_data[34][5] ), .B1(n22674), .B2(
        \xmem_data[35][5] ), .ZN(n12962) );
  AOI22_X1 U17101 ( .A1(n29437), .A2(\xmem_data[36][5] ), .B1(n25383), .B2(
        \xmem_data[37][5] ), .ZN(n12961) );
  AOI22_X1 U17102 ( .A1(n23764), .A2(\xmem_data[38][5] ), .B1(n22718), .B2(
        \xmem_data[39][5] ), .ZN(n12960) );
  NAND4_X1 U17103 ( .A1(n12963), .A2(n12962), .A3(n12961), .A4(n12960), .ZN(
        n12979) );
  AOI22_X1 U17104 ( .A1(n23777), .A2(\xmem_data[40][5] ), .B1(n23776), .B2(
        \xmem_data[41][5] ), .ZN(n12967) );
  AOI22_X1 U17105 ( .A1(n28061), .A2(\xmem_data[42][5] ), .B1(n23778), .B2(
        \xmem_data[43][5] ), .ZN(n12966) );
  AOI22_X1 U17106 ( .A1(n23780), .A2(\xmem_data[44][5] ), .B1(n23779), .B2(
        \xmem_data[45][5] ), .ZN(n12965) );
  AOI22_X1 U17107 ( .A1(n24467), .A2(\xmem_data[46][5] ), .B1(n23781), .B2(
        \xmem_data[47][5] ), .ZN(n12964) );
  NAND4_X1 U17108 ( .A1(n12967), .A2(n12966), .A3(n12965), .A4(n12964), .ZN(
        n12978) );
  AOI22_X1 U17109 ( .A1(n23753), .A2(\xmem_data[48][5] ), .B1(n30524), .B2(
        \xmem_data[49][5] ), .ZN(n12971) );
  AOI22_X1 U17110 ( .A1(n3380), .A2(\xmem_data[50][5] ), .B1(n24525), .B2(
        \xmem_data[51][5] ), .ZN(n12970) );
  AOI22_X1 U17111 ( .A1(n23754), .A2(\xmem_data[52][5] ), .B1(n28501), .B2(
        \xmem_data[53][5] ), .ZN(n12969) );
  AOI22_X1 U17112 ( .A1(n23756), .A2(\xmem_data[54][5] ), .B1(n3222), .B2(
        \xmem_data[55][5] ), .ZN(n12968) );
  NAND4_X1 U17113 ( .A1(n12971), .A2(n12970), .A3(n12969), .A4(n12968), .ZN(
        n12977) );
  AOI22_X1 U17114 ( .A1(n23770), .A2(\xmem_data[56][5] ), .B1(n23769), .B2(
        \xmem_data[57][5] ), .ZN(n12975) );
  AOI22_X1 U17115 ( .A1(n24697), .A2(\xmem_data[58][5] ), .B1(n31275), .B2(
        \xmem_data[59][5] ), .ZN(n12974) );
  AOI22_X1 U17116 ( .A1(n3280), .A2(\xmem_data[60][5] ), .B1(n3231), .B2(
        \xmem_data[61][5] ), .ZN(n12973) );
  AOI22_X1 U17117 ( .A1(n27447), .A2(\xmem_data[62][5] ), .B1(n20982), .B2(
        \xmem_data[63][5] ), .ZN(n12972) );
  NAND4_X1 U17118 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12976) );
  OR4_X1 U17119 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12980) );
  AND2_X1 U17120 ( .A1(n12980), .A2(n23790), .ZN(n13013) );
  AOI22_X1 U17121 ( .A1(n29065), .A2(\xmem_data[24][5] ), .B1(n30534), .B2(
        \xmem_data[25][5] ), .ZN(n12981) );
  AOI22_X1 U17122 ( .A1(n23813), .A2(\xmem_data[30][5] ), .B1(n13475), .B2(
        \xmem_data[31][5] ), .ZN(n12983) );
  NAND2_X1 U17123 ( .A1(n3280), .A2(\xmem_data[28][5] ), .ZN(n12982) );
  NAND2_X1 U17124 ( .A1(n12983), .A2(n12982), .ZN(n12986) );
  AOI22_X1 U17125 ( .A1(n23812), .A2(\xmem_data[26][5] ), .B1(n23811), .B2(
        \xmem_data[27][5] ), .ZN(n12984) );
  INV_X1 U17126 ( .A(n12984), .ZN(n12985) );
  OR3_X1 U17127 ( .A1(n12987), .A2(n12986), .A3(n12985), .ZN(n12993) );
  AOI22_X1 U17128 ( .A1(n23792), .A2(\xmem_data[0][5] ), .B1(n24212), .B2(
        \xmem_data[1][5] ), .ZN(n12991) );
  AOI22_X1 U17129 ( .A1(n29310), .A2(\xmem_data[2][5] ), .B1(n23793), .B2(
        \xmem_data[3][5] ), .ZN(n12990) );
  AOI22_X1 U17130 ( .A1(n30543), .A2(\xmem_data[4][5] ), .B1(n3208), .B2(
        \xmem_data[5][5] ), .ZN(n12989) );
  AOI22_X1 U17131 ( .A1(n23717), .A2(\xmem_data[6][5] ), .B1(n23796), .B2(
        \xmem_data[7][5] ), .ZN(n12988) );
  NAND4_X1 U17132 ( .A1(n12991), .A2(n12990), .A3(n12989), .A4(n12988), .ZN(
        n12992) );
  OR2_X1 U17133 ( .A1(n12993), .A2(n12992), .ZN(n13009) );
  AND2_X1 U17134 ( .A1(n29124), .A2(\xmem_data[18][5] ), .ZN(n12995) );
  AND2_X1 U17135 ( .A1(n3219), .A2(\xmem_data[23][5] ), .ZN(n12994) );
  NOR2_X1 U17136 ( .A1(n12995), .A2(n12994), .ZN(n12998) );
  NAND2_X1 U17137 ( .A1(n20769), .A2(\xmem_data[17][5] ), .ZN(n12997) );
  AOI22_X1 U17138 ( .A1(n30864), .A2(\xmem_data[20][5] ), .B1(n25360), .B2(
        \xmem_data[21][5] ), .ZN(n12996) );
  NOR2_X1 U17139 ( .A1(n13000), .A2(n12999), .ZN(n13007) );
  AOI22_X1 U17140 ( .A1(n23802), .A2(\xmem_data[8][5] ), .B1(n23801), .B2(
        \xmem_data[9][5] ), .ZN(n13004) );
  AOI22_X1 U17141 ( .A1(n3205), .A2(\xmem_data[10][5] ), .B1(n30898), .B2(
        \xmem_data[11][5] ), .ZN(n13003) );
  AOI22_X1 U17142 ( .A1(n28955), .A2(\xmem_data[12][5] ), .B1(n23723), .B2(
        \xmem_data[13][5] ), .ZN(n13002) );
  AOI22_X1 U17143 ( .A1(n24685), .A2(\xmem_data[14][5] ), .B1(n17049), .B2(
        \xmem_data[15][5] ), .ZN(n13001) );
  NAND2_X1 U17144 ( .A1(n20708), .A2(\xmem_data[16][5] ), .ZN(n13006) );
  NAND2_X1 U17145 ( .A1(n24562), .A2(\xmem_data[22][5] ), .ZN(n13005) );
  NAND4_X1 U17146 ( .A1(n13007), .A2(n3811), .A3(n13006), .A4(n13005), .ZN(
        n13008) );
  NOR2_X1 U17147 ( .A1(n13009), .A2(n13008), .ZN(n13011) );
  NAND2_X1 U17148 ( .A1(n28307), .A2(\xmem_data[29][5] ), .ZN(n13010) );
  AOI21_X1 U17149 ( .B1(n13011), .B2(n13010), .A(n22877), .ZN(n13012) );
  AOI22_X1 U17150 ( .A1(n23802), .A2(\xmem_data[8][6] ), .B1(n23801), .B2(
        \xmem_data[9][6] ), .ZN(n13019) );
  AOI22_X1 U17151 ( .A1(n3177), .A2(\xmem_data[10][6] ), .B1(n30598), .B2(
        \xmem_data[11][6] ), .ZN(n13018) );
  AOI22_X1 U17152 ( .A1(n23780), .A2(\xmem_data[12][6] ), .B1(n30599), .B2(
        \xmem_data[13][6] ), .ZN(n13017) );
  AOI22_X1 U17153 ( .A1(n30497), .A2(\xmem_data[14][6] ), .B1(n31256), .B2(
        \xmem_data[15][6] ), .ZN(n13016) );
  NAND4_X1 U17154 ( .A1(n13019), .A2(n13018), .A3(n13017), .A4(n13016), .ZN(
        n13039) );
  AOI22_X1 U17155 ( .A1(n29725), .A2(\xmem_data[16][6] ), .B1(n17050), .B2(
        \xmem_data[17][6] ), .ZN(n13023) );
  AOI22_X1 U17156 ( .A1(n27500), .A2(\xmem_data[18][6] ), .B1(n21309), .B2(
        \xmem_data[19][6] ), .ZN(n13022) );
  AOI22_X1 U17157 ( .A1(n3350), .A2(\xmem_data[20][6] ), .B1(n28501), .B2(
        \xmem_data[21][6] ), .ZN(n13021) );
  AOI22_X1 U17158 ( .A1(n20576), .A2(\xmem_data[22][6] ), .B1(n3218), .B2(
        \xmem_data[23][6] ), .ZN(n13020) );
  NAND4_X1 U17159 ( .A1(n13023), .A2(n13022), .A3(n13021), .A4(n13020), .ZN(
        n13038) );
  AOI22_X1 U17160 ( .A1(n23792), .A2(\xmem_data[0][6] ), .B1(n14998), .B2(
        \xmem_data[1][6] ), .ZN(n13027) );
  AOI22_X1 U17161 ( .A1(n28980), .A2(\xmem_data[2][6] ), .B1(n23793), .B2(
        \xmem_data[3][6] ), .ZN(n13026) );
  AOI22_X1 U17162 ( .A1(n27945), .A2(\xmem_data[4][6] ), .B1(n3207), .B2(
        \xmem_data[5][6] ), .ZN(n13025) );
  AOI22_X1 U17163 ( .A1(n21007), .A2(\xmem_data[6][6] ), .B1(n23796), .B2(
        \xmem_data[7][6] ), .ZN(n13024) );
  NAND4_X1 U17164 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n13037) );
  AOI22_X1 U17165 ( .A1(n23812), .A2(\xmem_data[26][6] ), .B1(n23811), .B2(
        \xmem_data[27][6] ), .ZN(n13035) );
  AOI22_X1 U17166 ( .A1(n24139), .A2(\xmem_data[24][6] ), .B1(n27869), .B2(
        \xmem_data[25][6] ), .ZN(n13028) );
  INV_X1 U17167 ( .A(n13028), .ZN(n13033) );
  AND2_X1 U17168 ( .A1(n3280), .A2(\xmem_data[28][6] ), .ZN(n13032) );
  NAND2_X1 U17169 ( .A1(n13475), .A2(\xmem_data[31][6] ), .ZN(n13030) );
  NAND2_X1 U17170 ( .A1(n23813), .A2(\xmem_data[30][6] ), .ZN(n13029) );
  NAND2_X1 U17171 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  NOR3_X1 U17172 ( .A1(n13033), .A2(n13032), .A3(n13031), .ZN(n13034) );
  NAND2_X1 U17173 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NOR4_X1 U17174 ( .A1(n13039), .A2(n13038), .A3(n13037), .A4(n13036), .ZN(
        n13041) );
  NAND2_X1 U17175 ( .A1(n23771), .A2(\xmem_data[29][6] ), .ZN(n13040) );
  AOI21_X1 U17176 ( .B1(n13041), .B2(n13040), .A(n22877), .ZN(n13042) );
  INV_X1 U17177 ( .A(n13042), .ZN(n13110) );
  AOI22_X1 U17178 ( .A1(n23730), .A2(\xmem_data[112][6] ), .B1(n24122), .B2(
        \xmem_data[113][6] ), .ZN(n13046) );
  AOI22_X1 U17179 ( .A1(n27959), .A2(\xmem_data[114][6] ), .B1(n28037), .B2(
        \xmem_data[115][6] ), .ZN(n13045) );
  AOI22_X1 U17180 ( .A1(n23732), .A2(\xmem_data[116][6] ), .B1(n23731), .B2(
        \xmem_data[117][6] ), .ZN(n13044) );
  AOI22_X1 U17181 ( .A1(n23734), .A2(\xmem_data[118][6] ), .B1(n3221), .B2(
        \xmem_data[119][6] ), .ZN(n13043) );
  NAND4_X1 U17182 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13063) );
  AOI22_X1 U17183 ( .A1(n23722), .A2(\xmem_data[104][6] ), .B1(n24165), .B2(
        \xmem_data[105][6] ), .ZN(n13050) );
  AOI22_X1 U17184 ( .A1(n27952), .A2(\xmem_data[106][6] ), .B1(n27951), .B2(
        \xmem_data[107][6] ), .ZN(n13049) );
  AOI22_X1 U17185 ( .A1(n23724), .A2(\xmem_data[108][6] ), .B1(n23723), .B2(
        \xmem_data[109][6] ), .ZN(n13048) );
  AOI22_X1 U17186 ( .A1(n30497), .A2(\xmem_data[110][6] ), .B1(n23725), .B2(
        \xmem_data[111][6] ), .ZN(n13047) );
  NAND4_X1 U17187 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13061) );
  AOI22_X1 U17188 ( .A1(n23740), .A2(\xmem_data[120][6] ), .B1(n23739), .B2(
        \xmem_data[121][6] ), .ZN(n13054) );
  AOI22_X1 U17189 ( .A1(n23741), .A2(\xmem_data[122][6] ), .B1(n20559), .B2(
        \xmem_data[123][6] ), .ZN(n13053) );
  AOI22_X1 U17190 ( .A1(n23742), .A2(\xmem_data[124][6] ), .B1(n28045), .B2(
        \xmem_data[125][6] ), .ZN(n13052) );
  AOI22_X1 U17191 ( .A1(n27447), .A2(\xmem_data[126][6] ), .B1(n13475), .B2(
        \xmem_data[127][6] ), .ZN(n13051) );
  NAND4_X1 U17192 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13060) );
  AOI22_X1 U17193 ( .A1(n24640), .A2(\xmem_data[96][6] ), .B1(n30552), .B2(
        \xmem_data[97][6] ), .ZN(n13058) );
  AOI22_X1 U17194 ( .A1(n28298), .A2(\xmem_data[98][6] ), .B1(n23715), .B2(
        \xmem_data[99][6] ), .ZN(n13057) );
  AOI22_X1 U17195 ( .A1(n25607), .A2(\xmem_data[100][6] ), .B1(n23716), .B2(
        \xmem_data[101][6] ), .ZN(n13056) );
  AOI22_X1 U17196 ( .A1(n23717), .A2(\xmem_data[102][6] ), .B1(n25715), .B2(
        \xmem_data[103][6] ), .ZN(n13055) );
  NAND4_X1 U17197 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n13055), .ZN(
        n13059) );
  OR3_X1 U17198 ( .A1(n13061), .A2(n13060), .A3(n13059), .ZN(n13062) );
  OAI21_X1 U17199 ( .B1(n13063), .B2(n13062), .A(n23751), .ZN(n13109) );
  AOI22_X1 U17200 ( .A1(n23753), .A2(\xmem_data[48][6] ), .B1(n21059), .B2(
        \xmem_data[49][6] ), .ZN(n13067) );
  AOI22_X1 U17201 ( .A1(n3380), .A2(\xmem_data[50][6] ), .B1(n29118), .B2(
        \xmem_data[51][6] ), .ZN(n13066) );
  AOI22_X1 U17202 ( .A1(n23754), .A2(\xmem_data[52][6] ), .B1(n31347), .B2(
        \xmem_data[53][6] ), .ZN(n13065) );
  AOI22_X1 U17203 ( .A1(n23756), .A2(\xmem_data[54][6] ), .B1(n3218), .B2(
        \xmem_data[55][6] ), .ZN(n13064) );
  NAND4_X1 U17204 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13084) );
  AOI22_X1 U17205 ( .A1(n23777), .A2(\xmem_data[40][6] ), .B1(n23776), .B2(
        \xmem_data[41][6] ), .ZN(n13071) );
  AOI22_X1 U17206 ( .A1(n28385), .A2(\xmem_data[42][6] ), .B1(n23778), .B2(
        \xmem_data[43][6] ), .ZN(n13070) );
  AOI22_X1 U17207 ( .A1(n23780), .A2(\xmem_data[44][6] ), .B1(n23779), .B2(
        \xmem_data[45][6] ), .ZN(n13069) );
  AOI22_X1 U17208 ( .A1(n20818), .A2(\xmem_data[46][6] ), .B1(n23781), .B2(
        \xmem_data[47][6] ), .ZN(n13068) );
  NAND4_X1 U17209 ( .A1(n13071), .A2(n13070), .A3(n13069), .A4(n13068), .ZN(
        n13082) );
  AOI22_X1 U17210 ( .A1(n23770), .A2(\xmem_data[56][6] ), .B1(n23769), .B2(
        \xmem_data[57][6] ), .ZN(n13075) );
  AOI22_X1 U17211 ( .A1(n22666), .A2(\xmem_data[58][6] ), .B1(n22711), .B2(
        \xmem_data[59][6] ), .ZN(n13074) );
  AOI22_X1 U17212 ( .A1(n30698), .A2(\xmem_data[60][6] ), .B1(n31252), .B2(
        \xmem_data[61][6] ), .ZN(n13073) );
  AOI22_X1 U17213 ( .A1(n27447), .A2(\xmem_data[62][6] ), .B1(n24590), .B2(
        \xmem_data[63][6] ), .ZN(n13072) );
  NAND4_X1 U17214 ( .A1(n13075), .A2(n13074), .A3(n13073), .A4(n13072), .ZN(
        n13081) );
  AOI22_X1 U17215 ( .A1(n23762), .A2(\xmem_data[32][6] ), .B1(n23761), .B2(
        \xmem_data[33][6] ), .ZN(n13079) );
  AOI22_X1 U17216 ( .A1(n23763), .A2(\xmem_data[34][6] ), .B1(n27912), .B2(
        \xmem_data[35][6] ), .ZN(n13078) );
  AOI22_X1 U17217 ( .A1(n3466), .A2(\xmem_data[36][6] ), .B1(n20938), .B2(
        \xmem_data[37][6] ), .ZN(n13077) );
  AOI22_X1 U17218 ( .A1(n23764), .A2(\xmem_data[38][6] ), .B1(n25398), .B2(
        \xmem_data[39][6] ), .ZN(n13076) );
  NAND4_X1 U17219 ( .A1(n13079), .A2(n13078), .A3(n13077), .A4(n13076), .ZN(
        n13080) );
  OR3_X1 U17220 ( .A1(n13082), .A2(n13081), .A3(n13080), .ZN(n13083) );
  OAI21_X1 U17221 ( .B1(n13084), .B2(n13083), .A(n23790), .ZN(n13108) );
  AOI22_X1 U17222 ( .A1(n23753), .A2(\xmem_data[80][6] ), .B1(n22727), .B2(
        \xmem_data[81][6] ), .ZN(n13089) );
  AOI22_X1 U17223 ( .A1(n17030), .A2(\xmem_data[82][6] ), .B1(n24470), .B2(
        \xmem_data[83][6] ), .ZN(n13088) );
  AOI22_X1 U17224 ( .A1(n23754), .A2(\xmem_data[84][6] ), .B1(n3247), .B2(
        \xmem_data[85][6] ), .ZN(n13087) );
  AND2_X1 U17225 ( .A1(n3218), .A2(\xmem_data[87][6] ), .ZN(n13085) );
  AOI21_X1 U17226 ( .B1(n23756), .B2(\xmem_data[86][6] ), .A(n13085), .ZN(
        n13086) );
  NAND4_X1 U17227 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13106) );
  AOI22_X1 U17228 ( .A1(n23777), .A2(\xmem_data[72][6] ), .B1(n23776), .B2(
        \xmem_data[73][6] ), .ZN(n13093) );
  AOI22_X1 U17229 ( .A1(n25575), .A2(\xmem_data[74][6] ), .B1(n23778), .B2(
        \xmem_data[75][6] ), .ZN(n13092) );
  AOI22_X1 U17230 ( .A1(n23780), .A2(\xmem_data[76][6] ), .B1(n23779), .B2(
        \xmem_data[77][6] ), .ZN(n13091) );
  AOI22_X1 U17231 ( .A1(n25582), .A2(\xmem_data[78][6] ), .B1(n23781), .B2(
        \xmem_data[79][6] ), .ZN(n13090) );
  NAND4_X1 U17232 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        n13104) );
  AOI22_X1 U17233 ( .A1(n23770), .A2(\xmem_data[88][6] ), .B1(n23769), .B2(
        \xmem_data[89][6] ), .ZN(n13097) );
  AOI22_X1 U17234 ( .A1(n20969), .A2(\xmem_data[90][6] ), .B1(n25616), .B2(
        \xmem_data[91][6] ), .ZN(n13096) );
  AOI22_X1 U17235 ( .A1(n3374), .A2(\xmem_data[92][6] ), .B1(n28045), .B2(
        \xmem_data[93][6] ), .ZN(n13095) );
  AOI22_X1 U17236 ( .A1(n27447), .A2(\xmem_data[94][6] ), .B1(n20546), .B2(
        \xmem_data[95][6] ), .ZN(n13094) );
  NAND4_X1 U17237 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        n13103) );
  AOI22_X1 U17238 ( .A1(n23762), .A2(\xmem_data[64][6] ), .B1(n23761), .B2(
        \xmem_data[65][6] ), .ZN(n13101) );
  AOI22_X1 U17239 ( .A1(n23763), .A2(n20682), .B1(n25458), .B2(
        \xmem_data[67][6] ), .ZN(n13100) );
  AOI22_X1 U17240 ( .A1(n24545), .A2(\xmem_data[68][6] ), .B1(n25574), .B2(
        \xmem_data[69][6] ), .ZN(n13099) );
  AOI22_X1 U17241 ( .A1(n23764), .A2(\xmem_data[70][6] ), .B1(n16989), .B2(
        \xmem_data[71][6] ), .ZN(n13098) );
  NAND4_X1 U17242 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        n13102) );
  OR3_X1 U17243 ( .A1(n13104), .A2(n13103), .A3(n13102), .ZN(n13105) );
  OAI21_X1 U17244 ( .B1(n13106), .B2(n13105), .A(n23713), .ZN(n13107) );
  XNOR2_X1 U17245 ( .A(n33055), .B(\fmem_data[4][5] ), .ZN(n31822) );
  XOR2_X1 U17246 ( .A(\fmem_data[25][2] ), .B(\fmem_data[25][3] ), .Z(n13111)
         );
  AOI22_X1 U17247 ( .A1(n24470), .A2(\xmem_data[104][7] ), .B1(n27813), .B2(
        \xmem_data[105][7] ), .ZN(n13115) );
  BUF_X1 U17248 ( .A(n13468), .Z(n29173) );
  AOI22_X1 U17249 ( .A1(n29173), .A2(\xmem_data[106][7] ), .B1(n20518), .B2(
        \xmem_data[107][7] ), .ZN(n13114) );
  AOI22_X1 U17250 ( .A1(n3220), .A2(\xmem_data[108][7] ), .B1(n29065), .B2(
        \xmem_data[109][7] ), .ZN(n13113) );
  BUF_X1 U17251 ( .A(n14990), .Z(n29174) );
  AOI22_X1 U17252 ( .A1(n20500), .A2(\xmem_data[110][7] ), .B1(n29174), .B2(
        \xmem_data[111][7] ), .ZN(n13112) );
  NAND4_X1 U17253 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        n13126) );
  BUF_X1 U17254 ( .A(n14927), .Z(n29181) );
  BUF_X1 U17255 ( .A(n14991), .Z(n27396) );
  AOI22_X1 U17256 ( .A1(n29181), .A2(\xmem_data[112][7] ), .B1(n27396), .B2(
        \xmem_data[113][7] ), .ZN(n13119) );
  AOI22_X1 U17257 ( .A1(n31252), .A2(\xmem_data[114][7] ), .B1(n28972), .B2(
        \xmem_data[115][7] ), .ZN(n13118) );
  BUF_X1 U17258 ( .A(n14997), .Z(n29179) );
  AOI22_X1 U17259 ( .A1(n29180), .A2(\xmem_data[116][7] ), .B1(n29179), .B2(
        \xmem_data[117][7] ), .ZN(n13117) );
  AOI22_X1 U17260 ( .A1(n22702), .A2(\xmem_data[118][7] ), .B1(n29310), .B2(
        \xmem_data[119][7] ), .ZN(n13116) );
  NAND4_X1 U17261 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13125) );
  AOI22_X1 U17262 ( .A1(n27536), .A2(\xmem_data[120][7] ), .B1(n20776), .B2(
        \xmem_data[121][7] ), .ZN(n13123) );
  BUF_X1 U17263 ( .A(n13188), .Z(n29188) );
  AOI22_X1 U17264 ( .A1(n29188), .A2(\xmem_data[122][7] ), .B1(n24133), .B2(
        \xmem_data[123][7] ), .ZN(n13122) );
  AOI22_X1 U17265 ( .A1(n24459), .A2(\xmem_data[124][7] ), .B1(n30872), .B2(
        \xmem_data[125][7] ), .ZN(n13121) );
  BUF_X1 U17266 ( .A(n14913), .Z(n29190) );
  AOI22_X1 U17267 ( .A1(n29190), .A2(\xmem_data[126][7] ), .B1(n3205), .B2(
        \xmem_data[127][7] ), .ZN(n13120) );
  NAND4_X1 U17268 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13120), .ZN(
        n13124) );
  OR3_X1 U17269 ( .A1(n13126), .A2(n13125), .A3(n13124), .ZN(n13136) );
  AOI22_X1 U17270 ( .A1(n28494), .A2(\xmem_data[96][7] ), .B1(n30311), .B2(
        \xmem_data[97][7] ), .ZN(n13131) );
  AOI22_X1 U17271 ( .A1(n28098), .A2(\xmem_data[98][7] ), .B1(n31316), .B2(
        \xmem_data[99][7] ), .ZN(n13130) );
  AOI22_X1 U17272 ( .A1(n28328), .A2(\xmem_data[100][7] ), .B1(n27717), .B2(
        \xmem_data[101][7] ), .ZN(n13129) );
  AOI22_X1 U17273 ( .A1(n28035), .A2(\xmem_data[102][7] ), .B1(n28038), .B2(
        \xmem_data[103][7] ), .ZN(n13128) );
  NAND4_X1 U17274 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13135) );
  NAND2_X1 U17275 ( .A1(n37190), .A2(n13132), .ZN(n13133) );
  INV_X1 U17276 ( .A(n13133), .ZN(n13134) );
  AOI22_X1 U17277 ( .A1(load_xaddr_val[5]), .A2(n13133), .B1(n13134), .B2(
        n4499), .ZN(n13207) );
  AOI22_X1 U17278 ( .A1(n13134), .A2(n39040), .B1(n14909), .B2(n13133), .ZN(
        n13181) );
  AND2_X1 U17279 ( .A1(n13207), .A2(n13181), .ZN(n29171) );
  OAI21_X1 U17280 ( .B1(n13136), .B2(n13135), .A(n29171), .ZN(n13212) );
  BUF_X1 U17281 ( .A(n14973), .Z(n29089) );
  AOI22_X1 U17282 ( .A1(n29089), .A2(\xmem_data[32][7] ), .B1(n3307), .B2(
        \xmem_data[33][7] ), .ZN(n13140) );
  BUF_X1 U17283 ( .A(n14914), .Z(n27365) );
  AOI22_X1 U17284 ( .A1(n27365), .A2(\xmem_data[34][7] ), .B1(n20782), .B2(
        \xmem_data[35][7] ), .ZN(n13139) );
  BUF_X1 U17285 ( .A(n14919), .Z(n29086) );
  AOI22_X1 U17286 ( .A1(n29086), .A2(\xmem_data[36][7] ), .B1(n30674), .B2(
        \xmem_data[37][7] ), .ZN(n13138) );
  AOI22_X1 U17287 ( .A1(n30498), .A2(\xmem_data[38][7] ), .B1(n27564), .B2(
        \xmem_data[39][7] ), .ZN(n13137) );
  NAND4_X1 U17288 ( .A1(n13140), .A2(n13139), .A3(n13138), .A4(n13137), .ZN(
        n13157) );
  AOI22_X1 U17289 ( .A1(n12471), .A2(\xmem_data[40][7] ), .B1(n30864), .B2(
        \xmem_data[41][7] ), .ZN(n13144) );
  AOI22_X1 U17290 ( .A1(n14875), .A2(\xmem_data[42][7] ), .B1(n23756), .B2(
        \xmem_data[43][7] ), .ZN(n13143) );
  AOI22_X1 U17291 ( .A1(n3221), .A2(\xmem_data[44][7] ), .B1(n25448), .B2(
        \xmem_data[45][7] ), .ZN(n13142) );
  BUF_X1 U17292 ( .A(n14989), .Z(n29095) );
  AOI22_X1 U17293 ( .A1(n29095), .A2(\xmem_data[46][7] ), .B1(n25490), .B2(
        \xmem_data[47][7] ), .ZN(n13141) );
  NAND4_X1 U17294 ( .A1(n13144), .A2(n13143), .A3(n13142), .A4(n13141), .ZN(
        n13156) );
  BUF_X1 U17295 ( .A(n14890), .Z(n29104) );
  BUF_X1 U17296 ( .A(n14991), .Z(n29157) );
  AOI22_X1 U17297 ( .A1(n29104), .A2(\xmem_data[48][7] ), .B1(n29157), .B2(
        \xmem_data[49][7] ), .ZN(n13148) );
  AOI22_X1 U17298 ( .A1(n29103), .A2(\xmem_data[50][7] ), .B1(n27447), .B2(
        \xmem_data[51][7] ), .ZN(n13147) );
  AOI22_X1 U17299 ( .A1(n28415), .A2(\xmem_data[52][7] ), .B1(n17064), .B2(
        \xmem_data[53][7] ), .ZN(n13146) );
  BUF_X1 U17300 ( .A(n13436), .Z(n29109) );
  AOI22_X1 U17301 ( .A1(n24132), .A2(\xmem_data[54][7] ), .B1(n29109), .B2(
        \xmem_data[55][7] ), .ZN(n13145) );
  NAND4_X1 U17302 ( .A1(n13148), .A2(n13147), .A3(n13146), .A4(n13145), .ZN(
        n13155) );
  AOI22_X1 U17303 ( .A1(n25383), .A2(\xmem_data[58][7] ), .B1(n25635), .B2(
        \xmem_data[59][7] ), .ZN(n13153) );
  AOI22_X1 U17304 ( .A1(n30544), .A2(\xmem_data[60][7] ), .B1(n24115), .B2(
        \xmem_data[61][7] ), .ZN(n13152) );
  BUF_X1 U17305 ( .A(n3324), .Z(n29100) );
  BUF_X1 U17306 ( .A(n13481), .Z(n29101) );
  AOI22_X1 U17307 ( .A1(n17002), .A2(\xmem_data[63][7] ), .B1(
        \xmem_data[62][7] ), .B2(n29101), .ZN(n13151) );
  AOI22_X1 U17308 ( .A1(n25458), .A2(\xmem_data[56][7] ), .B1(n29437), .B2(
        \xmem_data[57][7] ), .ZN(n13150) );
  NAND4_X1 U17309 ( .A1(n13153), .A2(n13152), .A3(n13151), .A4(n13150), .ZN(
        n13154) );
  OR4_X1 U17310 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13158) );
  INV_X1 U17311 ( .A(n13181), .ZN(n13206) );
  AND2_X1 U17312 ( .A1(n13206), .A2(n13207), .ZN(n29145) );
  NAND2_X1 U17313 ( .A1(n13158), .A2(n29145), .ZN(n13211) );
  AND2_X1 U17314 ( .A1(n30589), .A2(\xmem_data[10][7] ), .ZN(n13159) );
  AOI21_X1 U17315 ( .B1(n27902), .B2(\xmem_data[11][7] ), .A(n13159), .ZN(
        n13163) );
  AOI22_X1 U17316 ( .A1(n29118), .A2(\xmem_data[8][7] ), .B1(n23732), .B2(
        \xmem_data[9][7] ), .ZN(n13162) );
  AOI22_X1 U17317 ( .A1(n3219), .A2(\xmem_data[12][7] ), .B1(n25612), .B2(
        \xmem_data[13][7] ), .ZN(n13161) );
  AOI22_X1 U17318 ( .A1(n25562), .A2(\xmem_data[14][7] ), .B1(n28083), .B2(
        \xmem_data[15][7] ), .ZN(n13160) );
  NAND4_X1 U17319 ( .A1(n13163), .A2(n13162), .A3(n13161), .A4(n13160), .ZN(
        n13180) );
  AOI22_X1 U17320 ( .A1(n17001), .A2(\xmem_data[0][7] ), .B1(n3269), .B2(
        \xmem_data[1][7] ), .ZN(n13167) );
  AOI22_X1 U17321 ( .A1(n27365), .A2(\xmem_data[2][7] ), .B1(n24685), .B2(
        \xmem_data[3][7] ), .ZN(n13166) );
  BUF_X1 U17322 ( .A(n14919), .Z(n29136) );
  AOI22_X1 U17323 ( .A1(n29136), .A2(\xmem_data[4][7] ), .B1(n21060), .B2(
        \xmem_data[5][7] ), .ZN(n13165) );
  BUF_X1 U17324 ( .A(n13457), .Z(n29125) );
  BUF_X1 U17325 ( .A(n31263), .Z(n29124) );
  AOI22_X1 U17326 ( .A1(n29125), .A2(\xmem_data[6][7] ), .B1(n29124), .B2(
        \xmem_data[7][7] ), .ZN(n13164) );
  NAND4_X1 U17327 ( .A1(n13167), .A2(n13166), .A3(n13165), .A4(n13164), .ZN(
        n13179) );
  AOI22_X1 U17328 ( .A1(n20993), .A2(\xmem_data[16][7] ), .B1(n29157), .B2(
        \xmem_data[17][7] ), .ZN(n13172) );
  AOI22_X1 U17329 ( .A1(n23771), .A2(\xmem_data[18][7] ), .B1(n27447), .B2(
        \xmem_data[19][7] ), .ZN(n13171) );
  AOI22_X1 U17330 ( .A1(n13475), .A2(\xmem_data[20][7] ), .B1(n22738), .B2(
        \xmem_data[21][7] ), .ZN(n13170) );
  AOI22_X1 U17331 ( .A1(n13168), .A2(\xmem_data[22][7] ), .B1(n20541), .B2(
        \xmem_data[23][7] ), .ZN(n13169) );
  NAND4_X1 U17332 ( .A1(n13172), .A2(n13171), .A3(n13170), .A4(n13169), .ZN(
        n13178) );
  AOI22_X1 U17333 ( .A1(n23715), .A2(\xmem_data[24][7] ), .B1(n30948), .B2(
        \xmem_data[25][7] ), .ZN(n13176) );
  AOI22_X1 U17334 ( .A1(n3207), .A2(\xmem_data[26][7] ), .B1(n24547), .B2(
        \xmem_data[27][7] ), .ZN(n13175) );
  AOI22_X1 U17335 ( .A1(n27518), .A2(\xmem_data[28][7] ), .B1(n28994), .B2(
        \xmem_data[29][7] ), .ZN(n13174) );
  AOI22_X1 U17336 ( .A1(n28380), .A2(\xmem_data[30][7] ), .B1(n29100), .B2(
        \xmem_data[31][7] ), .ZN(n13173) );
  NAND4_X1 U17337 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13177) );
  OR4_X1 U17338 ( .A1(n13180), .A2(n13179), .A3(n13178), .A4(n13177), .ZN(
        n13182) );
  NOR2_X1 U17339 ( .A1(n13207), .A2(n13181), .ZN(n29143) );
  NAND2_X1 U17340 ( .A1(n13182), .A2(n29143), .ZN(n13210) );
  AND2_X1 U17341 ( .A1(n25360), .A2(\xmem_data[74][7] ), .ZN(n13183) );
  AOI21_X1 U17342 ( .B1(n24443), .B2(\xmem_data[75][7] ), .A(n13183), .ZN(
        n13187) );
  AOI22_X1 U17343 ( .A1(n20578), .A2(\xmem_data[72][7] ), .B1(n3412), .B2(
        \xmem_data[73][7] ), .ZN(n13186) );
  AOI22_X1 U17344 ( .A1(n3218), .A2(\xmem_data[76][7] ), .B1(n31368), .B2(
        \xmem_data[77][7] ), .ZN(n13185) );
  AOI22_X1 U17345 ( .A1(n29095), .A2(\xmem_data[78][7] ), .B1(n20969), .B2(
        \xmem_data[79][7] ), .ZN(n13184) );
  NAND4_X1 U17346 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13205) );
  AOI22_X1 U17347 ( .A1(n28052), .A2(\xmem_data[88][7] ), .B1(n29396), .B2(
        \xmem_data[89][7] ), .ZN(n13192) );
  BUF_X1 U17348 ( .A(n13188), .Z(n29162) );
  AOI22_X1 U17349 ( .A1(n29162), .A2(\xmem_data[90][7] ), .B1(n25573), .B2(
        \xmem_data[91][7] ), .ZN(n13191) );
  AOI22_X1 U17350 ( .A1(n21006), .A2(\xmem_data[92][7] ), .B1(n31255), .B2(
        \xmem_data[93][7] ), .ZN(n13190) );
  AOI22_X1 U17351 ( .A1(n29101), .A2(\xmem_data[94][7] ), .B1(n24190), .B2(
        \xmem_data[95][7] ), .ZN(n13189) );
  NAND4_X1 U17352 ( .A1(n13192), .A2(n13191), .A3(n13190), .A4(n13189), .ZN(
        n13204) );
  AOI22_X1 U17353 ( .A1(n29104), .A2(\xmem_data[80][7] ), .B1(n27396), .B2(
        \xmem_data[81][7] ), .ZN(n13196) );
  AOI22_X1 U17354 ( .A1(n29103), .A2(\xmem_data[82][7] ), .B1(n30551), .B2(
        \xmem_data[83][7] ), .ZN(n13195) );
  AOI22_X1 U17355 ( .A1(n3358), .A2(\xmem_data[84][7] ), .B1(n29179), .B2(
        \xmem_data[85][7] ), .ZN(n13194) );
  AOI22_X1 U17356 ( .A1(n28375), .A2(\xmem_data[86][7] ), .B1(n29109), .B2(
        \xmem_data[87][7] ), .ZN(n13193) );
  NAND4_X1 U17357 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n13193), .ZN(
        n13203) );
  AOI22_X1 U17358 ( .A1(n29089), .A2(\xmem_data[64][7] ), .B1(n25636), .B2(
        \xmem_data[65][7] ), .ZN(n13201) );
  BUF_X1 U17359 ( .A(n14914), .Z(n29126) );
  BUF_X1 U17360 ( .A(n13486), .Z(n29151) );
  AOI22_X1 U17361 ( .A1(n29126), .A2(\xmem_data[66][7] ), .B1(n29151), .B2(
        \xmem_data[67][7] ), .ZN(n13200) );
  AND2_X1 U17362 ( .A1(n29086), .A2(\xmem_data[68][7] ), .ZN(n13197) );
  AOI21_X1 U17363 ( .B1(n29298), .B2(\xmem_data[69][7] ), .A(n13197), .ZN(
        n13199) );
  AOI22_X1 U17364 ( .A1(n27957), .A2(\xmem_data[70][7] ), .B1(n17056), .B2(
        \xmem_data[71][7] ), .ZN(n13198) );
  NAND4_X1 U17365 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        n13202) );
  OR4_X1 U17366 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13208) );
  NOR2_X1 U17367 ( .A1(n13207), .A2(n13206), .ZN(n29201) );
  NAND2_X1 U17368 ( .A1(n13208), .A2(n29201), .ZN(n13209) );
  XNOR2_X1 U17369 ( .A(n35326), .B(\fmem_data[25][3] ), .ZN(n33060) );
  INV_X1 U17370 ( .A(n13213), .ZN(n23922) );
  XNOR2_X1 U17371 ( .A(n31885), .B(\fmem_data[5][5] ), .ZN(n30435) );
  AOI22_X1 U17372 ( .A1(n3357), .A2(\xmem_data[96][6] ), .B1(n23792), .B2(
        \xmem_data[97][6] ), .ZN(n13217) );
  AOI22_X1 U17373 ( .A1(n22675), .A2(\xmem_data[98][6] ), .B1(n3176), .B2(
        \xmem_data[99][6] ), .ZN(n13216) );
  AOI22_X1 U17374 ( .A1(n22674), .A2(\xmem_data[100][6] ), .B1(n28752), .B2(
        \xmem_data[101][6] ), .ZN(n13215) );
  AOI22_X1 U17375 ( .A1(n22677), .A2(\xmem_data[102][6] ), .B1(n22676), .B2(
        \xmem_data[103][6] ), .ZN(n13214) );
  NAND4_X1 U17376 ( .A1(n13217), .A2(n13216), .A3(n13215), .A4(n13214), .ZN(
        n13220) );
  AOI22_X1 U17377 ( .A1(n25527), .A2(\xmem_data[112][6] ), .B1(n20577), .B2(
        \xmem_data[113][6] ), .ZN(n13218) );
  INV_X1 U17378 ( .A(n13218), .ZN(n13219) );
  NOR2_X1 U17379 ( .A1(n13220), .A2(n13219), .ZN(n13235) );
  AOI22_X1 U17380 ( .A1(n20568), .A2(\xmem_data[118][6] ), .B1(n25508), .B2(
        \xmem_data[119][6] ), .ZN(n13234) );
  AOI22_X1 U17381 ( .A1(n3219), .A2(\xmem_data[120][6] ), .B1(n29422), .B2(
        \xmem_data[121][6] ), .ZN(n13224) );
  AOI22_X1 U17382 ( .A1(n22667), .A2(\xmem_data[122][6] ), .B1(n22666), .B2(
        \xmem_data[123][6] ), .ZN(n13223) );
  AOI22_X1 U17383 ( .A1(n22669), .A2(\xmem_data[124][6] ), .B1(n22668), .B2(
        \xmem_data[125][6] ), .ZN(n13222) );
  AOI22_X1 U17384 ( .A1(n3231), .A2(\xmem_data[126][6] ), .B1(n28374), .B2(
        \xmem_data[127][6] ), .ZN(n13221) );
  NAND4_X1 U17385 ( .A1(n13224), .A2(n13223), .A3(n13222), .A4(n13221), .ZN(
        n13228) );
  AOI22_X1 U17386 ( .A1(n28366), .A2(\xmem_data[116][6] ), .B1(n3424), .B2(
        \xmem_data[117][6] ), .ZN(n13226) );
  AOI22_X1 U17387 ( .A1(n28329), .A2(\xmem_data[114][6] ), .B1(n27500), .B2(
        \xmem_data[115][6] ), .ZN(n13225) );
  NAND2_X1 U17388 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  NOR2_X1 U17389 ( .A1(n13228), .A2(n13227), .ZN(n13233) );
  AOI22_X1 U17390 ( .A1(n25398), .A2(\xmem_data[104][6] ), .B1(n22682), .B2(
        \xmem_data[105][6] ), .ZN(n13232) );
  AOI22_X1 U17391 ( .A1(n20941), .A2(\xmem_data[106][6] ), .B1(n22683), .B2(
        \xmem_data[107][6] ), .ZN(n13231) );
  AOI22_X1 U17392 ( .A1(n14882), .A2(\xmem_data[108][6] ), .B1(n30645), .B2(
        \xmem_data[109][6] ), .ZN(n13230) );
  AOI22_X1 U17393 ( .A1(n22685), .A2(\xmem_data[110][6] ), .B1(n22684), .B2(
        \xmem_data[111][6] ), .ZN(n13229) );
  NAND4_X1 U17394 ( .A1(n13235), .A2(n13234), .A3(n13233), .A4(n3744), .ZN(
        n13236) );
  NAND2_X1 U17395 ( .A1(n13236), .A2(n22698), .ZN(n13309) );
  AOI22_X1 U17396 ( .A1(n22701), .A2(\xmem_data[32][6] ), .B1(n31327), .B2(
        \xmem_data[33][6] ), .ZN(n13240) );
  AOI22_X1 U17397 ( .A1(n22702), .A2(\xmem_data[34][6] ), .B1(n28980), .B2(
        \xmem_data[35][6] ), .ZN(n13239) );
  AOI22_X1 U17398 ( .A1(n22703), .A2(\xmem_data[36][6] ), .B1(n25607), .B2(
        \xmem_data[37][6] ), .ZN(n13238) );
  AOI22_X1 U17399 ( .A1(n3213), .A2(\xmem_data[38][6] ), .B1(n20800), .B2(
        \xmem_data[39][6] ), .ZN(n13237) );
  NAND4_X1 U17400 ( .A1(n13240), .A2(n13239), .A3(n13238), .A4(n13237), .ZN(
        n13257) );
  AOI22_X1 U17401 ( .A1(n22718), .A2(\xmem_data[40][6] ), .B1(n22717), .B2(
        \xmem_data[41][6] ), .ZN(n13244) );
  AOI22_X1 U17402 ( .A1(n29318), .A2(\xmem_data[42][6] ), .B1(n30849), .B2(
        \xmem_data[43][6] ), .ZN(n13243) );
  AOI22_X1 U17403 ( .A1(n29089), .A2(\xmem_data[44][6] ), .B1(n3329), .B2(
        \xmem_data[45][6] ), .ZN(n13242) );
  AOI22_X1 U17404 ( .A1(n24223), .A2(\xmem_data[46][6] ), .B1(n22719), .B2(
        \xmem_data[47][6] ), .ZN(n13241) );
  NAND4_X1 U17405 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13256) );
  AOI22_X1 U17406 ( .A1(n27526), .A2(\xmem_data[48][6] ), .B1(n20985), .B2(
        \xmem_data[49][6] ), .ZN(n13249) );
  AOI22_X1 U17407 ( .A1(n22727), .A2(\xmem_data[50][6] ), .B1(n25686), .B2(
        \xmem_data[51][6] ), .ZN(n13248) );
  AOI22_X1 U17408 ( .A1(n22729), .A2(\xmem_data[52][6] ), .B1(n22728), .B2(
        \xmem_data[53][6] ), .ZN(n13247) );
  AND2_X1 U17409 ( .A1(n22753), .A2(\xmem_data[54][6] ), .ZN(n13245) );
  AOI21_X1 U17410 ( .B1(n28044), .B2(\xmem_data[55][6] ), .A(n13245), .ZN(
        n13246) );
  NAND4_X1 U17411 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        n13255) );
  AOI22_X1 U17412 ( .A1(n3222), .A2(\xmem_data[56][6] ), .B1(n22708), .B2(
        \xmem_data[57][6] ), .ZN(n13253) );
  AOI22_X1 U17413 ( .A1(n22710), .A2(\xmem_data[58][6] ), .B1(n22709), .B2(
        \xmem_data[59][6] ), .ZN(n13252) );
  AOI22_X1 U17414 ( .A1(n22711), .A2(\xmem_data[60][6] ), .B1(n3126), .B2(
        \xmem_data[61][6] ), .ZN(n13251) );
  AOI22_X1 U17415 ( .A1(n24657), .A2(\xmem_data[62][6] ), .B1(n22712), .B2(
        \xmem_data[63][6] ), .ZN(n13250) );
  NAND4_X1 U17416 ( .A1(n13253), .A2(n13252), .A3(n13251), .A4(n13250), .ZN(
        n13254) );
  OR4_X1 U17417 ( .A1(n13257), .A2(n13256), .A3(n13255), .A4(n13254), .ZN(
        n13258) );
  NAND2_X1 U17418 ( .A1(n13258), .A2(n22735), .ZN(n13308) );
  AOI22_X1 U17419 ( .A1(n29136), .A2(\xmem_data[80][6] ), .B1(n20770), .B2(
        \xmem_data[81][6] ), .ZN(n13270) );
  AOI22_X1 U17420 ( .A1(n22729), .A2(\xmem_data[84][6] ), .B1(n22728), .B2(
        \xmem_data[85][6] ), .ZN(n13259) );
  INV_X1 U17421 ( .A(n13259), .ZN(n13262) );
  AOI22_X1 U17422 ( .A1(n22727), .A2(\xmem_data[82][6] ), .B1(n28354), .B2(
        \xmem_data[83][6] ), .ZN(n13260) );
  INV_X1 U17423 ( .A(n13260), .ZN(n13261) );
  NOR2_X1 U17424 ( .A1(n13262), .A2(n13261), .ZN(n13269) );
  AND2_X1 U17425 ( .A1(n25442), .A2(\xmem_data[86][6] ), .ZN(n13263) );
  AOI21_X1 U17426 ( .B1(n24532), .B2(\xmem_data[87][6] ), .A(n13263), .ZN(
        n13268) );
  AOI22_X1 U17427 ( .A1(n3217), .A2(\xmem_data[88][6] ), .B1(n22708), .B2(
        \xmem_data[89][6] ), .ZN(n13267) );
  AOI22_X1 U17428 ( .A1(n22710), .A2(\xmem_data[90][6] ), .B1(n22709), .B2(
        \xmem_data[91][6] ), .ZN(n13266) );
  AOI22_X1 U17429 ( .A1(n22711), .A2(\xmem_data[92][6] ), .B1(n3375), .B2(
        \xmem_data[93][6] ), .ZN(n13265) );
  AOI22_X1 U17430 ( .A1(n25450), .A2(\xmem_data[94][6] ), .B1(n22712), .B2(
        \xmem_data[95][6] ), .ZN(n13264) );
  NAND4_X1 U17431 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n3745), .ZN(
        n13282) );
  AOI22_X1 U17432 ( .A1(n22718), .A2(\xmem_data[72][6] ), .B1(n22717), .B2(
        \xmem_data[73][6] ), .ZN(n13274) );
  AOI22_X1 U17433 ( .A1(n28301), .A2(\xmem_data[74][6] ), .B1(n21010), .B2(
        \xmem_data[75][6] ), .ZN(n13273) );
  AOI22_X1 U17434 ( .A1(n25581), .A2(\xmem_data[76][6] ), .B1(n3329), .B2(
        \xmem_data[77][6] ), .ZN(n13272) );
  AOI22_X1 U17435 ( .A1(n24622), .A2(\xmem_data[78][6] ), .B1(n22719), .B2(
        \xmem_data[79][6] ), .ZN(n13271) );
  NAND4_X1 U17436 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13280) );
  AOI22_X1 U17437 ( .A1(n22701), .A2(\xmem_data[64][6] ), .B1(n24556), .B2(
        \xmem_data[65][6] ), .ZN(n13278) );
  AOI22_X1 U17438 ( .A1(n22702), .A2(n20682), .B1(n25567), .B2(
        \xmem_data[67][6] ), .ZN(n13277) );
  AOI22_X1 U17439 ( .A1(n22703), .A2(\xmem_data[68][6] ), .B1(n3158), .B2(
        \xmem_data[69][6] ), .ZN(n13276) );
  AOI22_X1 U17440 ( .A1(n28335), .A2(\xmem_data[70][6] ), .B1(n29010), .B2(
        \xmem_data[71][6] ), .ZN(n13275) );
  NAND4_X1 U17441 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13279) );
  OR2_X1 U17442 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  OAI21_X1 U17443 ( .B1(n13282), .B2(n13281), .A(n22663), .ZN(n13307) );
  AND2_X1 U17444 ( .A1(n22751), .A2(\xmem_data[16][6] ), .ZN(n13283) );
  AOI21_X1 U17445 ( .B1(n29725), .B2(\xmem_data[17][6] ), .A(n13283), .ZN(
        n13287) );
  AOI22_X1 U17446 ( .A1(n16999), .A2(\xmem_data[18][6] ), .B1(n28076), .B2(
        \xmem_data[19][6] ), .ZN(n13286) );
  AOI22_X1 U17447 ( .A1(n22752), .A2(\xmem_data[20][6] ), .B1(n25443), .B2(
        \xmem_data[21][6] ), .ZN(n13285) );
  AOI22_X1 U17448 ( .A1(n22753), .A2(\xmem_data[22][6] ), .B1(n29064), .B2(
        \xmem_data[23][6] ), .ZN(n13284) );
  NAND4_X1 U17449 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13288) );
  AOI22_X1 U17450 ( .A1(n22739), .A2(\xmem_data[0][6] ), .B1(n22738), .B2(
        \xmem_data[1][6] ), .ZN(n13292) );
  AOI22_X1 U17451 ( .A1(n22740), .A2(\xmem_data[2][6] ), .B1(n28298), .B2(
        \xmem_data[3][6] ), .ZN(n13291) );
  AOI22_X1 U17452 ( .A1(n22741), .A2(\xmem_data[4][6] ), .B1(n29315), .B2(
        \xmem_data[5][6] ), .ZN(n13290) );
  AOI22_X1 U17453 ( .A1(n22742), .A2(\xmem_data[6][6] ), .B1(n28096), .B2(
        \xmem_data[7][6] ), .ZN(n13289) );
  NAND4_X1 U17454 ( .A1(n13292), .A2(n13291), .A3(n13290), .A4(n13289), .ZN(
        n13304) );
  AOI22_X1 U17455 ( .A1(n25581), .A2(\xmem_data[12][6] ), .B1(n20950), .B2(
        \xmem_data[13][6] ), .ZN(n13296) );
  AOI22_X1 U17456 ( .A1(n28983), .A2(\xmem_data[14][6] ), .B1(n20734), .B2(
        \xmem_data[15][6] ), .ZN(n13295) );
  AOI22_X1 U17457 ( .A1(n27918), .A2(\xmem_data[8][6] ), .B1(n31255), .B2(
        \xmem_data[9][6] ), .ZN(n13294) );
  AOI22_X1 U17458 ( .A1(n28428), .A2(\xmem_data[11][6] ), .B1(
        \xmem_data[10][6] ), .B2(n29238), .ZN(n13293) );
  NAND4_X1 U17459 ( .A1(n13296), .A2(n13295), .A3(n13294), .A4(n13293), .ZN(
        n13303) );
  AOI22_X1 U17460 ( .A1(n22759), .A2(\xmem_data[28][6] ), .B1(n30710), .B2(
        \xmem_data[29][6] ), .ZN(n13297) );
  INV_X1 U17461 ( .A(n13297), .ZN(n13302) );
  AOI22_X1 U17462 ( .A1(n3222), .A2(\xmem_data[24][6] ), .B1(n29288), .B2(
        \xmem_data[25][6] ), .ZN(n13300) );
  AOI22_X1 U17463 ( .A1(n20598), .A2(\xmem_data[26][6] ), .B1(n22758), .B2(
        \xmem_data[27][6] ), .ZN(n13299) );
  NAND2_X1 U17464 ( .A1(n16974), .A2(\xmem_data[31][6] ), .ZN(n13298) );
  NAND3_X1 U17465 ( .A1(n13300), .A2(n13299), .A3(n13298), .ZN(n13301) );
  OAI21_X1 U17466 ( .B1(n3982), .B2(n13305), .A(n22768), .ZN(n13306) );
  AOI22_X1 U17467 ( .A1(n3172), .A2(\xmem_data[96][5] ), .B1(n23725), .B2(
        \xmem_data[97][5] ), .ZN(n13313) );
  AOI22_X1 U17468 ( .A1(n28036), .A2(\xmem_data[98][5] ), .B1(n28035), .B2(
        \xmem_data[99][5] ), .ZN(n13312) );
  AOI22_X1 U17469 ( .A1(n28038), .A2(\xmem_data[100][5] ), .B1(n28037), .B2(
        \xmem_data[101][5] ), .ZN(n13311) );
  AOI22_X1 U17470 ( .A1(n28039), .A2(\xmem_data[102][5] ), .B1(n28501), .B2(
        \xmem_data[103][5] ), .ZN(n13310) );
  NAND4_X1 U17471 ( .A1(n13313), .A2(n13312), .A3(n13311), .A4(n13310), .ZN(
        n13329) );
  AOI22_X1 U17472 ( .A1(n28044), .A2(\xmem_data[104][5] ), .B1(n3221), .B2(
        \xmem_data[105][5] ), .ZN(n13317) );
  AOI22_X1 U17473 ( .A1(n31368), .A2(\xmem_data[106][5] ), .B1(n25509), .B2(
        \xmem_data[107][5] ), .ZN(n13316) );
  AOI22_X1 U17474 ( .A1(n25449), .A2(\xmem_data[108][5] ), .B1(n21068), .B2(
        \xmem_data[109][5] ), .ZN(n13315) );
  AOI22_X1 U17475 ( .A1(n3375), .A2(\xmem_data[110][5] ), .B1(n28343), .B2(
        \xmem_data[111][5] ), .ZN(n13314) );
  NAND4_X1 U17476 ( .A1(n13317), .A2(n13316), .A3(n13315), .A4(n13314), .ZN(
        n13328) );
  AOI22_X1 U17477 ( .A1(n28050), .A2(\xmem_data[112][5] ), .B1(n28481), .B2(
        \xmem_data[113][5] ), .ZN(n13321) );
  AOI22_X1 U17478 ( .A1(n28051), .A2(\xmem_data[114][5] ), .B1(n21075), .B2(
        \xmem_data[115][5] ), .ZN(n13320) );
  AOI22_X1 U17479 ( .A1(n27515), .A2(\xmem_data[116][5] ), .B1(n28052), .B2(
        \xmem_data[117][5] ), .ZN(n13319) );
  AOI22_X1 U17480 ( .A1(n27517), .A2(\xmem_data[118][5] ), .B1(n30542), .B2(
        \xmem_data[119][5] ), .ZN(n13318) );
  NAND4_X1 U17481 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13327) );
  AOI22_X1 U17482 ( .A1(n28059), .A2(\xmem_data[120][5] ), .B1(n28058), .B2(
        \xmem_data[121][5] ), .ZN(n13325) );
  AOI22_X1 U17483 ( .A1(n29012), .A2(\xmem_data[122][5] ), .B1(n25576), .B2(
        \xmem_data[123][5] ), .ZN(n13324) );
  AOI22_X1 U17484 ( .A1(n28061), .A2(\xmem_data[124][5] ), .B1(n28060), .B2(
        \xmem_data[125][5] ), .ZN(n13323) );
  AOI22_X1 U17485 ( .A1(n24623), .A2(\xmem_data[126][5] ), .B1(n28062), .B2(
        \xmem_data[127][5] ), .ZN(n13322) );
  NAND4_X1 U17486 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13326) );
  OR4_X1 U17487 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13351) );
  AOI22_X1 U17488 ( .A1(n14976), .A2(\xmem_data[64][5] ), .B1(n28468), .B2(
        \xmem_data[65][5] ), .ZN(n13333) );
  AOI22_X1 U17489 ( .A1(n30257), .A2(\xmem_data[66][5] ), .B1(n29248), .B2(
        \xmem_data[67][5] ), .ZN(n13332) );
  AOI22_X1 U17490 ( .A1(n28076), .A2(\xmem_data[68][5] ), .B1(n28075), .B2(
        \xmem_data[69][5] ), .ZN(n13331) );
  AOI22_X1 U17491 ( .A1(n3434), .A2(\xmem_data[70][5] ), .B1(n3247), .B2(
        \xmem_data[71][5] ), .ZN(n13330) );
  NAND4_X1 U17492 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n13349) );
  AOI22_X1 U17493 ( .A1(n28082), .A2(\xmem_data[72][5] ), .B1(n3220), .B2(
        \xmem_data[73][5] ), .ZN(n13337) );
  AOI22_X1 U17494 ( .A1(n30964), .A2(\xmem_data[74][5] ), .B1(n23769), .B2(
        \xmem_data[75][5] ), .ZN(n13336) );
  AOI22_X1 U17495 ( .A1(n28083), .A2(\xmem_data[76][5] ), .B1(n13444), .B2(
        \xmem_data[77][5] ), .ZN(n13335) );
  AOI22_X1 U17496 ( .A1(n28084), .A2(\xmem_data[78][5] ), .B1(n25492), .B2(
        \xmem_data[79][5] ), .ZN(n13334) );
  NAND4_X1 U17497 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13348) );
  AOI22_X1 U17498 ( .A1(n27551), .A2(\xmem_data[80][5] ), .B1(n13475), .B2(
        \xmem_data[81][5] ), .ZN(n13341) );
  AOI22_X1 U17499 ( .A1(n28089), .A2(\xmem_data[82][5] ), .B1(n24212), .B2(
        \xmem_data[83][5] ), .ZN(n13340) );
  AOI22_X1 U17500 ( .A1(n28980), .A2(\xmem_data[84][5] ), .B1(n28090), .B2(
        \xmem_data[85][5] ), .ZN(n13339) );
  AOI22_X1 U17501 ( .A1(n20776), .A2(\xmem_data[86][5] ), .B1(n27864), .B2(
        \xmem_data[87][5] ), .ZN(n13338) );
  NAND4_X1 U17502 ( .A1(n13341), .A2(n13340), .A3(n13339), .A4(n13338), .ZN(
        n13347) );
  AOI22_X1 U17503 ( .A1(n28096), .A2(\xmem_data[88][5] ), .B1(n31355), .B2(
        \xmem_data[89][5] ), .ZN(n13345) );
  AOI22_X1 U17504 ( .A1(n28994), .A2(\xmem_data[90][5] ), .B1(n28097), .B2(
        \xmem_data[91][5] ), .ZN(n13344) );
  AOI22_X1 U17505 ( .A1(n21010), .A2(\xmem_data[92][5] ), .B1(n21051), .B2(
        \xmem_data[93][5] ), .ZN(n13343) );
  AOI22_X1 U17506 ( .A1(n17004), .A2(\xmem_data[94][5] ), .B1(n28098), .B2(
        \xmem_data[95][5] ), .ZN(n13342) );
  NAND4_X1 U17507 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13346) );
  OR4_X1 U17508 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13350) );
  AOI22_X1 U17509 ( .A1(n28071), .A2(n13351), .B1(n28033), .B2(n13350), .ZN(
        n13405) );
  AOI22_X1 U17510 ( .A1(n28059), .A2(\xmem_data[24][5] ), .B1(n28492), .B2(
        \xmem_data[25][5] ), .ZN(n13355) );
  AOI22_X1 U17511 ( .A1(n30893), .A2(\xmem_data[26][5] ), .B1(n13481), .B2(
        \xmem_data[27][5] ), .ZN(n13354) );
  AOI22_X1 U17512 ( .A1(n27974), .A2(\xmem_data[28][5] ), .B1(n30495), .B2(
        \xmem_data[29][5] ), .ZN(n13353) );
  AOI22_X1 U17513 ( .A1(n3330), .A2(\xmem_data[30][5] ), .B1(n27975), .B2(
        \xmem_data[31][5] ), .ZN(n13352) );
  NAND4_X1 U17514 ( .A1(n13355), .A2(n13354), .A3(n13353), .A4(n13352), .ZN(
        n13361) );
  AOI22_X1 U17515 ( .A1(n25582), .A2(\xmem_data[0][5] ), .B1(n27981), .B2(
        \xmem_data[1][5] ), .ZN(n13359) );
  AOI22_X1 U17516 ( .A1(n23730), .A2(\xmem_data[2][5] ), .B1(n30524), .B2(
        \xmem_data[3][5] ), .ZN(n13358) );
  AOI22_X1 U17517 ( .A1(n28076), .A2(\xmem_data[4][5] ), .B1(n20489), .B2(
        \xmem_data[5][5] ), .ZN(n13357) );
  AOI22_X1 U17518 ( .A1(n3449), .A2(\xmem_data[6][5] ), .B1(n29173), .B2(
        \xmem_data[7][5] ), .ZN(n13356) );
  NAND4_X1 U17519 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        n13360) );
  OR2_X1 U17520 ( .A1(n13361), .A2(n13360), .ZN(n13378) );
  NAND2_X1 U17521 ( .A1(n28044), .A2(\xmem_data[8][5] ), .ZN(n13363) );
  NAND2_X1 U17522 ( .A1(n3218), .A2(\xmem_data[9][5] ), .ZN(n13362) );
  NAND2_X1 U17523 ( .A1(n13363), .A2(n13362), .ZN(n13367) );
  AOI22_X1 U17524 ( .A1(n28475), .A2(\xmem_data[12][5] ), .B1(n27994), .B2(
        \xmem_data[13][5] ), .ZN(n13365) );
  NAND2_X1 U17525 ( .A1(n3138), .A2(\xmem_data[14][5] ), .ZN(n13364) );
  NAND2_X1 U17526 ( .A1(n13365), .A2(n13364), .ZN(n13366) );
  NOR2_X1 U17527 ( .A1(n13367), .A2(n13366), .ZN(n13376) );
  AOI22_X1 U17528 ( .A1(n30607), .A2(\xmem_data[16][5] ), .B1(n27988), .B2(
        \xmem_data[17][5] ), .ZN(n13371) );
  AOI22_X1 U17529 ( .A1(n29179), .A2(\xmem_data[18][5] ), .B1(n28515), .B2(
        \xmem_data[19][5] ), .ZN(n13370) );
  AOI22_X1 U17530 ( .A1(n13436), .A2(\xmem_data[20][5] ), .B1(n23793), .B2(
        \xmem_data[21][5] ), .ZN(n13369) );
  AOI22_X1 U17531 ( .A1(n23795), .A2(\xmem_data[22][5] ), .B1(n27989), .B2(
        \xmem_data[23][5] ), .ZN(n13368) );
  NAND4_X1 U17532 ( .A1(n13371), .A2(n13370), .A3(n13369), .A4(n13368), .ZN(
        n13374) );
  AOI22_X1 U17533 ( .A1(n20805), .A2(\xmem_data[10][5] ), .B1(n24695), .B2(
        \xmem_data[11][5] ), .ZN(n13372) );
  NOR2_X1 U17534 ( .A1(n13374), .A2(n13373), .ZN(n13375) );
  NAND2_X1 U17535 ( .A1(n13376), .A2(n13375), .ZN(n13377) );
  NOR2_X1 U17536 ( .A1(n13378), .A2(n13377), .ZN(n13380) );
  NAND2_X1 U17537 ( .A1(n31252), .A2(\xmem_data[15][5] ), .ZN(n13379) );
  AOI21_X1 U17538 ( .B1(n13380), .B2(n13379), .A(n24043), .ZN(n13403) );
  AOI22_X1 U17539 ( .A1(n3172), .A2(\xmem_data[32][5] ), .B1(n27981), .B2(
        \xmem_data[33][5] ), .ZN(n13384) );
  AOI22_X1 U17540 ( .A1(n30901), .A2(\xmem_data[34][5] ), .B1(n30524), .B2(
        \xmem_data[35][5] ), .ZN(n13383) );
  AOI22_X1 U17541 ( .A1(n28076), .A2(\xmem_data[36][5] ), .B1(n28075), .B2(
        \xmem_data[37][5] ), .ZN(n13382) );
  AOI22_X1 U17542 ( .A1(n3434), .A2(\xmem_data[38][5] ), .B1(n3247), .B2(
        \xmem_data[39][5] ), .ZN(n13381) );
  NAND4_X1 U17543 ( .A1(n13384), .A2(n13383), .A3(n13382), .A4(n13381), .ZN(
        n13400) );
  AOI22_X1 U17544 ( .A1(n28082), .A2(\xmem_data[40][5] ), .B1(n3219), .B2(
        \xmem_data[41][5] ), .ZN(n13388) );
  AOI22_X1 U17545 ( .A1(n27445), .A2(\xmem_data[42][5] ), .B1(n23739), .B2(
        \xmem_data[43][5] ), .ZN(n13387) );
  AOI22_X1 U17546 ( .A1(n28083), .A2(\xmem_data[44][5] ), .B1(n28509), .B2(
        \xmem_data[45][5] ), .ZN(n13386) );
  AOI22_X1 U17547 ( .A1(n28084), .A2(\xmem_data[46][5] ), .B1(n25450), .B2(
        \xmem_data[47][5] ), .ZN(n13385) );
  NAND4_X1 U17548 ( .A1(n13388), .A2(n13387), .A3(n13386), .A4(n13385), .ZN(
        n13399) );
  AOI22_X1 U17549 ( .A1(n27551), .A2(\xmem_data[48][5] ), .B1(n13475), .B2(
        \xmem_data[49][5] ), .ZN(n13392) );
  AOI22_X1 U17550 ( .A1(n28089), .A2(\xmem_data[50][5] ), .B1(n27535), .B2(
        \xmem_data[51][5] ), .ZN(n13391) );
  AOI22_X1 U17551 ( .A1(n13436), .A2(\xmem_data[52][5] ), .B1(n28090), .B2(
        \xmem_data[53][5] ), .ZN(n13390) );
  AOI22_X1 U17552 ( .A1(n28091), .A2(\xmem_data[54][5] ), .B1(n3208), .B2(
        \xmem_data[55][5] ), .ZN(n13389) );
  NAND4_X1 U17553 ( .A1(n13392), .A2(n13391), .A3(n13390), .A4(n13389), .ZN(
        n13398) );
  AOI22_X1 U17554 ( .A1(n28096), .A2(\xmem_data[56][5] ), .B1(n31355), .B2(
        \xmem_data[57][5] ), .ZN(n13396) );
  AOI22_X1 U17555 ( .A1(n25400), .A2(\xmem_data[58][5] ), .B1(n28097), .B2(
        \xmem_data[59][5] ), .ZN(n13395) );
  AOI22_X1 U17556 ( .A1(n3177), .A2(\xmem_data[60][5] ), .B1(n28429), .B2(
        \xmem_data[61][5] ), .ZN(n13394) );
  AOI22_X1 U17557 ( .A1(n25636), .A2(\xmem_data[62][5] ), .B1(n28098), .B2(
        \xmem_data[63][5] ), .ZN(n13393) );
  NAND4_X1 U17558 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        n13397) );
  OR4_X1 U17559 ( .A1(n13400), .A2(n13399), .A3(n13398), .A4(n13397), .ZN(
        n13401) );
  AND2_X1 U17560 ( .A1(n13401), .A2(n28107), .ZN(n13402) );
  NOR2_X1 U17561 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  XOR2_X1 U17562 ( .A(\fmem_data[22][5] ), .B(\fmem_data[22][4] ), .Z(n13406)
         );
  AOI22_X1 U17563 ( .A1(n29661), .A2(\xmem_data[32][3] ), .B1(n3247), .B2(
        \xmem_data[33][3] ), .ZN(n13410) );
  BUF_X1 U17564 ( .A(n29064), .Z(n24562) );
  AOI22_X1 U17565 ( .A1(n24562), .A2(\xmem_data[34][3] ), .B1(n3221), .B2(
        \xmem_data[35][3] ), .ZN(n13409) );
  BUF_X1 U17566 ( .A(n14988), .Z(n24563) );
  AOI22_X1 U17567 ( .A1(n24563), .A2(\xmem_data[36][3] ), .B1(n29255), .B2(
        \xmem_data[37][3] ), .ZN(n13408) );
  BUF_X1 U17568 ( .A(n14926), .Z(n24565) );
  BUF_X1 U17569 ( .A(n14927), .Z(n24564) );
  AOI22_X1 U17570 ( .A1(n24565), .A2(\xmem_data[38][3] ), .B1(n24564), .B2(
        \xmem_data[39][3] ), .ZN(n13407) );
  NAND4_X1 U17571 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13428) );
  BUF_X1 U17572 ( .A(n15011), .Z(n24553) );
  AOI22_X1 U17573 ( .A1(n3344), .A2(\xmem_data[40][3] ), .B1(n24553), .B2(
        \xmem_data[41][3] ), .ZN(n13414) );
  BUF_X1 U17574 ( .A(n31276), .Z(n24554) );
  AOI22_X1 U17575 ( .A1(n24554), .A2(\xmem_data[42][3] ), .B1(n29180), .B2(
        \xmem_data[43][3] ), .ZN(n13413) );
  BUF_X1 U17576 ( .A(n14997), .Z(n24556) );
  BUF_X1 U17577 ( .A(n13435), .Z(n24555) );
  AOI22_X1 U17578 ( .A1(n24556), .A2(\xmem_data[44][3] ), .B1(n24555), .B2(
        \xmem_data[45][3] ), .ZN(n13412) );
  AOI22_X1 U17579 ( .A1(n16986), .A2(\xmem_data[46][3] ), .B1(n24160), .B2(
        \xmem_data[47][3] ), .ZN(n13411) );
  NAND4_X1 U17580 ( .A1(n13414), .A2(n13413), .A3(n13412), .A4(n13411), .ZN(
        n13427) );
  BUF_X1 U17581 ( .A(n3464), .Z(n24545) );
  AOI22_X1 U17582 ( .A1(n24545), .A2(\xmem_data[48][3] ), .B1(n31269), .B2(
        \xmem_data[49][3] ), .ZN(n13419) );
  BUF_X1 U17583 ( .A(n14937), .Z(n24547) );
  BUF_X1 U17584 ( .A(n13415), .Z(n24546) );
  AOI22_X1 U17585 ( .A1(n24547), .A2(\xmem_data[50][3] ), .B1(n24546), .B2(
        \xmem_data[51][3] ), .ZN(n13418) );
  AOI22_X1 U17586 ( .A1(n25678), .A2(\xmem_data[52][3] ), .B1(n24460), .B2(
        \xmem_data[53][3] ), .ZN(n13417) );
  BUF_X1 U17587 ( .A(n3324), .Z(n24548) );
  AOI22_X1 U17588 ( .A1(n24548), .A2(\xmem_data[54][3] ), .B1(n29281), .B2(
        \xmem_data[55][3] ), .ZN(n13416) );
  NAND4_X1 U17589 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        n13426) );
  BUF_X1 U17590 ( .A(n14974), .Z(n24571) );
  BUF_X1 U17591 ( .A(n14914), .Z(n24570) );
  AOI22_X1 U17592 ( .A1(n24571), .A2(\xmem_data[56][3] ), .B1(n24570), .B2(
        \xmem_data[57][3] ), .ZN(n13424) );
  BUF_X1 U17593 ( .A(n14976), .Z(n24572) );
  AOI22_X1 U17594 ( .A1(n24572), .A2(\xmem_data[58][3] ), .B1(n21057), .B2(
        \xmem_data[59][3] ), .ZN(n13423) );
  AOI22_X1 U17595 ( .A1(n27852), .A2(\xmem_data[60][3] ), .B1(n16999), .B2(
        \xmem_data[61][3] ), .ZN(n13422) );
  BUF_X1 U17596 ( .A(n28947), .Z(n24573) );
  AOI22_X1 U17597 ( .A1(n29124), .A2(\xmem_data[62][3] ), .B1(n24573), .B2(
        \xmem_data[63][3] ), .ZN(n13421) );
  NAND4_X1 U17598 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n13421), .ZN(
        n13425) );
  OR4_X1 U17599 ( .A1(n13428), .A2(n13427), .A3(n13426), .A4(n13425), .ZN(
        n13434) );
  INV_X1 U17600 ( .A(n13467), .ZN(n13496) );
  MUX2_X1 U17601 ( .A(n37191), .B(n4499), .S(n13432), .Z(n13433) );
  INV_X1 U17602 ( .A(n13433), .ZN(n13497) );
  BUF_X1 U17603 ( .A(n29064), .Z(n24443) );
  BUF_X1 U17604 ( .A(n13435), .Z(n24448) );
  AOI22_X1 U17605 ( .A1(n27944), .A2(\xmem_data[12][3] ), .B1(n24448), .B2(
        \xmem_data[13][3] ), .ZN(n13439) );
  AOI22_X1 U17606 ( .A1(n17041), .A2(\xmem_data[14][3] ), .B1(n24160), .B2(
        \xmem_data[15][3] ), .ZN(n13438) );
  BUF_X1 U17607 ( .A(n25604), .Z(n24450) );
  AOI22_X1 U17608 ( .A1(n24450), .A2(\xmem_data[10][3] ), .B1(n27863), .B2(
        \xmem_data[11][3] ), .ZN(n13437) );
  BUF_X1 U17609 ( .A(n13468), .Z(n24439) );
  AOI22_X1 U17610 ( .A1(n22728), .A2(\xmem_data[0][3] ), .B1(n24439), .B2(
        \xmem_data[1][3] ), .ZN(n13440) );
  INV_X1 U17611 ( .A(n13440), .ZN(n13441) );
  BUF_X1 U17612 ( .A(n14974), .Z(n24466) );
  AOI22_X1 U17613 ( .A1(n3338), .A2(\xmem_data[24][3] ), .B1(n28098), .B2(
        \xmem_data[25][3] ), .ZN(n13443) );
  AOI22_X1 U17614 ( .A1(n24632), .A2(\xmem_data[4][3] ), .B1(n20500), .B2(
        \xmem_data[5][3] ), .ZN(n13442) );
  BUF_X1 U17615 ( .A(n14990), .Z(n24438) );
  AOI22_X1 U17616 ( .A1(n24438), .A2(\xmem_data[6][3] ), .B1(n17061), .B2(
        \xmem_data[7][3] ), .ZN(n13446) );
  BUF_X1 U17617 ( .A(n13486), .Z(n24467) );
  AOI22_X1 U17618 ( .A1(n24467), .A2(\xmem_data[26][3] ), .B1(n23725), .B2(
        \xmem_data[27][3] ), .ZN(n13445) );
  NAND2_X1 U17619 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NOR2_X1 U17620 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  NAND4_X1 U17621 ( .A1(n13451), .A2(n3907), .A3(n13450), .A4(n13449), .ZN(
        n13463) );
  BUF_X1 U17622 ( .A(n3464), .Z(n24458) );
  BUF_X1 U17623 ( .A(n14936), .Z(n24457) );
  AOI22_X1 U17624 ( .A1(n24458), .A2(\xmem_data[16][3] ), .B1(n24457), .B2(
        \xmem_data[17][3] ), .ZN(n13456) );
  BUF_X1 U17625 ( .A(n14912), .Z(n24459) );
  AOI22_X1 U17626 ( .A1(n24133), .A2(\xmem_data[18][3] ), .B1(n24459), .B2(
        \xmem_data[19][3] ), .ZN(n13455) );
  BUF_X1 U17627 ( .A(n13452), .Z(n24460) );
  AOI22_X1 U17628 ( .A1(n30893), .A2(\xmem_data[20][3] ), .B1(n24460), .B2(
        \xmem_data[21][3] ), .ZN(n13454) );
  BUF_X1 U17629 ( .A(n14972), .Z(n24461) );
  AOI22_X1 U17630 ( .A1(n3178), .A2(\xmem_data[22][3] ), .B1(n30955), .B2(
        \xmem_data[23][3] ), .ZN(n13453) );
  NAND4_X1 U17631 ( .A1(n13456), .A2(n13455), .A3(n13454), .A4(n13453), .ZN(
        n13461) );
  BUF_X1 U17632 ( .A(n13457), .Z(n24468) );
  NAND2_X1 U17633 ( .A1(n24468), .A2(\xmem_data[29][3] ), .ZN(n13459) );
  BUF_X1 U17634 ( .A(n28947), .Z(n24470) );
  NAND2_X1 U17635 ( .A1(n24470), .A2(\xmem_data[31][3] ), .ZN(n13458) );
  NAND4_X1 U17636 ( .A1(n3556), .A2(n13459), .A3(n13458), .A4(n4001), .ZN(
        n13460) );
  OR2_X1 U17637 ( .A1(n13461), .A2(n13460), .ZN(n13462) );
  NOR2_X1 U17638 ( .A1(n13463), .A2(n13462), .ZN(n13464) );
  NOR2_X1 U17639 ( .A1(n13497), .A2(n13467), .ZN(n22180) );
  AOI21_X1 U17640 ( .B1(n27878), .B2(n13464), .A(n22298), .ZN(n13466) );
  NAND2_X1 U17641 ( .A1(n13464), .A2(n39034), .ZN(n13465) );
  NAND2_X1 U17642 ( .A1(n13466), .A2(n13465), .ZN(n13521) );
  AND2_X1 U17643 ( .A1(n13497), .A2(n13467), .ZN(n24542) );
  AOI22_X1 U17644 ( .A1(n3449), .A2(\xmem_data[96][3] ), .B1(n28501), .B2(
        \xmem_data[97][3] ), .ZN(n13473) );
  BUF_X1 U17645 ( .A(n29064), .Z(n24532) );
  AOI22_X1 U17646 ( .A1(n24532), .A2(\xmem_data[98][3] ), .B1(n3220), .B2(
        \xmem_data[99][3] ), .ZN(n13472) );
  BUF_X1 U17647 ( .A(n14988), .Z(n24533) );
  AOI22_X1 U17648 ( .A1(n24533), .A2(\xmem_data[100][3] ), .B1(n20500), .B2(
        \xmem_data[101][3] ), .ZN(n13471) );
  BUF_X1 U17649 ( .A(n14926), .Z(n24534) );
  AOI22_X1 U17650 ( .A1(n24534), .A2(\xmem_data[102][3] ), .B1(n30550), .B2(
        \xmem_data[103][3] ), .ZN(n13470) );
  NAND4_X1 U17651 ( .A1(n13473), .A2(n13472), .A3(n13471), .A4(n13470), .ZN(
        n13495) );
  AOI22_X1 U17652 ( .A1(n3375), .A2(\xmem_data[104][3] ), .B1(n29103), .B2(
        \xmem_data[105][3] ), .ZN(n13480) );
  AOI22_X1 U17653 ( .A1(n25604), .A2(\xmem_data[106][3] ), .B1(n29307), .B2(
        \xmem_data[107][3] ), .ZN(n13479) );
  BUF_X1 U17654 ( .A(n14934), .Z(n24516) );
  AOI22_X1 U17655 ( .A1(n20545), .A2(\xmem_data[108][3] ), .B1(n24516), .B2(
        \xmem_data[109][3] ), .ZN(n13478) );
  AOI22_X1 U17656 ( .A1(n28298), .A2(\xmem_data[110][3] ), .B1(n23793), .B2(
        \xmem_data[111][3] ), .ZN(n13477) );
  NAND4_X1 U17657 ( .A1(n13480), .A2(n13479), .A3(n13478), .A4(n13477), .ZN(
        n13494) );
  AOI22_X1 U17658 ( .A1(n30892), .A2(\xmem_data[112][3] ), .B1(n27864), .B2(
        \xmem_data[113][3] ), .ZN(n13485) );
  AOI22_X1 U17659 ( .A1(n24509), .A2(\xmem_data[114][3] ), .B1(n27518), .B2(
        \xmem_data[115][3] ), .ZN(n13484) );
  BUF_X1 U17660 ( .A(n13481), .Z(n24510) );
  AOI22_X1 U17661 ( .A1(n23777), .A2(\xmem_data[116][3] ), .B1(n24510), .B2(
        \xmem_data[117][3] ), .ZN(n13483) );
  BUF_X1 U17662 ( .A(n14881), .Z(n24511) );
  AOI22_X1 U17663 ( .A1(n24511), .A2(\xmem_data[118][3] ), .B1(n21051), .B2(
        \xmem_data[119][3] ), .ZN(n13482) );
  NAND4_X1 U17664 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n13493) );
  BUF_X1 U17665 ( .A(n14974), .Z(n24522) );
  BUF_X1 U17666 ( .A(n14914), .Z(n24521) );
  AOI22_X1 U17667 ( .A1(n24522), .A2(\xmem_data[120][3] ), .B1(n24521), .B2(
        \xmem_data[121][3] ), .ZN(n13491) );
  BUF_X1 U17668 ( .A(n13486), .Z(n24523) );
  AOI22_X1 U17669 ( .A1(n3209), .A2(\xmem_data[122][3] ), .B1(n28500), .B2(
        \xmem_data[123][3] ), .ZN(n13490) );
  BUF_X1 U17670 ( .A(n13487), .Z(n24524) );
  AOI22_X1 U17671 ( .A1(n20952), .A2(\xmem_data[124][3] ), .B1(n24524), .B2(
        \xmem_data[125][3] ), .ZN(n13489) );
  BUF_X1 U17672 ( .A(n31263), .Z(n24526) );
  AOI22_X1 U17673 ( .A1(n24526), .A2(\xmem_data[126][3] ), .B1(n24525), .B2(
        \xmem_data[127][3] ), .ZN(n13488) );
  NAND4_X1 U17674 ( .A1(n13491), .A2(n13490), .A3(n13489), .A4(n13488), .ZN(
        n13492) );
  OR4_X1 U17675 ( .A1(n13495), .A2(n13494), .A3(n13493), .A4(n13492), .ZN(
        n13519) );
  NOR2_X1 U17676 ( .A1(n13497), .A2(n13496), .ZN(n24581) );
  AOI22_X1 U17677 ( .A1(n30864), .A2(\xmem_data[64][3] ), .B1(n29253), .B2(
        \xmem_data[65][3] ), .ZN(n13501) );
  AOI22_X1 U17678 ( .A1(n24532), .A2(\xmem_data[66][3] ), .B1(n3220), .B2(
        \xmem_data[67][3] ), .ZN(n13500) );
  AOI22_X1 U17679 ( .A1(n24533), .A2(\xmem_data[68][3] ), .B1(n23739), .B2(
        \xmem_data[69][3] ), .ZN(n13499) );
  AOI22_X1 U17680 ( .A1(n24534), .A2(\xmem_data[70][3] ), .B1(n28372), .B2(
        \xmem_data[71][3] ), .ZN(n13498) );
  NAND4_X1 U17681 ( .A1(n13501), .A2(n13500), .A3(n13499), .A4(n13498), .ZN(
        n13517) );
  AOI22_X1 U17682 ( .A1(n28344), .A2(\xmem_data[72][3] ), .B1(n27446), .B2(
        \xmem_data[73][3] ), .ZN(n13505) );
  AOI22_X1 U17683 ( .A1(n28972), .A2(\xmem_data[74][3] ), .B1(n25481), .B2(
        \xmem_data[75][3] ), .ZN(n13504) );
  AOI22_X1 U17684 ( .A1(n23762), .A2(\xmem_data[76][3] ), .B1(n24516), .B2(
        \xmem_data[77][3] ), .ZN(n13503) );
  AOI22_X1 U17685 ( .A1(n3176), .A2(\xmem_data[78][3] ), .B1(n14935), .B2(
        \xmem_data[79][3] ), .ZN(n13502) );
  NAND4_X1 U17686 ( .A1(n13505), .A2(n13504), .A3(n13503), .A4(n13502), .ZN(
        n13516) );
  AOI22_X1 U17687 ( .A1(n30892), .A2(\xmem_data[80][3] ), .B1(n3213), .B2(
        \xmem_data[81][3] ), .ZN(n13509) );
  AOI22_X1 U17688 ( .A1(n24509), .A2(\xmem_data[82][3] ), .B1(n24707), .B2(
        \xmem_data[83][3] ), .ZN(n13508) );
  AOI22_X1 U17689 ( .A1(n29239), .A2(\xmem_data[84][3] ), .B1(n24510), .B2(
        \xmem_data[85][3] ), .ZN(n13507) );
  AOI22_X1 U17690 ( .A1(n24511), .A2(\xmem_data[86][3] ), .B1(n25679), .B2(
        \xmem_data[87][3] ), .ZN(n13506) );
  NAND4_X1 U17691 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        n13515) );
  AOI22_X1 U17692 ( .A1(n24522), .A2(\xmem_data[88][3] ), .B1(n24521), .B2(
        \xmem_data[89][3] ), .ZN(n13513) );
  AOI22_X1 U17693 ( .A1(n3209), .A2(\xmem_data[90][3] ), .B1(n17049), .B2(
        \xmem_data[91][3] ), .ZN(n13512) );
  AOI22_X1 U17694 ( .A1(n30674), .A2(\xmem_data[92][3] ), .B1(n24524), .B2(
        \xmem_data[93][3] ), .ZN(n13511) );
  AOI22_X1 U17695 ( .A1(n24526), .A2(\xmem_data[94][3] ), .B1(n24525), .B2(
        \xmem_data[95][3] ), .ZN(n13510) );
  NAND4_X1 U17696 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        n13514) );
  OR4_X1 U17697 ( .A1(n13517), .A2(n13516), .A3(n13515), .A4(n13514), .ZN(
        n13518) );
  AOI22_X1 U17698 ( .A1(n24542), .A2(n13519), .B1(n24581), .B2(n13518), .ZN(
        n13520) );
  AOI22_X1 U17699 ( .A1(n3318), .A2(\xmem_data[96][2] ), .B1(n27437), .B2(
        \xmem_data[97][2] ), .ZN(n13525) );
  AOI22_X1 U17700 ( .A1(n24532), .A2(\xmem_data[98][2] ), .B1(n3222), .B2(
        \xmem_data[99][2] ), .ZN(n13524) );
  AOI22_X1 U17701 ( .A1(n24533), .A2(\xmem_data[100][2] ), .B1(n20500), .B2(
        \xmem_data[101][2] ), .ZN(n13523) );
  AOI22_X1 U17702 ( .A1(n24534), .A2(\xmem_data[102][2] ), .B1(n25486), .B2(
        \xmem_data[103][2] ), .ZN(n13522) );
  NAND4_X1 U17703 ( .A1(n13525), .A2(n13524), .A3(n13523), .A4(n13522), .ZN(
        n13541) );
  AOI22_X1 U17704 ( .A1(n3345), .A2(\xmem_data[104][2] ), .B1(n28045), .B2(
        \xmem_data[105][2] ), .ZN(n13529) );
  AOI22_X1 U17705 ( .A1(n30885), .A2(\xmem_data[106][2] ), .B1(n24158), .B2(
        \xmem_data[107][2] ), .ZN(n13528) );
  AOI22_X1 U17706 ( .A1(n22738), .A2(\xmem_data[108][2] ), .B1(n24516), .B2(
        \xmem_data[109][2] ), .ZN(n13527) );
  AOI22_X1 U17707 ( .A1(n3176), .A2(\xmem_data[110][2] ), .B1(n28052), .B2(
        \xmem_data[111][2] ), .ZN(n13526) );
  NAND4_X1 U17708 ( .A1(n13529), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13540) );
  AOI22_X1 U17709 ( .A1(n20718), .A2(\xmem_data[112][2] ), .B1(n3212), .B2(
        \xmem_data[113][2] ), .ZN(n13533) );
  AOI22_X1 U17710 ( .A1(n24509), .A2(\xmem_data[114][2] ), .B1(n24459), .B2(
        \xmem_data[115][2] ), .ZN(n13532) );
  AOI22_X1 U17711 ( .A1(n14971), .A2(\xmem_data[116][2] ), .B1(n24510), .B2(
        \xmem_data[117][2] ), .ZN(n13531) );
  AOI22_X1 U17712 ( .A1(n24511), .A2(\xmem_data[118][2] ), .B1(n28291), .B2(
        \xmem_data[119][2] ), .ZN(n13530) );
  NAND4_X1 U17713 ( .A1(n13533), .A2(n13532), .A3(n13531), .A4(n13530), .ZN(
        n13539) );
  AOI22_X1 U17714 ( .A1(n24522), .A2(\xmem_data[120][2] ), .B1(n24521), .B2(
        \xmem_data[121][2] ), .ZN(n13537) );
  AOI22_X1 U17715 ( .A1(n3209), .A2(\xmem_data[122][2] ), .B1(n17049), .B2(
        \xmem_data[123][2] ), .ZN(n13536) );
  AOI22_X1 U17716 ( .A1(n20577), .A2(\xmem_data[124][2] ), .B1(n24524), .B2(
        \xmem_data[125][2] ), .ZN(n13535) );
  AOI22_X1 U17717 ( .A1(n24526), .A2(\xmem_data[126][2] ), .B1(n24525), .B2(
        \xmem_data[127][2] ), .ZN(n13534) );
  NAND4_X1 U17718 ( .A1(n13537), .A2(n13536), .A3(n13535), .A4(n13534), .ZN(
        n13538) );
  OR4_X1 U17719 ( .A1(n13541), .A2(n13540), .A3(n13539), .A4(n13538), .ZN(
        n13563) );
  AOI22_X1 U17720 ( .A1(n3153), .A2(\xmem_data[64][2] ), .B1(n27437), .B2(
        \xmem_data[65][2] ), .ZN(n13545) );
  AOI22_X1 U17721 ( .A1(n24532), .A2(\xmem_data[66][2] ), .B1(n3221), .B2(
        \xmem_data[67][2] ), .ZN(n13544) );
  AOI22_X1 U17722 ( .A1(n24533), .A2(\xmem_data[68][2] ), .B1(n27507), .B2(
        \xmem_data[69][2] ), .ZN(n13543) );
  AOI22_X1 U17723 ( .A1(n24534), .A2(\xmem_data[70][2] ), .B1(n29104), .B2(
        \xmem_data[71][2] ), .ZN(n13542) );
  NAND4_X1 U17724 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13561) );
  AOI22_X1 U17725 ( .A1(n16973), .A2(\xmem_data[72][2] ), .B1(n25514), .B2(
        \xmem_data[73][2] ), .ZN(n13549) );
  AOI22_X1 U17726 ( .A1(n27551), .A2(\xmem_data[74][2] ), .B1(n25481), .B2(
        \xmem_data[75][2] ), .ZN(n13548) );
  AOI22_X1 U17727 ( .A1(n29403), .A2(\xmem_data[76][2] ), .B1(n24516), .B2(
        \xmem_data[77][2] ), .ZN(n13547) );
  AOI22_X1 U17728 ( .A1(n28298), .A2(\xmem_data[78][2] ), .B1(n24160), .B2(
        \xmem_data[79][2] ), .ZN(n13546) );
  NAND4_X1 U17729 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13560) );
  AOI22_X1 U17730 ( .A1(n24213), .A2(\xmem_data[80][2] ), .B1(n3208), .B2(
        \xmem_data[81][2] ), .ZN(n13553) );
  AOI22_X1 U17731 ( .A1(n24509), .A2(\xmem_data[82][2] ), .B1(n21006), .B2(
        \xmem_data[83][2] ), .ZN(n13552) );
  AOI22_X1 U17732 ( .A1(n20730), .A2(\xmem_data[84][2] ), .B1(n24510), .B2(
        \xmem_data[85][2] ), .ZN(n13551) );
  AOI22_X1 U17733 ( .A1(n24511), .A2(\xmem_data[86][2] ), .B1(n30898), .B2(
        \xmem_data[87][2] ), .ZN(n13550) );
  NAND4_X1 U17734 ( .A1(n13553), .A2(n13552), .A3(n13551), .A4(n13550), .ZN(
        n13559) );
  AOI22_X1 U17735 ( .A1(n24522), .A2(\xmem_data[88][2] ), .B1(n24521), .B2(
        \xmem_data[89][2] ), .ZN(n13557) );
  AOI22_X1 U17736 ( .A1(n3209), .A2(\xmem_data[90][2] ), .B1(n27981), .B2(
        \xmem_data[91][2] ), .ZN(n13556) );
  AOI22_X1 U17737 ( .A1(n24687), .A2(\xmem_data[92][2] ), .B1(n24524), .B2(
        \xmem_data[93][2] ), .ZN(n13555) );
  AOI22_X1 U17738 ( .A1(n24526), .A2(\xmem_data[94][2] ), .B1(n24525), .B2(
        \xmem_data[95][2] ), .ZN(n13554) );
  NAND4_X1 U17739 ( .A1(n13557), .A2(n13556), .A3(n13555), .A4(n13554), .ZN(
        n13558) );
  OR4_X1 U17740 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n13562) );
  AOI22_X1 U17741 ( .A1(n24542), .A2(n13563), .B1(n24581), .B2(n13562), .ZN(
        n13614) );
  NOR2_X1 U17742 ( .A1(n22298), .A2(n39037), .ZN(n13564) );
  NAND2_X1 U17743 ( .A1(n25450), .A2(n13564), .ZN(n13613) );
  AOI22_X1 U17744 ( .A1(n28973), .A2(\xmem_data[32][2] ), .B1(n24172), .B2(
        \xmem_data[33][2] ), .ZN(n13568) );
  AOI22_X1 U17745 ( .A1(n24562), .A2(\xmem_data[34][2] ), .B1(n3218), .B2(
        \xmem_data[35][2] ), .ZN(n13567) );
  AOI22_X1 U17746 ( .A1(n24563), .A2(\xmem_data[36][2] ), .B1(n13469), .B2(
        \xmem_data[37][2] ), .ZN(n13566) );
  AOI22_X1 U17747 ( .A1(n24565), .A2(\xmem_data[38][2] ), .B1(n24564), .B2(
        \xmem_data[39][2] ), .ZN(n13565) );
  NAND4_X1 U17748 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13584) );
  AOI22_X1 U17749 ( .A1(n3375), .A2(\xmem_data[40][2] ), .B1(n24553), .B2(
        \xmem_data[41][2] ), .ZN(n13572) );
  AOI22_X1 U17750 ( .A1(n24554), .A2(\xmem_data[42][2] ), .B1(n29307), .B2(
        \xmem_data[43][2] ), .ZN(n13571) );
  AOI22_X1 U17751 ( .A1(n24556), .A2(\xmem_data[44][2] ), .B1(n24555), .B2(
        \xmem_data[45][2] ), .ZN(n13570) );
  AOI22_X1 U17752 ( .A1(n16986), .A2(\xmem_data[46][2] ), .B1(n25671), .B2(
        \xmem_data[47][2] ), .ZN(n13569) );
  NAND4_X1 U17753 ( .A1(n13572), .A2(n13571), .A3(n13570), .A4(n13569), .ZN(
        n13583) );
  AOI22_X1 U17754 ( .A1(n24545), .A2(\xmem_data[48][2] ), .B1(n28335), .B2(
        \xmem_data[49][2] ), .ZN(n13576) );
  AOI22_X1 U17755 ( .A1(n24547), .A2(\xmem_data[50][2] ), .B1(n24546), .B2(
        \xmem_data[51][2] ), .ZN(n13575) );
  AOI22_X1 U17756 ( .A1(n31255), .A2(\xmem_data[52][2] ), .B1(n25399), .B2(
        \xmem_data[53][2] ), .ZN(n13574) );
  AOI22_X1 U17757 ( .A1(n24548), .A2(\xmem_data[54][2] ), .B1(n31361), .B2(
        \xmem_data[55][2] ), .ZN(n13573) );
  NAND4_X1 U17758 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13582) );
  AOI22_X1 U17759 ( .A1(n24571), .A2(\xmem_data[56][2] ), .B1(n24570), .B2(
        \xmem_data[57][2] ), .ZN(n13580) );
  AOI22_X1 U17760 ( .A1(n24572), .A2(\xmem_data[58][2] ), .B1(n25359), .B2(
        \xmem_data[59][2] ), .ZN(n13579) );
  AOI22_X1 U17761 ( .A1(n20770), .A2(\xmem_data[60][2] ), .B1(n30498), .B2(
        \xmem_data[61][2] ), .ZN(n13578) );
  AOI22_X1 U17762 ( .A1(n20827), .A2(\xmem_data[62][2] ), .B1(n24573), .B2(
        \xmem_data[63][2] ), .ZN(n13577) );
  NAND4_X1 U17763 ( .A1(n13580), .A2(n13579), .A3(n13578), .A4(n13577), .ZN(
        n13581) );
  OR4_X1 U17764 ( .A1(n13584), .A2(n13583), .A3(n13582), .A4(n13581), .ZN(
        n13611) );
  AOI22_X1 U17765 ( .A1(n30744), .A2(\xmem_data[12][2] ), .B1(n24448), .B2(
        \xmem_data[13][2] ), .ZN(n13591) );
  AOI22_X1 U17766 ( .A1(n30614), .A2(\xmem_data[14][2] ), .B1(n30541), .B2(
        \xmem_data[15][2] ), .ZN(n13585) );
  INV_X1 U17767 ( .A(n13585), .ZN(n13589) );
  AOI22_X1 U17768 ( .A1(n24450), .A2(\xmem_data[10][2] ), .B1(n30854), .B2(
        \xmem_data[11][2] ), .ZN(n13587) );
  NAND2_X1 U17769 ( .A1(n28308), .A2(\xmem_data[8][2] ), .ZN(n13586) );
  NAND2_X1 U17770 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  NOR2_X1 U17771 ( .A1(n13589), .A2(n13588), .ZN(n13590) );
  NAND2_X1 U17772 ( .A1(n13591), .A2(n13590), .ZN(n13602) );
  AOI22_X1 U17773 ( .A1(n24458), .A2(\xmem_data[16][2] ), .B1(n24457), .B2(
        \xmem_data[17][2] ), .ZN(n13595) );
  AOI22_X1 U17774 ( .A1(n24133), .A2(\xmem_data[18][2] ), .B1(n24459), .B2(
        \xmem_data[19][2] ), .ZN(n13594) );
  AOI22_X1 U17775 ( .A1(n29410), .A2(\xmem_data[20][2] ), .B1(n24460), .B2(
        \xmem_data[21][2] ), .ZN(n13593) );
  AOI22_X1 U17776 ( .A1(n3178), .A2(\xmem_data[22][2] ), .B1(n25364), .B2(
        \xmem_data[23][2] ), .ZN(n13592) );
  NAND4_X1 U17777 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13601) );
  AOI22_X1 U17778 ( .A1(n24630), .A2(\xmem_data[0][2] ), .B1(n24439), .B2(
        \xmem_data[1][2] ), .ZN(n13599) );
  AOI22_X1 U17779 ( .A1(n24443), .A2(\xmem_data[2][2] ), .B1(n3222), .B2(
        \xmem_data[3][2] ), .ZN(n13598) );
  AOI22_X1 U17780 ( .A1(n24696), .A2(\xmem_data[4][2] ), .B1(n28476), .B2(
        \xmem_data[5][2] ), .ZN(n13597) );
  AOI22_X1 U17781 ( .A1(n24438), .A2(\xmem_data[6][2] ), .B1(n29181), .B2(
        \xmem_data[7][2] ), .ZN(n13596) );
  NAND4_X1 U17782 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13600) );
  OR3_X1 U17783 ( .A1(n13602), .A2(n13601), .A3(n13600), .ZN(n13608) );
  AOI22_X1 U17784 ( .A1(n3338), .A2(\xmem_data[24][2] ), .B1(n25583), .B2(
        \xmem_data[25][2] ), .ZN(n13606) );
  AOI22_X1 U17785 ( .A1(n24467), .A2(\xmem_data[26][2] ), .B1(n27526), .B2(
        \xmem_data[27][2] ), .ZN(n13605) );
  AOI22_X1 U17786 ( .A1(n24687), .A2(\xmem_data[28][2] ), .B1(n24468), .B2(
        \xmem_data[29][2] ), .ZN(n13604) );
  AOI22_X1 U17787 ( .A1(n27500), .A2(\xmem_data[30][2] ), .B1(n24470), .B2(
        \xmem_data[31][2] ), .ZN(n13603) );
  NAND4_X1 U17788 ( .A1(n13606), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        n13607) );
  NOR2_X1 U17789 ( .A1(n13608), .A2(n13607), .ZN(n13609) );
  INV_X1 U17790 ( .A(n22180), .ZN(n22298) );
  NOR2_X1 U17791 ( .A1(n13609), .A2(n22298), .ZN(n13610) );
  AOI21_X1 U17792 ( .B1(n13611), .B2(n24508), .A(n13610), .ZN(n13612) );
  NAND3_X1 U17793 ( .A1(n13614), .A2(n13613), .A3(n13612), .ZN(n32005) );
  XNOR2_X1 U17794 ( .A(n32005), .B(\fmem_data[16][7] ), .ZN(n17851) );
  XOR2_X1 U17795 ( .A(\fmem_data[16][6] ), .B(\fmem_data[16][7] ), .Z(n13615)
         );
  AOI22_X1 U17796 ( .A1(n28291), .A2(\xmem_data[0][3] ), .B1(n30686), .B2(
        \xmem_data[1][3] ), .ZN(n13619) );
  AOI22_X1 U17797 ( .A1(n27365), .A2(\xmem_data[2][3] ), .B1(n25526), .B2(
        \xmem_data[3][3] ), .ZN(n13618) );
  AOI22_X1 U17798 ( .A1(n29136), .A2(\xmem_data[4][3] ), .B1(n29657), .B2(
        \xmem_data[5][3] ), .ZN(n13617) );
  AOI22_X1 U17799 ( .A1(n29125), .A2(\xmem_data[6][3] ), .B1(n29124), .B2(
        \xmem_data[7][3] ), .ZN(n13616) );
  AND4_X1 U17800 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13635) );
  AOI22_X1 U17801 ( .A1(n29118), .A2(\xmem_data[8][3] ), .B1(n28164), .B2(
        \xmem_data[9][3] ), .ZN(n13623) );
  AOI22_X1 U17802 ( .A1(n3247), .A2(\xmem_data[10][3] ), .B1(n28082), .B2(
        \xmem_data[11][3] ), .ZN(n13622) );
  AOI22_X1 U17803 ( .A1(n3221), .A2(\xmem_data[12][3] ), .B1(n29422), .B2(
        \xmem_data[13][3] ), .ZN(n13621) );
  AOI22_X1 U17804 ( .A1(n25562), .A2(\xmem_data[14][3] ), .B1(n29257), .B2(
        \xmem_data[15][3] ), .ZN(n13620) );
  AND4_X1 U17805 ( .A1(n13623), .A2(n13622), .A3(n13621), .A4(n13620), .ZN(
        n13634) );
  AOI22_X1 U17806 ( .A1(n24633), .A2(\xmem_data[16][3] ), .B1(n29350), .B2(
        \xmem_data[17][3] ), .ZN(n13627) );
  AOI22_X1 U17807 ( .A1(n28045), .A2(\xmem_data[18][3] ), .B1(n25670), .B2(
        \xmem_data[19][3] ), .ZN(n13626) );
  AOI22_X1 U17808 ( .A1(n30854), .A2(\xmem_data[20][3] ), .B1(n29591), .B2(
        \xmem_data[21][3] ), .ZN(n13625) );
  AOI22_X1 U17809 ( .A1(n24212), .A2(\xmem_data[22][3] ), .B1(n28334), .B2(
        \xmem_data[23][3] ), .ZN(n13624) );
  AND4_X1 U17810 ( .A1(n13627), .A2(n13626), .A3(n13625), .A4(n13624), .ZN(
        n13633) );
  AOI22_X1 U17811 ( .A1(n29279), .A2(\xmem_data[26][3] ), .B1(n29317), .B2(
        \xmem_data[27][3] ), .ZN(n13631) );
  AOI22_X1 U17812 ( .A1(n22703), .A2(\xmem_data[24][3] ), .B1(n29187), .B2(
        \xmem_data[25][3] ), .ZN(n13630) );
  AOI22_X1 U17813 ( .A1(n28492), .A2(\xmem_data[28][3] ), .B1(n28781), .B2(
        \xmem_data[29][3] ), .ZN(n13629) );
  AOI22_X1 U17814 ( .A1(n29190), .A2(\xmem_data[30][3] ), .B1(n17002), .B2(
        \xmem_data[31][3] ), .ZN(n13628) );
  AND4_X1 U17815 ( .A1(n13631), .A2(n13630), .A3(n13629), .A4(n13628), .ZN(
        n13632) );
  NAND4_X1 U17816 ( .A1(n13635), .A2(n13634), .A3(n13633), .A4(n13632), .ZN(
        n13636) );
  AOI22_X1 U17817 ( .A1(n25514), .A2(\xmem_data[82][3] ), .B1(n31276), .B2(
        \xmem_data[83][3] ), .ZN(n13662) );
  AOI22_X1 U17818 ( .A1(n27567), .A2(\xmem_data[70][3] ), .B1(n24688), .B2(
        \xmem_data[71][3] ), .ZN(n13641) );
  AOI22_X1 U17819 ( .A1(n29126), .A2(\xmem_data[66][3] ), .B1(n3209), .B2(
        \xmem_data[67][3] ), .ZN(n13640) );
  AOI22_X1 U17820 ( .A1(n28494), .A2(\xmem_data[64][3] ), .B1(n29324), .B2(
        \xmem_data[65][3] ), .ZN(n13639) );
  AND2_X1 U17821 ( .A1(n21057), .A2(\xmem_data[68][3] ), .ZN(n13637) );
  AOI21_X1 U17822 ( .B1(n27717), .B2(\xmem_data[69][3] ), .A(n13637), .ZN(
        n13638) );
  NAND4_X1 U17823 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13645) );
  AOI22_X1 U17824 ( .A1(n29181), .A2(\xmem_data[80][3] ), .B1(n29157), .B2(
        \xmem_data[81][3] ), .ZN(n13643) );
  AOI22_X1 U17825 ( .A1(n20775), .A2(\xmem_data[86][3] ), .B1(n30614), .B2(
        \xmem_data[87][3] ), .ZN(n13642) );
  NAND2_X1 U17826 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  AOI22_X1 U17827 ( .A1(n30861), .A2(\xmem_data[72][3] ), .B1(n28245), .B2(
        \xmem_data[73][3] ), .ZN(n13649) );
  AOI22_X1 U17828 ( .A1(n29173), .A2(\xmem_data[74][3] ), .B1(n28318), .B2(
        \xmem_data[75][3] ), .ZN(n13648) );
  AOI22_X1 U17829 ( .A1(n3220), .A2(\xmem_data[76][3] ), .B1(n29256), .B2(
        \xmem_data[77][3] ), .ZN(n13647) );
  AOI22_X1 U17830 ( .A1(n30963), .A2(\xmem_data[78][3] ), .B1(n29174), .B2(
        \xmem_data[79][3] ), .ZN(n13646) );
  AND4_X1 U17831 ( .A1(n13649), .A2(n13648), .A3(n13647), .A4(n13646), .ZN(
        n13658) );
  AOI22_X1 U17832 ( .A1(n29162), .A2(\xmem_data[90][3] ), .B1(n20585), .B2(
        \xmem_data[91][3] ), .ZN(n13653) );
  AOI22_X1 U17833 ( .A1(n24160), .A2(\xmem_data[88][3] ), .B1(n29187), .B2(
        \xmem_data[89][3] ), .ZN(n13652) );
  AOI22_X1 U17834 ( .A1(n29048), .A2(\xmem_data[92][3] ), .B1(n21050), .B2(
        \xmem_data[93][3] ), .ZN(n13651) );
  AOI22_X1 U17835 ( .A1(n29190), .A2(\xmem_data[94][3] ), .B1(n3205), .B2(
        \xmem_data[95][3] ), .ZN(n13650) );
  NAND4_X1 U17836 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13656) );
  AOI22_X1 U17837 ( .A1(n29180), .A2(\xmem_data[84][3] ), .B1(n29179), .B2(
        \xmem_data[85][3] ), .ZN(n13654) );
  INV_X1 U17838 ( .A(n13654), .ZN(n13655) );
  NOR2_X1 U17839 ( .A1(n13656), .A2(n13655), .ZN(n13657) );
  NAND2_X1 U17840 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  NOR2_X1 U17841 ( .A1(n3968), .A2(n13659), .ZN(n13661) );
  INV_X1 U17842 ( .A(n29201), .ZN(n13660) );
  AOI21_X1 U17843 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13714) );
  AOI22_X1 U17844 ( .A1(n28045), .A2(\xmem_data[114][3] ), .B1(n24554), .B2(
        \xmem_data[115][3] ), .ZN(n13686) );
  AOI22_X1 U17845 ( .A1(n24457), .A2(\xmem_data[122][3] ), .B1(n25573), .B2(
        \xmem_data[123][3] ), .ZN(n13666) );
  AOI22_X1 U17846 ( .A1(n22741), .A2(\xmem_data[120][3] ), .B1(n3464), .B2(
        \xmem_data[121][3] ), .ZN(n13665) );
  AOI22_X1 U17847 ( .A1(n29316), .A2(\xmem_data[124][3] ), .B1(n29410), .B2(
        \xmem_data[125][3] ), .ZN(n13664) );
  AOI22_X1 U17848 ( .A1(n29190), .A2(\xmem_data[126][3] ), .B1(n3206), .B2(
        \xmem_data[127][3] ), .ZN(n13663) );
  NAND4_X1 U17849 ( .A1(n13666), .A2(n13665), .A3(n13664), .A4(n13663), .ZN(
        n13683) );
  AOI22_X1 U17850 ( .A1(n29180), .A2(\xmem_data[116][3] ), .B1(n29179), .B2(
        \xmem_data[117][3] ), .ZN(n13681) );
  AOI22_X1 U17851 ( .A1(n31262), .A2(\xmem_data[104][3] ), .B1(n3413), .B2(
        \xmem_data[105][3] ), .ZN(n13670) );
  AOI22_X1 U17852 ( .A1(n29173), .A2(\xmem_data[106][3] ), .B1(n30503), .B2(
        \xmem_data[107][3] ), .ZN(n13669) );
  AOI22_X1 U17853 ( .A1(n3219), .A2(\xmem_data[108][3] ), .B1(n25612), .B2(
        \xmem_data[109][3] ), .ZN(n13668) );
  AOI22_X1 U17854 ( .A1(n25491), .A2(\xmem_data[110][3] ), .B1(n29174), .B2(
        \xmem_data[111][3] ), .ZN(n13667) );
  AND4_X1 U17855 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13680) );
  AOI22_X1 U17856 ( .A1(n25679), .A2(\xmem_data[96][3] ), .B1(n28461), .B2(
        \xmem_data[97][3] ), .ZN(n13674) );
  AOI22_X1 U17857 ( .A1(n29126), .A2(\xmem_data[98][3] ), .B1(n29151), .B2(
        \xmem_data[99][3] ), .ZN(n13673) );
  AOI22_X1 U17858 ( .A1(n28500), .A2(\xmem_data[100][3] ), .B1(n25684), .B2(
        \xmem_data[101][3] ), .ZN(n13672) );
  AOI22_X1 U17859 ( .A1(n20769), .A2(\xmem_data[102][3] ), .B1(n21061), .B2(
        \xmem_data[103][3] ), .ZN(n13671) );
  NAND4_X1 U17860 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13678) );
  AOI22_X1 U17861 ( .A1(n29181), .A2(\xmem_data[112][3] ), .B1(n30295), .B2(
        \xmem_data[113][3] ), .ZN(n13676) );
  AOI22_X1 U17862 ( .A1(n22675), .A2(\xmem_data[118][3] ), .B1(n30514), .B2(
        \xmem_data[119][3] ), .ZN(n13675) );
  NAND2_X1 U17863 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  NOR2_X1 U17864 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  NAND3_X1 U17865 ( .A1(n13681), .A2(n13680), .A3(n13679), .ZN(n13682) );
  NOR2_X1 U17866 ( .A1(n13683), .A2(n13682), .ZN(n13685) );
  INV_X1 U17867 ( .A(n29171), .ZN(n13684) );
  AOI21_X1 U17868 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13713) );
  AOI22_X1 U17869 ( .A1(n22739), .A2(\xmem_data[52][3] ), .B1(n30083), .B2(
        \xmem_data[53][3] ), .ZN(n13702) );
  AOI22_X1 U17870 ( .A1(n28366), .A2(\xmem_data[40][3] ), .B1(n28245), .B2(
        \xmem_data[41][3] ), .ZN(n13690) );
  AOI22_X1 U17871 ( .A1(n31347), .A2(\xmem_data[42][3] ), .B1(n24443), .B2(
        \xmem_data[43][3] ), .ZN(n13689) );
  AOI22_X1 U17872 ( .A1(n3217), .A2(\xmem_data[44][3] ), .B1(n27831), .B2(
        \xmem_data[45][3] ), .ZN(n13688) );
  AOI22_X1 U17873 ( .A1(n29095), .A2(\xmem_data[46][3] ), .B1(n3342), .B2(
        \xmem_data[47][3] ), .ZN(n13687) );
  AND4_X1 U17874 ( .A1(n13690), .A2(n13689), .A3(n13688), .A4(n13687), .ZN(
        n13701) );
  AOI22_X1 U17875 ( .A1(n29089), .A2(\xmem_data[32][3] ), .B1(n29816), .B2(
        \xmem_data[33][3] ), .ZN(n13695) );
  AOI22_X1 U17876 ( .A1(n29126), .A2(\xmem_data[34][3] ), .B1(n29151), .B2(
        \xmem_data[35][3] ), .ZN(n13694) );
  AND2_X1 U17877 ( .A1(n29086), .A2(\xmem_data[36][3] ), .ZN(n13691) );
  AOI21_X1 U17878 ( .B1(n28772), .B2(\xmem_data[37][3] ), .A(n13691), .ZN(
        n13693) );
  AOI22_X1 U17879 ( .A1(n16999), .A2(\xmem_data[38][3] ), .B1(n20827), .B2(
        \xmem_data[39][3] ), .ZN(n13692) );
  NAND4_X1 U17880 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13699) );
  AOI22_X1 U17881 ( .A1(n29104), .A2(\xmem_data[48][3] ), .B1(n3138), .B2(
        \xmem_data[49][3] ), .ZN(n13697) );
  AOI22_X1 U17882 ( .A1(n13168), .A2(\xmem_data[54][3] ), .B1(n29109), .B2(
        \xmem_data[55][3] ), .ZN(n13696) );
  NAND2_X1 U17883 ( .A1(n13697), .A2(n13696), .ZN(n13698) );
  NOR2_X1 U17884 ( .A1(n13699), .A2(n13698), .ZN(n13700) );
  AOI22_X1 U17885 ( .A1(n29188), .A2(\xmem_data[58][3] ), .B1(n17020), .B2(
        \xmem_data[59][3] ), .ZN(n13706) );
  AOI22_X1 U17886 ( .A1(n28090), .A2(\xmem_data[56][3] ), .B1(n29187), .B2(
        \xmem_data[57][3] ), .ZN(n13705) );
  AOI22_X1 U17887 ( .A1(n27518), .A2(\xmem_data[60][3] ), .B1(n28232), .B2(
        \xmem_data[61][3] ), .ZN(n13704) );
  AOI22_X1 U17888 ( .A1(n29101), .A2(\xmem_data[62][3] ), .B1(n28460), .B2(
        \xmem_data[63][3] ), .ZN(n13703) );
  NAND4_X1 U17889 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13709) );
  AOI22_X1 U17890 ( .A1(n29103), .A2(\xmem_data[50][3] ), .B1(n27910), .B2(
        \xmem_data[51][3] ), .ZN(n13707) );
  INV_X1 U17891 ( .A(n13707), .ZN(n13708) );
  NOR2_X1 U17892 ( .A1(n13709), .A2(n13708), .ZN(n13711) );
  INV_X1 U17893 ( .A(n29145), .ZN(n13710) );
  AOI21_X1 U17894 ( .B1(n3887), .B2(n13711), .A(n13710), .ZN(n13712) );
  AOI22_X1 U17895 ( .A1(n29118), .A2(\xmem_data[8][2] ), .B1(n28245), .B2(
        \xmem_data[9][2] ), .ZN(n13718) );
  AOI22_X1 U17896 ( .A1(n3247), .A2(\xmem_data[10][2] ), .B1(n28355), .B2(
        \xmem_data[11][2] ), .ZN(n13717) );
  AOI22_X1 U17897 ( .A1(n3217), .A2(\xmem_data[12][2] ), .B1(n29627), .B2(
        \xmem_data[13][2] ), .ZN(n13716) );
  AOI22_X1 U17898 ( .A1(n23739), .A2(\xmem_data[14][2] ), .B1(n22666), .B2(
        \xmem_data[15][2] ), .ZN(n13715) );
  NAND4_X1 U17899 ( .A1(n13718), .A2(n13717), .A3(n13716), .A4(n13715), .ZN(
        n13739) );
  AOI22_X1 U17900 ( .A1(n27536), .A2(\xmem_data[24][2] ), .B1(n24458), .B2(
        \xmem_data[25][2] ), .ZN(n13722) );
  AOI22_X1 U17901 ( .A1(n29188), .A2(\xmem_data[26][2] ), .B1(n25573), .B2(
        \xmem_data[27][2] ), .ZN(n13721) );
  AOI22_X1 U17902 ( .A1(n23796), .A2(\xmem_data[28][2] ), .B1(n29239), .B2(
        \xmem_data[29][2] ), .ZN(n13720) );
  AOI22_X1 U17903 ( .A1(n24510), .A2(\xmem_data[30][2] ), .B1(n20593), .B2(
        \xmem_data[31][2] ), .ZN(n13719) );
  AOI22_X1 U17904 ( .A1(n29306), .A2(\xmem_data[18][2] ), .B1(n27551), .B2(
        \xmem_data[19][2] ), .ZN(n13737) );
  NAND2_X1 U17905 ( .A1(n25628), .A2(\xmem_data[5][2] ), .ZN(n13724) );
  NAND2_X1 U17906 ( .A1(n29136), .A2(\xmem_data[4][2] ), .ZN(n13723) );
  NAND2_X1 U17907 ( .A1(n13724), .A2(n13723), .ZN(n13729) );
  AOI22_X1 U17908 ( .A1(n25716), .A2(\xmem_data[0][2] ), .B1(n3270), .B2(
        \xmem_data[1][2] ), .ZN(n13727) );
  AOI22_X1 U17909 ( .A1(n29126), .A2(\xmem_data[2][2] ), .B1(n29151), .B2(
        \xmem_data[3][2] ), .ZN(n13726) );
  AOI22_X1 U17910 ( .A1(n29125), .A2(\xmem_data[6][2] ), .B1(n29124), .B2(
        \xmem_data[7][2] ), .ZN(n13725) );
  NOR2_X1 U17911 ( .A1(n13729), .A2(n13728), .ZN(n13736) );
  AOI22_X1 U17912 ( .A1(n25456), .A2(\xmem_data[20][2] ), .B1(n31353), .B2(
        \xmem_data[21][2] ), .ZN(n13731) );
  AOI22_X1 U17913 ( .A1(n3256), .A2(\xmem_data[16][2] ), .B1(n27396), .B2(
        \xmem_data[17][2] ), .ZN(n13730) );
  NAND2_X1 U17914 ( .A1(n13731), .A2(n13730), .ZN(n13734) );
  AOI22_X1 U17915 ( .A1(n28515), .A2(\xmem_data[22][2] ), .B1(n20959), .B2(
        \xmem_data[23][2] ), .ZN(n13732) );
  INV_X1 U17916 ( .A(n13732), .ZN(n13733) );
  NOR2_X1 U17917 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NAND4_X1 U17918 ( .A1(n3832), .A2(n13737), .A3(n13736), .A4(n13735), .ZN(
        n13738) );
  OAI21_X1 U17919 ( .B1(n13739), .B2(n13738), .A(n29143), .ZN(n13813) );
  AOI22_X1 U17920 ( .A1(n20568), .A2(\xmem_data[42][2] ), .B1(n23756), .B2(
        \xmem_data[43][2] ), .ZN(n13743) );
  AOI22_X1 U17921 ( .A1(n22729), .A2(\xmem_data[40][2] ), .B1(n3318), .B2(
        \xmem_data[41][2] ), .ZN(n13742) );
  AOI22_X1 U17922 ( .A1(n3218), .A2(\xmem_data[44][2] ), .B1(n29431), .B2(
        \xmem_data[45][2] ), .ZN(n13741) );
  AOI22_X1 U17923 ( .A1(n29095), .A2(\xmem_data[46][2] ), .B1(n23812), .B2(
        \xmem_data[47][2] ), .ZN(n13740) );
  NAND4_X1 U17924 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13761) );
  AOI22_X1 U17925 ( .A1(n29089), .A2(\xmem_data[32][2] ), .B1(n30269), .B2(
        \xmem_data[33][2] ), .ZN(n13748) );
  AOI22_X1 U17926 ( .A1(n24622), .A2(\xmem_data[34][2] ), .B1(n27542), .B2(
        \xmem_data[35][2] ), .ZN(n13747) );
  AND2_X1 U17927 ( .A1(n29086), .A2(\xmem_data[36][2] ), .ZN(n13744) );
  AOI21_X1 U17928 ( .B1(n27568), .B2(\xmem_data[37][2] ), .A(n13744), .ZN(
        n13746) );
  AOI22_X1 U17929 ( .A1(n24468), .A2(\xmem_data[38][2] ), .B1(n25630), .B2(
        \xmem_data[39][2] ), .ZN(n13745) );
  NAND4_X1 U17930 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13759) );
  AOI22_X1 U17931 ( .A1(n24457), .A2(\xmem_data[58][2] ), .B1(n24214), .B2(
        \xmem_data[59][2] ), .ZN(n13752) );
  AOI22_X1 U17932 ( .A1(n25520), .A2(\xmem_data[60][2] ), .B1(n30950), .B2(
        \xmem_data[61][2] ), .ZN(n13751) );
  AOI22_X1 U17933 ( .A1(n24548), .A2(\xmem_data[63][2] ), .B1(
        \xmem_data[62][2] ), .B2(n29101), .ZN(n13750) );
  AOI22_X1 U17934 ( .A1(n27536), .A2(\xmem_data[56][2] ), .B1(n30666), .B2(
        \xmem_data[57][2] ), .ZN(n13749) );
  NAND4_X1 U17935 ( .A1(n13752), .A2(n13751), .A3(n13750), .A4(n13749), .ZN(
        n13758) );
  AOI22_X1 U17936 ( .A1(n24212), .A2(\xmem_data[54][2] ), .B1(n29109), .B2(
        \xmem_data[55][2] ), .ZN(n13756) );
  AOI22_X1 U17937 ( .A1(n29103), .A2(\xmem_data[50][2] ), .B1(n28050), .B2(
        \xmem_data[51][2] ), .ZN(n13755) );
  AOI22_X1 U17938 ( .A1(n28373), .A2(\xmem_data[52][2] ), .B1(n27514), .B2(
        \xmem_data[53][2] ), .ZN(n13754) );
  AOI22_X1 U17939 ( .A1(n29104), .A2(\xmem_data[48][2] ), .B1(n29157), .B2(
        \xmem_data[49][2] ), .ZN(n13753) );
  NAND4_X1 U17940 ( .A1(n13756), .A2(n13755), .A3(n13754), .A4(n13753), .ZN(
        n13757) );
  OR3_X1 U17941 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(n13760) );
  OAI21_X1 U17942 ( .B1(n13761), .B2(n13760), .A(n29145), .ZN(n13812) );
  AOI22_X1 U17943 ( .A1(n29009), .A2(\xmem_data[120][2] ), .B1(n27517), .B2(
        \xmem_data[121][2] ), .ZN(n13765) );
  AOI22_X1 U17944 ( .A1(n31269), .A2(\xmem_data[122][2] ), .B1(n25635), .B2(
        \xmem_data[123][2] ), .ZN(n13764) );
  AOI22_X1 U17945 ( .A1(n27518), .A2(\xmem_data[124][2] ), .B1(n20815), .B2(
        \xmem_data[125][2] ), .ZN(n13763) );
  AOI22_X1 U17946 ( .A1(n29190), .A2(\xmem_data[126][2] ), .B1(n3205), .B2(
        \xmem_data[127][2] ), .ZN(n13762) );
  AOI22_X1 U17947 ( .A1(n24555), .A2(\xmem_data[118][2] ), .B1(n25567), .B2(
        \xmem_data[119][2] ), .ZN(n13769) );
  AOI22_X1 U17948 ( .A1(n30877), .A2(\xmem_data[114][2] ), .B1(n27551), .B2(
        \xmem_data[115][2] ), .ZN(n13768) );
  AOI22_X1 U17949 ( .A1(n29180), .A2(\xmem_data[116][2] ), .B1(n29179), .B2(
        \xmem_data[117][2] ), .ZN(n13767) );
  AOI22_X1 U17950 ( .A1(n29181), .A2(\xmem_data[112][2] ), .B1(n27396), .B2(
        \xmem_data[113][2] ), .ZN(n13766) );
  AOI22_X1 U17951 ( .A1(n21051), .A2(\xmem_data[96][2] ), .B1(n30600), .B2(
        \xmem_data[97][2] ), .ZN(n13770) );
  INV_X1 U17952 ( .A(n13770), .ZN(n13774) );
  AOI22_X1 U17953 ( .A1(n31344), .A2(\xmem_data[102][2] ), .B1(n20710), .B2(
        \xmem_data[103][2] ), .ZN(n13772) );
  AOI22_X1 U17954 ( .A1(n29126), .A2(\xmem_data[98][2] ), .B1(n20782), .B2(
        \xmem_data[99][2] ), .ZN(n13771) );
  NAND2_X1 U17955 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  NOR2_X1 U17956 ( .A1(n13774), .A2(n13773), .ZN(n13776) );
  AOI22_X1 U17957 ( .A1(n30496), .A2(\xmem_data[100][2] ), .B1(n21060), .B2(
        \xmem_data[101][2] ), .ZN(n13775) );
  NAND4_X1 U17958 ( .A1(n3829), .A2(n3535), .A3(n13776), .A4(n13775), .ZN(
        n13783) );
  AOI22_X1 U17959 ( .A1(n24470), .A2(\xmem_data[104][2] ), .B1(n3388), .B2(
        \xmem_data[105][2] ), .ZN(n13781) );
  AND2_X1 U17960 ( .A1(n29173), .A2(\xmem_data[106][2] ), .ZN(n13777) );
  AOI21_X1 U17961 ( .B1(n23734), .B2(\xmem_data[107][2] ), .A(n13777), .ZN(
        n13780) );
  AOI22_X1 U17962 ( .A1(n3219), .A2(\xmem_data[108][2] ), .B1(n24696), .B2(
        \xmem_data[109][2] ), .ZN(n13779) );
  AOI22_X1 U17963 ( .A1(n23739), .A2(\xmem_data[110][2] ), .B1(n29174), .B2(
        \xmem_data[111][2] ), .ZN(n13778) );
  NAND4_X1 U17964 ( .A1(n13781), .A2(n13780), .A3(n13779), .A4(n13778), .ZN(
        n13782) );
  OAI21_X1 U17965 ( .B1(n13783), .B2(n13782), .A(n29171), .ZN(n13811) );
  AOI22_X1 U17966 ( .A1(n21015), .A2(\xmem_data[86][2] ), .B1(n25710), .B2(
        \xmem_data[87][2] ), .ZN(n13785) );
  AOI22_X1 U17967 ( .A1(n29173), .A2(\xmem_data[74][2] ), .B1(
        \xmem_data[73][2] ), .B2(n3384), .ZN(n13784) );
  NAND2_X1 U17968 ( .A1(n13784), .A2(n13785), .ZN(n13788) );
  AOI22_X1 U17969 ( .A1(n25581), .A2(\xmem_data[64][2] ), .B1(n31315), .B2(
        \xmem_data[65][2] ), .ZN(n13786) );
  INV_X1 U17970 ( .A(n13786), .ZN(n13787) );
  NOR2_X1 U17971 ( .A1(n13788), .A2(n13787), .ZN(n13797) );
  AOI22_X1 U17972 ( .A1(n20488), .A2(\xmem_data[68][2] ), .B1(n29383), .B2(
        \xmem_data[69][2] ), .ZN(n13796) );
  AOI22_X1 U17973 ( .A1(n23734), .A2(\xmem_data[75][2] ), .B1(n28037), .B2(
        \xmem_data[72][2] ), .ZN(n13795) );
  AOI22_X1 U17974 ( .A1(n20769), .A2(\xmem_data[70][2] ), .B1(n25408), .B2(
        \xmem_data[71][2] ), .ZN(n13789) );
  INV_X1 U17975 ( .A(n13789), .ZN(n13793) );
  AOI22_X1 U17976 ( .A1(n23739), .A2(\xmem_data[78][2] ), .B1(n29174), .B2(
        \xmem_data[79][2] ), .ZN(n13791) );
  AOI22_X1 U17977 ( .A1(n27365), .A2(\xmem_data[66][2] ), .B1(n27847), .B2(
        \xmem_data[67][2] ), .ZN(n13790) );
  NAND2_X1 U17978 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  NOR2_X1 U17979 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  NAND4_X1 U17980 ( .A1(n13797), .A2(n13796), .A3(n13795), .A4(n13794), .ZN(
        n13809) );
  AOI22_X1 U17981 ( .A1(n30541), .A2(\xmem_data[88][2] ), .B1(n3466), .B2(
        \xmem_data[89][2] ), .ZN(n13801) );
  AOI22_X1 U17982 ( .A1(n29162), .A2(\xmem_data[90][2] ), .B1(n25635), .B2(
        \xmem_data[91][2] ), .ZN(n13800) );
  AOI22_X1 U17983 ( .A1(n25398), .A2(\xmem_data[92][2] ), .B1(n20730), .B2(
        \xmem_data[93][2] ), .ZN(n13799) );
  AOI22_X1 U17984 ( .A1(n29190), .A2(\xmem_data[94][2] ), .B1(n3206), .B2(
        \xmem_data[95][2] ), .ZN(n13798) );
  NAND4_X1 U17985 ( .A1(n13801), .A2(n13800), .A3(n13799), .A4(n13798), .ZN(
        n13807) );
  AOI22_X1 U17986 ( .A1(n29180), .A2(\xmem_data[84][2] ), .B1(n29179), .B2(
        \xmem_data[85][2] ), .ZN(n13805) );
  AOI22_X1 U17987 ( .A1(n28045), .A2(\xmem_data[82][2] ), .B1(n27447), .B2(
        \xmem_data[83][2] ), .ZN(n13804) );
  AOI22_X1 U17988 ( .A1(n29181), .A2(\xmem_data[80][2] ), .B1(n27396), .B2(
        \xmem_data[81][2] ), .ZN(n13803) );
  AOI22_X1 U17989 ( .A1(n3221), .A2(\xmem_data[76][2] ), .B1(n29256), .B2(
        \xmem_data[77][2] ), .ZN(n13802) );
  NAND4_X1 U17990 ( .A1(n13805), .A2(n13804), .A3(n13803), .A4(n13802), .ZN(
        n13806) );
  OR2_X1 U17991 ( .A1(n13807), .A2(n13806), .ZN(n13808) );
  OAI21_X1 U17992 ( .B1(n13809), .B2(n13808), .A(n29201), .ZN(n13810) );
  XNOR2_X1 U17993 ( .A(n32513), .B(\fmem_data[25][7] ), .ZN(n30394) );
  XOR2_X1 U17994 ( .A(\fmem_data[25][6] ), .B(\fmem_data[25][7] ), .Z(n13814)
         );
  OAI22_X1 U17995 ( .A1(n33247), .A2(n35745), .B1(n30394), .B2(n35744), .ZN(
        n19510) );
  NAND2_X1 U17996 ( .A1(n25425), .A2(\xmem_data[4][5] ), .ZN(n13826) );
  AOI22_X1 U17997 ( .A1(n14976), .A2(\xmem_data[16][5] ), .B1(n28500), .B2(
        \xmem_data[17][5] ), .ZN(n13818) );
  AOI22_X1 U17998 ( .A1(n25628), .A2(\xmem_data[18][5] ), .B1(n30498), .B2(
        \xmem_data[19][5] ), .ZN(n13817) );
  AOI22_X1 U17999 ( .A1(n25630), .A2(\xmem_data[20][5] ), .B1(n25629), .B2(
        \xmem_data[21][5] ), .ZN(n13816) );
  AOI22_X1 U18000 ( .A1(n25624), .A2(\xmem_data[22][5] ), .B1(n3247), .B2(
        \xmem_data[23][5] ), .ZN(n13815) );
  NAND4_X1 U18001 ( .A1(n13818), .A2(n13817), .A3(n13816), .A4(n13815), .ZN(
        n13824) );
  AOI22_X1 U18002 ( .A1(n29451), .A2(\xmem_data[2][5] ), .B1(n25605), .B2(
        \xmem_data[3][5] ), .ZN(n13822) );
  AOI22_X1 U18003 ( .A1(n3158), .A2(\xmem_data[6][5] ), .B1(n29162), .B2(
        \xmem_data[7][5] ), .ZN(n13820) );
  AOI22_X1 U18004 ( .A1(n25606), .A2(\xmem_data[5][5] ), .B1(\xmem_data[1][5] ), .B2(n20546), .ZN(n13819) );
  AND2_X1 U18005 ( .A1(n13820), .A2(n13819), .ZN(n13821) );
  NAND2_X1 U18006 ( .A1(n13822), .A2(n13821), .ZN(n13823) );
  NOR2_X1 U18007 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  NAND2_X1 U18008 ( .A1(n13826), .A2(n13825), .ZN(n13844) );
  NAND2_X1 U18009 ( .A1(n28364), .A2(\xmem_data[24][5] ), .ZN(n13828) );
  NAND2_X1 U18010 ( .A1(n3222), .A2(\xmem_data[25][5] ), .ZN(n13827) );
  NAND2_X1 U18011 ( .A1(n13828), .A2(n13827), .ZN(n13833) );
  AOI22_X1 U18012 ( .A1(n25617), .A2(\xmem_data[28][5] ), .B1(n25616), .B2(
        \xmem_data[29][5] ), .ZN(n13831) );
  NAND2_X1 U18013 ( .A1(n25604), .A2(\xmem_data[0][5] ), .ZN(n13830) );
  NAND2_X1 U18014 ( .A1(n30295), .A2(\xmem_data[30][5] ), .ZN(n13829) );
  NAND3_X1 U18015 ( .A1(n13831), .A2(n13830), .A3(n13829), .ZN(n13832) );
  NOR2_X1 U18016 ( .A1(n13833), .A2(n13832), .ZN(n13842) );
  AOI22_X1 U18017 ( .A1(n25635), .A2(\xmem_data[8][5] ), .B1(n30544), .B2(
        \xmem_data[9][5] ), .ZN(n13837) );
  AOI22_X1 U18018 ( .A1(n30309), .A2(\xmem_data[10][5] ), .B1(n31360), .B2(
        \xmem_data[11][5] ), .ZN(n13836) );
  AOI22_X1 U18019 ( .A1(n25632), .A2(\xmem_data[12][5] ), .B1(n25581), .B2(
        \xmem_data[13][5] ), .ZN(n13835) );
  AOI22_X1 U18020 ( .A1(n25636), .A2(\xmem_data[14][5] ), .B1(n20949), .B2(
        \xmem_data[15][5] ), .ZN(n13834) );
  NAND4_X1 U18021 ( .A1(n13837), .A2(n13836), .A3(n13835), .A4(n13834), .ZN(
        n13840) );
  AOI22_X1 U18022 ( .A1(n25612), .A2(\xmem_data[26][5] ), .B1(n25562), .B2(
        \xmem_data[27][5] ), .ZN(n13838) );
  OR2_X1 U18023 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  AOI21_X1 U18024 ( .B1(n28045), .B2(\xmem_data[31][5] ), .A(n13845), .ZN(
        n13911) );
  AOI22_X1 U18025 ( .A1(n25707), .A2(\xmem_data[32][5] ), .B1(n3358), .B2(
        \xmem_data[33][5] ), .ZN(n13849) );
  AOI22_X1 U18026 ( .A1(n25708), .A2(\xmem_data[34][5] ), .B1(n13168), .B2(
        \xmem_data[35][5] ), .ZN(n13848) );
  AOI22_X1 U18027 ( .A1(n29023), .A2(\xmem_data[36][5] ), .B1(n25709), .B2(
        \xmem_data[37][5] ), .ZN(n13847) );
  AOI22_X1 U18028 ( .A1(n21048), .A2(\xmem_data[38][5] ), .B1(n20938), .B2(
        \xmem_data[39][5] ), .ZN(n13846) );
  NAND4_X1 U18029 ( .A1(n13849), .A2(n13848), .A3(n13847), .A4(n13846), .ZN(
        n13865) );
  AOI22_X1 U18030 ( .A1(n22676), .A2(\xmem_data[40][5] ), .B1(n25715), .B2(
        \xmem_data[41][5] ), .ZN(n13853) );
  AOI22_X1 U18031 ( .A1(n23777), .A2(\xmem_data[42][5] ), .B1(n24460), .B2(
        \xmem_data[43][5] ), .ZN(n13852) );
  AOI22_X1 U18032 ( .A1(n24190), .A2(\xmem_data[44][5] ), .B1(n28429), .B2(
        \xmem_data[45][5] ), .ZN(n13851) );
  AOI22_X1 U18033 ( .A1(n25718), .A2(\xmem_data[46][5] ), .B1(n24521), .B2(
        \xmem_data[47][5] ), .ZN(n13850) );
  NAND4_X1 U18034 ( .A1(n13853), .A2(n13852), .A3(n13851), .A4(n13850), .ZN(
        n13864) );
  AOI22_X1 U18035 ( .A1(n25582), .A2(\xmem_data[48][5] ), .B1(n25723), .B2(
        \xmem_data[49][5] ), .ZN(n13857) );
  AOI22_X1 U18036 ( .A1(n20952), .A2(\xmem_data[50][5] ), .B1(n25528), .B2(
        \xmem_data[51][5] ), .ZN(n13856) );
  AOI22_X1 U18037 ( .A1(n25724), .A2(\xmem_data[52][5] ), .B1(n28317), .B2(
        \xmem_data[53][5] ), .ZN(n13855) );
  AOI22_X1 U18038 ( .A1(n25725), .A2(\xmem_data[54][5] ), .B1(n30863), .B2(
        \xmem_data[55][5] ), .ZN(n13854) );
  NAND4_X1 U18039 ( .A1(n13857), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        n13863) );
  AOI22_X1 U18040 ( .A1(n25730), .A2(\xmem_data[56][5] ), .B1(n3220), .B2(
        \xmem_data[57][5] ), .ZN(n13861) );
  AOI22_X1 U18041 ( .A1(n25731), .A2(\xmem_data[58][5] ), .B1(n31367), .B2(
        \xmem_data[59][5] ), .ZN(n13860) );
  AOI22_X1 U18042 ( .A1(n20725), .A2(\xmem_data[60][5] ), .B1(n27550), .B2(
        \xmem_data[61][5] ), .ZN(n13859) );
  AOI22_X1 U18043 ( .A1(n25732), .A2(\xmem_data[62][5] ), .B1(n23771), .B2(
        \xmem_data[63][5] ), .ZN(n13858) );
  NAND4_X1 U18044 ( .A1(n13861), .A2(n13860), .A3(n13859), .A4(n13858), .ZN(
        n13862) );
  OR4_X1 U18045 ( .A1(n13865), .A2(n13864), .A3(n13863), .A4(n13862), .ZN(
        n13866) );
  NAND2_X1 U18046 ( .A1(n13866), .A2(n25741), .ZN(n13910) );
  AOI22_X1 U18047 ( .A1(n25670), .A2(\xmem_data[96][5] ), .B1(n25456), .B2(
        \xmem_data[97][5] ), .ZN(n13870) );
  AOI22_X1 U18048 ( .A1(n25708), .A2(\xmem_data[98][5] ), .B1(n24639), .B2(
        \xmem_data[99][5] ), .ZN(n13869) );
  AOI22_X1 U18049 ( .A1(n17041), .A2(\xmem_data[100][5] ), .B1(n25671), .B2(
        \xmem_data[101][5] ), .ZN(n13868) );
  AOI22_X1 U18050 ( .A1(n25672), .A2(\xmem_data[102][5] ), .B1(n22742), .B2(
        \xmem_data[103][5] ), .ZN(n13867) );
  NAND4_X1 U18051 ( .A1(n13870), .A2(n13869), .A3(n13868), .A4(n13867), .ZN(
        n13886) );
  AOI22_X1 U18052 ( .A1(n13149), .A2(\xmem_data[104][5] ), .B1(n25677), .B2(
        \xmem_data[105][5] ), .ZN(n13874) );
  AOI22_X1 U18053 ( .A1(n25678), .A2(\xmem_data[106][5] ), .B1(n24510), .B2(
        \xmem_data[107][5] ), .ZN(n13873) );
  AOI22_X1 U18054 ( .A1(n27524), .A2(\xmem_data[108][5] ), .B1(n30598), .B2(
        \xmem_data[109][5] ), .ZN(n13872) );
  AOI22_X1 U18055 ( .A1(n3151), .A2(\xmem_data[110][5] ), .B1(n24223), .B2(
        \xmem_data[111][5] ), .ZN(n13871) );
  NAND4_X1 U18056 ( .A1(n13874), .A2(n13873), .A3(n13872), .A4(n13871), .ZN(
        n13885) );
  AOI22_X1 U18057 ( .A1(n24166), .A2(\xmem_data[112][5] ), .B1(n22751), .B2(
        \xmem_data[113][5] ), .ZN(n13878) );
  AOI22_X1 U18058 ( .A1(n25684), .A2(\xmem_data[114][5] ), .B1(n27567), .B2(
        \xmem_data[115][5] ), .ZN(n13877) );
  AOI22_X1 U18059 ( .A1(n25686), .A2(\xmem_data[116][5] ), .B1(n25685), .B2(
        \xmem_data[117][5] ), .ZN(n13876) );
  AOI22_X1 U18060 ( .A1(n28973), .A2(\xmem_data[118][5] ), .B1(n25687), .B2(
        \xmem_data[119][5] ), .ZN(n13875) );
  NAND4_X1 U18061 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13875), .ZN(
        n13884) );
  AOI22_X1 U18062 ( .A1(n25692), .A2(\xmem_data[120][5] ), .B1(n3222), .B2(
        \xmem_data[121][5] ), .ZN(n13882) );
  AOI22_X1 U18063 ( .A1(n25693), .A2(\xmem_data[122][5] ), .B1(n25562), .B2(
        \xmem_data[123][5] ), .ZN(n13881) );
  AOI22_X1 U18064 ( .A1(n25694), .A2(\xmem_data[124][5] ), .B1(n31275), .B2(
        \xmem_data[125][5] ), .ZN(n13880) );
  AOI22_X1 U18065 ( .A1(n29350), .A2(\xmem_data[126][5] ), .B1(n3231), .B2(
        \xmem_data[127][5] ), .ZN(n13879) );
  NAND4_X1 U18066 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13883) );
  OR4_X1 U18067 ( .A1(n13886), .A2(n13885), .A3(n13884), .A4(n13883), .ZN(
        n13908) );
  AOI22_X1 U18068 ( .A1(n25707), .A2(\xmem_data[64][5] ), .B1(n20546), .B2(
        \xmem_data[65][5] ), .ZN(n13890) );
  AOI22_X1 U18069 ( .A1(n25708), .A2(\xmem_data[66][5] ), .B1(n24159), .B2(
        \xmem_data[67][5] ), .ZN(n13889) );
  AOI22_X1 U18070 ( .A1(n28980), .A2(\xmem_data[68][5] ), .B1(n25709), .B2(
        \xmem_data[69][5] ), .ZN(n13888) );
  AOI22_X1 U18071 ( .A1(n25672), .A2(\xmem_data[70][5] ), .B1(n27454), .B2(
        \xmem_data[71][5] ), .ZN(n13887) );
  NAND4_X1 U18072 ( .A1(n13890), .A2(n13889), .A3(n13888), .A4(n13887), .ZN(
        n13906) );
  AOI22_X1 U18073 ( .A1(n20585), .A2(\xmem_data[72][5] ), .B1(n25715), .B2(
        \xmem_data[73][5] ), .ZN(n13894) );
  AOI22_X1 U18074 ( .A1(n17044), .A2(\xmem_data[74][5] ), .B1(n29280), .B2(
        \xmem_data[75][5] ), .ZN(n13893) );
  AOI22_X1 U18075 ( .A1(n28460), .A2(\xmem_data[76][5] ), .B1(n20816), .B2(
        \xmem_data[77][5] ), .ZN(n13892) );
  AOI22_X1 U18076 ( .A1(n25718), .A2(\xmem_data[78][5] ), .B1(n23723), .B2(
        \xmem_data[79][5] ), .ZN(n13891) );
  NAND4_X1 U18077 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n13905) );
  AOI22_X1 U18078 ( .A1(n27542), .A2(\xmem_data[80][5] ), .B1(n25723), .B2(
        \xmem_data[81][5] ), .ZN(n13898) );
  AOI22_X1 U18079 ( .A1(n20770), .A2(\xmem_data[82][5] ), .B1(n24524), .B2(
        \xmem_data[83][5] ), .ZN(n13897) );
  AOI22_X1 U18080 ( .A1(n25724), .A2(\xmem_data[84][5] ), .B1(n24573), .B2(
        \xmem_data[85][5] ), .ZN(n13896) );
  AOI22_X1 U18081 ( .A1(n25725), .A2(\xmem_data[86][5] ), .B1(n25485), .B2(
        \xmem_data[87][5] ), .ZN(n13895) );
  NAND4_X1 U18082 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        n13904) );
  AOI22_X1 U18083 ( .A1(n25730), .A2(\xmem_data[88][5] ), .B1(n3220), .B2(
        \xmem_data[89][5] ), .ZN(n13902) );
  AOI22_X1 U18084 ( .A1(n25731), .A2(\xmem_data[90][5] ), .B1(n28319), .B2(
        \xmem_data[91][5] ), .ZN(n13901) );
  AOI22_X1 U18085 ( .A1(n27938), .A2(\xmem_data[92][5] ), .B1(n31275), .B2(
        \xmem_data[93][5] ), .ZN(n13900) );
  AOI22_X1 U18086 ( .A1(n25732), .A2(\xmem_data[94][5] ), .B1(n25514), .B2(
        \xmem_data[95][5] ), .ZN(n13899) );
  NAND4_X1 U18087 ( .A1(n13902), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13903) );
  OR4_X1 U18088 ( .A1(n13906), .A2(n13905), .A3(n13904), .A4(n13903), .ZN(
        n13907) );
  AOI22_X1 U18089 ( .A1(n25706), .A2(n13908), .B1(n25704), .B2(n13907), .ZN(
        n13909) );
  XNOR2_X1 U18090 ( .A(n30451), .B(\fmem_data[6][7] ), .ZN(n34930) );
  AOI22_X1 U18091 ( .A1(n29849), .A2(\xmem_data[32][7] ), .B1(n29848), .B2(
        \xmem_data[33][7] ), .ZN(n13916) );
  AOI22_X1 U18092 ( .A1(n29851), .A2(\xmem_data[34][7] ), .B1(n29850), .B2(
        \xmem_data[35][7] ), .ZN(n13915) );
  AOI22_X1 U18093 ( .A1(n29853), .A2(\xmem_data[36][7] ), .B1(n29852), .B2(
        \xmem_data[37][7] ), .ZN(n13914) );
  AOI22_X1 U18094 ( .A1(n29855), .A2(\xmem_data[38][7] ), .B1(n29854), .B2(
        \xmem_data[39][7] ), .ZN(n13913) );
  NAND4_X1 U18095 ( .A1(n13916), .A2(n13915), .A3(n13914), .A4(n13913), .ZN(
        n13932) );
  AOI22_X1 U18096 ( .A1(n29860), .A2(\xmem_data[40][7] ), .B1(n29976), .B2(
        \xmem_data[41][7] ), .ZN(n13920) );
  AOI22_X1 U18097 ( .A1(n29978), .A2(\xmem_data[42][7] ), .B1(n3195), .B2(
        \xmem_data[43][7] ), .ZN(n13919) );
  AOI22_X1 U18098 ( .A1(n29980), .A2(\xmem_data[44][7] ), .B1(n29979), .B2(
        \xmem_data[45][7] ), .ZN(n13918) );
  AOI22_X1 U18099 ( .A1(n29982), .A2(\xmem_data[46][7] ), .B1(n29981), .B2(
        \xmem_data[47][7] ), .ZN(n13917) );
  NAND4_X1 U18100 ( .A1(n13920), .A2(n13919), .A3(n13918), .A4(n13917), .ZN(
        n13931) );
  AOI22_X1 U18101 ( .A1(n29866), .A2(\xmem_data[48][7] ), .B1(n29865), .B2(
        \xmem_data[49][7] ), .ZN(n13924) );
  AOI22_X1 U18102 ( .A1(n29868), .A2(\xmem_data[50][7] ), .B1(n29867), .B2(
        \xmem_data[51][7] ), .ZN(n13923) );
  AOI22_X1 U18103 ( .A1(n29870), .A2(\xmem_data[52][7] ), .B1(n29869), .B2(
        \xmem_data[53][7] ), .ZN(n13922) );
  AOI22_X1 U18104 ( .A1(n29871), .A2(\xmem_data[54][7] ), .B1(n29993), .B2(
        \xmem_data[55][7] ), .ZN(n13921) );
  NAND4_X1 U18105 ( .A1(n13924), .A2(n13923), .A3(n13922), .A4(n13921), .ZN(
        n13930) );
  AOI22_X1 U18106 ( .A1(n29877), .A2(\xmem_data[56][7] ), .B1(n29876), .B2(
        \xmem_data[57][7] ), .ZN(n13928) );
  AOI22_X1 U18107 ( .A1(n29879), .A2(\xmem_data[58][7] ), .B1(n29878), .B2(
        \xmem_data[59][7] ), .ZN(n13927) );
  AOI22_X1 U18108 ( .A1(n29881), .A2(\xmem_data[60][7] ), .B1(n29880), .B2(
        \xmem_data[61][7] ), .ZN(n13926) );
  AOI22_X1 U18109 ( .A1(n29883), .A2(\xmem_data[62][7] ), .B1(n29882), .B2(
        \xmem_data[63][7] ), .ZN(n13925) );
  NAND4_X1 U18110 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n13929) );
  OR4_X1 U18111 ( .A1(n13932), .A2(n13931), .A3(n13930), .A4(n13929), .ZN(
        n13954) );
  AOI22_X1 U18112 ( .A1(n29893), .A2(\xmem_data[0][7] ), .B1(n29892), .B2(
        \xmem_data[1][7] ), .ZN(n13936) );
  AOI22_X1 U18113 ( .A1(n29895), .A2(\xmem_data[2][7] ), .B1(n29894), .B2(
        \xmem_data[3][7] ), .ZN(n13935) );
  AOI22_X1 U18114 ( .A1(n29897), .A2(\xmem_data[4][7] ), .B1(n29896), .B2(
        \xmem_data[5][7] ), .ZN(n13934) );
  AOI22_X1 U18115 ( .A1(n29899), .A2(\xmem_data[6][7] ), .B1(n29898), .B2(
        \xmem_data[7][7] ), .ZN(n13933) );
  NAND4_X1 U18116 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n13933), .ZN(
        n13952) );
  AOI22_X1 U18117 ( .A1(n29904), .A2(\xmem_data[8][7] ), .B1(n29942), .B2(
        \xmem_data[9][7] ), .ZN(n13940) );
  AOI22_X1 U18118 ( .A1(n29943), .A2(\xmem_data[10][7] ), .B1(n3196), .B2(
        \xmem_data[11][7] ), .ZN(n13939) );
  AOI22_X1 U18119 ( .A1(n29945), .A2(\xmem_data[12][7] ), .B1(n29906), .B2(
        \xmem_data[13][7] ), .ZN(n13938) );
  AOI22_X1 U18120 ( .A1(n29947), .A2(\xmem_data[14][7] ), .B1(n29908), .B2(
        \xmem_data[15][7] ), .ZN(n13937) );
  NAND4_X1 U18121 ( .A1(n13940), .A2(n13939), .A3(n13938), .A4(n13937), .ZN(
        n13951) );
  AOI22_X1 U18122 ( .A1(n29917), .A2(\xmem_data[18][7] ), .B1(n29916), .B2(
        \xmem_data[19][7] ), .ZN(n13944) );
  AOI22_X1 U18123 ( .A1(n29915), .A2(\xmem_data[16][7] ), .B1(n29914), .B2(
        \xmem_data[17][7] ), .ZN(n13943) );
  AOI22_X1 U18124 ( .A1(n29921), .A2(\xmem_data[22][7] ), .B1(n29920), .B2(
        \xmem_data[23][7] ), .ZN(n13942) );
  AOI22_X1 U18125 ( .A1(n29918), .A2(\xmem_data[21][7] ), .B1(n29919), .B2(
        \xmem_data[20][7] ), .ZN(n13941) );
  NAND4_X1 U18126 ( .A1(n13944), .A2(n13943), .A3(n13942), .A4(n13941), .ZN(
        n13950) );
  AOI22_X1 U18127 ( .A1(n3243), .A2(\xmem_data[24][7] ), .B1(n3242), .B2(
        \xmem_data[25][7] ), .ZN(n13948) );
  AOI22_X1 U18128 ( .A1(n3235), .A2(\xmem_data[26][7] ), .B1(n3238), .B2(
        \xmem_data[27][7] ), .ZN(n13947) );
  AOI22_X1 U18129 ( .A1(n3236), .A2(\xmem_data[28][7] ), .B1(n3225), .B2(
        \xmem_data[29][7] ), .ZN(n13946) );
  AOI22_X1 U18130 ( .A1(n3237), .A2(\xmem_data[30][7] ), .B1(n3234), .B2(
        \xmem_data[31][7] ), .ZN(n13945) );
  NAND4_X1 U18131 ( .A1(n13948), .A2(n13947), .A3(n13946), .A4(n13945), .ZN(
        n13949) );
  AOI22_X1 U18132 ( .A1(n29937), .A2(n13954), .B1(n29935), .B2(n13953), .ZN(
        n14001) );
  AOI22_X1 U18133 ( .A1(n29966), .A2(\xmem_data[96][7] ), .B1(n29965), .B2(
        \xmem_data[97][7] ), .ZN(n13958) );
  AOI22_X1 U18134 ( .A1(n29968), .A2(\xmem_data[98][7] ), .B1(n29967), .B2(
        \xmem_data[99][7] ), .ZN(n13957) );
  AOI22_X1 U18135 ( .A1(n29969), .A2(\xmem_data[100][7] ), .B1(n29896), .B2(
        \xmem_data[101][7] ), .ZN(n13956) );
  AOI22_X1 U18136 ( .A1(n29971), .A2(\xmem_data[102][7] ), .B1(n29970), .B2(
        \xmem_data[103][7] ), .ZN(n13955) );
  NAND4_X1 U18137 ( .A1(n13958), .A2(n13957), .A3(n13956), .A4(n13955), .ZN(
        n13974) );
  AOI22_X1 U18138 ( .A1(n29977), .A2(\xmem_data[104][7] ), .B1(n29976), .B2(
        \xmem_data[105][7] ), .ZN(n13962) );
  AOI22_X1 U18139 ( .A1(n29905), .A2(\xmem_data[106][7] ), .B1(n3195), .B2(
        \xmem_data[107][7] ), .ZN(n13961) );
  AOI22_X1 U18140 ( .A1(n29907), .A2(\xmem_data[108][7] ), .B1(n29906), .B2(
        \xmem_data[109][7] ), .ZN(n13960) );
  AOI22_X1 U18141 ( .A1(n29909), .A2(\xmem_data[110][7] ), .B1(n29908), .B2(
        \xmem_data[111][7] ), .ZN(n13959) );
  NAND4_X1 U18142 ( .A1(n13962), .A2(n13961), .A3(n13960), .A4(n13959), .ZN(
        n13973) );
  AOI22_X1 U18143 ( .A1(n29988), .A2(\xmem_data[112][7] ), .B1(n29987), .B2(
        \xmem_data[113][7] ), .ZN(n13966) );
  AOI22_X1 U18144 ( .A1(n29990), .A2(\xmem_data[114][7] ), .B1(n29989), .B2(
        \xmem_data[115][7] ), .ZN(n13965) );
  AOI22_X1 U18145 ( .A1(n29992), .A2(\xmem_data[116][7] ), .B1(n29991), .B2(
        \xmem_data[117][7] ), .ZN(n13964) );
  AOI22_X1 U18146 ( .A1(n29994), .A2(\xmem_data[118][7] ), .B1(n29952), .B2(
        \xmem_data[119][7] ), .ZN(n13963) );
  NAND4_X1 U18147 ( .A1(n13966), .A2(n13965), .A3(n13964), .A4(n13963), .ZN(
        n13972) );
  AOI22_X1 U18148 ( .A1(n3243), .A2(\xmem_data[120][7] ), .B1(n3242), .B2(
        \xmem_data[121][7] ), .ZN(n13970) );
  AOI22_X1 U18149 ( .A1(n3235), .A2(\xmem_data[122][7] ), .B1(n3238), .B2(
        \xmem_data[123][7] ), .ZN(n13969) );
  AOI22_X1 U18150 ( .A1(n3236), .A2(\xmem_data[124][7] ), .B1(n3225), .B2(
        \xmem_data[125][7] ), .ZN(n13968) );
  AOI22_X1 U18151 ( .A1(n3237), .A2(\xmem_data[126][7] ), .B1(n3234), .B2(
        \xmem_data[127][7] ), .ZN(n13967) );
  NAND4_X1 U18152 ( .A1(n13970), .A2(n13969), .A3(n13968), .A4(n13967), .ZN(
        n13971) );
  OR4_X1 U18153 ( .A1(n13974), .A2(n13973), .A3(n13972), .A4(n13971), .ZN(
        n13999) );
  AOI22_X1 U18154 ( .A1(n29860), .A2(\xmem_data[72][7] ), .B1(n29942), .B2(
        \xmem_data[73][7] ), .ZN(n13978) );
  AOI22_X1 U18155 ( .A1(n29943), .A2(\xmem_data[74][7] ), .B1(n3195), .B2(
        \xmem_data[75][7] ), .ZN(n13977) );
  AOI22_X1 U18156 ( .A1(n29945), .A2(\xmem_data[76][7] ), .B1(n29944), .B2(
        \xmem_data[77][7] ), .ZN(n13976) );
  AOI22_X1 U18157 ( .A1(n29947), .A2(\xmem_data[78][7] ), .B1(n29946), .B2(
        \xmem_data[79][7] ), .ZN(n13975) );
  NAND4_X1 U18158 ( .A1(n13978), .A2(n13977), .A3(n13976), .A4(n13975), .ZN(
        n13984) );
  AOI22_X1 U18159 ( .A1(n29866), .A2(\xmem_data[80][7] ), .B1(n29865), .B2(
        \xmem_data[81][7] ), .ZN(n13982) );
  AOI22_X1 U18160 ( .A1(n29868), .A2(\xmem_data[82][7] ), .B1(n29867), .B2(
        \xmem_data[83][7] ), .ZN(n13981) );
  AOI22_X1 U18161 ( .A1(n29870), .A2(\xmem_data[84][7] ), .B1(n29869), .B2(
        \xmem_data[85][7] ), .ZN(n13980) );
  AOI22_X1 U18162 ( .A1(n29871), .A2(\xmem_data[86][7] ), .B1(n29952), .B2(
        \xmem_data[87][7] ), .ZN(n13979) );
  NAND4_X1 U18163 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13983) );
  AOI22_X1 U18164 ( .A1(n29877), .A2(\xmem_data[88][7] ), .B1(n29876), .B2(
        \xmem_data[89][7] ), .ZN(n13988) );
  AOI22_X1 U18165 ( .A1(n29879), .A2(\xmem_data[90][7] ), .B1(n29878), .B2(
        \xmem_data[91][7] ), .ZN(n13987) );
  AOI22_X1 U18166 ( .A1(n29881), .A2(\xmem_data[92][7] ), .B1(n29880), .B2(
        \xmem_data[93][7] ), .ZN(n13986) );
  AOI22_X1 U18167 ( .A1(n29883), .A2(\xmem_data[94][7] ), .B1(n29882), .B2(
        \xmem_data[95][7] ), .ZN(n13985) );
  NAND4_X1 U18168 ( .A1(n13988), .A2(n13987), .A3(n13986), .A4(n13985), .ZN(
        n13994) );
  AOI22_X1 U18169 ( .A1(n29849), .A2(\xmem_data[64][7] ), .B1(n29848), .B2(
        \xmem_data[65][7] ), .ZN(n13992) );
  AOI22_X1 U18170 ( .A1(n29851), .A2(\xmem_data[66][7] ), .B1(n29850), .B2(
        \xmem_data[67][7] ), .ZN(n13991) );
  AOI22_X1 U18171 ( .A1(n29853), .A2(\xmem_data[68][7] ), .B1(n29852), .B2(
        \xmem_data[69][7] ), .ZN(n13990) );
  AOI22_X1 U18172 ( .A1(n29855), .A2(\xmem_data[70][7] ), .B1(n29854), .B2(
        \xmem_data[71][7] ), .ZN(n13989) );
  NAND4_X1 U18173 ( .A1(n13992), .A2(n13991), .A3(n13990), .A4(n13989), .ZN(
        n13993) );
  XNOR2_X1 U18174 ( .A(n35280), .B(\fmem_data[1][5] ), .ZN(n34940) );
  AOI22_X1 U18175 ( .A1(n29849), .A2(\xmem_data[32][6] ), .B1(n29848), .B2(
        \xmem_data[33][6] ), .ZN(n14005) );
  AOI22_X1 U18176 ( .A1(n29851), .A2(\xmem_data[34][6] ), .B1(n29850), .B2(
        \xmem_data[35][6] ), .ZN(n14004) );
  AOI22_X1 U18177 ( .A1(n29853), .A2(\xmem_data[36][6] ), .B1(n29852), .B2(
        \xmem_data[37][6] ), .ZN(n14003) );
  AOI22_X1 U18178 ( .A1(n29855), .A2(\xmem_data[38][6] ), .B1(n29854), .B2(
        \xmem_data[39][6] ), .ZN(n14002) );
  NAND4_X1 U18179 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14021) );
  AOI22_X1 U18180 ( .A1(n29860), .A2(\xmem_data[40][6] ), .B1(n29976), .B2(
        \xmem_data[41][6] ), .ZN(n14009) );
  AOI22_X1 U18181 ( .A1(n29978), .A2(\xmem_data[42][6] ), .B1(n3195), .B2(
        \xmem_data[43][6] ), .ZN(n14008) );
  AOI22_X1 U18182 ( .A1(n29980), .A2(\xmem_data[44][6] ), .B1(n29944), .B2(
        \xmem_data[45][6] ), .ZN(n14007) );
  AOI22_X1 U18183 ( .A1(n29982), .A2(\xmem_data[46][6] ), .B1(n29946), .B2(
        \xmem_data[47][6] ), .ZN(n14006) );
  NAND4_X1 U18184 ( .A1(n14009), .A2(n14008), .A3(n14007), .A4(n14006), .ZN(
        n14020) );
  AOI22_X1 U18185 ( .A1(n29866), .A2(\xmem_data[48][6] ), .B1(n29865), .B2(
        \xmem_data[49][6] ), .ZN(n14013) );
  AOI22_X1 U18186 ( .A1(n29868), .A2(\xmem_data[50][6] ), .B1(n29867), .B2(
        \xmem_data[51][6] ), .ZN(n14012) );
  AOI22_X1 U18187 ( .A1(n29870), .A2(\xmem_data[52][6] ), .B1(n29869), .B2(
        \xmem_data[53][6] ), .ZN(n14011) );
  AOI22_X1 U18188 ( .A1(n29871), .A2(\xmem_data[54][6] ), .B1(n29920), .B2(
        \xmem_data[55][6] ), .ZN(n14010) );
  NAND4_X1 U18189 ( .A1(n14013), .A2(n14012), .A3(n14011), .A4(n14010), .ZN(
        n14019) );
  AOI22_X1 U18190 ( .A1(n29877), .A2(\xmem_data[56][6] ), .B1(n29876), .B2(
        \xmem_data[57][6] ), .ZN(n14017) );
  AOI22_X1 U18191 ( .A1(n29879), .A2(\xmem_data[58][6] ), .B1(n29878), .B2(
        \xmem_data[59][6] ), .ZN(n14016) );
  AOI22_X1 U18192 ( .A1(n29881), .A2(\xmem_data[60][6] ), .B1(n29880), .B2(
        \xmem_data[61][6] ), .ZN(n14015) );
  AOI22_X1 U18193 ( .A1(n29883), .A2(\xmem_data[62][6] ), .B1(n29882), .B2(
        \xmem_data[63][6] ), .ZN(n14014) );
  NAND4_X1 U18194 ( .A1(n14017), .A2(n14016), .A3(n14015), .A4(n14014), .ZN(
        n14018) );
  OR4_X1 U18195 ( .A1(n14021), .A2(n14020), .A3(n14019), .A4(n14018), .ZN(
        n14043) );
  AOI22_X1 U18196 ( .A1(n29893), .A2(\xmem_data[0][6] ), .B1(n29892), .B2(
        \xmem_data[1][6] ), .ZN(n14025) );
  AOI22_X1 U18197 ( .A1(n29895), .A2(\xmem_data[2][6] ), .B1(n29894), .B2(
        \xmem_data[3][6] ), .ZN(n14024) );
  AOI22_X1 U18198 ( .A1(n29897), .A2(\xmem_data[4][6] ), .B1(n29896), .B2(
        \xmem_data[5][6] ), .ZN(n14023) );
  AOI22_X1 U18199 ( .A1(n29899), .A2(\xmem_data[6][6] ), .B1(n29898), .B2(
        \xmem_data[7][6] ), .ZN(n14022) );
  NAND4_X1 U18200 ( .A1(n14025), .A2(n14024), .A3(n14023), .A4(n14022), .ZN(
        n14041) );
  AOI22_X1 U18201 ( .A1(n29904), .A2(\xmem_data[8][6] ), .B1(n29976), .B2(
        \xmem_data[9][6] ), .ZN(n14029) );
  AOI22_X1 U18202 ( .A1(n29978), .A2(\xmem_data[10][6] ), .B1(n3196), .B2(
        \xmem_data[11][6] ), .ZN(n14028) );
  AOI22_X1 U18203 ( .A1(n29980), .A2(\xmem_data[12][6] ), .B1(n29979), .B2(
        \xmem_data[13][6] ), .ZN(n14027) );
  AOI22_X1 U18204 ( .A1(n29982), .A2(\xmem_data[14][6] ), .B1(n29981), .B2(
        \xmem_data[15][6] ), .ZN(n14026) );
  NAND4_X1 U18205 ( .A1(n14029), .A2(n14028), .A3(n14027), .A4(n14026), .ZN(
        n14040) );
  AOI22_X1 U18206 ( .A1(n29915), .A2(\xmem_data[16][6] ), .B1(n29914), .B2(
        \xmem_data[17][6] ), .ZN(n14033) );
  AOI22_X1 U18207 ( .A1(n29917), .A2(\xmem_data[18][6] ), .B1(n29916), .B2(
        \xmem_data[19][6] ), .ZN(n14032) );
  AOI22_X1 U18208 ( .A1(n29919), .A2(\xmem_data[20][6] ), .B1(n29918), .B2(
        \xmem_data[21][6] ), .ZN(n14031) );
  AOI22_X1 U18209 ( .A1(n29921), .A2(\xmem_data[22][6] ), .B1(n29952), .B2(
        \xmem_data[23][6] ), .ZN(n14030) );
  NAND4_X1 U18210 ( .A1(n14033), .A2(n14032), .A3(n14031), .A4(n14030), .ZN(
        n14039) );
  AOI22_X1 U18211 ( .A1(n3243), .A2(\xmem_data[24][6] ), .B1(n3242), .B2(
        \xmem_data[25][6] ), .ZN(n14037) );
  AOI22_X1 U18212 ( .A1(n3235), .A2(\xmem_data[26][6] ), .B1(n3238), .B2(
        \xmem_data[27][6] ), .ZN(n14036) );
  AOI22_X1 U18213 ( .A1(n3236), .A2(\xmem_data[28][6] ), .B1(n3225), .B2(
        \xmem_data[29][6] ), .ZN(n14035) );
  AOI22_X1 U18214 ( .A1(n3237), .A2(\xmem_data[30][6] ), .B1(n3234), .B2(
        \xmem_data[31][6] ), .ZN(n14034) );
  NAND4_X1 U18215 ( .A1(n14037), .A2(n14036), .A3(n14035), .A4(n14034), .ZN(
        n14038) );
  OR4_X1 U18216 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14042) );
  AOI22_X1 U18217 ( .A1(n29937), .A2(n14043), .B1(n29935), .B2(n14042), .ZN(
        n14087) );
  AOI22_X1 U18218 ( .A1(n29966), .A2(\xmem_data[96][6] ), .B1(n29965), .B2(
        \xmem_data[97][6] ), .ZN(n14047) );
  AOI22_X1 U18219 ( .A1(n29968), .A2(\xmem_data[98][6] ), .B1(n29967), .B2(
        \xmem_data[99][6] ), .ZN(n14046) );
  AOI22_X1 U18220 ( .A1(n29969), .A2(\xmem_data[100][6] ), .B1(n29896), .B2(
        \xmem_data[101][6] ), .ZN(n14045) );
  AOI22_X1 U18221 ( .A1(n29971), .A2(\xmem_data[102][6] ), .B1(n29970), .B2(
        \xmem_data[103][6] ), .ZN(n14044) );
  NAND4_X1 U18222 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        n14063) );
  AOI22_X1 U18223 ( .A1(n29977), .A2(\xmem_data[104][6] ), .B1(n29976), .B2(
        \xmem_data[105][6] ), .ZN(n14051) );
  AOI22_X1 U18224 ( .A1(n29905), .A2(\xmem_data[106][6] ), .B1(n3196), .B2(
        \xmem_data[107][6] ), .ZN(n14050) );
  AOI22_X1 U18225 ( .A1(n29907), .A2(\xmem_data[108][6] ), .B1(n29979), .B2(
        \xmem_data[109][6] ), .ZN(n14049) );
  AOI22_X1 U18226 ( .A1(n29909), .A2(\xmem_data[110][6] ), .B1(n29981), .B2(
        \xmem_data[111][6] ), .ZN(n14048) );
  NAND4_X1 U18227 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14062) );
  AOI22_X1 U18228 ( .A1(n29988), .A2(\xmem_data[112][6] ), .B1(n29987), .B2(
        \xmem_data[113][6] ), .ZN(n14055) );
  AOI22_X1 U18229 ( .A1(n29990), .A2(\xmem_data[114][6] ), .B1(n29989), .B2(
        \xmem_data[115][6] ), .ZN(n14054) );
  AOI22_X1 U18230 ( .A1(n29992), .A2(\xmem_data[116][6] ), .B1(n29991), .B2(
        \xmem_data[117][6] ), .ZN(n14053) );
  AOI22_X1 U18231 ( .A1(n29994), .A2(\xmem_data[118][6] ), .B1(n29993), .B2(
        \xmem_data[119][6] ), .ZN(n14052) );
  NAND4_X1 U18232 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14061) );
  AOI22_X1 U18233 ( .A1(n3243), .A2(\xmem_data[120][6] ), .B1(n3242), .B2(
        \xmem_data[121][6] ), .ZN(n14059) );
  AOI22_X1 U18234 ( .A1(n3235), .A2(\xmem_data[122][6] ), .B1(n3238), .B2(
        \xmem_data[123][6] ), .ZN(n14058) );
  AOI22_X1 U18235 ( .A1(n3236), .A2(\xmem_data[124][6] ), .B1(n3225), .B2(
        \xmem_data[125][6] ), .ZN(n14057) );
  AOI22_X1 U18236 ( .A1(n3237), .A2(\xmem_data[126][6] ), .B1(n3234), .B2(
        \xmem_data[127][6] ), .ZN(n14056) );
  NAND4_X1 U18237 ( .A1(n14059), .A2(n14058), .A3(n14057), .A4(n14056), .ZN(
        n14060) );
  OR4_X1 U18238 ( .A1(n14063), .A2(n14062), .A3(n14061), .A4(n14060), .ZN(
        n14085) );
  AOI22_X1 U18239 ( .A1(n29849), .A2(\xmem_data[64][6] ), .B1(n29848), .B2(
        \xmem_data[65][6] ), .ZN(n14067) );
  AOI22_X1 U18240 ( .A1(n29851), .A2(n20682), .B1(n29850), .B2(
        \xmem_data[67][6] ), .ZN(n14066) );
  AOI22_X1 U18241 ( .A1(n29853), .A2(\xmem_data[68][6] ), .B1(n29852), .B2(
        \xmem_data[69][6] ), .ZN(n14065) );
  AOI22_X1 U18242 ( .A1(n29855), .A2(\xmem_data[70][6] ), .B1(n29854), .B2(
        \xmem_data[71][6] ), .ZN(n14064) );
  NAND4_X1 U18243 ( .A1(n14067), .A2(n14066), .A3(n14065), .A4(n14064), .ZN(
        n14083) );
  AOI22_X1 U18244 ( .A1(n29860), .A2(\xmem_data[72][6] ), .B1(n29976), .B2(
        \xmem_data[73][6] ), .ZN(n14071) );
  AOI22_X1 U18245 ( .A1(n29905), .A2(\xmem_data[74][6] ), .B1(n3195), .B2(
        \xmem_data[75][6] ), .ZN(n14070) );
  AOI22_X1 U18246 ( .A1(n29907), .A2(\xmem_data[76][6] ), .B1(n29906), .B2(
        \xmem_data[77][6] ), .ZN(n14069) );
  AOI22_X1 U18247 ( .A1(n29909), .A2(\xmem_data[78][6] ), .B1(n29908), .B2(
        \xmem_data[79][6] ), .ZN(n14068) );
  NAND4_X1 U18248 ( .A1(n14071), .A2(n14070), .A3(n14069), .A4(n14068), .ZN(
        n14082) );
  AOI22_X1 U18249 ( .A1(n29866), .A2(\xmem_data[80][6] ), .B1(n29865), .B2(
        \xmem_data[81][6] ), .ZN(n14075) );
  AOI22_X1 U18250 ( .A1(n29868), .A2(\xmem_data[82][6] ), .B1(n29867), .B2(
        \xmem_data[83][6] ), .ZN(n14074) );
  AOI22_X1 U18251 ( .A1(n29870), .A2(\xmem_data[84][6] ), .B1(n29869), .B2(
        \xmem_data[85][6] ), .ZN(n14073) );
  AOI22_X1 U18252 ( .A1(n29871), .A2(\xmem_data[86][6] ), .B1(n29993), .B2(
        \xmem_data[87][6] ), .ZN(n14072) );
  NAND4_X1 U18253 ( .A1(n14075), .A2(n14074), .A3(n14073), .A4(n14072), .ZN(
        n14081) );
  AOI22_X1 U18254 ( .A1(n29877), .A2(\xmem_data[88][6] ), .B1(n29876), .B2(
        \xmem_data[89][6] ), .ZN(n14079) );
  AOI22_X1 U18255 ( .A1(n29879), .A2(\xmem_data[90][6] ), .B1(n29878), .B2(
        \xmem_data[91][6] ), .ZN(n14078) );
  AOI22_X1 U18256 ( .A1(n29881), .A2(\xmem_data[92][6] ), .B1(n29880), .B2(
        \xmem_data[93][6] ), .ZN(n14077) );
  AOI22_X1 U18257 ( .A1(n29883), .A2(\xmem_data[94][6] ), .B1(n29882), .B2(
        \xmem_data[95][6] ), .ZN(n14076) );
  NAND4_X1 U18258 ( .A1(n14079), .A2(n14078), .A3(n14077), .A4(n14076), .ZN(
        n14080) );
  OR4_X1 U18259 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14084) );
  AOI22_X1 U18260 ( .A1(n30007), .A2(n14085), .B1(n30009), .B2(n14084), .ZN(
        n14086) );
  AOI22_X1 U18261 ( .A1(n27568), .A2(\xmem_data[0][7] ), .B1(n27567), .B2(
        \xmem_data[1][7] ), .ZN(n14092) );
  AOI22_X1 U18262 ( .A1(n27564), .A2(\xmem_data[2][7] ), .B1(n27563), .B2(
        \xmem_data[3][7] ), .ZN(n14091) );
  AOI22_X1 U18263 ( .A1(n28039), .A2(\xmem_data[4][7] ), .B1(n28501), .B2(
        \xmem_data[5][7] ), .ZN(n14090) );
  AND2_X1 U18264 ( .A1(n3219), .A2(\xmem_data[7][7] ), .ZN(n14088) );
  AOI21_X1 U18265 ( .B1(n27439), .B2(\xmem_data[6][7] ), .A(n14088), .ZN(
        n14089) );
  NAND4_X1 U18266 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14116) );
  AOI22_X1 U18267 ( .A1(n27516), .A2(\xmem_data[21][7] ), .B1(
        \xmem_data[20][7] ), .B2(n3465), .ZN(n14093) );
  INV_X1 U18268 ( .A(n14093), .ZN(n14099) );
  AOI22_X1 U18269 ( .A1(n27453), .A2(\xmem_data[16][7] ), .B1(n27535), .B2(
        \xmem_data[17][7] ), .ZN(n14095) );
  AOI22_X1 U18270 ( .A1(n20800), .A2(\xmem_data[22][7] ), .B1(n20505), .B2(
        \xmem_data[23][7] ), .ZN(n14094) );
  NAND2_X1 U18271 ( .A1(n14095), .A2(n14094), .ZN(n14098) );
  AOI22_X1 U18272 ( .A1(n28980), .A2(\xmem_data[18][7] ), .B1(n27536), .B2(
        \xmem_data[19][7] ), .ZN(n14096) );
  INV_X1 U18273 ( .A(n14096), .ZN(n14097) );
  AOI22_X1 U18274 ( .A1(n21069), .A2(\xmem_data[10][7] ), .B1(n27550), .B2(
        \xmem_data[11][7] ), .ZN(n14100) );
  AOI22_X1 U18275 ( .A1(n28428), .A2(\xmem_data[26][7] ), .B1(n23778), .B2(
        \xmem_data[27][7] ), .ZN(n14101) );
  INV_X1 U18276 ( .A(n14101), .ZN(n14106) );
  AOI22_X1 U18277 ( .A1(n27542), .A2(\xmem_data[30][7] ), .B1(n28979), .B2(
        \xmem_data[31][7] ), .ZN(n14104) );
  AOI22_X1 U18278 ( .A1(n23802), .A2(\xmem_data[24][7] ), .B1(n13452), .B2(
        \xmem_data[25][7] ), .ZN(n14103) );
  AOI22_X1 U18279 ( .A1(n25636), .A2(\xmem_data[28][7] ), .B1(n14975), .B2(
        \xmem_data[29][7] ), .ZN(n14102) );
  NAND3_X1 U18280 ( .A1(n14104), .A2(n14103), .A3(n14102), .ZN(n14105) );
  NOR3_X1 U18281 ( .A1(n14107), .A2(n14106), .A3(n14105), .ZN(n14114) );
  AOI22_X1 U18282 ( .A1(n27551), .A2(\xmem_data[14][7] ), .B1(n20982), .B2(
        \xmem_data[15][7] ), .ZN(n14108) );
  INV_X1 U18283 ( .A(n14108), .ZN(n14112) );
  AND2_X1 U18284 ( .A1(n29231), .A2(\xmem_data[12][7] ), .ZN(n14111) );
  AOI22_X1 U18285 ( .A1(n29698), .A2(\xmem_data[8][7] ), .B1(n20992), .B2(
        \xmem_data[9][7] ), .ZN(n14109) );
  INV_X1 U18286 ( .A(n14109), .ZN(n14110) );
  NOR3_X1 U18287 ( .A1(n14112), .A2(n14111), .A3(n14110), .ZN(n14113) );
  NAND2_X1 U18288 ( .A1(n14114), .A2(n14113), .ZN(n14115) );
  NOR3_X1 U18289 ( .A1(n14116), .A2(n3918), .A3(n14115), .ZN(n14118) );
  NAND2_X1 U18290 ( .A1(n25450), .A2(\xmem_data[13][7] ), .ZN(n14117) );
  AOI21_X1 U18291 ( .B1(n14118), .B2(n14117), .A(n27573), .ZN(n14119) );
  INV_X1 U18292 ( .A(n14119), .ZN(n14187) );
  AOI22_X1 U18293 ( .A1(n29383), .A2(\xmem_data[96][7] ), .B1(n27435), .B2(
        \xmem_data[97][7] ), .ZN(n14123) );
  AOI22_X1 U18294 ( .A1(n27436), .A2(\xmem_data[98][7] ), .B1(n3203), .B2(
        \xmem_data[99][7] ), .ZN(n14122) );
  AOI22_X1 U18295 ( .A1(n3384), .A2(\xmem_data[100][7] ), .B1(n27437), .B2(
        \xmem_data[101][7] ), .ZN(n14121) );
  AOI22_X1 U18296 ( .A1(n27439), .A2(\xmem_data[102][7] ), .B1(n3219), .B2(
        \xmem_data[103][7] ), .ZN(n14120) );
  NAND4_X1 U18297 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14140) );
  AOI22_X1 U18298 ( .A1(n27453), .A2(\xmem_data[112][7] ), .B1(n27452), .B2(
        \xmem_data[113][7] ), .ZN(n14127) );
  AOI22_X1 U18299 ( .A1(n3175), .A2(\xmem_data[114][7] ), .B1(n29046), .B2(
        \xmem_data[115][7] ), .ZN(n14126) );
  AOI22_X1 U18300 ( .A1(n30543), .A2(\xmem_data[116][7] ), .B1(n27454), .B2(
        \xmem_data[117][7] ), .ZN(n14125) );
  AOI22_X1 U18301 ( .A1(n14937), .A2(\xmem_data[118][7] ), .B1(n28492), .B2(
        \xmem_data[119][7] ), .ZN(n14124) );
  NAND4_X1 U18302 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14138) );
  AOI22_X1 U18303 ( .A1(n29239), .A2(\xmem_data[120][7] ), .B1(n27460), .B2(
        \xmem_data[121][7] ), .ZN(n14131) );
  AOI22_X1 U18304 ( .A1(n27462), .A2(\xmem_data[122][7] ), .B1(n27461), .B2(
        \xmem_data[123][7] ), .ZN(n14130) );
  AOI22_X1 U18305 ( .A1(n3271), .A2(\xmem_data[124][7] ), .B1(n20781), .B2(
        \xmem_data[125][7] ), .ZN(n14129) );
  AOI22_X1 U18306 ( .A1(n3209), .A2(\xmem_data[126][7] ), .B1(n27463), .B2(
        \xmem_data[127][7] ), .ZN(n14128) );
  NAND4_X1 U18307 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14137) );
  AOI22_X1 U18308 ( .A1(n27445), .A2(\xmem_data[104][7] ), .B1(n27444), .B2(
        \xmem_data[105][7] ), .ZN(n14135) );
  AOI22_X1 U18309 ( .A1(n20994), .A2(\xmem_data[106][7] ), .B1(n28342), .B2(
        \xmem_data[107][7] ), .ZN(n14134) );
  AOI22_X1 U18310 ( .A1(n3344), .A2(\xmem_data[108][7] ), .B1(n27446), .B2(
        \xmem_data[109][7] ), .ZN(n14133) );
  AOI22_X1 U18311 ( .A1(n27447), .A2(\xmem_data[110][7] ), .B1(n24590), .B2(
        \xmem_data[111][7] ), .ZN(n14132) );
  NAND4_X1 U18312 ( .A1(n14135), .A2(n14134), .A3(n14133), .A4(n14132), .ZN(
        n14136) );
  OR3_X1 U18313 ( .A1(n14138), .A2(n14137), .A3(n14136), .ZN(n14139) );
  OAI21_X1 U18314 ( .B1(n14140), .B2(n14139), .A(n27496), .ZN(n14186) );
  AOI22_X1 U18315 ( .A1(n27498), .A2(\xmem_data[32][7] ), .B1(n24524), .B2(
        \xmem_data[33][7] ), .ZN(n14144) );
  AOI22_X1 U18316 ( .A1(n27500), .A2(\xmem_data[34][7] ), .B1(n27499), .B2(
        \xmem_data[35][7] ), .ZN(n14143) );
  AOI22_X1 U18317 ( .A1(n3317), .A2(\xmem_data[36][7] ), .B1(n27501), .B2(
        \xmem_data[37][7] ), .ZN(n14142) );
  AOI22_X1 U18318 ( .A1(n27502), .A2(\xmem_data[38][7] ), .B1(n3222), .B2(
        \xmem_data[39][7] ), .ZN(n14141) );
  NAND4_X1 U18319 ( .A1(n14144), .A2(n14143), .A3(n14142), .A4(n14141), .ZN(
        n14161) );
  AOI22_X1 U18320 ( .A1(n28302), .A2(\xmem_data[56][7] ), .B1(n27523), .B2(
        \xmem_data[57][7] ), .ZN(n14148) );
  AOI22_X1 U18321 ( .A1(n27524), .A2(\xmem_data[58][7] ), .B1(n30898), .B2(
        \xmem_data[59][7] ), .ZN(n14147) );
  AOI22_X1 U18322 ( .A1(n20732), .A2(\xmem_data[60][7] ), .B1(n27525), .B2(
        \xmem_data[61][7] ), .ZN(n14146) );
  AOI22_X1 U18323 ( .A1(n31316), .A2(\xmem_data[62][7] ), .B1(n27526), .B2(
        \xmem_data[63][7] ), .ZN(n14145) );
  NAND4_X1 U18324 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        n14159) );
  AOI22_X1 U18325 ( .A1(n27514), .A2(\xmem_data[48][7] ), .B1(n27513), .B2(
        \xmem_data[49][7] ), .ZN(n14152) );
  AOI22_X1 U18326 ( .A1(n27515), .A2(\xmem_data[50][7] ), .B1(n21076), .B2(
        \xmem_data[51][7] ), .ZN(n14151) );
  AOI22_X1 U18327 ( .A1(n30543), .A2(\xmem_data[52][7] ), .B1(n27516), .B2(
        \xmem_data[53][7] ), .ZN(n14150) );
  AOI22_X1 U18328 ( .A1(n13149), .A2(\xmem_data[54][7] ), .B1(n27518), .B2(
        \xmem_data[55][7] ), .ZN(n14149) );
  NAND4_X1 U18329 ( .A1(n14152), .A2(n14151), .A3(n14150), .A4(n14149), .ZN(
        n14158) );
  AOI22_X1 U18330 ( .A1(n22708), .A2(\xmem_data[40][7] ), .B1(n27507), .B2(
        \xmem_data[41][7] ), .ZN(n14156) );
  AOI22_X1 U18331 ( .A1(n29027), .A2(\xmem_data[42][7] ), .B1(n13444), .B2(
        \xmem_data[43][7] ), .ZN(n14155) );
  AOI22_X1 U18332 ( .A1(n30295), .A2(\xmem_data[44][7] ), .B1(n28510), .B2(
        \xmem_data[45][7] ), .ZN(n14154) );
  AOI22_X1 U18333 ( .A1(n27508), .A2(\xmem_data[46][7] ), .B1(n27943), .B2(
        \xmem_data[47][7] ), .ZN(n14153) );
  NAND4_X1 U18334 ( .A1(n14156), .A2(n14155), .A3(n14154), .A4(n14153), .ZN(
        n14157) );
  OAI21_X1 U18335 ( .B1(n14161), .B2(n14160), .A(n27577), .ZN(n14185) );
  AOI22_X1 U18336 ( .A1(n27498), .A2(\xmem_data[64][7] ), .B1(n20769), .B2(
        \xmem_data[65][7] ), .ZN(n14166) );
  AOI22_X1 U18337 ( .A1(n27500), .A2(\xmem_data[66][7] ), .B1(n27499), .B2(
        \xmem_data[67][7] ), .ZN(n14165) );
  AOI22_X1 U18338 ( .A1(n25624), .A2(\xmem_data[68][7] ), .B1(n27501), .B2(
        \xmem_data[69][7] ), .ZN(n14164) );
  AND2_X1 U18339 ( .A1(n3220), .A2(\xmem_data[71][7] ), .ZN(n14162) );
  AOI21_X1 U18340 ( .B1(n27502), .B2(\xmem_data[70][7] ), .A(n14162), .ZN(
        n14163) );
  NAND4_X1 U18341 ( .A1(n14166), .A2(n14165), .A3(n14164), .A4(n14163), .ZN(
        n14183) );
  AOI22_X1 U18342 ( .A1(n29319), .A2(\xmem_data[88][7] ), .B1(n27523), .B2(
        \xmem_data[89][7] ), .ZN(n14170) );
  AOI22_X1 U18343 ( .A1(n27524), .A2(\xmem_data[90][7] ), .B1(n27951), .B2(
        \xmem_data[91][7] ), .ZN(n14169) );
  AOI22_X1 U18344 ( .A1(n20732), .A2(\xmem_data[92][7] ), .B1(n27525), .B2(
        \xmem_data[93][7] ), .ZN(n14168) );
  AOI22_X1 U18345 ( .A1(n3209), .A2(\xmem_data[94][7] ), .B1(n27526), .B2(
        \xmem_data[95][7] ), .ZN(n14167) );
  NAND4_X1 U18346 ( .A1(n14170), .A2(n14169), .A3(n14168), .A4(n14167), .ZN(
        n14181) );
  AOI22_X1 U18347 ( .A1(n27818), .A2(\xmem_data[84][7] ), .B1(n27516), .B2(
        \xmem_data[85][7] ), .ZN(n14174) );
  AOI22_X1 U18348 ( .A1(n27515), .A2(\xmem_data[82][7] ), .B1(n29271), .B2(
        \xmem_data[83][7] ), .ZN(n14173) );
  AOI22_X1 U18349 ( .A1(n27514), .A2(\xmem_data[80][7] ), .B1(n27513), .B2(
        \xmem_data[81][7] ), .ZN(n14172) );
  AOI22_X1 U18350 ( .A1(n29010), .A2(\xmem_data[86][7] ), .B1(n27518), .B2(
        \xmem_data[87][7] ), .ZN(n14171) );
  NAND4_X1 U18351 ( .A1(n14174), .A2(n14173), .A3(n14172), .A4(n14171), .ZN(
        n14180) );
  AOI22_X1 U18352 ( .A1(n27831), .A2(\xmem_data[72][7] ), .B1(n27507), .B2(
        \xmem_data[73][7] ), .ZN(n14178) );
  AOI22_X1 U18353 ( .A1(n29174), .A2(\xmem_data[74][7] ), .B1(n13444), .B2(
        \xmem_data[75][7] ), .ZN(n14177) );
  AOI22_X1 U18354 ( .A1(n28084), .A2(\xmem_data[76][7] ), .B1(n27446), .B2(
        \xmem_data[77][7] ), .ZN(n14176) );
  AOI22_X1 U18355 ( .A1(n27508), .A2(\xmem_data[78][7] ), .B1(n27943), .B2(
        \xmem_data[79][7] ), .ZN(n14175) );
  NAND4_X1 U18356 ( .A1(n14178), .A2(n14177), .A3(n14176), .A4(n14175), .ZN(
        n14179) );
  OR3_X1 U18357 ( .A1(n14181), .A2(n14180), .A3(n14179), .ZN(n14182) );
  OAI21_X1 U18358 ( .B1(n14183), .B2(n14182), .A(n27494), .ZN(n14184) );
  XOR2_X1 U18359 ( .A(\fmem_data[20][3] ), .B(\fmem_data[20][2] ), .Z(n14188)
         );
  AOI22_X1 U18360 ( .A1(n29055), .A2(\xmem_data[48][7] ), .B1(n29054), .B2(
        \xmem_data[49][7] ), .ZN(n14192) );
  AOI22_X1 U18361 ( .A1(n24167), .A2(\xmem_data[50][7] ), .B1(n24166), .B2(
        \xmem_data[51][7] ), .ZN(n14191) );
  AOI22_X1 U18362 ( .A1(n21057), .A2(\xmem_data[52][7] ), .B1(n29820), .B2(
        \xmem_data[53][7] ), .ZN(n14190) );
  AOI22_X1 U18363 ( .A1(n27435), .A2(\xmem_data[54][7] ), .B1(n29057), .B2(
        \xmem_data[55][7] ), .ZN(n14189) );
  NAND4_X1 U18364 ( .A1(n14192), .A2(n14191), .A3(n14190), .A4(n14189), .ZN(
        n14193) );
  NAND2_X1 U18365 ( .A1(n14193), .A2(n29078), .ZN(n14217) );
  AOI22_X1 U18366 ( .A1(n25442), .A2(\xmem_data[90][7] ), .B1(n20991), .B2(
        \xmem_data[91][7] ), .ZN(n14197) );
  AOI22_X1 U18367 ( .A1(n28317), .A2(\xmem_data[88][7] ), .B1(n21308), .B2(
        \xmem_data[89][7] ), .ZN(n14196) );
  AOI22_X1 U18368 ( .A1(n3222), .A2(\xmem_data[92][7] ), .B1(n29065), .B2(
        \xmem_data[93][7] ), .ZN(n14195) );
  AOI22_X1 U18369 ( .A1(n20723), .A2(\xmem_data[94][7] ), .B1(n24697), .B2(
        \xmem_data[95][7] ), .ZN(n14194) );
  NAND4_X1 U18370 ( .A1(n14197), .A2(n14196), .A3(n14195), .A4(n14194), .ZN(
        n14198) );
  NAND2_X1 U18371 ( .A1(n14198), .A2(n29041), .ZN(n14216) );
  AOI22_X1 U18372 ( .A1(n23731), .A2(\xmem_data[26][7] ), .B1(n24443), .B2(
        \xmem_data[27][7] ), .ZN(n14202) );
  AOI22_X1 U18373 ( .A1(n25561), .A2(\xmem_data[24][7] ), .B1(n3333), .B2(
        \xmem_data[25][7] ), .ZN(n14201) );
  AOI22_X1 U18374 ( .A1(n3219), .A2(\xmem_data[28][7] ), .B1(n27831), .B2(
        \xmem_data[29][7] ), .ZN(n14200) );
  AOI22_X1 U18375 ( .A1(n28508), .A2(\xmem_data[30][7] ), .B1(n27904), .B2(
        \xmem_data[31][7] ), .ZN(n14199) );
  NAND4_X1 U18376 ( .A1(n14202), .A2(n14201), .A3(n14200), .A4(n14199), .ZN(
        n14203) );
  NAND2_X1 U18377 ( .A1(n14203), .A2(n29002), .ZN(n14215) );
  AOI22_X1 U18378 ( .A1(n29009), .A2(\xmem_data[104][7] ), .B1(n29008), .B2(
        \xmem_data[105][7] ), .ZN(n14207) );
  AOI22_X1 U18379 ( .A1(n3212), .A2(\xmem_data[106][7] ), .B1(n29010), .B2(
        \xmem_data[107][7] ), .ZN(n14206) );
  AOI22_X1 U18380 ( .A1(n24459), .A2(\xmem_data[108][7] ), .B1(n29012), .B2(
        \xmem_data[109][7] ), .ZN(n14205) );
  AOI22_X1 U18381 ( .A1(n20941), .A2(\xmem_data[110][7] ), .B1(n28428), .B2(
        \xmem_data[111][7] ), .ZN(n14204) );
  NAND4_X1 U18382 ( .A1(n14207), .A2(n14206), .A3(n14205), .A4(n14204), .ZN(
        n14213) );
  AOI22_X1 U18383 ( .A1(n24564), .A2(\xmem_data[32][7] ), .B1(n28344), .B2(
        \xmem_data[33][7] ), .ZN(n14211) );
  AOI22_X1 U18384 ( .A1(n28510), .A2(\xmem_data[34][7] ), .B1(n28972), .B2(
        \xmem_data[35][7] ), .ZN(n14210) );
  AOI22_X1 U18385 ( .A1(n28373), .A2(\xmem_data[36][7] ), .B1(n22738), .B2(
        \xmem_data[37][7] ), .ZN(n14209) );
  AOI22_X1 U18386 ( .A1(n29232), .A2(\xmem_data[38][7] ), .B1(n28334), .B2(
        \xmem_data[39][7] ), .ZN(n14208) );
  NAND4_X1 U18387 ( .A1(n14211), .A2(n14210), .A3(n14209), .A4(n14208), .ZN(
        n14212) );
  AOI22_X1 U18388 ( .A1(n14213), .A2(n28968), .B1(n14212), .B2(n29078), .ZN(
        n14214) );
  NAND4_X1 U18389 ( .A1(n14217), .A2(n14216), .A3(n14215), .A4(n14214), .ZN(
        n14287) );
  AOI22_X1 U18390 ( .A1(n30861), .A2(\xmem_data[56][7] ), .B1(n28164), .B2(
        \xmem_data[57][7] ), .ZN(n14221) );
  AOI22_X1 U18391 ( .A1(n29173), .A2(\xmem_data[58][7] ), .B1(n27902), .B2(
        \xmem_data[59][7] ), .ZN(n14220) );
  AOI22_X1 U18392 ( .A1(n3217), .A2(\xmem_data[60][7] ), .B1(n29065), .B2(
        \xmem_data[61][7] ), .ZN(n14219) );
  AOI22_X1 U18393 ( .A1(n28508), .A2(\xmem_data[62][7] ), .B1(n27904), .B2(
        \xmem_data[63][7] ), .ZN(n14218) );
  NAND4_X1 U18394 ( .A1(n14221), .A2(n14220), .A3(n14219), .A4(n14218), .ZN(
        n14222) );
  NAND2_X1 U18395 ( .A1(n14222), .A2(n29078), .ZN(n14229) );
  AOI22_X1 U18396 ( .A1(n21309), .A2(\xmem_data[120][7] ), .B1(n25624), .B2(
        \xmem_data[121][7] ), .ZN(n14226) );
  AOI22_X1 U18397 ( .A1(n30589), .A2(\xmem_data[122][7] ), .B1(n25413), .B2(
        \xmem_data[123][7] ), .ZN(n14225) );
  AOI22_X1 U18398 ( .A1(n3222), .A2(\xmem_data[124][7] ), .B1(n29026), .B2(
        \xmem_data[125][7] ), .ZN(n14224) );
  AOI22_X1 U18399 ( .A1(n29028), .A2(\xmem_data[126][7] ), .B1(n29027), .B2(
        \xmem_data[127][7] ), .ZN(n14223) );
  NAND4_X1 U18400 ( .A1(n14226), .A2(n14225), .A3(n14224), .A4(n14223), .ZN(
        n14227) );
  NAND2_X1 U18401 ( .A1(n14227), .A2(n28968), .ZN(n14228) );
  NAND2_X1 U18402 ( .A1(n14229), .A2(n14228), .ZN(n14286) );
  AOI22_X1 U18403 ( .A1(n25581), .A2(\xmem_data[16][7] ), .B1(n30645), .B2(
        \xmem_data[17][7] ), .ZN(n14233) );
  AOI22_X1 U18404 ( .A1(n28983), .A2(\xmem_data[18][7] ), .B1(n24467), .B2(
        \xmem_data[19][7] ), .ZN(n14232) );
  AOI22_X1 U18405 ( .A1(n28979), .A2(\xmem_data[20][7] ), .B1(n20708), .B2(
        \xmem_data[21][7] ), .ZN(n14231) );
  AOI22_X1 U18406 ( .A1(n24468), .A2(\xmem_data[22][7] ), .B1(n17030), .B2(
        \xmem_data[23][7] ), .ZN(n14230) );
  NAND4_X1 U18407 ( .A1(n14233), .A2(n14232), .A3(n14231), .A4(n14230), .ZN(
        n14234) );
  NAND2_X1 U18408 ( .A1(n14234), .A2(n29002), .ZN(n14258) );
  AOI22_X1 U18409 ( .A1(n25415), .A2(\xmem_data[64][7] ), .B1(n29567), .B2(
        \xmem_data[65][7] ), .ZN(n14238) );
  AOI22_X1 U18410 ( .A1(n29045), .A2(\xmem_data[66][7] ), .B1(n25422), .B2(
        \xmem_data[67][7] ), .ZN(n14237) );
  AOI22_X1 U18411 ( .A1(n29180), .A2(\xmem_data[68][7] ), .B1(n17064), .B2(
        \xmem_data[69][7] ), .ZN(n14236) );
  AOI22_X1 U18412 ( .A1(n27513), .A2(\xmem_data[70][7] ), .B1(n27913), .B2(
        \xmem_data[71][7] ), .ZN(n14235) );
  NAND4_X1 U18413 ( .A1(n14238), .A2(n14237), .A3(n14236), .A4(n14235), .ZN(
        n14244) );
  AOI22_X1 U18414 ( .A1(n30513), .A2(\xmem_data[8][7] ), .B1(n3157), .B2(
        \xmem_data[9][7] ), .ZN(n14242) );
  AOI22_X1 U18415 ( .A1(n28993), .A2(\xmem_data[10][7] ), .B1(n24593), .B2(
        \xmem_data[11][7] ), .ZN(n14241) );
  AOI22_X1 U18416 ( .A1(n25715), .A2(\xmem_data[12][7] ), .B1(n28994), .B2(
        \xmem_data[13][7] ), .ZN(n14240) );
  AOI22_X1 U18417 ( .A1(n28380), .A2(\xmem_data[14][7] ), .B1(n3204), .B2(
        \xmem_data[15][7] ), .ZN(n14239) );
  NAND4_X1 U18418 ( .A1(n14242), .A2(n14241), .A3(n14240), .A4(n14239), .ZN(
        n14243) );
  AOI22_X1 U18419 ( .A1(n14244), .A2(n29041), .B1(n14243), .B2(n29002), .ZN(
        n14257) );
  AOI22_X1 U18420 ( .A1(n20559), .A2(\xmem_data[0][7] ), .B1(n28952), .B2(
        \xmem_data[1][7] ), .ZN(n14248) );
  AOI22_X1 U18421 ( .A1(n25450), .A2(\xmem_data[2][7] ), .B1(n24638), .B2(
        \xmem_data[3][7] ), .ZN(n14247) );
  AOI22_X1 U18422 ( .A1(n22701), .A2(\xmem_data[4][7] ), .B1(n23792), .B2(
        \xmem_data[5][7] ), .ZN(n14246) );
  AOI22_X1 U18423 ( .A1(n28345), .A2(\xmem_data[6][7] ), .B1(n25710), .B2(
        \xmem_data[7][7] ), .ZN(n14245) );
  NAND4_X1 U18424 ( .A1(n14248), .A2(n14247), .A3(n14246), .A4(n14245), .ZN(
        n14249) );
  NAND2_X1 U18425 ( .A1(n14249), .A2(n29002), .ZN(n14256) );
  AOI22_X1 U18426 ( .A1(n24140), .A2(\xmem_data[96][7] ), .B1(n3374), .B2(
        \xmem_data[97][7] ), .ZN(n14253) );
  AOI22_X1 U18427 ( .A1(n29045), .A2(\xmem_data[98][7] ), .B1(n27447), .B2(
        \xmem_data[99][7] ), .ZN(n14252) );
  AOI22_X1 U18428 ( .A1(n3357), .A2(\xmem_data[100][7] ), .B1(n28089), .B2(
        \xmem_data[101][7] ), .ZN(n14251) );
  AOI22_X1 U18429 ( .A1(n22740), .A2(\xmem_data[102][7] ), .B1(n30891), .B2(
        \xmem_data[103][7] ), .ZN(n14250) );
  NAND4_X1 U18430 ( .A1(n14253), .A2(n14252), .A3(n14251), .A4(n14250), .ZN(
        n14254) );
  NAND2_X1 U18431 ( .A1(n14254), .A2(n28968), .ZN(n14255) );
  NAND4_X1 U18432 ( .A1(n14258), .A2(n14257), .A3(n14256), .A4(n14255), .ZN(
        n14285) );
  AOI22_X1 U18433 ( .A1(n25716), .A2(\xmem_data[112][7] ), .B1(n28955), .B2(
        \xmem_data[113][7] ), .ZN(n14262) );
  AOI22_X1 U18434 ( .A1(n28983), .A2(\xmem_data[114][7] ), .B1(n3179), .B2(
        \xmem_data[115][7] ), .ZN(n14261) );
  AOI22_X1 U18435 ( .A1(n29017), .A2(\xmem_data[116][7] ), .B1(n20770), .B2(
        \xmem_data[117][7] ), .ZN(n14260) );
  AOI22_X1 U18436 ( .A1(n20951), .A2(\xmem_data[118][7] ), .B1(n30909), .B2(
        \xmem_data[119][7] ), .ZN(n14259) );
  NAND4_X1 U18437 ( .A1(n14262), .A2(n14261), .A3(n14260), .A4(n14259), .ZN(
        n14263) );
  NAND2_X1 U18438 ( .A1(n14263), .A2(n28968), .ZN(n14283) );
  AOI22_X1 U18439 ( .A1(n14975), .A2(\xmem_data[82][7] ), .B1(n20552), .B2(
        \xmem_data[83][7] ), .ZN(n14267) );
  AOI22_X1 U18440 ( .A1(n29055), .A2(\xmem_data[80][7] ), .B1(n29054), .B2(
        \xmem_data[81][7] ), .ZN(n14266) );
  AOI22_X1 U18441 ( .A1(n24524), .A2(\xmem_data[86][7] ), .B1(n29057), .B2(
        \xmem_data[87][7] ), .ZN(n14265) );
  NAND4_X1 U18442 ( .A1(n14268), .A2(n14267), .A3(n14266), .A4(n14265), .ZN(
        n14269) );
  NAND2_X1 U18443 ( .A1(n14269), .A2(n29041), .ZN(n14282) );
  AOI22_X1 U18444 ( .A1(n29046), .A2(\xmem_data[72][7] ), .B1(n30666), .B2(
        \xmem_data[73][7] ), .ZN(n14273) );
  AOI22_X1 U18445 ( .A1(n3213), .A2(\xmem_data[74][7] ), .B1(n13149), .B2(
        \xmem_data[75][7] ), .ZN(n14272) );
  AOI22_X1 U18446 ( .A1(n29048), .A2(\xmem_data[76][7] ), .B1(n29047), .B2(
        \xmem_data[77][7] ), .ZN(n14271) );
  AOI22_X1 U18447 ( .A1(n29049), .A2(\xmem_data[78][7] ), .B1(n28428), .B2(
        \xmem_data[79][7] ), .ZN(n14270) );
  NAND4_X1 U18448 ( .A1(n14273), .A2(n14272), .A3(n14271), .A4(n14270), .ZN(
        n14274) );
  NAND2_X1 U18449 ( .A1(n14274), .A2(n29041), .ZN(n14281) );
  AOI22_X1 U18450 ( .A1(n29046), .A2(\xmem_data[40][7] ), .B1(n29437), .B2(
        \xmem_data[41][7] ), .ZN(n14278) );
  AOI22_X1 U18451 ( .A1(n25383), .A2(\xmem_data[42][7] ), .B1(n20585), .B2(
        \xmem_data[43][7] ), .ZN(n14277) );
  AOI22_X1 U18452 ( .A1(n29048), .A2(\xmem_data[44][7] ), .B1(n29047), .B2(
        \xmem_data[45][7] ), .ZN(n14276) );
  AOI22_X1 U18453 ( .A1(n29049), .A2(\xmem_data[46][7] ), .B1(n30849), .B2(
        \xmem_data[47][7] ), .ZN(n14275) );
  NAND4_X1 U18454 ( .A1(n14278), .A2(n14277), .A3(n14276), .A4(n14275), .ZN(
        n14279) );
  NAND2_X1 U18455 ( .A1(n14279), .A2(n29078), .ZN(n14280) );
  NAND4_X1 U18456 ( .A1(n14283), .A2(n14282), .A3(n14281), .A4(n14280), .ZN(
        n14284) );
  XNOR2_X1 U18457 ( .A(n35338), .B(\fmem_data[9][3] ), .ZN(n33044) );
  INV_X1 U18458 ( .A(n14288), .ZN(n23599) );
  AOI22_X1 U18459 ( .A1(n22708), .A2(\xmem_data[32][5] ), .B1(n30963), .B2(
        \xmem_data[33][5] ), .ZN(n14292) );
  AOI22_X1 U18460 ( .A1(n20994), .A2(\xmem_data[34][5] ), .B1(n31275), .B2(
        \xmem_data[35][5] ), .ZN(n14291) );
  AOI22_X1 U18461 ( .A1(n22668), .A2(\xmem_data[36][5] ), .B1(n25450), .B2(
        \xmem_data[37][5] ), .ZN(n14290) );
  AOI22_X1 U18462 ( .A1(n31321), .A2(\xmem_data[38][5] ), .B1(n13475), .B2(
        \xmem_data[39][5] ), .ZN(n14289) );
  NAND4_X1 U18463 ( .A1(n14292), .A2(n14291), .A3(n14290), .A4(n14289), .ZN(
        n14308) );
  AOI22_X1 U18464 ( .A1(n31327), .A2(\xmem_data[40][5] ), .B1(n31326), .B2(
        \xmem_data[41][5] ), .ZN(n14296) );
  AOI22_X1 U18465 ( .A1(n29272), .A2(\xmem_data[42][5] ), .B1(n25572), .B2(
        \xmem_data[43][5] ), .ZN(n14295) );
  AOI22_X1 U18466 ( .A1(n31328), .A2(\xmem_data[44][5] ), .B1(n23716), .B2(
        \xmem_data[45][5] ), .ZN(n14294) );
  AOI22_X1 U18467 ( .A1(n31330), .A2(\xmem_data[46][5] ), .B1(n31329), .B2(
        \xmem_data[47][5] ), .ZN(n14293) );
  NAND4_X1 U18468 ( .A1(n14296), .A2(n14295), .A3(n14294), .A4(n14293), .ZN(
        n14307) );
  AOI22_X1 U18469 ( .A1(n20730), .A2(\xmem_data[48][5] ), .B1(n23776), .B2(
        \xmem_data[49][5] ), .ZN(n14300) );
  AOI22_X1 U18470 ( .A1(n20731), .A2(\xmem_data[50][5] ), .B1(n28429), .B2(
        \xmem_data[51][5] ), .ZN(n14299) );
  AOI22_X1 U18471 ( .A1(n31315), .A2(\xmem_data[52][5] ), .B1(n31314), .B2(
        \xmem_data[53][5] ), .ZN(n14298) );
  AOI22_X1 U18472 ( .A1(n31316), .A2(\xmem_data[54][5] ), .B1(n25406), .B2(
        \xmem_data[55][5] ), .ZN(n14297) );
  NAND4_X1 U18473 ( .A1(n14300), .A2(n14299), .A3(n14298), .A4(n14297), .ZN(
        n14306) );
  AOI22_X1 U18474 ( .A1(n31308), .A2(\xmem_data[56][5] ), .B1(n20769), .B2(
        \xmem_data[57][5] ), .ZN(n14304) );
  AOI22_X1 U18475 ( .A1(n24607), .A2(\xmem_data[58][5] ), .B1(n31309), .B2(
        \xmem_data[59][5] ), .ZN(n14303) );
  AOI22_X1 U18476 ( .A1(n3245), .A2(\xmem_data[60][5] ), .B1(n3247), .B2(
        \xmem_data[61][5] ), .ZN(n14302) );
  AOI22_X1 U18477 ( .A1(n30962), .A2(\xmem_data[62][5] ), .B1(n3218), .B2(
        \xmem_data[63][5] ), .ZN(n14301) );
  NAND4_X1 U18478 ( .A1(n14304), .A2(n14303), .A3(n14302), .A4(n14301), .ZN(
        n14305) );
  OR4_X1 U18479 ( .A1(n14308), .A2(n14307), .A3(n14306), .A4(n14305), .ZN(
        n14310) );
  NOR2_X1 U18480 ( .A1(n31041), .A2(n39026), .ZN(n14309) );
  AOI21_X1 U18481 ( .B1(n14310), .B2(n31340), .A(n3899), .ZN(n14382) );
  AOI22_X1 U18482 ( .A1(n31345), .A2(\xmem_data[120][5] ), .B1(n31344), .B2(
        \xmem_data[121][5] ), .ZN(n14314) );
  AOI22_X1 U18483 ( .A1(n24688), .A2(\xmem_data[122][5] ), .B1(n31346), .B2(
        \xmem_data[123][5] ), .ZN(n14313) );
  AOI22_X1 U18484 ( .A1(n3352), .A2(\xmem_data[124][5] ), .B1(n31347), .B2(
        \xmem_data[125][5] ), .ZN(n14312) );
  AOI22_X1 U18485 ( .A1(n31348), .A2(\xmem_data[126][5] ), .B1(n3221), .B2(
        \xmem_data[127][5] ), .ZN(n14311) );
  NAND4_X1 U18486 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        n14331) );
  AOI22_X1 U18487 ( .A1(n31353), .A2(\xmem_data[104][5] ), .B1(n30552), .B2(
        \xmem_data[105][5] ), .ZN(n14318) );
  AOI22_X1 U18488 ( .A1(n27913), .A2(\xmem_data[106][5] ), .B1(n14999), .B2(
        \xmem_data[107][5] ), .ZN(n14317) );
  AOI22_X1 U18489 ( .A1(n30948), .A2(\xmem_data[108][5] ), .B1(n3212), .B2(
        \xmem_data[109][5] ), .ZN(n14316) );
  AOI22_X1 U18490 ( .A1(n23717), .A2(\xmem_data[110][5] ), .B1(n31355), .B2(
        \xmem_data[111][5] ), .ZN(n14315) );
  NAND4_X1 U18491 ( .A1(n14318), .A2(n14317), .A3(n14316), .A4(n14315), .ZN(
        n14329) );
  AOI22_X1 U18492 ( .A1(n30309), .A2(\xmem_data[112][5] ), .B1(n31360), .B2(
        \xmem_data[113][5] ), .ZN(n14322) );
  AOI22_X1 U18493 ( .A1(n25717), .A2(\xmem_data[114][5] ), .B1(n31361), .B2(
        \xmem_data[115][5] ), .ZN(n14321) );
  AOI22_X1 U18494 ( .A1(n25401), .A2(\xmem_data[116][5] ), .B1(n31362), .B2(
        \xmem_data[117][5] ), .ZN(n14320) );
  AOI22_X1 U18495 ( .A1(n20734), .A2(\xmem_data[118][5] ), .B1(n23725), .B2(
        \xmem_data[119][5] ), .ZN(n14319) );
  NAND4_X1 U18496 ( .A1(n14322), .A2(n14321), .A3(n14320), .A4(n14319), .ZN(
        n14328) );
  AOI22_X1 U18497 ( .A1(n31368), .A2(\xmem_data[96][5] ), .B1(n31367), .B2(
        \xmem_data[97][5] ), .ZN(n14326) );
  AOI22_X1 U18498 ( .A1(n20725), .A2(\xmem_data[98][5] ), .B1(n29104), .B2(
        \xmem_data[99][5] ), .ZN(n14325) );
  AOI22_X1 U18499 ( .A1(n3344), .A2(\xmem_data[100][5] ), .B1(n24657), .B2(
        \xmem_data[101][5] ), .ZN(n14324) );
  AOI22_X1 U18500 ( .A1(n25422), .A2(\xmem_data[102][5] ), .B1(n14933), .B2(
        \xmem_data[103][5] ), .ZN(n14323) );
  NAND4_X1 U18501 ( .A1(n14326), .A2(n14325), .A3(n14324), .A4(n14323), .ZN(
        n14327) );
  AOI22_X1 U18502 ( .A1(n31308), .A2(\xmem_data[88][5] ), .B1(n30900), .B2(
        \xmem_data[89][5] ), .ZN(n14335) );
  AOI22_X1 U18503 ( .A1(n20827), .A2(\xmem_data[90][5] ), .B1(n31309), .B2(
        \xmem_data[91][5] ), .ZN(n14334) );
  AOI22_X1 U18504 ( .A1(n28973), .A2(\xmem_data[92][5] ), .B1(n29253), .B2(
        \xmem_data[93][5] ), .ZN(n14333) );
  AOI22_X1 U18505 ( .A1(n20991), .A2(\xmem_data[94][5] ), .B1(n3220), .B2(
        \xmem_data[95][5] ), .ZN(n14332) );
  NAND4_X1 U18506 ( .A1(n14335), .A2(n14334), .A3(n14333), .A4(n14332), .ZN(
        n14352) );
  AOI22_X1 U18507 ( .A1(n29319), .A2(\xmem_data[80][5] ), .B1(n23801), .B2(
        \xmem_data[81][5] ), .ZN(n14339) );
  AOI22_X1 U18508 ( .A1(n30557), .A2(\xmem_data[82][5] ), .B1(n25581), .B2(
        \xmem_data[83][5] ), .ZN(n14338) );
  AOI22_X1 U18509 ( .A1(n31315), .A2(\xmem_data[84][5] ), .B1(n31314), .B2(
        \xmem_data[85][5] ), .ZN(n14337) );
  AOI22_X1 U18510 ( .A1(n31316), .A2(\xmem_data[86][5] ), .B1(n28292), .B2(
        \xmem_data[87][5] ), .ZN(n14336) );
  NAND4_X1 U18511 ( .A1(n14339), .A2(n14338), .A3(n14337), .A4(n14336), .ZN(
        n14350) );
  AOI22_X1 U18512 ( .A1(n24533), .A2(\xmem_data[64][5] ), .B1(n28476), .B2(
        \xmem_data[65][5] ), .ZN(n14343) );
  AOI22_X1 U18513 ( .A1(n20725), .A2(\xmem_data[66][5] ), .B1(n22759), .B2(
        \xmem_data[67][5] ), .ZN(n14342) );
  AOI22_X1 U18514 ( .A1(n3281), .A2(\xmem_data[68][5] ), .B1(n25492), .B2(
        \xmem_data[69][5] ), .ZN(n14341) );
  AOI22_X1 U18515 ( .A1(n31321), .A2(\xmem_data[70][5] ), .B1(n13475), .B2(
        \xmem_data[71][5] ), .ZN(n14340) );
  NAND4_X1 U18516 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n14340), .ZN(
        n14349) );
  AOI22_X1 U18517 ( .A1(n31327), .A2(\xmem_data[72][5] ), .B1(n31326), .B2(
        \xmem_data[73][5] ), .ZN(n14347) );
  AOI22_X1 U18518 ( .A1(n29023), .A2(\xmem_data[74][5] ), .B1(n25382), .B2(
        \xmem_data[75][5] ), .ZN(n14346) );
  AOI22_X1 U18519 ( .A1(n31328), .A2(\xmem_data[76][5] ), .B1(n3207), .B2(
        \xmem_data[77][5] ), .ZN(n14345) );
  AOI22_X1 U18520 ( .A1(n31330), .A2(\xmem_data[78][5] ), .B1(n31329), .B2(
        \xmem_data[79][5] ), .ZN(n14344) );
  NAND4_X1 U18521 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14348) );
  AOI22_X1 U18522 ( .A1(n31255), .A2(\xmem_data[16][5] ), .B1(n31254), .B2(
        \xmem_data[17][5] ), .ZN(n14356) );
  AOI22_X1 U18523 ( .A1(n24548), .A2(\xmem_data[18][5] ), .B1(n25364), .B2(
        \xmem_data[19][5] ), .ZN(n14355) );
  AOI22_X1 U18524 ( .A1(n30269), .A2(\xmem_data[20][5] ), .B1(n31362), .B2(
        \xmem_data[21][5] ), .ZN(n14354) );
  AOI22_X1 U18525 ( .A1(n30497), .A2(\xmem_data[22][5] ), .B1(n31256), .B2(
        \xmem_data[23][5] ), .ZN(n14353) );
  NAND4_X1 U18526 ( .A1(n14356), .A2(n14355), .A3(n14354), .A4(n14353), .ZN(
        n14359) );
  AOI22_X1 U18527 ( .A1(n3387), .A2(\xmem_data[28][5] ), .B1(n22753), .B2(
        \xmem_data[29][5] ), .ZN(n14357) );
  NOR2_X1 U18528 ( .A1(n14359), .A2(n14358), .ZN(n14363) );
  AOI22_X1 U18529 ( .A1(n25354), .A2(\xmem_data[30][5] ), .B1(n3219), .B2(
        \xmem_data[31][5] ), .ZN(n14362) );
  AOI22_X1 U18530 ( .A1(n3380), .A2(\xmem_data[26][5] ), .B1(n31262), .B2(
        \xmem_data[27][5] ), .ZN(n14361) );
  AOI22_X1 U18531 ( .A1(n23753), .A2(\xmem_data[24][5] ), .B1(n31261), .B2(
        \xmem_data[25][5] ), .ZN(n14360) );
  AOI22_X1 U18532 ( .A1(n29565), .A2(\xmem_data[0][5] ), .B1(n30963), .B2(
        \xmem_data[1][5] ), .ZN(n14370) );
  AOI22_X1 U18533 ( .A1(n17010), .A2(\xmem_data[2][5] ), .B1(n31275), .B2(
        \xmem_data[3][5] ), .ZN(n14364) );
  INV_X1 U18534 ( .A(n14364), .ZN(n14368) );
  AOI22_X1 U18535 ( .A1(n31276), .A2(\xmem_data[6][5] ), .B1(n27943), .B2(
        \xmem_data[7][5] ), .ZN(n14366) );
  NAND2_X1 U18536 ( .A1(n3375), .A2(\xmem_data[4][5] ), .ZN(n14365) );
  NAND2_X1 U18537 ( .A1(n14366), .A2(n14365), .ZN(n14367) );
  NOR2_X1 U18538 ( .A1(n14368), .A2(n14367), .ZN(n14369) );
  NAND2_X1 U18539 ( .A1(n14370), .A2(n14369), .ZN(n14376) );
  AOI22_X1 U18540 ( .A1(n28233), .A2(\xmem_data[8][5] ), .B1(n24448), .B2(
        \xmem_data[9][5] ), .ZN(n14374) );
  AOI22_X1 U18541 ( .A1(n31268), .A2(\xmem_data[10][5] ), .B1(n25382), .B2(
        \xmem_data[11][5] ), .ZN(n14373) );
  AOI22_X1 U18542 ( .A1(n31354), .A2(\xmem_data[12][5] ), .B1(n31269), .B2(
        \xmem_data[13][5] ), .ZN(n14372) );
  AOI22_X1 U18543 ( .A1(n27919), .A2(\xmem_data[14][5] ), .B1(n31270), .B2(
        \xmem_data[15][5] ), .ZN(n14371) );
  NAND4_X1 U18544 ( .A1(n14374), .A2(n14373), .A3(n14372), .A4(n14371), .ZN(
        n14375) );
  OR2_X1 U18545 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  XOR2_X1 U18546 ( .A(\fmem_data[12][4] ), .B(\fmem_data[12][5] ), .Z(n14383)
         );
  AOI22_X1 U18547 ( .A1(n31345), .A2(\xmem_data[120][6] ), .B1(n31344), .B2(
        \xmem_data[121][6] ), .ZN(n14388) );
  AOI22_X1 U18548 ( .A1(n27564), .A2(\xmem_data[122][6] ), .B1(n31346), .B2(
        \xmem_data[123][6] ), .ZN(n14387) );
  AOI22_X1 U18549 ( .A1(n3434), .A2(\xmem_data[124][6] ), .B1(n31347), .B2(
        \xmem_data[125][6] ), .ZN(n14386) );
  AND2_X1 U18550 ( .A1(n3220), .A2(\xmem_data[127][6] ), .ZN(n14384) );
  AOI21_X1 U18551 ( .B1(n31348), .B2(\xmem_data[126][6] ), .A(n14384), .ZN(
        n14385) );
  NAND4_X1 U18552 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14405) );
  AOI22_X1 U18553 ( .A1(n25425), .A2(\xmem_data[106][6] ), .B1(n25671), .B2(
        \xmem_data[107][6] ), .ZN(n14392) );
  AOI22_X1 U18554 ( .A1(n31353), .A2(\xmem_data[104][6] ), .B1(n28345), .B2(
        \xmem_data[105][6] ), .ZN(n14391) );
  AOI22_X1 U18555 ( .A1(n29317), .A2(\xmem_data[110][6] ), .B1(n31355), .B2(
        \xmem_data[111][6] ), .ZN(n14390) );
  AOI22_X1 U18556 ( .A1(n31269), .A2(\xmem_data[109][6] ), .B1(
        \xmem_data[108][6] ), .B2(n25461), .ZN(n14389) );
  NAND4_X1 U18557 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n14403) );
  AOI22_X1 U18558 ( .A1(n16990), .A2(\xmem_data[112][6] ), .B1(n31360), .B2(
        \xmem_data[113][6] ), .ZN(n14396) );
  AOI22_X1 U18559 ( .A1(n21010), .A2(\xmem_data[114][6] ), .B1(n31361), .B2(
        \xmem_data[115][6] ), .ZN(n14395) );
  AOI22_X1 U18560 ( .A1(n25401), .A2(\xmem_data[116][6] ), .B1(n31362), .B2(
        \xmem_data[117][6] ), .ZN(n14394) );
  AOI22_X1 U18561 ( .A1(n24685), .A2(\xmem_data[118][6] ), .B1(n20733), .B2(
        \xmem_data[119][6] ), .ZN(n14393) );
  NAND4_X1 U18562 ( .A1(n14396), .A2(n14395), .A3(n14394), .A4(n14393), .ZN(
        n14402) );
  AOI22_X1 U18563 ( .A1(n31368), .A2(\xmem_data[96][6] ), .B1(n31367), .B2(
        \xmem_data[97][6] ), .ZN(n14400) );
  AOI22_X1 U18564 ( .A1(n20725), .A2(\xmem_data[98][6] ), .B1(n22759), .B2(
        \xmem_data[99][6] ), .ZN(n14399) );
  AOI22_X1 U18565 ( .A1(n21074), .A2(\xmem_data[100][6] ), .B1(n29103), .B2(
        \xmem_data[101][6] ), .ZN(n14398) );
  AOI22_X1 U18566 ( .A1(n25422), .A2(\xmem_data[102][6] ), .B1(n27943), .B2(
        \xmem_data[103][6] ), .ZN(n14397) );
  NAND4_X1 U18567 ( .A1(n14400), .A2(n14399), .A3(n14398), .A4(n14397), .ZN(
        n14401) );
  OR3_X1 U18568 ( .A1(n14403), .A2(n14402), .A3(n14401), .ZN(n14404) );
  OR2_X1 U18569 ( .A1(n14405), .A2(n14404), .ZN(n14427) );
  AOI22_X1 U18570 ( .A1(n29494), .A2(\xmem_data[64][6] ), .B1(n23769), .B2(
        \xmem_data[65][6] ), .ZN(n14409) );
  AOI22_X1 U18571 ( .A1(n29174), .A2(\xmem_data[66][6] ), .B1(n24633), .B2(
        \xmem_data[67][6] ), .ZN(n14408) );
  AOI22_X1 U18572 ( .A1(n3375), .A2(\xmem_data[68][6] ), .B1(n25492), .B2(
        \xmem_data[69][6] ), .ZN(n14407) );
  AOI22_X1 U18573 ( .A1(n31321), .A2(\xmem_data[70][6] ), .B1(n29180), .B2(
        \xmem_data[71][6] ), .ZN(n14406) );
  NAND4_X1 U18574 ( .A1(n14409), .A2(n14408), .A3(n14407), .A4(n14406), .ZN(
        n14425) );
  AOI22_X1 U18575 ( .A1(n31327), .A2(\xmem_data[72][6] ), .B1(n31326), .B2(
        \xmem_data[73][6] ), .ZN(n14413) );
  AOI22_X1 U18576 ( .A1(n29272), .A2(\xmem_data[74][6] ), .B1(n22741), .B2(
        \xmem_data[75][6] ), .ZN(n14412) );
  AOI22_X1 U18577 ( .A1(n31328), .A2(\xmem_data[76][6] ), .B1(n20543), .B2(
        \xmem_data[77][6] ), .ZN(n14411) );
  AOI22_X1 U18578 ( .A1(n31330), .A2(\xmem_data[78][6] ), .B1(n31329), .B2(
        \xmem_data[79][6] ), .ZN(n14410) );
  NAND4_X1 U18579 ( .A1(n14413), .A2(n14412), .A3(n14411), .A4(n14410), .ZN(
        n14424) );
  AOI22_X1 U18580 ( .A1(n17044), .A2(\xmem_data[80][6] ), .B1(n29190), .B2(
        \xmem_data[81][6] ), .ZN(n14417) );
  AOI22_X1 U18581 ( .A1(n25521), .A2(\xmem_data[82][6] ), .B1(n20506), .B2(
        \xmem_data[83][6] ), .ZN(n14416) );
  AOI22_X1 U18582 ( .A1(n31315), .A2(\xmem_data[84][6] ), .B1(n31314), .B2(
        \xmem_data[85][6] ), .ZN(n14415) );
  AOI22_X1 U18583 ( .A1(n31316), .A2(\xmem_data[86][6] ), .B1(n25406), .B2(
        \xmem_data[87][6] ), .ZN(n14414) );
  NAND4_X1 U18584 ( .A1(n14417), .A2(n14416), .A3(n14415), .A4(n14414), .ZN(
        n14423) );
  AOI22_X1 U18585 ( .A1(n31308), .A2(\xmem_data[88][6] ), .B1(n20769), .B2(
        \xmem_data[89][6] ), .ZN(n14421) );
  AOI22_X1 U18586 ( .A1(n25358), .A2(\xmem_data[90][6] ), .B1(n31309), .B2(
        \xmem_data[91][6] ), .ZN(n14420) );
  AOI22_X1 U18587 ( .A1(n3317), .A2(\xmem_data[92][6] ), .B1(n28501), .B2(
        \xmem_data[93][6] ), .ZN(n14419) );
  AOI22_X1 U18588 ( .A1(n30906), .A2(\xmem_data[94][6] ), .B1(n3217), .B2(
        \xmem_data[95][6] ), .ZN(n14418) );
  NAND4_X1 U18589 ( .A1(n14421), .A2(n14420), .A3(n14419), .A4(n14418), .ZN(
        n14422) );
  OR4_X1 U18590 ( .A1(n14425), .A2(n14424), .A3(n14423), .A4(n14422), .ZN(
        n14426) );
  AOI22_X1 U18591 ( .A1(n31376), .A2(n14427), .B1(n31342), .B2(n14426), .ZN(
        n14471) );
  AOI22_X1 U18592 ( .A1(n29422), .A2(\xmem_data[32][6] ), .B1(n28508), .B2(
        \xmem_data[33][6] ), .ZN(n14431) );
  AOI22_X1 U18593 ( .A1(n24697), .A2(\xmem_data[34][6] ), .B1(n30882), .B2(
        \xmem_data[35][6] ), .ZN(n14430) );
  AOI22_X1 U18594 ( .A1(n30710), .A2(\xmem_data[36][6] ), .B1(n27547), .B2(
        \xmem_data[37][6] ), .ZN(n14429) );
  AOI22_X1 U18595 ( .A1(n31321), .A2(\xmem_data[38][6] ), .B1(n3357), .B2(
        \xmem_data[39][6] ), .ZN(n14428) );
  NAND4_X1 U18596 ( .A1(n14431), .A2(n14430), .A3(n14429), .A4(n14428), .ZN(
        n14447) );
  AOI22_X1 U18597 ( .A1(n31327), .A2(\xmem_data[40][6] ), .B1(n31326), .B2(
        \xmem_data[41][6] ), .ZN(n14435) );
  AOI22_X1 U18598 ( .A1(n3176), .A2(\xmem_data[42][6] ), .B1(n25458), .B2(
        \xmem_data[43][6] ), .ZN(n14434) );
  AOI22_X1 U18599 ( .A1(n31328), .A2(\xmem_data[44][6] ), .B1(n28335), .B2(
        \xmem_data[45][6] ), .ZN(n14433) );
  AOI22_X1 U18600 ( .A1(n31330), .A2(\xmem_data[46][6] ), .B1(n31329), .B2(
        \xmem_data[47][6] ), .ZN(n14432) );
  NAND4_X1 U18601 ( .A1(n14435), .A2(n14434), .A3(n14433), .A4(n14432), .ZN(
        n14446) );
  AOI22_X1 U18602 ( .A1(n29239), .A2(\xmem_data[48][6] ), .B1(n28380), .B2(
        \xmem_data[49][6] ), .ZN(n14439) );
  AOI22_X1 U18603 ( .A1(n20731), .A2(\xmem_data[50][6] ), .B1(n21009), .B2(
        \xmem_data[51][6] ), .ZN(n14438) );
  AOI22_X1 U18604 ( .A1(n31315), .A2(\xmem_data[52][6] ), .B1(n31314), .B2(
        \xmem_data[53][6] ), .ZN(n14437) );
  AOI22_X1 U18605 ( .A1(n31316), .A2(\xmem_data[54][6] ), .B1(n11008), .B2(
        \xmem_data[55][6] ), .ZN(n14436) );
  NAND4_X1 U18606 ( .A1(n14439), .A2(n14438), .A3(n14437), .A4(n14436), .ZN(
        n14445) );
  AOI22_X1 U18607 ( .A1(n31308), .A2(\xmem_data[56][6] ), .B1(n20769), .B2(
        \xmem_data[57][6] ), .ZN(n14443) );
  AOI22_X1 U18608 ( .A1(n25630), .A2(\xmem_data[58][6] ), .B1(n31309), .B2(
        \xmem_data[59][6] ), .ZN(n14442) );
  AOI22_X1 U18609 ( .A1(n3334), .A2(\xmem_data[60][6] ), .B1(n3247), .B2(
        \xmem_data[61][6] ), .ZN(n14441) );
  AOI22_X1 U18610 ( .A1(n28044), .A2(\xmem_data[62][6] ), .B1(n3218), .B2(
        \xmem_data[63][6] ), .ZN(n14440) );
  NAND4_X1 U18611 ( .A1(n14443), .A2(n14442), .A3(n14441), .A4(n14440), .ZN(
        n14444) );
  OR4_X1 U18612 ( .A1(n14447), .A2(n14446), .A3(n14445), .A4(n14444), .ZN(
        n14469) );
  AOI22_X1 U18613 ( .A1(n29422), .A2(\xmem_data[0][6] ), .B1(n20500), .B2(
        \xmem_data[1][6] ), .ZN(n14451) );
  AOI22_X1 U18614 ( .A1(n27904), .A2(\xmem_data[2][6] ), .B1(n31275), .B2(
        \xmem_data[3][6] ), .ZN(n14450) );
  AOI22_X1 U18615 ( .A1(n29231), .A2(\xmem_data[4][6] ), .B1(n29306), .B2(
        \xmem_data[5][6] ), .ZN(n14449) );
  AOI22_X1 U18616 ( .A1(n31276), .A2(\xmem_data[6][6] ), .B1(n3357), .B2(
        \xmem_data[7][6] ), .ZN(n14448) );
  NAND4_X1 U18617 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        n14467) );
  AOI22_X1 U18618 ( .A1(n30943), .A2(\xmem_data[8][6] ), .B1(n28416), .B2(
        \xmem_data[9][6] ), .ZN(n14455) );
  AOI22_X1 U18619 ( .A1(n31268), .A2(\xmem_data[10][6] ), .B1(n23715), .B2(
        \xmem_data[11][6] ), .ZN(n14454) );
  AOI22_X1 U18620 ( .A1(n31354), .A2(\xmem_data[12][6] ), .B1(n31269), .B2(
        \xmem_data[13][6] ), .ZN(n14453) );
  AOI22_X1 U18621 ( .A1(n13149), .A2(\xmem_data[14][6] ), .B1(n31270), .B2(
        \xmem_data[15][6] ), .ZN(n14452) );
  NAND4_X1 U18622 ( .A1(n14455), .A2(n14454), .A3(n14453), .A4(n14452), .ZN(
        n14466) );
  AOI22_X1 U18623 ( .A1(n31255), .A2(\xmem_data[16][6] ), .B1(n31254), .B2(
        \xmem_data[17][6] ), .ZN(n14459) );
  AOI22_X1 U18624 ( .A1(n3206), .A2(\xmem_data[18][6] ), .B1(n25581), .B2(
        \xmem_data[19][6] ), .ZN(n14458) );
  AOI22_X1 U18625 ( .A1(n28461), .A2(\xmem_data[20][6] ), .B1(n28098), .B2(
        \xmem_data[21][6] ), .ZN(n14457) );
  AOI22_X1 U18626 ( .A1(n20734), .A2(\xmem_data[22][6] ), .B1(n31256), .B2(
        \xmem_data[23][6] ), .ZN(n14456) );
  NAND4_X1 U18627 ( .A1(n14459), .A2(n14458), .A3(n14457), .A4(n14456), .ZN(
        n14465) );
  AOI22_X1 U18628 ( .A1(n25684), .A2(\xmem_data[24][6] ), .B1(n31261), .B2(
        \xmem_data[25][6] ), .ZN(n14463) );
  AOI22_X1 U18629 ( .A1(n31263), .A2(\xmem_data[26][6] ), .B1(n31262), .B2(
        \xmem_data[27][6] ), .ZN(n14462) );
  AOI22_X1 U18630 ( .A1(n30864), .A2(\xmem_data[28][6] ), .B1(n27437), .B2(
        \xmem_data[29][6] ), .ZN(n14461) );
  AOI22_X1 U18631 ( .A1(n30962), .A2(\xmem_data[30][6] ), .B1(n3221), .B2(
        \xmem_data[31][6] ), .ZN(n14460) );
  NAND4_X1 U18632 ( .A1(n14463), .A2(n14462), .A3(n14461), .A4(n14460), .ZN(
        n14464) );
  OR4_X1 U18633 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14468) );
  AOI22_X1 U18634 ( .A1(n31340), .A2(n14469), .B1(n31284), .B2(n14468), .ZN(
        n14470) );
  XNOR2_X1 U18635 ( .A(n31663), .B(\fmem_data[12][5] ), .ZN(n33372) );
  OAI22_X1 U18636 ( .A1(n30472), .A2(n33973), .B1(n33372), .B2(n33975), .ZN(
        n23598) );
  XOR2_X1 U18637 ( .A(\fmem_data[16][3] ), .B(\fmem_data[16][2] ), .Z(n14472)
         );
  AOI22_X1 U18638 ( .A1(n24450), .A2(\xmem_data[10][7] ), .B1(n22701), .B2(
        \xmem_data[11][7] ), .ZN(n14476) );
  NAND2_X1 U18639 ( .A1(n30698), .A2(\xmem_data[8][7] ), .ZN(n14475) );
  NAND2_X1 U18640 ( .A1(n14476), .A2(n14475), .ZN(n14480) );
  NAND2_X1 U18641 ( .A1(n28772), .A2(\xmem_data[28][7] ), .ZN(n14478) );
  NAND2_X1 U18642 ( .A1(n24468), .A2(\xmem_data[29][7] ), .ZN(n14477) );
  NAND2_X1 U18643 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  NOR2_X1 U18644 ( .A1(n14480), .A2(n14479), .ZN(n14500) );
  AOI22_X1 U18645 ( .A1(n24458), .A2(\xmem_data[16][7] ), .B1(n24457), .B2(
        \xmem_data[17][7] ), .ZN(n14484) );
  AOI22_X1 U18646 ( .A1(n24133), .A2(\xmem_data[18][7] ), .B1(n24459), .B2(
        \xmem_data[19][7] ), .ZN(n14483) );
  AOI22_X1 U18647 ( .A1(n28232), .A2(\xmem_data[20][7] ), .B1(n24460), .B2(
        \xmem_data[21][7] ), .ZN(n14482) );
  AOI22_X1 U18648 ( .A1(n3178), .A2(\xmem_data[22][7] ), .B1(n20506), .B2(
        \xmem_data[23][7] ), .ZN(n14481) );
  AOI22_X1 U18649 ( .A1(n3222), .A2(\xmem_data[3][7] ), .B1(n29124), .B2(
        \xmem_data[30][7] ), .ZN(n14487) );
  AOI22_X1 U18650 ( .A1(n3334), .A2(\xmem_data[0][7] ), .B1(n24439), .B2(
        \xmem_data[1][7] ), .ZN(n14486) );
  AOI22_X1 U18651 ( .A1(n22708), .A2(\xmem_data[4][7] ), .B1(n25491), .B2(
        \xmem_data[5][7] ), .ZN(n14485) );
  AOI22_X1 U18652 ( .A1(n24467), .A2(\xmem_data[26][7] ), .B1(n31256), .B2(
        \xmem_data[27][7] ), .ZN(n14489) );
  AOI22_X1 U18653 ( .A1(n24438), .A2(\xmem_data[6][7] ), .B1(n30882), .B2(
        \xmem_data[7][7] ), .ZN(n14488) );
  NAND2_X1 U18654 ( .A1(n14489), .A2(n14488), .ZN(n14490) );
  NOR2_X1 U18655 ( .A1(n14491), .A2(n14490), .ZN(n14499) );
  AOI22_X1 U18656 ( .A1(n25710), .A2(\xmem_data[14][7] ), .B1(n23715), .B2(
        \xmem_data[15][7] ), .ZN(n14492) );
  INV_X1 U18657 ( .A(n14492), .ZN(n14496) );
  AOI22_X1 U18658 ( .A1(n27911), .A2(\xmem_data[12][7] ), .B1(n24448), .B2(
        \xmem_data[13][7] ), .ZN(n14494) );
  AOI22_X1 U18659 ( .A1(n3338), .A2(\xmem_data[24][7] ), .B1(n28098), .B2(
        \xmem_data[25][7] ), .ZN(n14493) );
  NAND2_X1 U18660 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  NOR2_X1 U18661 ( .A1(n14496), .A2(n14495), .ZN(n14498) );
  NAND2_X1 U18662 ( .A1(n29045), .A2(\xmem_data[9][7] ), .ZN(n14497) );
  NAND4_X1 U18663 ( .A1(n14501), .A2(n14500), .A3(n3522), .A4(n3917), .ZN(
        n14502) );
  NAND2_X1 U18664 ( .A1(n14502), .A2(n22180), .ZN(n14572) );
  AOI22_X1 U18665 ( .A1(n24556), .A2(\xmem_data[44][7] ), .B1(n24555), .B2(
        \xmem_data[45][7] ), .ZN(n14504) );
  AOI22_X1 U18666 ( .A1(n22717), .A2(\xmem_data[52][7] ), .B1(n14913), .B2(
        \xmem_data[53][7] ), .ZN(n14503) );
  NAND2_X1 U18667 ( .A1(n14504), .A2(n14503), .ZN(n14510) );
  AOI22_X1 U18668 ( .A1(n27913), .A2(\xmem_data[46][7] ), .B1(n24597), .B2(
        \xmem_data[47][7] ), .ZN(n14505) );
  INV_X1 U18669 ( .A(n14505), .ZN(n14509) );
  AOI22_X1 U18670 ( .A1(n24547), .A2(\xmem_data[50][7] ), .B1(n24546), .B2(
        \xmem_data[51][7] ), .ZN(n14507) );
  AOI22_X1 U18671 ( .A1(n3280), .A2(\xmem_data[40][7] ), .B1(n24553), .B2(
        \xmem_data[41][7] ), .ZN(n14506) );
  NAND2_X1 U18672 ( .A1(n14507), .A2(n14506), .ZN(n14508) );
  AOI22_X1 U18673 ( .A1(n16980), .A2(\xmem_data[32][7] ), .B1(n31347), .B2(
        \xmem_data[33][7] ), .ZN(n14514) );
  AOI22_X1 U18674 ( .A1(n24562), .A2(\xmem_data[34][7] ), .B1(n3219), .B2(
        \xmem_data[35][7] ), .ZN(n14513) );
  AOI22_X1 U18675 ( .A1(n24563), .A2(\xmem_data[36][7] ), .B1(n24695), .B2(
        \xmem_data[37][7] ), .ZN(n14512) );
  AOI22_X1 U18676 ( .A1(n24565), .A2(\xmem_data[38][7] ), .B1(n24564), .B2(
        \xmem_data[39][7] ), .ZN(n14511) );
  NAND4_X1 U18677 ( .A1(n14514), .A2(n14513), .A3(n14512), .A4(n14511), .ZN(
        n14525) );
  AOI22_X1 U18678 ( .A1(n24571), .A2(\xmem_data[56][7] ), .B1(n24570), .B2(
        \xmem_data[57][7] ), .ZN(n14519) );
  AOI22_X1 U18679 ( .A1(n24572), .A2(\xmem_data[58][7] ), .B1(n21057), .B2(
        \xmem_data[59][7] ), .ZN(n14518) );
  AOI22_X1 U18680 ( .A1(n17051), .A2(\xmem_data[60][7] ), .B1(n28035), .B2(
        \xmem_data[61][7] ), .ZN(n14517) );
  AND2_X1 U18681 ( .A1(n29057), .A2(\xmem_data[62][7] ), .ZN(n14515) );
  AOI21_X1 U18682 ( .B1(n24573), .B2(\xmem_data[63][7] ), .A(n14515), .ZN(
        n14516) );
  NAND4_X1 U18683 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14516), .ZN(
        n14524) );
  AOI22_X1 U18684 ( .A1(n24545), .A2(\xmem_data[48][7] ), .B1(n27516), .B2(
        \xmem_data[49][7] ), .ZN(n14522) );
  AOI22_X1 U18685 ( .A1(n24554), .A2(\xmem_data[42][7] ), .B1(n3357), .B2(
        \xmem_data[43][7] ), .ZN(n14521) );
  AOI22_X1 U18686 ( .A1(n3326), .A2(\xmem_data[54][7] ), .B1(n21051), .B2(
        \xmem_data[55][7] ), .ZN(n14520) );
  NAND3_X1 U18687 ( .A1(n14522), .A2(n14521), .A3(n14520), .ZN(n14523) );
  OR4_X1 U18688 ( .A1(n3971), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14526) );
  NAND2_X1 U18689 ( .A1(n14526), .A2(n24508), .ZN(n14571) );
  AOI22_X1 U18690 ( .A1(n3449), .A2(\xmem_data[96][7] ), .B1(n20711), .B2(
        \xmem_data[97][7] ), .ZN(n14530) );
  AOI22_X1 U18691 ( .A1(n24532), .A2(\xmem_data[98][7] ), .B1(n3217), .B2(
        \xmem_data[99][7] ), .ZN(n14529) );
  AOI22_X1 U18692 ( .A1(n24533), .A2(\xmem_data[100][7] ), .B1(n29028), .B2(
        \xmem_data[101][7] ), .ZN(n14528) );
  AOI22_X1 U18693 ( .A1(n24534), .A2(\xmem_data[102][7] ), .B1(n24633), .B2(
        \xmem_data[103][7] ), .ZN(n14527) );
  NAND4_X1 U18694 ( .A1(n14530), .A2(n14529), .A3(n14528), .A4(n14527), .ZN(
        n14546) );
  AOI22_X1 U18695 ( .A1(n24522), .A2(\xmem_data[120][7] ), .B1(n24521), .B2(
        \xmem_data[121][7] ), .ZN(n14534) );
  AOI22_X1 U18696 ( .A1(n3209), .A2(\xmem_data[122][7] ), .B1(n29136), .B2(
        \xmem_data[123][7] ), .ZN(n14533) );
  AOI22_X1 U18697 ( .A1(n21060), .A2(\xmem_data[124][7] ), .B1(n24524), .B2(
        \xmem_data[125][7] ), .ZN(n14532) );
  AOI22_X1 U18698 ( .A1(n24526), .A2(\xmem_data[126][7] ), .B1(n24525), .B2(
        \xmem_data[127][7] ), .ZN(n14531) );
  NAND4_X1 U18699 ( .A1(n14534), .A2(n14533), .A3(n14532), .A4(n14531), .ZN(
        n14545) );
  AOI22_X1 U18700 ( .A1(n30543), .A2(\xmem_data[112][7] ), .B1(n15000), .B2(
        \xmem_data[113][7] ), .ZN(n14538) );
  AOI22_X1 U18701 ( .A1(n24509), .A2(\xmem_data[114][7] ), .B1(n25398), .B2(
        \xmem_data[115][7] ), .ZN(n14537) );
  AOI22_X1 U18702 ( .A1(n30872), .A2(\xmem_data[116][7] ), .B1(n24510), .B2(
        \xmem_data[117][7] ), .ZN(n14536) );
  AOI22_X1 U18703 ( .A1(n24511), .A2(\xmem_data[118][7] ), .B1(n23778), .B2(
        \xmem_data[119][7] ), .ZN(n14535) );
  NAND4_X1 U18704 ( .A1(n14538), .A2(n14537), .A3(n14536), .A4(n14535), .ZN(
        n14544) );
  AOI22_X1 U18705 ( .A1(n25732), .A2(\xmem_data[104][7] ), .B1(n25514), .B2(
        \xmem_data[105][7] ), .ZN(n14542) );
  AOI22_X1 U18706 ( .A1(n25422), .A2(\xmem_data[106][7] ), .B1(n29307), .B2(
        \xmem_data[107][7] ), .ZN(n14541) );
  AOI22_X1 U18707 ( .A1(n23762), .A2(\xmem_data[108][7] ), .B1(n24516), .B2(
        \xmem_data[109][7] ), .ZN(n14540) );
  AOI22_X1 U18708 ( .A1(n3175), .A2(\xmem_data[110][7] ), .B1(n29309), .B2(
        \xmem_data[111][7] ), .ZN(n14539) );
  NAND4_X1 U18709 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        n14543) );
  OR4_X1 U18710 ( .A1(n14546), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        n14547) );
  NAND2_X1 U18711 ( .A1(n14547), .A2(n24542), .ZN(n14570) );
  AOI22_X1 U18712 ( .A1(n3413), .A2(\xmem_data[64][7] ), .B1(n28501), .B2(
        \xmem_data[65][7] ), .ZN(n14551) );
  AOI22_X1 U18713 ( .A1(n24562), .A2(\xmem_data[66][7] ), .B1(n3220), .B2(
        \xmem_data[67][7] ), .ZN(n14550) );
  AOI22_X1 U18714 ( .A1(n24563), .A2(\xmem_data[68][7] ), .B1(n20787), .B2(
        \xmem_data[69][7] ), .ZN(n14549) );
  AOI22_X1 U18715 ( .A1(n24565), .A2(\xmem_data[70][7] ), .B1(n24564), .B2(
        \xmem_data[71][7] ), .ZN(n14548) );
  NAND4_X1 U18716 ( .A1(n14551), .A2(n14550), .A3(n14549), .A4(n14548), .ZN(
        n14567) );
  AOI22_X1 U18717 ( .A1(n24571), .A2(\xmem_data[88][7] ), .B1(n24570), .B2(
        \xmem_data[89][7] ), .ZN(n14555) );
  AOI22_X1 U18718 ( .A1(n24572), .A2(\xmem_data[90][7] ), .B1(n29247), .B2(
        \xmem_data[91][7] ), .ZN(n14554) );
  AOI22_X1 U18719 ( .A1(n25628), .A2(\xmem_data[92][7] ), .B1(n25528), .B2(
        \xmem_data[93][7] ), .ZN(n14553) );
  AOI22_X1 U18720 ( .A1(n20710), .A2(\xmem_data[94][7] ), .B1(n24573), .B2(
        \xmem_data[95][7] ), .ZN(n14552) );
  NAND4_X1 U18721 ( .A1(n14555), .A2(n14554), .A3(n14553), .A4(n14552), .ZN(
        n14566) );
  AOI22_X1 U18722 ( .A1(n24545), .A2(\xmem_data[80][7] ), .B1(n27516), .B2(
        \xmem_data[81][7] ), .ZN(n14559) );
  AOI22_X1 U18723 ( .A1(n24547), .A2(\xmem_data[82][7] ), .B1(n24546), .B2(
        \xmem_data[83][7] ), .ZN(n14558) );
  AOI22_X1 U18724 ( .A1(n27825), .A2(\xmem_data[84][7] ), .B1(n30871), .B2(
        \xmem_data[85][7] ), .ZN(n14557) );
  AOI22_X1 U18725 ( .A1(n24190), .A2(\xmem_data[86][7] ), .B1(n25679), .B2(
        \xmem_data[87][7] ), .ZN(n14556) );
  NAND4_X1 U18726 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14556), .ZN(
        n14565) );
  AOI22_X1 U18727 ( .A1(n30295), .A2(\xmem_data[72][7] ), .B1(n24553), .B2(
        \xmem_data[73][7] ), .ZN(n14563) );
  AOI22_X1 U18728 ( .A1(n24554), .A2(\xmem_data[74][7] ), .B1(n29180), .B2(
        \xmem_data[75][7] ), .ZN(n14562) );
  AOI22_X1 U18729 ( .A1(n24556), .A2(\xmem_data[76][7] ), .B1(n24555), .B2(
        \xmem_data[77][7] ), .ZN(n14561) );
  AOI22_X1 U18730 ( .A1(n28334), .A2(\xmem_data[78][7] ), .B1(n25382), .B2(
        \xmem_data[79][7] ), .ZN(n14560) );
  NAND4_X1 U18731 ( .A1(n14563), .A2(n14562), .A3(n14561), .A4(n14560), .ZN(
        n14564) );
  OR4_X1 U18732 ( .A1(n14567), .A2(n14566), .A3(n14565), .A4(n14564), .ZN(
        n14568) );
  NAND2_X1 U18733 ( .A1(n14568), .A2(n24581), .ZN(n14569) );
  XNOR2_X1 U18734 ( .A(n35397), .B(\fmem_data[16][3] ), .ZN(n30380) );
  AOI21_X1 U18735 ( .B1(n34501), .B2(n34499), .A(n30380), .ZN(n14573) );
  INV_X1 U18736 ( .A(n14573), .ZN(n34871) );
  AOI22_X1 U18737 ( .A1(n23779), .A2(\xmem_data[26][5] ), .B1(n30525), .B2(
        \xmem_data[27][5] ), .ZN(n14574) );
  INV_X1 U18738 ( .A(n14574), .ZN(n14576) );
  AND2_X1 U18739 ( .A1(n30496), .A2(\xmem_data[28][5] ), .ZN(n14575) );
  NOR2_X1 U18740 ( .A1(n14576), .A2(n14575), .ZN(n14580) );
  AOI22_X1 U18741 ( .A1(n25716), .A2(\xmem_data[24][5] ), .B1(n30645), .B2(
        \xmem_data[25][5] ), .ZN(n14579) );
  AOI22_X1 U18742 ( .A1(n30498), .A2(\xmem_data[30][5] ), .B1(n25358), .B2(
        \xmem_data[31][5] ), .ZN(n14578) );
  NAND2_X1 U18743 ( .A1(n20708), .A2(\xmem_data[29][5] ), .ZN(n14577) );
  NAND4_X1 U18744 ( .A1(n14580), .A2(n14579), .A3(n14578), .A4(n14577), .ZN(
        n14594) );
  AOI22_X1 U18745 ( .A1(n25481), .A2(\xmem_data[12][5] ), .B1(n28743), .B2(
        \xmem_data[13][5] ), .ZN(n14587) );
  AOI22_X1 U18746 ( .A1(n25486), .A2(\xmem_data[8][5] ), .B1(n22668), .B2(
        \xmem_data[9][5] ), .ZN(n14581) );
  INV_X1 U18747 ( .A(n14581), .ZN(n14585) );
  AOI22_X1 U18748 ( .A1(n20775), .A2(\xmem_data[14][5] ), .B1(n13436), .B2(
        \xmem_data[15][5] ), .ZN(n14583) );
  NAND2_X1 U18749 ( .A1(n25422), .A2(\xmem_data[11][5] ), .ZN(n14582) );
  NAND2_X1 U18750 ( .A1(n14583), .A2(n14582), .ZN(n14584) );
  NOR2_X1 U18751 ( .A1(n14585), .A2(n14584), .ZN(n14586) );
  NAND2_X1 U18752 ( .A1(n14587), .A2(n14586), .ZN(n14593) );
  AOI22_X1 U18753 ( .A1(n25572), .A2(\xmem_data[16][5] ), .B1(n25672), .B2(
        \xmem_data[17][5] ), .ZN(n14591) );
  AOI22_X1 U18754 ( .A1(n3208), .A2(\xmem_data[18][5] ), .B1(n28096), .B2(
        \xmem_data[19][5] ), .ZN(n14590) );
  AOI22_X1 U18755 ( .A1(n28427), .A2(\xmem_data[20][5] ), .B1(n17044), .B2(
        \xmem_data[21][5] ), .ZN(n14589) );
  AOI22_X1 U18756 ( .A1(n30545), .A2(\xmem_data[22][5] ), .B1(n24511), .B2(
        \xmem_data[23][5] ), .ZN(n14588) );
  NAND4_X1 U18757 ( .A1(n14591), .A2(n14590), .A3(n14589), .A4(n14588), .ZN(
        n14592) );
  OR3_X1 U18758 ( .A1(n14594), .A2(n14593), .A3(n14592), .ZN(n14600) );
  AOI22_X1 U18759 ( .A1(n25485), .A2(\xmem_data[2][5] ), .B1(n28355), .B2(
        \xmem_data[3][5] ), .ZN(n14598) );
  AOI22_X1 U18760 ( .A1(n21309), .A2(\xmem_data[0][5] ), .B1(n28718), .B2(
        \xmem_data[1][5] ), .ZN(n14597) );
  AOI22_X1 U18761 ( .A1(n3221), .A2(\xmem_data[4][5] ), .B1(n27708), .B2(
        \xmem_data[5][5] ), .ZN(n14596) );
  AOI22_X1 U18762 ( .A1(n25491), .A2(\xmem_data[6][5] ), .B1(n25490), .B2(
        \xmem_data[7][5] ), .ZN(n14595) );
  NAND4_X1 U18763 ( .A1(n14598), .A2(n14597), .A3(n14596), .A4(n14595), .ZN(
        n14599) );
  NOR2_X1 U18764 ( .A1(n14600), .A2(n14599), .ZN(n14602) );
  NAND2_X1 U18765 ( .A1(n25492), .A2(\xmem_data[10][5] ), .ZN(n14601) );
  AOI21_X1 U18766 ( .B1(n14602), .B2(n14601), .A(n25505), .ZN(n14603) );
  INV_X1 U18767 ( .A(n14603), .ZN(n14669) );
  AOI22_X1 U18768 ( .A1(n25561), .A2(\xmem_data[96][5] ), .B1(n16980), .B2(
        \xmem_data[97][5] ), .ZN(n14607) );
  AOI22_X1 U18769 ( .A1(n27501), .A2(\xmem_data[98][5] ), .B1(n25508), .B2(
        \xmem_data[99][5] ), .ZN(n14606) );
  AOI22_X1 U18770 ( .A1(n3217), .A2(\xmem_data[100][5] ), .B1(n24632), .B2(
        \xmem_data[101][5] ), .ZN(n14605) );
  AOI22_X1 U18771 ( .A1(n25509), .A2(\xmem_data[102][5] ), .B1(n23741), .B2(
        \xmem_data[103][5] ), .ZN(n14604) );
  NAND4_X1 U18772 ( .A1(n14607), .A2(n14606), .A3(n14605), .A4(n14604), .ZN(
        n14623) );
  AOI22_X1 U18773 ( .A1(n28509), .A2(\xmem_data[104][5] ), .B1(n27905), .B2(
        \xmem_data[105][5] ), .ZN(n14611) );
  AOI22_X1 U18774 ( .A1(n25514), .A2(\xmem_data[106][5] ), .B1(n25422), .B2(
        \xmem_data[107][5] ), .ZN(n14610) );
  AOI22_X1 U18775 ( .A1(n22739), .A2(\xmem_data[108][5] ), .B1(n31327), .B2(
        \xmem_data[109][5] ), .ZN(n14609) );
  AOI22_X1 U18776 ( .A1(n27535), .A2(\xmem_data[110][5] ), .B1(n29272), .B2(
        \xmem_data[111][5] ), .ZN(n14608) );
  NAND4_X1 U18777 ( .A1(n14611), .A2(n14610), .A3(n14609), .A4(n14608), .ZN(
        n14622) );
  AOI22_X1 U18778 ( .A1(n25572), .A2(\xmem_data[112][5] ), .B1(n25519), .B2(
        \xmem_data[113][5] ), .ZN(n14615) );
  AOI22_X1 U18779 ( .A1(n27864), .A2(\xmem_data[114][5] ), .B1(n24509), .B2(
        \xmem_data[115][5] ), .ZN(n14614) );
  AOI22_X1 U18780 ( .A1(n25520), .A2(\xmem_data[116][5] ), .B1(n30872), .B2(
        \xmem_data[117][5] ), .ZN(n14613) );
  AOI22_X1 U18781 ( .A1(n27460), .A2(\xmem_data[118][5] ), .B1(n25521), .B2(
        \xmem_data[119][5] ), .ZN(n14612) );
  NAND4_X1 U18782 ( .A1(n14615), .A2(n14614), .A3(n14613), .A4(n14612), .ZN(
        n14621) );
  AOI22_X1 U18783 ( .A1(n24117), .A2(\xmem_data[120][5] ), .B1(n29324), .B2(
        \xmem_data[121][5] ), .ZN(n14619) );
  AOI22_X1 U18784 ( .A1(n14975), .A2(\xmem_data[122][5] ), .B1(n25526), .B2(
        \xmem_data[123][5] ), .ZN(n14618) );
  AOI22_X1 U18785 ( .A1(n25527), .A2(\xmem_data[124][5] ), .B1(n17051), .B2(
        \xmem_data[125][5] ), .ZN(n14617) );
  AOI22_X1 U18786 ( .A1(n25528), .A2(\xmem_data[126][5] ), .B1(n25724), .B2(
        \xmem_data[127][5] ), .ZN(n14616) );
  NAND4_X1 U18787 ( .A1(n14619), .A2(n14618), .A3(n14617), .A4(n14616), .ZN(
        n14620) );
  OR4_X1 U18788 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        n14645) );
  AOI22_X1 U18789 ( .A1(n25561), .A2(\xmem_data[64][5] ), .B1(n3305), .B2(
        \xmem_data[65][5] ), .ZN(n14627) );
  AOI22_X1 U18790 ( .A1(n14983), .A2(\xmem_data[66][5] ), .B1(n24562), .B2(
        \xmem_data[67][5] ), .ZN(n14626) );
  AOI22_X1 U18791 ( .A1(n3221), .A2(\xmem_data[68][5] ), .B1(n25693), .B2(
        \xmem_data[69][5] ), .ZN(n14625) );
  AOI22_X1 U18792 ( .A1(n25562), .A2(\xmem_data[70][5] ), .B1(n3341), .B2(
        \xmem_data[71][5] ), .ZN(n14624) );
  NAND4_X1 U18793 ( .A1(n14627), .A2(n14626), .A3(n14625), .A4(n14624), .ZN(
        n14643) );
  AOI22_X1 U18794 ( .A1(n25616), .A2(\xmem_data[72][5] ), .B1(n29350), .B2(
        \xmem_data[73][5] ), .ZN(n14631) );
  AOI22_X1 U18795 ( .A1(n24553), .A2(\xmem_data[74][5] ), .B1(n27447), .B2(
        \xmem_data[75][5] ), .ZN(n14630) );
  AOI22_X1 U18796 ( .A1(n28373), .A2(\xmem_data[76][5] ), .B1(n27453), .B2(
        \xmem_data[77][5] ), .ZN(n14629) );
  AOI22_X1 U18797 ( .A1(n27452), .A2(\xmem_data[78][5] ), .B1(n25567), .B2(
        \xmem_data[79][5] ), .ZN(n14628) );
  NAND4_X1 U18798 ( .A1(n14631), .A2(n14630), .A3(n14629), .A4(n14628), .ZN(
        n14642) );
  AOI22_X1 U18799 ( .A1(n24597), .A2(\xmem_data[80][5] ), .B1(n21048), .B2(
        \xmem_data[81][5] ), .ZN(n14635) );
  AOI22_X1 U18800 ( .A1(n25574), .A2(\xmem_data[82][5] ), .B1(n25573), .B2(
        \xmem_data[83][5] ), .ZN(n14634) );
  AOI22_X1 U18801 ( .A1(n25398), .A2(\xmem_data[84][5] ), .B1(n30617), .B2(
        \xmem_data[85][5] ), .ZN(n14633) );
  AOI22_X1 U18802 ( .A1(n25576), .A2(\xmem_data[86][5] ), .B1(n25575), .B2(
        \xmem_data[87][5] ), .ZN(n14632) );
  NAND4_X1 U18803 ( .A1(n14635), .A2(n14634), .A3(n14633), .A4(n14632), .ZN(
        n14641) );
  AOI22_X1 U18804 ( .A1(n25581), .A2(\xmem_data[88][5] ), .B1(n24623), .B2(
        \xmem_data[89][5] ), .ZN(n14639) );
  AOI22_X1 U18805 ( .A1(n25583), .A2(\xmem_data[90][5] ), .B1(n25582), .B2(
        \xmem_data[91][5] ), .ZN(n14638) );
  AOI22_X1 U18806 ( .A1(n28468), .A2(\xmem_data[92][5] ), .B1(n25584), .B2(
        \xmem_data[93][5] ), .ZN(n14637) );
  AOI22_X1 U18807 ( .A1(n20769), .A2(\xmem_data[94][5] ), .B1(n17030), .B2(
        \xmem_data[95][5] ), .ZN(n14636) );
  NAND4_X1 U18808 ( .A1(n14639), .A2(n14638), .A3(n14637), .A4(n14636), .ZN(
        n14640) );
  OR4_X1 U18809 ( .A1(n14643), .A2(n14642), .A3(n14641), .A4(n14640), .ZN(
        n14644) );
  AOI22_X1 U18810 ( .A1(n25560), .A2(n14645), .B1(n25558), .B2(n14644), .ZN(
        n14668) );
  AOI22_X1 U18811 ( .A1(n25561), .A2(\xmem_data[32][5] ), .B1(n3153), .B2(
        \xmem_data[33][5] ), .ZN(n14649) );
  AOI22_X1 U18812 ( .A1(n23731), .A2(\xmem_data[34][5] ), .B1(n28318), .B2(
        \xmem_data[35][5] ), .ZN(n14648) );
  AOI22_X1 U18813 ( .A1(n3219), .A2(\xmem_data[36][5] ), .B1(n30593), .B2(
        \xmem_data[37][5] ), .ZN(n14647) );
  AOI22_X1 U18814 ( .A1(n25562), .A2(\xmem_data[38][5] ), .B1(n3342), .B2(
        \xmem_data[39][5] ), .ZN(n14646) );
  NAND4_X1 U18815 ( .A1(n14649), .A2(n14648), .A3(n14647), .A4(n14646), .ZN(
        n14665) );
  AOI22_X1 U18816 ( .A1(n23811), .A2(\xmem_data[40][5] ), .B1(n3131), .B2(
        \xmem_data[41][5] ), .ZN(n14653) );
  AOI22_X1 U18817 ( .A1(n3231), .A2(\xmem_data[42][5] ), .B1(n28050), .B2(
        \xmem_data[43][5] ), .ZN(n14652) );
  AOI22_X1 U18818 ( .A1(n29180), .A2(\xmem_data[44][5] ), .B1(n28346), .B2(
        \xmem_data[45][5] ), .ZN(n14651) );
  AOI22_X1 U18819 ( .A1(n24516), .A2(\xmem_data[46][5] ), .B1(n25567), .B2(
        \xmem_data[47][5] ), .ZN(n14650) );
  NAND4_X1 U18820 ( .A1(n14653), .A2(n14652), .A3(n14651), .A4(n14650), .ZN(
        n14664) );
  AOI22_X1 U18821 ( .A1(n27536), .A2(\xmem_data[48][5] ), .B1(n21048), .B2(
        \xmem_data[49][5] ), .ZN(n14657) );
  AOI22_X1 U18822 ( .A1(n25574), .A2(\xmem_data[50][5] ), .B1(n25573), .B2(
        \xmem_data[51][5] ), .ZN(n14656) );
  AOI22_X1 U18823 ( .A1(n16989), .A2(\xmem_data[52][5] ), .B1(n29410), .B2(
        \xmem_data[53][5] ), .ZN(n14655) );
  AOI22_X1 U18824 ( .A1(n25576), .A2(\xmem_data[54][5] ), .B1(n25575), .B2(
        \xmem_data[55][5] ), .ZN(n14654) );
  NAND4_X1 U18825 ( .A1(n14657), .A2(n14656), .A3(n14655), .A4(n14654), .ZN(
        n14663) );
  AOI22_X1 U18826 ( .A1(n20816), .A2(\xmem_data[56][5] ), .B1(n24571), .B2(
        \xmem_data[57][5] ), .ZN(n14661) );
  AOI22_X1 U18827 ( .A1(n25583), .A2(\xmem_data[58][5] ), .B1(n25582), .B2(
        \xmem_data[59][5] ), .ZN(n14660) );
  AOI22_X1 U18828 ( .A1(n27463), .A2(\xmem_data[60][5] ), .B1(n25584), .B2(
        \xmem_data[61][5] ), .ZN(n14659) );
  AOI22_X1 U18829 ( .A1(n31261), .A2(\xmem_data[62][5] ), .B1(n27959), .B2(
        \xmem_data[63][5] ), .ZN(n14658) );
  NAND4_X1 U18830 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        n14662) );
  OR4_X1 U18831 ( .A1(n14665), .A2(n14664), .A3(n14663), .A4(n14662), .ZN(
        n14666) );
  NAND2_X1 U18832 ( .A1(n14666), .A2(n25593), .ZN(n14667) );
  AOI22_X1 U18833 ( .A1(n20489), .A2(\xmem_data[96][6] ), .B1(n3142), .B2(
        \xmem_data[97][6] ), .ZN(n14674) );
  AOI22_X1 U18834 ( .A1(n24172), .A2(\xmem_data[98][6] ), .B1(n25508), .B2(
        \xmem_data[99][6] ), .ZN(n14673) );
  AOI22_X1 U18835 ( .A1(n3222), .A2(\xmem_data[100][6] ), .B1(n25731), .B2(
        \xmem_data[101][6] ), .ZN(n14672) );
  AOI22_X1 U18836 ( .A1(n25509), .A2(\xmem_data[102][6] ), .B1(n20994), .B2(
        \xmem_data[103][6] ), .ZN(n14671) );
  NAND4_X1 U18837 ( .A1(n14674), .A2(n14673), .A3(n14672), .A4(n14671), .ZN(
        n14690) );
  AOI22_X1 U18838 ( .A1(n28509), .A2(\xmem_data[104][6] ), .B1(n30710), .B2(
        \xmem_data[105][6] ), .ZN(n14678) );
  AOI22_X1 U18839 ( .A1(n25514), .A2(\xmem_data[106][6] ), .B1(n16974), .B2(
        \xmem_data[107][6] ), .ZN(n14677) );
  AOI22_X1 U18840 ( .A1(n22701), .A2(\xmem_data[108][6] ), .B1(n25457), .B2(
        \xmem_data[109][6] ), .ZN(n14676) );
  AOI22_X1 U18841 ( .A1(n24516), .A2(\xmem_data[110][6] ), .B1(n28298), .B2(
        \xmem_data[111][6] ), .ZN(n14675) );
  NAND4_X1 U18842 ( .A1(n14678), .A2(n14677), .A3(n14676), .A4(n14675), .ZN(
        n14689) );
  AOI22_X1 U18843 ( .A1(n25572), .A2(\xmem_data[112][6] ), .B1(n25519), .B2(
        \xmem_data[113][6] ), .ZN(n14682) );
  AOI22_X1 U18844 ( .A1(n3213), .A2(\xmem_data[114][6] ), .B1(n17020), .B2(
        \xmem_data[115][6] ), .ZN(n14681) );
  AOI22_X1 U18845 ( .A1(n25520), .A2(\xmem_data[116][6] ), .B1(n29239), .B2(
        \xmem_data[117][6] ), .ZN(n14680) );
  AOI22_X1 U18846 ( .A1(n29101), .A2(\xmem_data[118][6] ), .B1(n25521), .B2(
        \xmem_data[119][6] ), .ZN(n14679) );
  NAND4_X1 U18847 ( .A1(n14682), .A2(n14681), .A3(n14680), .A4(n14679), .ZN(
        n14688) );
  AOI22_X1 U18848 ( .A1(n24222), .A2(\xmem_data[120][6] ), .B1(n3328), .B2(
        \xmem_data[121][6] ), .ZN(n14686) );
  AOI22_X1 U18849 ( .A1(n20507), .A2(\xmem_data[122][6] ), .B1(n25526), .B2(
        \xmem_data[123][6] ), .ZN(n14685) );
  AOI22_X1 U18850 ( .A1(n25527), .A2(\xmem_data[124][6] ), .B1(n25684), .B2(
        \xmem_data[125][6] ), .ZN(n14684) );
  AOI22_X1 U18851 ( .A1(n25528), .A2(\xmem_data[126][6] ), .B1(n24526), .B2(
        \xmem_data[127][6] ), .ZN(n14683) );
  NAND4_X1 U18852 ( .A1(n14686), .A2(n14685), .A3(n14684), .A4(n14683), .ZN(
        n14687) );
  OR4_X1 U18853 ( .A1(n14690), .A2(n14689), .A3(n14688), .A4(n14687), .ZN(
        n14713) );
  AOI22_X1 U18854 ( .A1(n25561), .A2(\xmem_data[64][6] ), .B1(n3229), .B2(
        \xmem_data[65][6] ), .ZN(n14694) );
  AOI22_X1 U18855 ( .A1(n29286), .A2(\xmem_data[66][6] ), .B1(n28082), .B2(
        \xmem_data[67][6] ), .ZN(n14693) );
  AOI22_X1 U18856 ( .A1(n3222), .A2(\xmem_data[68][6] ), .B1(n29256), .B2(
        \xmem_data[69][6] ), .ZN(n14692) );
  AOI22_X1 U18857 ( .A1(n25562), .A2(\xmem_data[70][6] ), .B1(n3340), .B2(
        \xmem_data[71][6] ), .ZN(n14691) );
  NAND4_X1 U18858 ( .A1(n14694), .A2(n14693), .A3(n14692), .A4(n14691), .ZN(
        n14711) );
  AOI22_X1 U18859 ( .A1(n22669), .A2(\xmem_data[72][6] ), .B1(n28952), .B2(
        \xmem_data[73][6] ), .ZN(n14698) );
  AOI22_X1 U18860 ( .A1(n31252), .A2(\xmem_data[74][6] ), .B1(n23813), .B2(
        \xmem_data[75][6] ), .ZN(n14697) );
  AOI22_X1 U18861 ( .A1(n14996), .A2(\xmem_data[76][6] ), .B1(n24640), .B2(
        \xmem_data[77][6] ), .ZN(n14696) );
  AOI22_X1 U18862 ( .A1(n24212), .A2(\xmem_data[78][6] ), .B1(n25567), .B2(
        \xmem_data[79][6] ), .ZN(n14695) );
  NAND4_X1 U18863 ( .A1(n14698), .A2(n14697), .A3(n14696), .A4(n14695), .ZN(
        n14710) );
  AOI22_X1 U18864 ( .A1(n25572), .A2(\xmem_data[80][6] ), .B1(n28336), .B2(
        \xmem_data[81][6] ), .ZN(n14702) );
  AOI22_X1 U18865 ( .A1(n25574), .A2(\xmem_data[82][6] ), .B1(n25573), .B2(
        \xmem_data[83][6] ), .ZN(n14701) );
  AOI22_X1 U18866 ( .A1(n25398), .A2(\xmem_data[84][6] ), .B1(n21050), .B2(
        \xmem_data[85][6] ), .ZN(n14700) );
  AOI22_X1 U18867 ( .A1(n25576), .A2(\xmem_data[86][6] ), .B1(n25575), .B2(
        \xmem_data[87][6] ), .ZN(n14699) );
  NAND4_X1 U18868 ( .A1(n14702), .A2(n14701), .A3(n14700), .A4(n14699), .ZN(
        n14709) );
  AOI22_X1 U18869 ( .A1(n25679), .A2(\xmem_data[88][6] ), .B1(n20950), .B2(
        \xmem_data[89][6] ), .ZN(n14707) );
  AOI22_X1 U18870 ( .A1(n25583), .A2(\xmem_data[90][6] ), .B1(n25582), .B2(
        \xmem_data[91][6] ), .ZN(n14706) );
  AND2_X1 U18871 ( .A1(n23725), .A2(\xmem_data[92][6] ), .ZN(n14703) );
  AOI21_X1 U18872 ( .B1(n25584), .B2(\xmem_data[93][6] ), .A(n14703), .ZN(
        n14705) );
  AOI22_X1 U18873 ( .A1(n30900), .A2(\xmem_data[94][6] ), .B1(n25686), .B2(
        \xmem_data[95][6] ), .ZN(n14704) );
  NAND4_X1 U18874 ( .A1(n14707), .A2(n14706), .A3(n14705), .A4(n14704), .ZN(
        n14708) );
  OR4_X1 U18875 ( .A1(n14711), .A2(n14710), .A3(n14709), .A4(n14708), .ZN(
        n14712) );
  AOI22_X1 U18876 ( .A1(n25560), .A2(n14713), .B1(n25558), .B2(n14712), .ZN(
        n14768) );
  AOI22_X1 U18877 ( .A1(n25561), .A2(\xmem_data[32][6] ), .B1(n25725), .B2(
        \xmem_data[33][6] ), .ZN(n14717) );
  AOI22_X1 U18878 ( .A1(n3247), .A2(\xmem_data[34][6] ), .B1(n20991), .B2(
        \xmem_data[35][6] ), .ZN(n14716) );
  AOI22_X1 U18879 ( .A1(n3217), .A2(\xmem_data[36][6] ), .B1(n28367), .B2(
        \xmem_data[37][6] ), .ZN(n14715) );
  AOI22_X1 U18880 ( .A1(n25562), .A2(\xmem_data[38][6] ), .B1(n3341), .B2(
        \xmem_data[39][6] ), .ZN(n14714) );
  NAND4_X1 U18881 ( .A1(n14717), .A2(n14716), .A3(n14715), .A4(n14714), .ZN(
        n14733) );
  AOI22_X1 U18882 ( .A1(n17061), .A2(\xmem_data[40][6] ), .B1(n29706), .B2(
        \xmem_data[41][6] ), .ZN(n14721) );
  AOI22_X1 U18883 ( .A1(n28045), .A2(\xmem_data[42][6] ), .B1(n28050), .B2(
        \xmem_data[43][6] ), .ZN(n14720) );
  AOI22_X1 U18884 ( .A1(n14933), .A2(\xmem_data[44][6] ), .B1(n30943), .B2(
        \xmem_data[45][6] ), .ZN(n14719) );
  AOI22_X1 U18885 ( .A1(n24212), .A2(\xmem_data[46][6] ), .B1(n25567), .B2(
        \xmem_data[47][6] ), .ZN(n14718) );
  NAND4_X1 U18886 ( .A1(n14721), .A2(n14720), .A3(n14719), .A4(n14718), .ZN(
        n14732) );
  AOI22_X1 U18887 ( .A1(n28517), .A2(\xmem_data[48][6] ), .B1(n28053), .B2(
        \xmem_data[49][6] ), .ZN(n14725) );
  AOI22_X1 U18888 ( .A1(n25574), .A2(\xmem_data[50][6] ), .B1(n25573), .B2(
        \xmem_data[51][6] ), .ZN(n14724) );
  AOI22_X1 U18889 ( .A1(n29048), .A2(\xmem_data[52][6] ), .B1(n17021), .B2(
        \xmem_data[53][6] ), .ZN(n14723) );
  AOI22_X1 U18890 ( .A1(n25576), .A2(\xmem_data[54][6] ), .B1(n25575), .B2(
        \xmem_data[55][6] ), .ZN(n14722) );
  NAND4_X1 U18891 ( .A1(n14725), .A2(n14724), .A3(n14723), .A4(n14722), .ZN(
        n14731) );
  AOI22_X1 U18892 ( .A1(n28462), .A2(\xmem_data[56][6] ), .B1(n30269), .B2(
        \xmem_data[57][6] ), .ZN(n14729) );
  AOI22_X1 U18893 ( .A1(n25583), .A2(\xmem_data[58][6] ), .B1(n25582), .B2(
        \xmem_data[59][6] ), .ZN(n14728) );
  AOI22_X1 U18894 ( .A1(n28292), .A2(\xmem_data[60][6] ), .B1(n25584), .B2(
        \xmem_data[61][6] ), .ZN(n14727) );
  AOI22_X1 U18895 ( .A1(n16999), .A2(\xmem_data[62][6] ), .B1(n20827), .B2(
        \xmem_data[63][6] ), .ZN(n14726) );
  NAND4_X1 U18896 ( .A1(n14729), .A2(n14728), .A3(n14727), .A4(n14726), .ZN(
        n14730) );
  OR4_X1 U18897 ( .A1(n14733), .A2(n14732), .A3(n14731), .A4(n14730), .ZN(
        n14734) );
  AOI22_X1 U18898 ( .A1(n25481), .A2(\xmem_data[12][6] ), .B1(n29591), .B2(
        \xmem_data[13][6] ), .ZN(n14735) );
  INV_X1 U18899 ( .A(n14735), .ZN(n14744) );
  AOI22_X1 U18900 ( .A1(n3207), .A2(\xmem_data[18][6] ), .B1(n30949), .B2(
        \xmem_data[19][6] ), .ZN(n14738) );
  AOI22_X1 U18901 ( .A1(n21059), .A2(\xmem_data[30][6] ), .B1(n27500), .B2(
        \xmem_data[31][6] ), .ZN(n14737) );
  AOI22_X1 U18902 ( .A1(n29281), .A2(\xmem_data[24][6] ), .B1(n29573), .B2(
        \xmem_data[25][6] ), .ZN(n14736) );
  AND2_X1 U18903 ( .A1(n30496), .A2(\xmem_data[28][6] ), .ZN(n14739) );
  AOI21_X1 U18904 ( .B1(n27717), .B2(\xmem_data[29][6] ), .A(n14739), .ZN(
        n14741) );
  AOI22_X1 U18905 ( .A1(n25629), .A2(\xmem_data[0][6] ), .B1(n24630), .B2(
        \xmem_data[1][6] ), .ZN(n14740) );
  NAND2_X1 U18906 ( .A1(n14741), .A2(n14740), .ZN(n14742) );
  NOR3_X1 U18907 ( .A1(n14744), .A2(n14743), .A3(n14742), .ZN(n14764) );
  AOI22_X1 U18908 ( .A1(n25486), .A2(\xmem_data[8][6] ), .B1(n30698), .B2(
        \xmem_data[9][6] ), .ZN(n14747) );
  AOI22_X1 U18909 ( .A1(n23761), .A2(\xmem_data[14][6] ), .B1(n30514), .B2(
        \xmem_data[15][6] ), .ZN(n14746) );
  NAND2_X1 U18910 ( .A1(n20961), .A2(\xmem_data[11][6] ), .ZN(n14745) );
  NAND3_X1 U18911 ( .A1(n14747), .A2(n14746), .A3(n14745), .ZN(n14762) );
  AOI22_X1 U18912 ( .A1(n3218), .A2(\xmem_data[4][6] ), .B1(n29627), .B2(
        \xmem_data[5][6] ), .ZN(n14751) );
  AOI22_X1 U18913 ( .A1(n20505), .A2(\xmem_data[20][6] ), .B1(n28781), .B2(
        \xmem_data[21][6] ), .ZN(n14750) );
  AOI22_X1 U18914 ( .A1(n24521), .A2(\xmem_data[26][6] ), .B1(n24606), .B2(
        \xmem_data[27][6] ), .ZN(n14749) );
  NAND2_X1 U18915 ( .A1(n30906), .A2(\xmem_data[3][6] ), .ZN(n14748) );
  NAND4_X1 U18916 ( .A1(n14751), .A2(n14750), .A3(n14749), .A4(n14748), .ZN(
        n14761) );
  AOI22_X1 U18917 ( .A1(n30545), .A2(\xmem_data[22][6] ), .B1(n30849), .B2(
        \xmem_data[23][6] ), .ZN(n14759) );
  AOI22_X1 U18918 ( .A1(n25709), .A2(\xmem_data[16][6] ), .B1(n25607), .B2(
        \xmem_data[17][6] ), .ZN(n14758) );
  AOI22_X1 U18919 ( .A1(n25491), .A2(\xmem_data[6][6] ), .B1(n25490), .B2(
        \xmem_data[7][6] ), .ZN(n14752) );
  INV_X1 U18920 ( .A(n14752), .ZN(n14756) );
  NAND2_X1 U18921 ( .A1(n25492), .A2(\xmem_data[10][6] ), .ZN(n14754) );
  NAND2_X1 U18922 ( .A1(n25485), .A2(\xmem_data[2][6] ), .ZN(n14753) );
  NAND2_X1 U18923 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  NOR2_X1 U18924 ( .A1(n14756), .A2(n14755), .ZN(n14757) );
  NOR3_X1 U18925 ( .A1(n14762), .A2(n14761), .A3(n14760), .ZN(n14763) );
  AOI21_X1 U18926 ( .B1(n14764), .B2(n14763), .A(n25505), .ZN(n14765) );
  INV_X1 U18927 ( .A(n14765), .ZN(n14766) );
  XNOR2_X1 U18928 ( .A(n31705), .B(\fmem_data[17][5] ), .ZN(n33126) );
  OAI22_X1 U18929 ( .A1(n30473), .A2(n34043), .B1(n34045), .B2(n33126), .ZN(
        n34870) );
  XNOR2_X1 U18930 ( .A(n34871), .B(n34870), .ZN(n14874) );
  XNOR2_X1 U18931 ( .A(n31247), .B(\fmem_data[11][7] ), .ZN(n23925) );
  AOI22_X1 U18932 ( .A1(n28765), .A2(\xmem_data[120][3] ), .B1(n3124), .B2(
        \xmem_data[121][3] ), .ZN(n14773) );
  AOI22_X1 U18933 ( .A1(n28719), .A2(\xmem_data[122][3] ), .B1(n28718), .B2(
        \xmem_data[123][3] ), .ZN(n14772) );
  AOI22_X1 U18934 ( .A1(n29788), .A2(\xmem_data[124][3] ), .B1(n29831), .B2(
        \xmem_data[125][3] ), .ZN(n14771) );
  AND2_X1 U18935 ( .A1(n28733), .A2(\xmem_data[127][3] ), .ZN(n14769) );
  AOI21_X1 U18936 ( .B1(n28700), .B2(\xmem_data[126][3] ), .A(n14769), .ZN(
        n14770) );
  NAND4_X1 U18937 ( .A1(n14773), .A2(n14772), .A3(n14771), .A4(n14770), .ZN(
        n14790) );
  AOI22_X1 U18938 ( .A1(n28740), .A2(\xmem_data[96][3] ), .B1(n30696), .B2(
        \xmem_data[97][3] ), .ZN(n14777) );
  AOI22_X1 U18939 ( .A1(n3244), .A2(\xmem_data[98][3] ), .B1(n3126), .B2(
        \xmem_data[99][3] ), .ZN(n14776) );
  AOI22_X1 U18940 ( .A1(n29801), .A2(\xmem_data[100][3] ), .B1(n28665), .B2(
        \xmem_data[101][3] ), .ZN(n14775) );
  AOI22_X1 U18941 ( .A1(n28744), .A2(\xmem_data[102][3] ), .B1(n28743), .B2(
        \xmem_data[103][3] ), .ZN(n14774) );
  NAND4_X1 U18942 ( .A1(n14777), .A2(n14776), .A3(n14775), .A4(n14774), .ZN(
        n14789) );
  AOI22_X1 U18943 ( .A1(n29363), .A2(\xmem_data[112][3] ), .B1(n29640), .B2(
        \xmem_data[113][3] ), .ZN(n14781) );
  AOI22_X1 U18944 ( .A1(n28720), .A2(\xmem_data[114][3] ), .B1(n29379), .B2(
        \xmem_data[115][3] ), .ZN(n14780) );
  AOI22_X1 U18945 ( .A1(n28725), .A2(\xmem_data[116][3] ), .B1(n28724), .B2(
        \xmem_data[117][3] ), .ZN(n14779) );
  AOI22_X1 U18946 ( .A1(n28727), .A2(\xmem_data[118][3] ), .B1(n25407), .B2(
        \xmem_data[119][3] ), .ZN(n14778) );
  NAND4_X1 U18947 ( .A1(n14781), .A2(n14780), .A3(n14779), .A4(n14778), .ZN(
        n14788) );
  AOI22_X1 U18948 ( .A1(n29769), .A2(\xmem_data[104][3] ), .B1(n30301), .B2(
        \xmem_data[105][3] ), .ZN(n14786) );
  AOI22_X1 U18949 ( .A1(n28753), .A2(\xmem_data[106][3] ), .B1(n29396), .B2(
        \xmem_data[107][3] ), .ZN(n14785) );
  AOI22_X1 U18950 ( .A1(n3162), .A2(\xmem_data[108][3] ), .B1(n3185), .B2(
        \xmem_data[109][3] ), .ZN(n14784) );
  AND2_X1 U18951 ( .A1(n28687), .A2(\xmem_data[111][3] ), .ZN(n14782) );
  AOI21_X1 U18952 ( .B1(n30070), .B2(\xmem_data[110][3] ), .A(n14782), .ZN(
        n14783) );
  NAND4_X1 U18953 ( .A1(n14786), .A2(n14785), .A3(n14784), .A4(n14783), .ZN(
        n14787) );
  NAND2_X1 U18954 ( .A1(n14791), .A2(n28762), .ZN(n14872) );
  NAND2_X1 U18955 ( .A1(n29790), .A2(\xmem_data[94][3] ), .ZN(n14793) );
  NAND2_X1 U18956 ( .A1(n28733), .A2(\xmem_data[95][3] ), .ZN(n14792) );
  NAND2_X1 U18957 ( .A1(n14793), .A2(n14792), .ZN(n14799) );
  AOI22_X1 U18958 ( .A1(n30766), .A2(\xmem_data[80][3] ), .B1(n30644), .B2(
        \xmem_data[81][3] ), .ZN(n14797) );
  AOI22_X1 U18959 ( .A1(n28720), .A2(\xmem_data[82][3] ), .B1(n3328), .B2(
        \xmem_data[83][3] ), .ZN(n14796) );
  AOI22_X1 U18960 ( .A1(n28725), .A2(\xmem_data[84][3] ), .B1(n28724), .B2(
        \xmem_data[85][3] ), .ZN(n14795) );
  AOI22_X1 U18961 ( .A1(n28727), .A2(\xmem_data[86][3] ), .B1(n31345), .B2(
        \xmem_data[87][3] ), .ZN(n14794) );
  NAND4_X1 U18962 ( .A1(n14797), .A2(n14796), .A3(n14795), .A4(n14794), .ZN(
        n14798) );
  NOR2_X1 U18963 ( .A1(n14799), .A2(n14798), .ZN(n14806) );
  AOI22_X1 U18964 ( .A1(n27741), .A2(\xmem_data[92][3] ), .B1(n27013), .B2(
        \xmem_data[93][3] ), .ZN(n14800) );
  INV_X1 U18965 ( .A(n14800), .ZN(n14804) );
  AOI22_X1 U18966 ( .A1(n28765), .A2(\xmem_data[88][3] ), .B1(n3124), .B2(
        \xmem_data[89][3] ), .ZN(n14802) );
  AOI22_X1 U18967 ( .A1(n28719), .A2(\xmem_data[90][3] ), .B1(n28718), .B2(
        \xmem_data[91][3] ), .ZN(n14801) );
  NAND2_X1 U18968 ( .A1(n14802), .A2(n14801), .ZN(n14803) );
  NOR2_X1 U18969 ( .A1(n14804), .A2(n14803), .ZN(n14805) );
  NAND2_X1 U18970 ( .A1(n14806), .A2(n14805), .ZN(n14822) );
  NAND2_X1 U18971 ( .A1(n29589), .A2(\xmem_data[69][3] ), .ZN(n14808) );
  NAND2_X1 U18972 ( .A1(n29590), .A2(\xmem_data[68][3] ), .ZN(n14807) );
  NAND2_X1 U18973 ( .A1(n14808), .A2(n14807), .ZN(n14815) );
  NAND2_X1 U18974 ( .A1(n28208), .A2(\xmem_data[65][3] ), .ZN(n14810) );
  NAND2_X1 U18975 ( .A1(n28740), .A2(\xmem_data[64][3] ), .ZN(n14809) );
  NAND2_X1 U18976 ( .A1(n14810), .A2(n14809), .ZN(n14814) );
  AOI22_X1 U18977 ( .A1(n3244), .A2(\xmem_data[66][3] ), .B1(n3126), .B2(
        \xmem_data[67][3] ), .ZN(n14812) );
  AOI22_X1 U18978 ( .A1(n28744), .A2(\xmem_data[70][3] ), .B1(n28743), .B2(
        \xmem_data[71][3] ), .ZN(n14811) );
  NAND2_X1 U18979 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  NOR3_X1 U18980 ( .A1(n14815), .A2(n14814), .A3(n14813), .ZN(n14820) );
  AOI22_X1 U18981 ( .A1(n28685), .A2(\xmem_data[72][3] ), .B1(n27753), .B2(
        \xmem_data[73][3] ), .ZN(n14819) );
  AOI22_X1 U18982 ( .A1(n28753), .A2(\xmem_data[74][3] ), .B1(n28516), .B2(
        \xmem_data[75][3] ), .ZN(n14818) );
  AOI22_X1 U18983 ( .A1(n3164), .A2(\xmem_data[76][3] ), .B1(n3188), .B2(
        \xmem_data[77][3] ), .ZN(n14817) );
  AOI22_X1 U18984 ( .A1(n30715), .A2(\xmem_data[78][3] ), .B1(n28754), .B2(
        \xmem_data[79][3] ), .ZN(n14816) );
  NAND2_X1 U18985 ( .A1(n14820), .A2(n3761), .ZN(n14821) );
  OAI21_X1 U18986 ( .B1(n14822), .B2(n14821), .A(n28662), .ZN(n14871) );
  AOI22_X1 U18987 ( .A1(n29647), .A2(\xmem_data[36][3] ), .B1(n29646), .B2(
        \xmem_data[37][3] ), .ZN(n14823) );
  INV_X1 U18988 ( .A(n14823), .ZN(n14830) );
  NAND2_X1 U18989 ( .A1(n28667), .A2(\xmem_data[33][3] ), .ZN(n14825) );
  NAND2_X1 U18990 ( .A1(n30280), .A2(\xmem_data[32][3] ), .ZN(n14824) );
  NAND2_X1 U18991 ( .A1(n14825), .A2(n14824), .ZN(n14829) );
  AOI22_X1 U18992 ( .A1(n28670), .A2(\xmem_data[34][3] ), .B1(n3140), .B2(
        \xmem_data[35][3] ), .ZN(n14827) );
  AOI22_X1 U18993 ( .A1(n28744), .A2(\xmem_data[38][3] ), .B1(n28671), .B2(
        \xmem_data[39][3] ), .ZN(n14826) );
  NAND2_X1 U18994 ( .A1(n14827), .A2(n14826), .ZN(n14828) );
  NOR3_X1 U18995 ( .A1(n14830), .A2(n14829), .A3(n14828), .ZN(n14846) );
  AOI22_X1 U18996 ( .A1(n29788), .A2(\xmem_data[60][3] ), .B1(n29672), .B2(
        \xmem_data[61][3] ), .ZN(n14831) );
  INV_X1 U18997 ( .A(n14831), .ZN(n14836) );
  AOI22_X1 U18998 ( .A1(n29628), .A2(\xmem_data[62][3] ), .B1(n30278), .B2(
        \xmem_data[63][3] ), .ZN(n14834) );
  AOI22_X1 U18999 ( .A1(n3227), .A2(\xmem_data[58][3] ), .B1(n28677), .B2(
        \xmem_data[59][3] ), .ZN(n14833) );
  AOI22_X1 U19000 ( .A1(n29829), .A2(\xmem_data[56][3] ), .B1(n27723), .B2(
        \xmem_data[57][3] ), .ZN(n14832) );
  NOR2_X1 U19001 ( .A1(n14836), .A2(n14835), .ZN(n14845) );
  AOI22_X1 U19002 ( .A1(n29769), .A2(\xmem_data[40][3] ), .B1(n28110), .B2(
        \xmem_data[41][3] ), .ZN(n14840) );
  AOI22_X1 U19003 ( .A1(n28686), .A2(\xmem_data[42][3] ), .B1(n3466), .B2(
        \xmem_data[43][3] ), .ZN(n14839) );
  AOI22_X1 U19004 ( .A1(n3168), .A2(\xmem_data[44][3] ), .B1(n3183), .B2(
        \xmem_data[45][3] ), .ZN(n14838) );
  AOI22_X1 U19005 ( .A1(n30062), .A2(\xmem_data[46][3] ), .B1(n28781), .B2(
        \xmem_data[47][3] ), .ZN(n14837) );
  AOI22_X1 U19006 ( .A1(n29722), .A2(\xmem_data[48][3] ), .B1(n29721), .B2(
        \xmem_data[49][3] ), .ZN(n14844) );
  AOI22_X1 U19007 ( .A1(n28702), .A2(\xmem_data[50][3] ), .B1(n28701), .B2(
        \xmem_data[51][3] ), .ZN(n14843) );
  AOI22_X1 U19008 ( .A1(n29724), .A2(\xmem_data[52][3] ), .B1(n28696), .B2(
        \xmem_data[53][3] ), .ZN(n14842) );
  AOI22_X1 U19009 ( .A1(n28681), .A2(\xmem_data[54][3] ), .B1(n28036), .B2(
        \xmem_data[55][3] ), .ZN(n14841) );
  NAND4_X1 U19010 ( .A1(n14846), .A2(n14845), .A3(n3795), .A4(n3517), .ZN(
        n14847) );
  NAND2_X1 U19011 ( .A1(n14847), .A2(n28713), .ZN(n14870) );
  AOI22_X1 U19012 ( .A1(n28787), .A2(\xmem_data[0][3] ), .B1(n29708), .B2(
        \xmem_data[1][3] ), .ZN(n14851) );
  AOI22_X1 U19013 ( .A1(n3244), .A2(\xmem_data[2][3] ), .B1(n3138), .B2(
        \xmem_data[3][3] ), .ZN(n14850) );
  AOI22_X1 U19014 ( .A1(n29705), .A2(\xmem_data[4][3] ), .B1(n30662), .B2(
        \xmem_data[5][3] ), .ZN(n14849) );
  AOI22_X1 U19015 ( .A1(n28788), .A2(\xmem_data[6][3] ), .B1(n30663), .B2(
        \xmem_data[7][3] ), .ZN(n14848) );
  AND4_X1 U19016 ( .A1(n14851), .A2(n14850), .A3(n14849), .A4(n14848), .ZN(
        n14867) );
  AOI22_X1 U19017 ( .A1(n30302), .A2(\xmem_data[8][3] ), .B1(n30193), .B2(
        \xmem_data[9][3] ), .ZN(n14855) );
  AOI22_X1 U19018 ( .A1(n28780), .A2(\xmem_data[10][3] ), .B1(n29237), .B2(
        \xmem_data[11][3] ), .ZN(n14854) );
  AOI22_X1 U19019 ( .A1(n3164), .A2(\xmem_data[12][3] ), .B1(n3187), .B2(
        \xmem_data[13][3] ), .ZN(n14853) );
  AOI22_X1 U19020 ( .A1(n30764), .A2(\xmem_data[14][3] ), .B1(n28687), .B2(
        \xmem_data[15][3] ), .ZN(n14852) );
  AND4_X1 U19021 ( .A1(n14855), .A2(n14854), .A3(n14853), .A4(n14852), .ZN(
        n14866) );
  AOI22_X1 U19022 ( .A1(n29488), .A2(\xmem_data[16][3] ), .B1(n29640), .B2(
        \xmem_data[17][3] ), .ZN(n14859) );
  AOI22_X1 U19023 ( .A1(n28702), .A2(\xmem_data[18][3] ), .B1(n29816), .B2(
        \xmem_data[19][3] ), .ZN(n14858) );
  AOI22_X1 U19024 ( .A1(n27716), .A2(\xmem_data[20][3] ), .B1(n27805), .B2(
        \xmem_data[21][3] ), .ZN(n14857) );
  AOI22_X1 U19025 ( .A1(n27806), .A2(\xmem_data[22][3] ), .B1(n28772), .B2(
        \xmem_data[23][3] ), .ZN(n14856) );
  AND4_X1 U19026 ( .A1(n14859), .A2(n14858), .A3(n14857), .A4(n14856), .ZN(
        n14865) );
  AOI22_X1 U19027 ( .A1(n28765), .A2(\xmem_data[24][3] ), .B1(n27723), .B2(
        \xmem_data[25][3] ), .ZN(n14863) );
  AOI22_X1 U19028 ( .A1(n3227), .A2(\xmem_data[26][3] ), .B1(n3153), .B2(
        \xmem_data[27][3] ), .ZN(n14862) );
  AOI22_X1 U19029 ( .A1(n29433), .A2(\xmem_data[28][3] ), .B1(n29432), .B2(
        \xmem_data[29][3] ), .ZN(n14861) );
  AOI22_X1 U19030 ( .A1(n29790), .A2(\xmem_data[30][3] ), .B1(n29832), .B2(
        \xmem_data[31][3] ), .ZN(n14860) );
  AND4_X1 U19031 ( .A1(n14863), .A2(n14862), .A3(n14861), .A4(n14860), .ZN(
        n14864) );
  NAND4_X1 U19032 ( .A1(n14867), .A2(n14866), .A3(n14865), .A4(n14864), .ZN(
        n14868) );
  NAND2_X1 U19033 ( .A1(n14868), .A2(n28794), .ZN(n14869) );
  NAND4_X2 U19034 ( .A1(n14872), .A2(n14871), .A3(n14870), .A4(n14869), .ZN(
        n32023) );
  XNOR2_X1 U19035 ( .A(n32023), .B(\fmem_data[11][7] ), .ZN(n24835) );
  XOR2_X1 U19036 ( .A(\fmem_data[11][6] ), .B(\fmem_data[11][7] ), .Z(n14873)
         );
  XNOR2_X1 U19037 ( .A(n14874), .B(n34869), .ZN(n18726) );
  AOI22_X1 U19038 ( .A1(n17003), .A2(\xmem_data[8][3] ), .B1(n30901), .B2(
        \xmem_data[9][3] ), .ZN(n14880) );
  AOI22_X1 U19039 ( .A1(n25388), .A2(\xmem_data[10][3] ), .B1(n28038), .B2(
        \xmem_data[11][3] ), .ZN(n14879) );
  AOI22_X1 U19040 ( .A1(n30908), .A2(\xmem_data[12][3] ), .B1(n29661), .B2(
        \xmem_data[13][3] ), .ZN(n14878) );
  AND2_X1 U19041 ( .A1(n25360), .A2(\xmem_data[14][3] ), .ZN(n14876) );
  AOI21_X1 U19042 ( .B1(n28503), .B2(\xmem_data[15][3] ), .A(n14876), .ZN(
        n14877) );
  NAND4_X1 U19043 ( .A1(n14880), .A2(n14879), .A3(n14878), .A4(n14877), .ZN(
        n14889) );
  BUF_X1 U19044 ( .A(n14912), .Z(n28427) );
  AOI22_X1 U19045 ( .A1(n28427), .A2(\xmem_data[0][3] ), .B1(n29410), .B2(
        \xmem_data[1][3] ), .ZN(n14887) );
  AOI22_X1 U19046 ( .A1(n30616), .A2(\xmem_data[2][3] ), .B1(n28428), .B2(
        \xmem_data[3][3] ), .ZN(n14886) );
  BUF_X1 U19047 ( .A(n14882), .Z(n28429) );
  AOI22_X1 U19048 ( .A1(n25581), .A2(\xmem_data[4][3] ), .B1(n30686), .B2(
        \xmem_data[5][3] ), .ZN(n14885) );
  AOI22_X1 U19049 ( .A1(n24167), .A2(\xmem_data[6][3] ), .B1(n14976), .B2(
        \xmem_data[7][3] ), .ZN(n14884) );
  NAND4_X1 U19050 ( .A1(n14887), .A2(n14886), .A3(n14885), .A4(n14884), .ZN(
        n14888) );
  OR2_X1 U19051 ( .A1(n14889), .A2(n14888), .ZN(n14906) );
  AOI22_X1 U19052 ( .A1(n3221), .A2(\xmem_data[16][3] ), .B1(n28137), .B2(
        \xmem_data[17][3] ), .ZN(n14897) );
  AOI22_X1 U19053 ( .A1(n3255), .A2(\xmem_data[20][3] ), .B1(n3374), .B2(
        \xmem_data[21][3] ), .ZN(n14891) );
  INV_X1 U19054 ( .A(n14891), .ZN(n14895) );
  AOI22_X1 U19055 ( .A1(n24207), .A2(\xmem_data[18][3] ), .B1(n3341), .B2(
        \xmem_data[19][3] ), .ZN(n14893) );
  NAND2_X1 U19056 ( .A1(n25422), .A2(\xmem_data[23][3] ), .ZN(n14892) );
  NAND2_X1 U19057 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  NOR2_X1 U19058 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  NAND2_X1 U19059 ( .A1(n14897), .A2(n14896), .ZN(n14904) );
  AOI22_X1 U19060 ( .A1(n27943), .A2(\xmem_data[24][3] ), .B1(n27944), .B2(
        \xmem_data[25][3] ), .ZN(n14902) );
  AOI22_X1 U19061 ( .A1(n28416), .A2(\xmem_data[26][3] ), .B1(n17041), .B2(
        \xmem_data[27][3] ), .ZN(n14901) );
  AOI22_X1 U19062 ( .A1(n25458), .A2(\xmem_data[28][3] ), .B1(n25672), .B2(
        \xmem_data[29][3] ), .ZN(n14900) );
  AOI22_X1 U19063 ( .A1(n27989), .A2(\xmem_data[30][3] ), .B1(n21007), .B2(
        \xmem_data[31][3] ), .ZN(n14899) );
  NAND4_X1 U19064 ( .A1(n14902), .A2(n14901), .A3(n14900), .A4(n14899), .ZN(
        n14903) );
  OR2_X1 U19065 ( .A1(n14904), .A2(n14903), .ZN(n14905) );
  NOR2_X1 U19066 ( .A1(n14906), .A2(n14905), .ZN(n14911) );
  NAND2_X1 U19067 ( .A1(n37190), .A2(n14907), .ZN(n14908) );
  INV_X1 U19068 ( .A(n14908), .ZN(n14910) );
  AOI22_X1 U19069 ( .A1(load_xaddr_val[5]), .A2(n14908), .B1(n14910), .B2(
        n4499), .ZN(n15009) );
  AOI22_X1 U19070 ( .A1(n14910), .A2(n39040), .B1(n14909), .B2(n14908), .ZN(
        n14967) );
  AOI22_X1 U19071 ( .A1(n28492), .A2(\xmem_data[96][3] ), .B1(n28687), .B2(
        \xmem_data[97][3] ), .ZN(n14918) );
  BUF_X1 U19072 ( .A(n14972), .Z(n28493) );
  AOI22_X1 U19073 ( .A1(n29190), .A2(\xmem_data[98][3] ), .B1(n28493), .B2(
        \xmem_data[99][3] ), .ZN(n14917) );
  BUF_X1 U19074 ( .A(n14973), .Z(n28494) );
  AOI22_X1 U19075 ( .A1(n28494), .A2(\xmem_data[100][3] ), .B1(n29816), .B2(
        \xmem_data[101][3] ), .ZN(n14916) );
  BUF_X1 U19076 ( .A(n14914), .Z(n28495) );
  AOI22_X1 U19077 ( .A1(n28495), .A2(\xmem_data[102][3] ), .B1(n20552), .B2(
        \xmem_data[103][3] ), .ZN(n14915) );
  NAND4_X1 U19078 ( .A1(n14918), .A2(n14917), .A3(n14916), .A4(n14915), .ZN(
        n14945) );
  AOI22_X1 U19079 ( .A1(n28500), .A2(\xmem_data[104][3] ), .B1(n30901), .B2(
        \xmem_data[105][3] ), .ZN(n14924) );
  AOI22_X1 U19080 ( .A1(n27567), .A2(\xmem_data[106][3] ), .B1(n28038), .B2(
        \xmem_data[107][3] ), .ZN(n14923) );
  AOI22_X1 U19081 ( .A1(n28075), .A2(\xmem_data[108][3] ), .B1(n3333), .B2(
        \xmem_data[109][3] ), .ZN(n14922) );
  BUF_X1 U19082 ( .A(n29064), .Z(n28503) );
  AND2_X1 U19083 ( .A1(n28501), .A2(\xmem_data[110][3] ), .ZN(n14920) );
  AOI21_X1 U19084 ( .B1(n28503), .B2(\xmem_data[111][3] ), .A(n14920), .ZN(
        n14921) );
  NAND4_X1 U19085 ( .A1(n14924), .A2(n14923), .A3(n14922), .A4(n14921), .ZN(
        n14944) );
  AOI22_X1 U19086 ( .A1(n3221), .A2(\xmem_data[112][3] ), .B1(n23770), .B2(
        \xmem_data[113][3] ), .ZN(n14932) );
  BUF_X1 U19087 ( .A(n14925), .Z(n28508) );
  AOI22_X1 U19088 ( .A1(n28508), .A2(\xmem_data[114][3] ), .B1(n3342), .B2(
        \xmem_data[115][3] ), .ZN(n14931) );
  BUF_X1 U19089 ( .A(n14927), .Z(n28509) );
  AOI22_X1 U19090 ( .A1(n28509), .A2(\xmem_data[116][3] ), .B1(n3128), .B2(
        \xmem_data[117][3] ), .ZN(n14930) );
  BUF_X1 U19091 ( .A(n14928), .Z(n28510) );
  AOI22_X1 U19092 ( .A1(n25450), .A2(\xmem_data[118][3] ), .B1(n28374), .B2(
        \xmem_data[119][3] ), .ZN(n14929) );
  NAND4_X1 U19093 ( .A1(n14932), .A2(n14931), .A3(n14930), .A4(n14929), .ZN(
        n14943) );
  AOI22_X1 U19094 ( .A1(n3358), .A2(\xmem_data[120][3] ), .B1(n31353), .B2(
        \xmem_data[121][3] ), .ZN(n14941) );
  AOI22_X1 U19095 ( .A1(n28515), .A2(\xmem_data[122][3] ), .B1(n27537), .B2(
        \xmem_data[123][3] ), .ZN(n14940) );
  BUF_X1 U19096 ( .A(n14935), .Z(n28517) );
  BUF_X1 U19097 ( .A(n29187), .Z(n28516) );
  AOI22_X1 U19098 ( .A1(n28517), .A2(\xmem_data[124][3] ), .B1(n3465), .B2(
        \xmem_data[125][3] ), .ZN(n14939) );
  AOI22_X1 U19099 ( .A1(n24457), .A2(\xmem_data[126][3] ), .B1(n28059), .B2(
        \xmem_data[127][3] ), .ZN(n14938) );
  NAND4_X1 U19100 ( .A1(n14941), .A2(n14940), .A3(n14939), .A4(n14938), .ZN(
        n14942) );
  OR4_X1 U19101 ( .A1(n14945), .A2(n14944), .A3(n14943), .A4(n14942), .ZN(
        n14969) );
  AND2_X1 U19102 ( .A1(n15009), .A2(n14967), .ZN(n28458) );
  AOI22_X1 U19103 ( .A1(n28492), .A2(\xmem_data[64][3] ), .B1(n17021), .B2(
        \xmem_data[65][3] ), .ZN(n14949) );
  AOI22_X1 U19104 ( .A1(n20941), .A2(\xmem_data[66][3] ), .B1(n28493), .B2(
        \xmem_data[67][3] ), .ZN(n14948) );
  AOI22_X1 U19105 ( .A1(n28494), .A2(\xmem_data[68][3] ), .B1(n28226), .B2(
        \xmem_data[69][3] ), .ZN(n14947) );
  AOI22_X1 U19106 ( .A1(n28495), .A2(\xmem_data[70][3] ), .B1(n25526), .B2(
        \xmem_data[71][3] ), .ZN(n14946) );
  NAND4_X1 U19107 ( .A1(n14949), .A2(n14948), .A3(n14947), .A4(n14946), .ZN(
        n14966) );
  AOI22_X1 U19108 ( .A1(n28500), .A2(\xmem_data[72][3] ), .B1(n29657), .B2(
        \xmem_data[73][3] ), .ZN(n14954) );
  AOI22_X1 U19109 ( .A1(n24468), .A2(\xmem_data[74][3] ), .B1(n30588), .B2(
        \xmem_data[75][3] ), .ZN(n14953) );
  AOI22_X1 U19110 ( .A1(n29328), .A2(\xmem_data[76][3] ), .B1(n29661), .B2(
        \xmem_data[77][3] ), .ZN(n14952) );
  AND2_X1 U19111 ( .A1(n28501), .A2(\xmem_data[78][3] ), .ZN(n14950) );
  AOI21_X1 U19112 ( .B1(n28503), .B2(\xmem_data[79][3] ), .A(n14950), .ZN(
        n14951) );
  NAND4_X1 U19113 ( .A1(n14954), .A2(n14953), .A3(n14952), .A4(n14951), .ZN(
        n14965) );
  AOI22_X1 U19114 ( .A1(n3218), .A2(\xmem_data[80][3] ), .B1(n23770), .B2(
        \xmem_data[81][3] ), .ZN(n14958) );
  AOI22_X1 U19115 ( .A1(n28508), .A2(\xmem_data[82][3] ), .B1(n3322), .B2(
        \xmem_data[83][3] ), .ZN(n14957) );
  AOI22_X1 U19116 ( .A1(n28509), .A2(\xmem_data[84][3] ), .B1(n3135), .B2(
        \xmem_data[85][3] ), .ZN(n14956) );
  AOI22_X1 U19117 ( .A1(n29306), .A2(\xmem_data[86][3] ), .B1(n28374), .B2(
        \xmem_data[87][3] ), .ZN(n14955) );
  NAND4_X1 U19118 ( .A1(n14958), .A2(n14957), .A3(n14956), .A4(n14955), .ZN(
        n14964) );
  AOI22_X1 U19119 ( .A1(n28517), .A2(\xmem_data[92][3] ), .B1(n3465), .B2(
        \xmem_data[93][3] ), .ZN(n14962) );
  AOI22_X1 U19120 ( .A1(n28515), .A2(\xmem_data[90][3] ), .B1(n29310), .B2(
        \xmem_data[91][3] ), .ZN(n14961) );
  AOI22_X1 U19121 ( .A1(n24590), .A2(\xmem_data[88][3] ), .B1(n17064), .B2(
        \xmem_data[89][3] ), .ZN(n14960) );
  AOI22_X1 U19122 ( .A1(n27989), .A2(\xmem_data[94][3] ), .B1(n27919), .B2(
        \xmem_data[95][3] ), .ZN(n14959) );
  NAND4_X1 U19123 ( .A1(n14962), .A2(n14961), .A3(n14960), .A4(n14959), .ZN(
        n14963) );
  OR4_X1 U19124 ( .A1(n14966), .A2(n14965), .A3(n14964), .A4(n14963), .ZN(
        n14968) );
  INV_X1 U19125 ( .A(n14967), .ZN(n15010) );
  NOR2_X1 U19126 ( .A1(n15009), .A2(n15010), .ZN(n28526) );
  AOI22_X1 U19127 ( .A1(n14969), .A2(n28458), .B1(n14968), .B2(n28526), .ZN(
        n15015) );
  AOI22_X1 U19128 ( .A1(n25520), .A2(\xmem_data[32][3] ), .B1(n25400), .B2(
        \xmem_data[33][3] ), .ZN(n14980) );
  AOI22_X1 U19129 ( .A1(n27523), .A2(\xmem_data[34][3] ), .B1(n24615), .B2(
        \xmem_data[35][3] ), .ZN(n14979) );
  BUF_X1 U19130 ( .A(n14973), .Z(n28462) );
  BUF_X1 U19131 ( .A(n14974), .Z(n28461) );
  AOI22_X1 U19132 ( .A1(n28462), .A2(\xmem_data[36][3] ), .B1(n28461), .B2(
        \xmem_data[37][3] ), .ZN(n14978) );
  AOI22_X1 U19133 ( .A1(n27975), .A2(\xmem_data[38][3] ), .B1(n20734), .B2(
        \xmem_data[39][3] ), .ZN(n14977) );
  NAND4_X1 U19134 ( .A1(n14980), .A2(n14979), .A3(n14978), .A4(n14977), .ZN(
        n15008) );
  BUF_X1 U19135 ( .A(n14982), .Z(n28467) );
  AOI22_X1 U19136 ( .A1(n28468), .A2(\xmem_data[40][3] ), .B1(n28467), .B2(
        \xmem_data[41][3] ), .ZN(n14987) );
  AOI22_X1 U19137 ( .A1(n28035), .A2(\xmem_data[42][3] ), .B1(n27959), .B2(
        \xmem_data[43][3] ), .ZN(n14986) );
  AOI22_X1 U19138 ( .A1(n30571), .A2(\xmem_data[44][3] ), .B1(n3449), .B2(
        \xmem_data[45][3] ), .ZN(n14985) );
  BUF_X1 U19139 ( .A(n29064), .Z(n28470) );
  AOI22_X1 U19140 ( .A1(n25360), .A2(\xmem_data[46][3] ), .B1(n28470), .B2(
        \xmem_data[47][3] ), .ZN(n14984) );
  NAND4_X1 U19141 ( .A1(n14987), .A2(n14986), .A3(n14985), .A4(n14984), .ZN(
        n15007) );
  AOI22_X1 U19142 ( .A1(n3222), .A2(\xmem_data[48][3] ), .B1(n27708), .B2(
        \xmem_data[49][3] ), .ZN(n14995) );
  BUF_X1 U19143 ( .A(n14989), .Z(n28476) );
  BUF_X1 U19144 ( .A(n14990), .Z(n28475) );
  AOI22_X1 U19145 ( .A1(n28476), .A2(\xmem_data[50][3] ), .B1(n28475), .B2(
        \xmem_data[51][3] ), .ZN(n14994) );
  AOI22_X1 U19146 ( .A1(n20806), .A2(\xmem_data[52][3] ), .B1(n28084), .B2(
        \xmem_data[53][3] ), .ZN(n14993) );
  AOI22_X1 U19147 ( .A1(n25514), .A2(\xmem_data[54][3] ), .B1(n23813), .B2(
        \xmem_data[55][3] ), .ZN(n14992) );
  NAND4_X1 U19148 ( .A1(n14995), .A2(n14994), .A3(n14993), .A4(n14992), .ZN(
        n15006) );
  BUF_X1 U19149 ( .A(n14996), .Z(n28481) );
  AOI22_X1 U19150 ( .A1(n28481), .A2(\xmem_data[56][3] ), .B1(n24556), .B2(
        \xmem_data[57][3] ), .ZN(n15004) );
  AOI22_X1 U19151 ( .A1(n14998), .A2(\xmem_data[58][3] ), .B1(n16986), .B2(
        \xmem_data[59][3] ), .ZN(n15003) );
  AOI22_X1 U19152 ( .A1(n20584), .A2(\xmem_data[60][3] ), .B1(n29807), .B2(
        \xmem_data[61][3] ), .ZN(n15002) );
  AOI22_X1 U19153 ( .A1(n30542), .A2(\xmem_data[62][3] ), .B1(n29010), .B2(
        \xmem_data[63][3] ), .ZN(n15001) );
  NAND4_X1 U19154 ( .A1(n15004), .A2(n15003), .A3(n15002), .A4(n15001), .ZN(
        n15005) );
  OR4_X1 U19155 ( .A1(n15008), .A2(n15007), .A3(n15006), .A4(n15005), .ZN(
        n15013) );
  AND2_X1 U19156 ( .A1(n15010), .A2(n15009), .ZN(n28490) );
  NOR2_X1 U19157 ( .A1(n15043), .A2(n39006), .ZN(n15012) );
  AOI21_X1 U19158 ( .B1(n15013), .B2(n28490), .A(n3890), .ZN(n15014) );
  XOR2_X1 U19159 ( .A(\fmem_data[29][7] ), .B(\fmem_data[29][6] ), .Z(n15016)
         );
  AOI22_X1 U19160 ( .A1(n28501), .A2(\xmem_data[14][4] ), .B1(n27439), .B2(
        \xmem_data[15][4] ), .ZN(n15027) );
  AOI22_X1 U19161 ( .A1(n25685), .A2(\xmem_data[12][4] ), .B1(n3414), .B2(
        \xmem_data[13][4] ), .ZN(n15017) );
  INV_X1 U19162 ( .A(n15017), .ZN(n15020) );
  AOI22_X1 U19163 ( .A1(n28329), .A2(\xmem_data[10][4] ), .B1(n25358), .B2(
        \xmem_data[11][4] ), .ZN(n15018) );
  INV_X1 U19164 ( .A(n15018), .ZN(n15019) );
  NOR2_X1 U19165 ( .A1(n15020), .A2(n15019), .ZN(n15026) );
  AOI22_X1 U19166 ( .A1(n27526), .A2(\xmem_data[8][4] ), .B1(n30674), .B2(
        \xmem_data[9][4] ), .ZN(n15025) );
  AOI22_X1 U19167 ( .A1(n28427), .A2(\xmem_data[0][4] ), .B1(n27825), .B2(
        \xmem_data[1][4] ), .ZN(n15024) );
  AOI22_X1 U19168 ( .A1(n23776), .A2(\xmem_data[2][4] ), .B1(n28428), .B2(
        \xmem_data[3][4] ), .ZN(n15023) );
  AOI22_X1 U19169 ( .A1(n20506), .A2(\xmem_data[4][4] ), .B1(n3329), .B2(
        \xmem_data[5][4] ), .ZN(n15022) );
  AOI22_X1 U19170 ( .A1(n20983), .A2(\xmem_data[6][4] ), .B1(n20552), .B2(
        \xmem_data[7][4] ), .ZN(n15021) );
  NAND4_X1 U19171 ( .A1(n15027), .A2(n15026), .A3(n15025), .A4(n3746), .ZN(
        n15042) );
  AOI22_X1 U19172 ( .A1(n3218), .A2(\xmem_data[16][4] ), .B1(n28137), .B2(
        \xmem_data[17][4] ), .ZN(n15034) );
  AOI22_X1 U19173 ( .A1(n3255), .A2(\xmem_data[20][4] ), .B1(n17063), .B2(
        \xmem_data[21][4] ), .ZN(n15028) );
  INV_X1 U19174 ( .A(n15028), .ZN(n15032) );
  AOI22_X1 U19175 ( .A1(n20787), .A2(\xmem_data[18][4] ), .B1(n24438), .B2(
        \xmem_data[19][4] ), .ZN(n15030) );
  NAND2_X1 U19176 ( .A1(n25422), .A2(\xmem_data[23][4] ), .ZN(n15029) );
  NAND2_X1 U19177 ( .A1(n15030), .A2(n15029), .ZN(n15031) );
  NOR2_X1 U19178 ( .A1(n15032), .A2(n15031), .ZN(n15033) );
  NAND2_X1 U19179 ( .A1(n15034), .A2(n15033), .ZN(n15040) );
  AOI22_X1 U19180 ( .A1(n25456), .A2(\xmem_data[24][4] ), .B1(n27911), .B2(
        \xmem_data[25][4] ), .ZN(n15038) );
  AOI22_X1 U19181 ( .A1(n28416), .A2(\xmem_data[26][4] ), .B1(n13436), .B2(
        \xmem_data[27][4] ), .ZN(n15037) );
  AOI22_X1 U19182 ( .A1(n25671), .A2(\xmem_data[28][4] ), .B1(n16988), .B2(
        \xmem_data[29][4] ), .ZN(n15036) );
  AOI22_X1 U19183 ( .A1(n29162), .A2(\xmem_data[30][4] ), .B1(n23717), .B2(
        \xmem_data[31][4] ), .ZN(n15035) );
  NAND4_X1 U19184 ( .A1(n15038), .A2(n15037), .A3(n15036), .A4(n15035), .ZN(
        n15039) );
  OR2_X1 U19185 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  NOR2_X1 U19186 ( .A1(n15042), .A2(n15041), .ZN(n15045) );
  NAND2_X1 U19187 ( .A1(n28045), .A2(\xmem_data[22][4] ), .ZN(n15044) );
  AOI21_X1 U19188 ( .B1(n15045), .B2(n15044), .A(n15043), .ZN(n15070) );
  AOI22_X1 U19189 ( .A1(n28468), .A2(\xmem_data[40][4] ), .B1(n28467), .B2(
        \xmem_data[41][4] ), .ZN(n15050) );
  AOI22_X1 U19190 ( .A1(n20769), .A2(\xmem_data[42][4] ), .B1(n25358), .B2(
        \xmem_data[43][4] ), .ZN(n15049) );
  AOI22_X1 U19191 ( .A1(n31262), .A2(\xmem_data[44][4] ), .B1(n24693), .B2(
        \xmem_data[45][4] ), .ZN(n15048) );
  AND2_X1 U19192 ( .A1(n25360), .A2(\xmem_data[46][4] ), .ZN(n15046) );
  AOI21_X1 U19193 ( .B1(n28470), .B2(\xmem_data[47][4] ), .A(n15046), .ZN(
        n15047) );
  NAND4_X1 U19194 ( .A1(n15050), .A2(n15049), .A3(n15048), .A4(n15047), .ZN(
        n15067) );
  AOI22_X1 U19195 ( .A1(n29316), .A2(\xmem_data[32][4] ), .B1(n16990), .B2(
        \xmem_data[33][4] ), .ZN(n15054) );
  AOI22_X1 U19196 ( .A1(n30515), .A2(\xmem_data[34][4] ), .B1(n24190), .B2(
        \xmem_data[35][4] ), .ZN(n15053) );
  AOI22_X1 U19197 ( .A1(n28462), .A2(\xmem_data[36][4] ), .B1(n28461), .B2(
        \xmem_data[37][4] ), .ZN(n15052) );
  AOI22_X1 U19198 ( .A1(n30599), .A2(\xmem_data[38][4] ), .B1(n29325), .B2(
        \xmem_data[39][4] ), .ZN(n15051) );
  NAND4_X1 U19199 ( .A1(n15054), .A2(n15053), .A3(n15052), .A4(n15051), .ZN(
        n15065) );
  AOI22_X1 U19200 ( .A1(n3221), .A2(\xmem_data[48][4] ), .B1(n24632), .B2(
        \xmem_data[49][4] ), .ZN(n15058) );
  AOI22_X1 U19201 ( .A1(n28476), .A2(\xmem_data[50][4] ), .B1(n28475), .B2(
        \xmem_data[51][4] ), .ZN(n15057) );
  AOI22_X1 U19202 ( .A1(n29181), .A2(\xmem_data[52][4] ), .B1(n3129), .B2(
        \xmem_data[53][4] ), .ZN(n15056) );
  AOI22_X1 U19203 ( .A1(n3231), .A2(\xmem_data[54][4] ), .B1(n27508), .B2(
        \xmem_data[55][4] ), .ZN(n15055) );
  NAND4_X1 U19204 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        n15064) );
  AOI22_X1 U19205 ( .A1(n28481), .A2(\xmem_data[56][4] ), .B1(n30943), .B2(
        \xmem_data[57][4] ), .ZN(n15062) );
  AOI22_X1 U19206 ( .A1(n21015), .A2(\xmem_data[58][4] ), .B1(n30891), .B2(
        \xmem_data[59][4] ), .ZN(n15061) );
  AOI22_X1 U19207 ( .A1(n25671), .A2(\xmem_data[60][4] ), .B1(n25607), .B2(
        \xmem_data[61][4] ), .ZN(n15060) );
  AOI22_X1 U19208 ( .A1(n24134), .A2(\xmem_data[62][4] ), .B1(n28096), .B2(
        \xmem_data[63][4] ), .ZN(n15059) );
  NAND4_X1 U19209 ( .A1(n15062), .A2(n15061), .A3(n15060), .A4(n15059), .ZN(
        n15063) );
  OR3_X1 U19210 ( .A1(n15065), .A2(n15064), .A3(n15063), .ZN(n15066) );
  OAI21_X1 U19211 ( .B1(n15067), .B2(n15066), .A(n28490), .ZN(n15068) );
  INV_X1 U19212 ( .A(n15068), .ZN(n15069) );
  NOR2_X1 U19213 ( .A1(n15070), .A2(n15069), .ZN(n15115) );
  AOI22_X1 U19214 ( .A1(n28492), .A2(\xmem_data[96][4] ), .B1(n23777), .B2(
        \xmem_data[97][4] ), .ZN(n15074) );
  AOI22_X1 U19215 ( .A1(n25435), .A2(\xmem_data[98][4] ), .B1(n28493), .B2(
        \xmem_data[99][4] ), .ZN(n15073) );
  AOI22_X1 U19216 ( .A1(n28494), .A2(\xmem_data[100][4] ), .B1(n25401), .B2(
        \xmem_data[101][4] ), .ZN(n15072) );
  AOI22_X1 U19217 ( .A1(n28495), .A2(\xmem_data[102][4] ), .B1(n3209), .B2(
        \xmem_data[103][4] ), .ZN(n15071) );
  NAND4_X1 U19218 ( .A1(n15074), .A2(n15073), .A3(n15072), .A4(n15071), .ZN(
        n15090) );
  AOI22_X1 U19219 ( .A1(n28500), .A2(\xmem_data[104][4] ), .B1(n29820), .B2(
        \xmem_data[105][4] ), .ZN(n15078) );
  AOI22_X1 U19220 ( .A1(n20951), .A2(\xmem_data[106][4] ), .B1(n20827), .B2(
        \xmem_data[107][4] ), .ZN(n15077) );
  AOI22_X1 U19221 ( .A1(n25561), .A2(\xmem_data[108][4] ), .B1(n23732), .B2(
        \xmem_data[109][4] ), .ZN(n15076) );
  AOI22_X1 U19222 ( .A1(n28501), .A2(\xmem_data[110][4] ), .B1(n28503), .B2(
        \xmem_data[111][4] ), .ZN(n15075) );
  NAND4_X1 U19223 ( .A1(n15078), .A2(n15077), .A3(n15076), .A4(n15075), .ZN(
        n15089) );
  AOI22_X1 U19224 ( .A1(n3220), .A2(\xmem_data[112][4] ), .B1(n27708), .B2(
        \xmem_data[113][4] ), .ZN(n15082) );
  AOI22_X1 U19225 ( .A1(n28508), .A2(\xmem_data[114][4] ), .B1(n3342), .B2(
        \xmem_data[115][4] ), .ZN(n15081) );
  AOI22_X1 U19226 ( .A1(n28509), .A2(\xmem_data[116][4] ), .B1(n3137), .B2(
        \xmem_data[117][4] ), .ZN(n15080) );
  AOI22_X1 U19227 ( .A1(n28045), .A2(\xmem_data[118][4] ), .B1(n28374), .B2(
        \xmem_data[119][4] ), .ZN(n15079) );
  NAND4_X1 U19228 ( .A1(n15082), .A2(n15081), .A3(n15080), .A4(n15079), .ZN(
        n15088) );
  AOI22_X1 U19229 ( .A1(n3358), .A2(\xmem_data[120][4] ), .B1(n31327), .B2(
        \xmem_data[121][4] ), .ZN(n15086) );
  AOI22_X1 U19230 ( .A1(n28515), .A2(\xmem_data[122][4] ), .B1(n16986), .B2(
        \xmem_data[123][4] ), .ZN(n15085) );
  AOI22_X1 U19231 ( .A1(n28517), .A2(\xmem_data[124][4] ), .B1(n30666), .B2(
        \xmem_data[125][4] ), .ZN(n15084) );
  AOI22_X1 U19232 ( .A1(n3208), .A2(\xmem_data[126][4] ), .B1(n30949), .B2(
        \xmem_data[127][4] ), .ZN(n15083) );
  NAND4_X1 U19233 ( .A1(n15086), .A2(n15085), .A3(n15084), .A4(n15083), .ZN(
        n15087) );
  OR4_X1 U19234 ( .A1(n15090), .A2(n15089), .A3(n15088), .A4(n15087), .ZN(
        n15113) );
  AOI22_X1 U19235 ( .A1(n27518), .A2(\xmem_data[64][4] ), .B1(n27825), .B2(
        \xmem_data[65][4] ), .ZN(n15094) );
  AOI22_X1 U19236 ( .A1(n30515), .A2(\xmem_data[66][4] ), .B1(n20593), .B2(
        \xmem_data[67][4] ), .ZN(n15093) );
  AOI22_X1 U19237 ( .A1(n28462), .A2(\xmem_data[68][4] ), .B1(n28461), .B2(
        \xmem_data[69][4] ), .ZN(n15092) );
  AOI22_X1 U19238 ( .A1(n31314), .A2(\xmem_data[70][4] ), .B1(n24685), .B2(
        \xmem_data[71][4] ), .ZN(n15091) );
  NAND4_X1 U19239 ( .A1(n15094), .A2(n15093), .A3(n15092), .A4(n15091), .ZN(
        n15111) );
  AOI22_X1 U19240 ( .A1(n28468), .A2(\xmem_data[72][4] ), .B1(n28467), .B2(
        \xmem_data[73][4] ), .ZN(n15099) );
  AOI22_X1 U19241 ( .A1(n27435), .A2(\xmem_data[74][4] ), .B1(n28038), .B2(
        \xmem_data[75][4] ), .ZN(n15098) );
  AOI22_X1 U19242 ( .A1(n22752), .A2(\xmem_data[76][4] ), .B1(n3433), .B2(
        \xmem_data[77][4] ), .ZN(n15097) );
  AND2_X1 U19243 ( .A1(n24439), .A2(\xmem_data[78][4] ), .ZN(n15095) );
  AOI21_X1 U19244 ( .B1(n28470), .B2(\xmem_data[79][4] ), .A(n15095), .ZN(
        n15096) );
  NAND4_X1 U19245 ( .A1(n15099), .A2(n15098), .A3(n15097), .A4(n15096), .ZN(
        n15110) );
  AOI22_X1 U19246 ( .A1(n3221), .A2(\xmem_data[80][4] ), .B1(n30593), .B2(
        \xmem_data[81][4] ), .ZN(n15103) );
  AOI22_X1 U19247 ( .A1(n28476), .A2(\xmem_data[82][4] ), .B1(n28475), .B2(
        \xmem_data[83][4] ), .ZN(n15102) );
  AOI22_X1 U19248 ( .A1(n28372), .A2(\xmem_data[84][4] ), .B1(n3282), .B2(
        \xmem_data[85][4] ), .ZN(n15101) );
  AOI22_X1 U19249 ( .A1(n28510), .A2(\xmem_data[86][4] ), .B1(n27551), .B2(
        \xmem_data[87][4] ), .ZN(n15100) );
  NAND4_X1 U19250 ( .A1(n15103), .A2(n15102), .A3(n15101), .A4(n15100), .ZN(
        n15109) );
  AOI22_X1 U19251 ( .A1(n28481), .A2(\xmem_data[88][4] ), .B1(n24157), .B2(
        \xmem_data[89][4] ), .ZN(n15107) );
  AOI22_X1 U19252 ( .A1(n28375), .A2(\xmem_data[90][4] ), .B1(n29023), .B2(
        \xmem_data[91][4] ), .ZN(n15106) );
  AOI22_X1 U19253 ( .A1(n20717), .A2(\xmem_data[92][4] ), .B1(n27755), .B2(
        \xmem_data[93][4] ), .ZN(n15105) );
  AOI22_X1 U19254 ( .A1(n28335), .A2(\xmem_data[94][4] ), .B1(n25434), .B2(
        \xmem_data[95][4] ), .ZN(n15104) );
  NAND4_X1 U19255 ( .A1(n15107), .A2(n15106), .A3(n15105), .A4(n15104), .ZN(
        n15108) );
  OR4_X1 U19256 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15112) );
  AOI22_X1 U19257 ( .A1(n28458), .A2(n15113), .B1(n28526), .B2(n15112), .ZN(
        n15114) );
  XNOR2_X1 U19258 ( .A(n32242), .B(\fmem_data[29][7] ), .ZN(n33128) );
  OAI22_X1 U19259 ( .A1(n30450), .A2(n35614), .B1(n33128), .B2(n35615), .ZN(
        n34880) );
  AOI22_X1 U19260 ( .A1(n30886), .A2(\xmem_data[6][3] ), .B1(n20958), .B2(
        \xmem_data[7][3] ), .ZN(n15116) );
  AOI22_X1 U19261 ( .A1(n23813), .A2(\xmem_data[4][3] ), .B1(n30854), .B2(
        \xmem_data[5][3] ), .ZN(n15118) );
  NAND2_X1 U19262 ( .A1(n30710), .A2(\xmem_data[2][3] ), .ZN(n15117) );
  NAND2_X1 U19263 ( .A1(n15118), .A2(n15117), .ZN(n15121) );
  AOI22_X1 U19264 ( .A1(n3341), .A2(\xmem_data[0][3] ), .B1(n29181), .B2(
        \xmem_data[1][3] ), .ZN(n15119) );
  INV_X1 U19265 ( .A(n15119), .ZN(n15120) );
  OR3_X1 U19266 ( .A1(n15122), .A2(n15121), .A3(n15120), .ZN(n15128) );
  AOI22_X1 U19267 ( .A1(n28980), .A2(\xmem_data[8][3] ), .B1(n24160), .B2(
        \xmem_data[9][3] ), .ZN(n15126) );
  AOI22_X1 U19268 ( .A1(n28231), .A2(\xmem_data[10][3] ), .B1(n30542), .B2(
        \xmem_data[11][3] ), .ZN(n15125) );
  AOI22_X1 U19269 ( .A1(n30949), .A2(\xmem_data[12][3] ), .B1(n31270), .B2(
        \xmem_data[13][3] ), .ZN(n15124) );
  AOI22_X1 U19270 ( .A1(n30872), .A2(\xmem_data[14][3] ), .B1(n30871), .B2(
        \xmem_data[15][3] ), .ZN(n15123) );
  NAND4_X1 U19271 ( .A1(n15126), .A2(n15125), .A3(n15124), .A4(n15123), .ZN(
        n15127) );
  NOR2_X1 U19272 ( .A1(n15128), .A2(n15127), .ZN(n15148) );
  AOI22_X1 U19273 ( .A1(n29254), .A2(\xmem_data[28][3] ), .B1(n3217), .B2(
        \xmem_data[29][3] ), .ZN(n15129) );
  INV_X1 U19274 ( .A(n15129), .ZN(n15146) );
  AOI22_X1 U19275 ( .A1(n23740), .A2(\xmem_data[30][3] ), .B1(n20500), .B2(
        \xmem_data[31][3] ), .ZN(n15130) );
  INV_X1 U19276 ( .A(n15130), .ZN(n15133) );
  AOI22_X1 U19277 ( .A1(n30864), .A2(\xmem_data[26][3] ), .B1(n30863), .B2(
        \xmem_data[27][3] ), .ZN(n15131) );
  INV_X1 U19278 ( .A(n15131), .ZN(n15132) );
  NOR2_X1 U19279 ( .A1(n15133), .A2(n15132), .ZN(n15135) );
  AOI22_X1 U19280 ( .A1(n30862), .A2(\xmem_data[24][3] ), .B1(n30861), .B2(
        \xmem_data[25][3] ), .ZN(n15134) );
  NAND2_X1 U19281 ( .A1(n15135), .A2(n15134), .ZN(n15145) );
  AOI22_X1 U19282 ( .A1(n20770), .A2(\xmem_data[22][3] ), .B1(n27567), .B2(
        \xmem_data[23][3] ), .ZN(n15143) );
  AOI22_X1 U19283 ( .A1(n30849), .A2(\xmem_data[16][3] ), .B1(n3372), .B2(
        \xmem_data[17][3] ), .ZN(n15136) );
  INV_X1 U19284 ( .A(n15136), .ZN(n15141) );
  AOI22_X1 U19285 ( .A1(n29325), .A2(\xmem_data[20][3] ), .B1(n31256), .B2(
        \xmem_data[21][3] ), .ZN(n15139) );
  NAND2_X1 U19286 ( .A1(n28045), .A2(\xmem_data[3][3] ), .ZN(n15138) );
  AOI22_X1 U19287 ( .A1(n29054), .A2(\xmem_data[18][3] ), .B1(n14975), .B2(
        \xmem_data[19][3] ), .ZN(n15137) );
  NOR2_X1 U19288 ( .A1(n15141), .A2(n15140), .ZN(n15142) );
  NAND2_X1 U19289 ( .A1(n15143), .A2(n15142), .ZN(n15144) );
  NOR3_X1 U19290 ( .A1(n15146), .A2(n15145), .A3(n15144), .ZN(n15147) );
  AOI21_X1 U19291 ( .B1(n15148), .B2(n15147), .A(n30879), .ZN(n15149) );
  INV_X1 U19292 ( .A(n15149), .ZN(n15216) );
  AOI22_X1 U19293 ( .A1(n22709), .A2(\xmem_data[64][3] ), .B1(n27994), .B2(
        \xmem_data[65][3] ), .ZN(n15153) );
  AOI22_X1 U19294 ( .A1(n3129), .A2(\xmem_data[66][3] ), .B1(n27547), .B2(
        \xmem_data[67][3] ), .ZN(n15152) );
  AOI22_X1 U19295 ( .A1(n27551), .A2(\xmem_data[68][3] ), .B1(n27943), .B2(
        \xmem_data[69][3] ), .ZN(n15151) );
  AOI22_X1 U19296 ( .A1(n30943), .A2(\xmem_data[70][3] ), .B1(n13168), .B2(
        \xmem_data[71][3] ), .ZN(n15150) );
  NAND4_X1 U19297 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        n15169) );
  AOI22_X1 U19298 ( .A1(n17041), .A2(\xmem_data[72][3] ), .B1(n29046), .B2(
        \xmem_data[73][3] ), .ZN(n15157) );
  AOI22_X1 U19299 ( .A1(n20718), .A2(\xmem_data[74][3] ), .B1(n13188), .B2(
        \xmem_data[75][3] ), .ZN(n15156) );
  AOI22_X1 U19300 ( .A1(n30949), .A2(\xmem_data[76][3] ), .B1(n31329), .B2(
        \xmem_data[77][3] ), .ZN(n15155) );
  AOI22_X1 U19301 ( .A1(n30950), .A2(\xmem_data[78][3] ), .B1(n29190), .B2(
        \xmem_data[79][3] ), .ZN(n15154) );
  NAND4_X1 U19302 ( .A1(n15157), .A2(n15156), .A3(n15155), .A4(n15154), .ZN(
        n15168) );
  AOI22_X1 U19303 ( .A1(n30956), .A2(\xmem_data[80][3] ), .B1(n30955), .B2(
        \xmem_data[81][3] ), .ZN(n15161) );
  AOI22_X1 U19304 ( .A1(n3270), .A2(\xmem_data[82][3] ), .B1(n20507), .B2(
        \xmem_data[83][3] ), .ZN(n15160) );
  AOI22_X1 U19305 ( .A1(n27542), .A2(\xmem_data[84][3] ), .B1(n29017), .B2(
        \xmem_data[85][3] ), .ZN(n15159) );
  AOI22_X1 U19306 ( .A1(n20567), .A2(\xmem_data[86][3] ), .B1(n31344), .B2(
        \xmem_data[87][3] ), .ZN(n15158) );
  NAND4_X1 U19307 ( .A1(n15161), .A2(n15160), .A3(n15159), .A4(n15158), .ZN(
        n15167) );
  AOI22_X1 U19308 ( .A1(n3380), .A2(\xmem_data[88][3] ), .B1(n27499), .B2(
        \xmem_data[89][3] ), .ZN(n15165) );
  AOI22_X1 U19309 ( .A1(n3333), .A2(\xmem_data[90][3] ), .B1(n30589), .B2(
        \xmem_data[91][3] ), .ZN(n15164) );
  AOI22_X1 U19310 ( .A1(n30962), .A2(\xmem_data[92][3] ), .B1(n3222), .B2(
        \xmem_data[93][3] ), .ZN(n15163) );
  AOI22_X1 U19311 ( .A1(n30964), .A2(\xmem_data[94][3] ), .B1(n30963), .B2(
        \xmem_data[95][3] ), .ZN(n15162) );
  NAND4_X1 U19312 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15166) );
  OR4_X1 U19313 ( .A1(n15169), .A2(n15168), .A3(n15167), .A4(n15166), .ZN(
        n15170) );
  NAND2_X1 U19314 ( .A1(n15170), .A2(n30974), .ZN(n15215) );
  AOI22_X1 U19315 ( .A1(n25449), .A2(\xmem_data[96][3] ), .B1(n28509), .B2(
        \xmem_data[97][3] ), .ZN(n15174) );
  AOI22_X1 U19316 ( .A1(n3128), .A2(\xmem_data[98][3] ), .B1(n28045), .B2(
        \xmem_data[99][3] ), .ZN(n15173) );
  AOI22_X1 U19317 ( .A1(n27551), .A2(\xmem_data[100][3] ), .B1(n27988), .B2(
        \xmem_data[101][3] ), .ZN(n15172) );
  AOI22_X1 U19318 ( .A1(n30943), .A2(\xmem_data[102][3] ), .B1(n13168), .B2(
        \xmem_data[103][3] ), .ZN(n15171) );
  NAND4_X1 U19319 ( .A1(n15174), .A2(n15173), .A3(n15172), .A4(n15171), .ZN(
        n15190) );
  AOI22_X1 U19320 ( .A1(n30614), .A2(\xmem_data[104][3] ), .B1(n14898), .B2(
        \xmem_data[105][3] ), .ZN(n15178) );
  AOI22_X1 U19321 ( .A1(n3121), .A2(\xmem_data[106][3] ), .B1(n29162), .B2(
        \xmem_data[107][3] ), .ZN(n15177) );
  AOI22_X1 U19322 ( .A1(n30949), .A2(\xmem_data[108][3] ), .B1(n31355), .B2(
        \xmem_data[109][3] ), .ZN(n15176) );
  AOI22_X1 U19323 ( .A1(n30950), .A2(\xmem_data[110][3] ), .B1(n29238), .B2(
        \xmem_data[111][3] ), .ZN(n15175) );
  NAND4_X1 U19324 ( .A1(n15178), .A2(n15177), .A3(n15176), .A4(n15175), .ZN(
        n15189) );
  AOI22_X1 U19325 ( .A1(n30956), .A2(\xmem_data[112][3] ), .B1(n30955), .B2(
        \xmem_data[113][3] ), .ZN(n15182) );
  AOI22_X1 U19326 ( .A1(n29816), .A2(\xmem_data[114][3] ), .B1(n14975), .B2(
        \xmem_data[115][3] ), .ZN(n15181) );
  AOI22_X1 U19327 ( .A1(n28293), .A2(\xmem_data[116][3] ), .B1(n22751), .B2(
        \xmem_data[117][3] ), .ZN(n15180) );
  AOI22_X1 U19328 ( .A1(n20952), .A2(\xmem_data[118][3] ), .B1(n25440), .B2(
        \xmem_data[119][3] ), .ZN(n15179) );
  NAND4_X1 U19329 ( .A1(n15182), .A2(n15181), .A3(n15180), .A4(n15179), .ZN(
        n15188) );
  AOI22_X1 U19330 ( .A1(n27925), .A2(\xmem_data[120][3] ), .B1(n25629), .B2(
        \xmem_data[121][3] ), .ZN(n15186) );
  AOI22_X1 U19331 ( .A1(n3333), .A2(\xmem_data[122][3] ), .B1(n30589), .B2(
        \xmem_data[123][3] ), .ZN(n15185) );
  AOI22_X1 U19332 ( .A1(n30962), .A2(\xmem_data[124][3] ), .B1(n3220), .B2(
        \xmem_data[125][3] ), .ZN(n15184) );
  AOI22_X1 U19333 ( .A1(n30964), .A2(\xmem_data[126][3] ), .B1(n30963), .B2(
        \xmem_data[127][3] ), .ZN(n15183) );
  NAND4_X1 U19334 ( .A1(n15186), .A2(n15185), .A3(n15184), .A4(n15183), .ZN(
        n15187) );
  OR4_X1 U19335 ( .A1(n15190), .A2(n15189), .A3(n15188), .A4(n15187), .ZN(
        n15191) );
  NAND2_X1 U19336 ( .A1(n15191), .A2(n30976), .ZN(n15214) );
  AOI22_X1 U19337 ( .A1(n30883), .A2(\xmem_data[32][3] ), .B1(n30882), .B2(
        \xmem_data[33][3] ), .ZN(n15195) );
  AOI22_X1 U19338 ( .A1(n25451), .A2(\xmem_data[34][3] ), .B1(n28045), .B2(
        \xmem_data[35][3] ), .ZN(n15194) );
  AOI22_X1 U19339 ( .A1(n30885), .A2(\xmem_data[36][3] ), .B1(n30884), .B2(
        \xmem_data[37][3] ), .ZN(n15193) );
  AOI22_X1 U19340 ( .A1(n30886), .A2(\xmem_data[38][3] ), .B1(n28345), .B2(
        \xmem_data[39][3] ), .ZN(n15192) );
  NAND4_X1 U19341 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15211) );
  AOI22_X1 U19342 ( .A1(n30891), .A2(\xmem_data[40][3] ), .B1(n20584), .B2(
        \xmem_data[41][3] ), .ZN(n15199) );
  AOI22_X1 U19343 ( .A1(n27455), .A2(\xmem_data[42][3] ), .B1(n31269), .B2(
        \xmem_data[43][3] ), .ZN(n15198) );
  AOI22_X1 U19344 ( .A1(n24708), .A2(\xmem_data[44][3] ), .B1(n28427), .B2(
        \xmem_data[45][3] ), .ZN(n15197) );
  AOI22_X1 U19345 ( .A1(n30893), .A2(\xmem_data[46][3] ), .B1(n20941), .B2(
        \xmem_data[47][3] ), .ZN(n15196) );
  NAND4_X1 U19346 ( .A1(n15199), .A2(n15198), .A3(n15197), .A4(n15196), .ZN(
        n15210) );
  AOI22_X1 U19347 ( .A1(n20593), .A2(\xmem_data[48][3] ), .B1(n30898), .B2(
        \xmem_data[49][3] ), .ZN(n15203) );
  AOI22_X1 U19348 ( .A1(n3302), .A2(\xmem_data[50][3] ), .B1(n30599), .B2(
        \xmem_data[51][3] ), .ZN(n15202) );
  AOI22_X1 U19349 ( .A1(n24572), .A2(\xmem_data[52][3] ), .B1(n28979), .B2(
        \xmem_data[53][3] ), .ZN(n15201) );
  AOI22_X1 U19350 ( .A1(n30901), .A2(\xmem_data[54][3] ), .B1(n30900), .B2(
        \xmem_data[55][3] ), .ZN(n15200) );
  NAND4_X1 U19351 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        n15209) );
  AOI22_X1 U19352 ( .A1(n30909), .A2(\xmem_data[56][3] ), .B1(n30908), .B2(
        \xmem_data[57][3] ), .ZN(n15207) );
  AOI22_X1 U19353 ( .A1(n3352), .A2(\xmem_data[58][3] ), .B1(n25360), .B2(
        \xmem_data[59][3] ), .ZN(n15206) );
  AOI22_X1 U19354 ( .A1(n30906), .A2(\xmem_data[60][3] ), .B1(n3218), .B2(
        \xmem_data[61][3] ), .ZN(n15205) );
  AOI22_X1 U19355 ( .A1(n28733), .A2(\xmem_data[62][3] ), .B1(n29095), .B2(
        \xmem_data[63][3] ), .ZN(n15204) );
  NAND4_X1 U19356 ( .A1(n15207), .A2(n15206), .A3(n15205), .A4(n15204), .ZN(
        n15208) );
  OR4_X1 U19357 ( .A1(n15211), .A2(n15210), .A3(n15209), .A4(n15208), .ZN(
        n15212) );
  NAND2_X1 U19358 ( .A1(n15212), .A2(n30918), .ZN(n15213) );
  XNOR2_X1 U19359 ( .A(n31451), .B(\fmem_data[10][7] ), .ZN(n30417) );
  XOR2_X1 U19360 ( .A(\fmem_data[10][6] ), .B(\fmem_data[10][7] ), .Z(n15217)
         );
  AOI22_X1 U19361 ( .A1(n30883), .A2(\xmem_data[32][4] ), .B1(n30882), .B2(
        \xmem_data[33][4] ), .ZN(n15221) );
  AOI22_X1 U19362 ( .A1(n16973), .A2(\xmem_data[34][4] ), .B1(n29045), .B2(
        \xmem_data[35][4] ), .ZN(n15220) );
  AOI22_X1 U19363 ( .A1(n30885), .A2(\xmem_data[36][4] ), .B1(n30884), .B2(
        \xmem_data[37][4] ), .ZN(n15219) );
  AOI22_X1 U19364 ( .A1(n30886), .A2(\xmem_data[38][4] ), .B1(n27452), .B2(
        \xmem_data[39][4] ), .ZN(n15218) );
  NAND4_X1 U19365 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        n15237) );
  AOI22_X1 U19366 ( .A1(n25710), .A2(\xmem_data[40][4] ), .B1(n22741), .B2(
        \xmem_data[41][4] ), .ZN(n15225) );
  AOI22_X1 U19367 ( .A1(n27517), .A2(\xmem_data[42][4] ), .B1(n24134), .B2(
        \xmem_data[43][4] ), .ZN(n15224) );
  AOI22_X1 U19368 ( .A1(n24214), .A2(\xmem_data[44][4] ), .B1(n22718), .B2(
        \xmem_data[45][4] ), .ZN(n15223) );
  AOI22_X1 U19369 ( .A1(n30893), .A2(\xmem_data[46][4] ), .B1(n24592), .B2(
        \xmem_data[47][4] ), .ZN(n15222) );
  NAND4_X1 U19370 ( .A1(n15225), .A2(n15224), .A3(n15223), .A4(n15222), .ZN(
        n15236) );
  AOI22_X1 U19371 ( .A1(n30899), .A2(\xmem_data[48][4] ), .B1(n30898), .B2(
        \xmem_data[49][4] ), .ZN(n15229) );
  AOI22_X1 U19372 ( .A1(n3302), .A2(\xmem_data[50][4] ), .B1(n24167), .B2(
        \xmem_data[51][4] ), .ZN(n15228) );
  AOI22_X1 U19373 ( .A1(n24467), .A2(\xmem_data[52][4] ), .B1(n11008), .B2(
        \xmem_data[53][4] ), .ZN(n15227) );
  AOI22_X1 U19374 ( .A1(n30901), .A2(\xmem_data[54][4] ), .B1(n30900), .B2(
        \xmem_data[55][4] ), .ZN(n15226) );
  NAND4_X1 U19375 ( .A1(n15229), .A2(n15228), .A3(n15227), .A4(n15226), .ZN(
        n15235) );
  AOI22_X1 U19376 ( .A1(n30909), .A2(\xmem_data[56][4] ), .B1(n30908), .B2(
        \xmem_data[57][4] ), .ZN(n15233) );
  AOI22_X1 U19377 ( .A1(n3351), .A2(\xmem_data[58][4] ), .B1(n25442), .B2(
        \xmem_data[59][4] ), .ZN(n15232) );
  AOI22_X1 U19378 ( .A1(n30906), .A2(\xmem_data[60][4] ), .B1(n3217), .B2(
        \xmem_data[61][4] ), .ZN(n15231) );
  AOI22_X1 U19379 ( .A1(n29494), .A2(\xmem_data[62][4] ), .B1(n23769), .B2(
        \xmem_data[63][4] ), .ZN(n15230) );
  NAND4_X1 U19380 ( .A1(n15233), .A2(n15232), .A3(n15231), .A4(n15230), .ZN(
        n15234) );
  OR4_X1 U19381 ( .A1(n15237), .A2(n15236), .A3(n15235), .A4(n15234), .ZN(
        n15238) );
  NAND2_X1 U19382 ( .A1(n15238), .A2(n30918), .ZN(n15308) );
  AOI22_X1 U19383 ( .A1(n28083), .A2(\xmem_data[96][4] ), .B1(n27994), .B2(
        \xmem_data[97][4] ), .ZN(n15242) );
  AOI22_X1 U19384 ( .A1(n3129), .A2(\xmem_data[98][4] ), .B1(n27547), .B2(
        \xmem_data[99][4] ), .ZN(n15241) );
  AOI22_X1 U19385 ( .A1(n27551), .A2(\xmem_data[100][4] ), .B1(n27988), .B2(
        \xmem_data[101][4] ), .ZN(n15240) );
  AOI22_X1 U19386 ( .A1(n30943), .A2(\xmem_data[102][4] ), .B1(n13168), .B2(
        \xmem_data[103][4] ), .ZN(n15239) );
  NAND4_X1 U19387 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        n15258) );
  AOI22_X1 U19388 ( .A1(n17041), .A2(\xmem_data[104][4] ), .B1(n14999), .B2(
        \xmem_data[105][4] ), .ZN(n15246) );
  AOI22_X1 U19389 ( .A1(n31328), .A2(\xmem_data[106][4] ), .B1(n13188), .B2(
        \xmem_data[107][4] ), .ZN(n15245) );
  AOI22_X1 U19390 ( .A1(n30949), .A2(\xmem_data[108][4] ), .B1(n25398), .B2(
        \xmem_data[109][4] ), .ZN(n15244) );
  AOI22_X1 U19391 ( .A1(n30950), .A2(\xmem_data[110][4] ), .B1(n29190), .B2(
        \xmem_data[111][4] ), .ZN(n15243) );
  NAND4_X1 U19392 ( .A1(n15246), .A2(n15245), .A3(n15244), .A4(n15243), .ZN(
        n15257) );
  AOI22_X1 U19393 ( .A1(n30956), .A2(\xmem_data[112][4] ), .B1(n30955), .B2(
        \xmem_data[113][4] ), .ZN(n15250) );
  AOI22_X1 U19394 ( .A1(n28461), .A2(\xmem_data[114][4] ), .B1(n22685), .B2(
        \xmem_data[115][4] ), .ZN(n15249) );
  AOI22_X1 U19395 ( .A1(n24685), .A2(\xmem_data[116][4] ), .B1(n31256), .B2(
        \xmem_data[117][4] ), .ZN(n15248) );
  AOI22_X1 U19396 ( .A1(n20770), .A2(\xmem_data[118][4] ), .B1(n21059), .B2(
        \xmem_data[119][4] ), .ZN(n15247) );
  NAND4_X1 U19397 ( .A1(n15250), .A2(n15249), .A3(n15248), .A4(n15247), .ZN(
        n15256) );
  AOI22_X1 U19398 ( .A1(n27564), .A2(\xmem_data[120][4] ), .B1(n28366), .B2(
        \xmem_data[121][4] ), .ZN(n15254) );
  AOI22_X1 U19399 ( .A1(n3332), .A2(\xmem_data[122][4] ), .B1(n28501), .B2(
        \xmem_data[123][4] ), .ZN(n15253) );
  AOI22_X1 U19400 ( .A1(n30962), .A2(\xmem_data[124][4] ), .B1(n3218), .B2(
        \xmem_data[125][4] ), .ZN(n15252) );
  AOI22_X1 U19401 ( .A1(n30964), .A2(\xmem_data[126][4] ), .B1(n30963), .B2(
        \xmem_data[127][4] ), .ZN(n15251) );
  NAND4_X1 U19402 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15255) );
  OR4_X1 U19403 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15259) );
  NAND2_X1 U19404 ( .A1(n15259), .A2(n30976), .ZN(n15307) );
  AOI22_X1 U19405 ( .A1(n30883), .A2(\xmem_data[64][4] ), .B1(n30882), .B2(
        \xmem_data[65][4] ), .ZN(n15263) );
  AOI22_X1 U19406 ( .A1(n24702), .A2(\xmem_data[66][4] ), .B1(n28343), .B2(
        \xmem_data[67][4] ), .ZN(n15262) );
  AOI22_X1 U19407 ( .A1(n30885), .A2(\xmem_data[68][4] ), .B1(n30884), .B2(
        \xmem_data[69][4] ), .ZN(n15261) );
  AOI22_X1 U19408 ( .A1(n30886), .A2(\xmem_data[70][4] ), .B1(n14998), .B2(
        \xmem_data[71][4] ), .ZN(n15260) );
  NAND4_X1 U19409 ( .A1(n15263), .A2(n15262), .A3(n15261), .A4(n15260), .ZN(
        n15280) );
  AOI22_X1 U19410 ( .A1(n30891), .A2(\xmem_data[72][4] ), .B1(n24160), .B2(
        \xmem_data[73][4] ), .ZN(n15267) );
  AOI22_X1 U19411 ( .A1(n29315), .A2(\xmem_data[74][4] ), .B1(n20586), .B2(
        \xmem_data[75][4] ), .ZN(n15266) );
  AOI22_X1 U19412 ( .A1(n23717), .A2(\xmem_data[76][4] ), .B1(n21006), .B2(
        \xmem_data[77][4] ), .ZN(n15265) );
  AOI22_X1 U19413 ( .A1(n30893), .A2(\xmem_data[78][4] ), .B1(n24592), .B2(
        \xmem_data[79][4] ), .ZN(n15264) );
  NAND4_X1 U19414 ( .A1(n15267), .A2(n15266), .A3(n15265), .A4(n15264), .ZN(
        n15279) );
  AOI22_X1 U19415 ( .A1(n25717), .A2(\xmem_data[80][4] ), .B1(n30898), .B2(
        \xmem_data[81][4] ), .ZN(n15272) );
  AOI22_X1 U19416 ( .A1(n3302), .A2(\xmem_data[82][4] ), .B1(n24521), .B2(
        \xmem_data[83][4] ), .ZN(n15271) );
  AOI22_X1 U19417 ( .A1(n25526), .A2(\xmem_data[84][4] ), .B1(n11008), .B2(
        \xmem_data[85][4] ), .ZN(n15270) );
  AND2_X1 U19418 ( .A1(n30900), .A2(\xmem_data[87][4] ), .ZN(n15268) );
  AOI21_X1 U19419 ( .B1(n30901), .B2(\xmem_data[86][4] ), .A(n15268), .ZN(
        n15269) );
  NAND4_X1 U19420 ( .A1(n15272), .A2(n15271), .A3(n15270), .A4(n15269), .ZN(
        n15278) );
  AOI22_X1 U19421 ( .A1(n30906), .A2(\xmem_data[92][4] ), .B1(n3218), .B2(
        \xmem_data[93][4] ), .ZN(n15276) );
  AOI22_X1 U19422 ( .A1(n3350), .A2(\xmem_data[90][4] ), .B1(n28501), .B2(
        \xmem_data[91][4] ), .ZN(n15275) );
  AOI22_X1 U19423 ( .A1(n30909), .A2(\xmem_data[88][4] ), .B1(n30908), .B2(
        \xmem_data[89][4] ), .ZN(n15274) );
  AOI22_X1 U19424 ( .A1(n24563), .A2(\xmem_data[94][4] ), .B1(n28319), .B2(
        \xmem_data[95][4] ), .ZN(n15273) );
  NAND4_X1 U19425 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15277) );
  OR4_X1 U19426 ( .A1(n15280), .A2(n15279), .A3(n15278), .A4(n15277), .ZN(
        n15281) );
  NAND2_X1 U19427 ( .A1(n15281), .A2(n30974), .ZN(n15306) );
  AOI22_X1 U19428 ( .A1(n30614), .A2(\xmem_data[8][4] ), .B1(n22703), .B2(
        \xmem_data[9][4] ), .ZN(n15285) );
  AOI22_X1 U19429 ( .A1(n27455), .A2(\xmem_data[10][4] ), .B1(n3208), .B2(
        \xmem_data[11][4] ), .ZN(n15284) );
  AOI22_X1 U19430 ( .A1(n29317), .A2(\xmem_data[12][4] ), .B1(n30544), .B2(
        \xmem_data[13][4] ), .ZN(n15283) );
  AOI22_X1 U19431 ( .A1(n30872), .A2(\xmem_data[14][4] ), .B1(n30871), .B2(
        \xmem_data[15][4] ), .ZN(n15282) );
  NAND4_X1 U19432 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15291) );
  AOI22_X1 U19433 ( .A1(n30862), .A2(\xmem_data[24][4] ), .B1(n30861), .B2(
        \xmem_data[25][4] ), .ZN(n15289) );
  AOI22_X1 U19434 ( .A1(n30864), .A2(\xmem_data[26][4] ), .B1(n30863), .B2(
        \xmem_data[27][4] ), .ZN(n15288) );
  AOI22_X1 U19435 ( .A1(n25692), .A2(\xmem_data[28][4] ), .B1(n3220), .B2(
        \xmem_data[29][4] ), .ZN(n15287) );
  AOI22_X1 U19436 ( .A1(n21067), .A2(\xmem_data[30][4] ), .B1(n23769), .B2(
        \xmem_data[31][4] ), .ZN(n15286) );
  NAND4_X1 U19437 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15290) );
  OR2_X1 U19438 ( .A1(n15291), .A2(n15290), .ZN(n15304) );
  AOI22_X1 U19439 ( .A1(n30849), .A2(\xmem_data[16][4] ), .B1(n27856), .B2(
        \xmem_data[17][4] ), .ZN(n15295) );
  AOI22_X1 U19440 ( .A1(n23724), .A2(\xmem_data[18][4] ), .B1(n14975), .B2(
        \xmem_data[19][4] ), .ZN(n15294) );
  AOI22_X1 U19441 ( .A1(n21058), .A2(\xmem_data[20][4] ), .B1(n27463), .B2(
        \xmem_data[21][4] ), .ZN(n15293) );
  AOI22_X1 U19442 ( .A1(n25684), .A2(\xmem_data[22][4] ), .B1(n31344), .B2(
        \xmem_data[23][4] ), .ZN(n15292) );
  NAND4_X1 U19443 ( .A1(n15295), .A2(n15294), .A3(n15293), .A4(n15292), .ZN(
        n15302) );
  AOI22_X1 U19444 ( .A1(n24157), .A2(\xmem_data[6][4] ), .B1(n13168), .B2(
        \xmem_data[7][4] ), .ZN(n15298) );
  AOI22_X1 U19445 ( .A1(n23813), .A2(\xmem_data[4][4] ), .B1(n30854), .B2(
        \xmem_data[5][4] ), .ZN(n15297) );
  AOI22_X1 U19446 ( .A1(n24697), .A2(\xmem_data[0][4] ), .B1(n13444), .B2(
        \xmem_data[1][4] ), .ZN(n15296) );
  NAND3_X1 U19447 ( .A1(n15298), .A2(n15297), .A3(n15296), .ZN(n15301) );
  AND2_X1 U19448 ( .A1(n3126), .A2(\xmem_data[2][4] ), .ZN(n15299) );
  AOI22_X1 U19449 ( .A1(n3222), .A2(\xmem_data[16][5] ), .B1(n29431), .B2(
        \xmem_data[17][5] ), .ZN(n15313) );
  AOI22_X1 U19450 ( .A1(n24140), .A2(\xmem_data[20][5] ), .B1(n28344), .B2(
        \xmem_data[21][5] ), .ZN(n15309) );
  AOI22_X1 U19451 ( .A1(n29255), .A2(\xmem_data[18][5] ), .B1(n3340), .B2(
        \xmem_data[19][5] ), .ZN(n15311) );
  NAND2_X1 U19452 ( .A1(n25422), .A2(\xmem_data[23][5] ), .ZN(n15310) );
  NAND2_X1 U19453 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  AOI22_X1 U19454 ( .A1(n28415), .A2(\xmem_data[24][5] ), .B1(n29451), .B2(
        \xmem_data[25][5] ), .ZN(n15317) );
  AOI22_X1 U19455 ( .A1(n28416), .A2(\xmem_data[26][5] ), .B1(n17041), .B2(
        \xmem_data[27][5] ), .ZN(n15316) );
  AOI22_X1 U19456 ( .A1(n30613), .A2(\xmem_data[28][5] ), .B1(n17018), .B2(
        \xmem_data[29][5] ), .ZN(n15315) );
  AOI22_X1 U19457 ( .A1(n3208), .A2(\xmem_data[30][5] ), .B1(n20542), .B2(
        \xmem_data[31][5] ), .ZN(n15314) );
  NAND4_X1 U19458 ( .A1(n15317), .A2(n15316), .A3(n15315), .A4(n15314), .ZN(
        n15318) );
  OR2_X1 U19459 ( .A1(n15319), .A2(n15318), .ZN(n15334) );
  AOI22_X1 U19460 ( .A1(n27437), .A2(\xmem_data[14][5] ), .B1(n30592), .B2(
        \xmem_data[15][5] ), .ZN(n15320) );
  INV_X1 U19461 ( .A(n15320), .ZN(n15333) );
  AOI22_X1 U19462 ( .A1(n3203), .A2(\xmem_data[12][5] ), .B1(n29661), .B2(
        \xmem_data[13][5] ), .ZN(n15323) );
  AND2_X1 U19463 ( .A1(n27526), .A2(\xmem_data[8][5] ), .ZN(n15321) );
  AOI21_X1 U19464 ( .B1(n30257), .B2(\xmem_data[9][5] ), .A(n15321), .ZN(
        n15322) );
  NAND2_X1 U19465 ( .A1(n15323), .A2(n15322), .ZN(n15331) );
  AOI22_X1 U19466 ( .A1(n28427), .A2(\xmem_data[0][5] ), .B1(n28687), .B2(
        \xmem_data[1][5] ), .ZN(n15327) );
  AOI22_X1 U19467 ( .A1(n27523), .A2(\xmem_data[2][5] ), .B1(n28428), .B2(
        \xmem_data[3][5] ), .ZN(n15326) );
  AOI22_X1 U19468 ( .A1(n21051), .A2(\xmem_data[4][5] ), .B1(n3330), .B2(
        \xmem_data[5][5] ), .ZN(n15325) );
  AOI22_X1 U19469 ( .A1(n28098), .A2(\xmem_data[6][5] ), .B1(n3171), .B2(
        \xmem_data[7][5] ), .ZN(n15324) );
  NAND4_X1 U19470 ( .A1(n15327), .A2(n15326), .A3(n15325), .A4(n15324), .ZN(
        n15330) );
  AOI22_X1 U19471 ( .A1(n25388), .A2(\xmem_data[10][5] ), .B1(n25358), .B2(
        \xmem_data[11][5] ), .ZN(n15328) );
  INV_X1 U19472 ( .A(n15328), .ZN(n15329) );
  OR3_X1 U19473 ( .A1(n15331), .A2(n15330), .A3(n15329), .ZN(n15332) );
  NOR3_X1 U19474 ( .A1(n15334), .A2(n15333), .A3(n15332), .ZN(n15336) );
  NAND2_X1 U19475 ( .A1(n25492), .A2(\xmem_data[22][5] ), .ZN(n15335) );
  AOI21_X1 U19476 ( .B1(n15336), .B2(n15335), .A(n15043), .ZN(n15337) );
  INV_X1 U19477 ( .A(n15337), .ZN(n15403) );
  AOI22_X1 U19478 ( .A1(n28492), .A2(\xmem_data[96][5] ), .B1(n25678), .B2(
        \xmem_data[97][5] ), .ZN(n15341) );
  AOI22_X1 U19479 ( .A1(n30616), .A2(\xmem_data[98][5] ), .B1(n28493), .B2(
        \xmem_data[99][5] ), .ZN(n15340) );
  AOI22_X1 U19480 ( .A1(n28494), .A2(\xmem_data[100][5] ), .B1(n31315), .B2(
        \xmem_data[101][5] ), .ZN(n15339) );
  AOI22_X1 U19481 ( .A1(n28495), .A2(\xmem_data[102][5] ), .B1(n28293), .B2(
        \xmem_data[103][5] ), .ZN(n15338) );
  NAND4_X1 U19482 ( .A1(n15341), .A2(n15340), .A3(n15339), .A4(n15338), .ZN(
        n15357) );
  AOI22_X1 U19483 ( .A1(n28500), .A2(\xmem_data[104][5] ), .B1(n28036), .B2(
        \xmem_data[105][5] ), .ZN(n15345) );
  AOI22_X1 U19484 ( .A1(n24468), .A2(\xmem_data[106][5] ), .B1(n17030), .B2(
        \xmem_data[107][5] ), .ZN(n15344) );
  AOI22_X1 U19485 ( .A1(n27499), .A2(\xmem_data[108][5] ), .B1(n3142), .B2(
        \xmem_data[109][5] ), .ZN(n15343) );
  AOI22_X1 U19486 ( .A1(n28501), .A2(\xmem_data[110][5] ), .B1(n28503), .B2(
        \xmem_data[111][5] ), .ZN(n15342) );
  NAND4_X1 U19487 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15356) );
  AOI22_X1 U19488 ( .A1(n3219), .A2(\xmem_data[112][5] ), .B1(n27445), .B2(
        \xmem_data[113][5] ), .ZN(n15349) );
  AOI22_X1 U19489 ( .A1(n28508), .A2(\xmem_data[114][5] ), .B1(n3342), .B2(
        \xmem_data[115][5] ), .ZN(n15348) );
  AOI22_X1 U19490 ( .A1(n28509), .A2(\xmem_data[116][5] ), .B1(n30710), .B2(
        \xmem_data[117][5] ), .ZN(n15347) );
  AOI22_X1 U19491 ( .A1(n25450), .A2(\xmem_data[118][5] ), .B1(n28374), .B2(
        \xmem_data[119][5] ), .ZN(n15346) );
  NAND4_X1 U19492 ( .A1(n15349), .A2(n15348), .A3(n15347), .A4(n15346), .ZN(
        n15355) );
  AOI22_X1 U19493 ( .A1(n14933), .A2(\xmem_data[120][5] ), .B1(n29451), .B2(
        \xmem_data[121][5] ), .ZN(n15353) );
  AOI22_X1 U19494 ( .A1(n28515), .A2(\xmem_data[122][5] ), .B1(n28334), .B2(
        \xmem_data[123][5] ), .ZN(n15352) );
  AOI22_X1 U19495 ( .A1(n28517), .A2(\xmem_data[124][5] ), .B1(n24213), .B2(
        \xmem_data[125][5] ), .ZN(n15351) );
  AOI22_X1 U19496 ( .A1(n27864), .A2(\xmem_data[126][5] ), .B1(n20800), .B2(
        \xmem_data[127][5] ), .ZN(n15350) );
  NAND4_X1 U19497 ( .A1(n15353), .A2(n15352), .A3(n15351), .A4(n15350), .ZN(
        n15354) );
  OR4_X1 U19498 ( .A1(n15357), .A2(n15356), .A3(n15355), .A4(n15354), .ZN(
        n15379) );
  AOI22_X1 U19499 ( .A1(n29048), .A2(\xmem_data[64][5] ), .B1(n30309), .B2(
        \xmem_data[65][5] ), .ZN(n15361) );
  AOI22_X1 U19500 ( .A1(n24592), .A2(\xmem_data[66][5] ), .B1(n29100), .B2(
        \xmem_data[67][5] ), .ZN(n15360) );
  AOI22_X1 U19501 ( .A1(n28462), .A2(\xmem_data[68][5] ), .B1(n28461), .B2(
        \xmem_data[69][5] ), .ZN(n15359) );
  AOI22_X1 U19502 ( .A1(n28062), .A2(\xmem_data[70][5] ), .B1(n29151), .B2(
        \xmem_data[71][5] ), .ZN(n15358) );
  NAND4_X1 U19503 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15377) );
  AOI22_X1 U19504 ( .A1(n28468), .A2(\xmem_data[72][5] ), .B1(n28467), .B2(
        \xmem_data[73][5] ), .ZN(n15365) );
  AOI22_X1 U19505 ( .A1(n20951), .A2(\xmem_data[74][5] ), .B1(n20986), .B2(
        \xmem_data[75][5] ), .ZN(n15364) );
  AOI22_X1 U19506 ( .A1(n30908), .A2(\xmem_data[76][5] ), .B1(n24630), .B2(
        \xmem_data[77][5] ), .ZN(n15363) );
  AOI22_X1 U19507 ( .A1(n29173), .A2(\xmem_data[78][5] ), .B1(n28470), .B2(
        \xmem_data[79][5] ), .ZN(n15362) );
  NAND4_X1 U19508 ( .A1(n15365), .A2(n15364), .A3(n15363), .A4(n15362), .ZN(
        n15376) );
  AOI22_X1 U19509 ( .A1(n3218), .A2(\xmem_data[80][5] ), .B1(n31368), .B2(
        \xmem_data[81][5] ), .ZN(n15369) );
  AOI22_X1 U19510 ( .A1(n28476), .A2(\xmem_data[82][5] ), .B1(n28475), .B2(
        \xmem_data[83][5] ), .ZN(n15368) );
  AOI22_X1 U19511 ( .A1(n17061), .A2(\xmem_data[84][5] ), .B1(n3374), .B2(
        \xmem_data[85][5] ), .ZN(n15367) );
  AOI22_X1 U19512 ( .A1(n29306), .A2(\xmem_data[86][5] ), .B1(n25422), .B2(
        \xmem_data[87][5] ), .ZN(n15366) );
  NAND4_X1 U19513 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15375) );
  AOI22_X1 U19514 ( .A1(n28481), .A2(\xmem_data[88][5] ), .B1(n27453), .B2(
        \xmem_data[89][5] ), .ZN(n15373) );
  AOI22_X1 U19515 ( .A1(n24212), .A2(\xmem_data[90][5] ), .B1(n25425), .B2(
        \xmem_data[91][5] ), .ZN(n15372) );
  AOI22_X1 U19516 ( .A1(n25709), .A2(\xmem_data[92][5] ), .B1(n31354), .B2(
        \xmem_data[93][5] ), .ZN(n15371) );
  AOI22_X1 U19517 ( .A1(n24134), .A2(\xmem_data[94][5] ), .B1(n17020), .B2(
        \xmem_data[95][5] ), .ZN(n15370) );
  NAND4_X1 U19518 ( .A1(n15373), .A2(n15372), .A3(n15371), .A4(n15370), .ZN(
        n15374) );
  OR4_X1 U19519 ( .A1(n15377), .A2(n15376), .A3(n15375), .A4(n15374), .ZN(
        n15378) );
  AOI22_X1 U19520 ( .A1(n28458), .A2(n15379), .B1(n28526), .B2(n15378), .ZN(
        n15402) );
  AOI22_X1 U19521 ( .A1(n13415), .A2(\xmem_data[32][5] ), .B1(n28754), .B2(
        \xmem_data[33][5] ), .ZN(n15383) );
  AOI22_X1 U19522 ( .A1(n29190), .A2(\xmem_data[34][5] ), .B1(n24220), .B2(
        \xmem_data[35][5] ), .ZN(n15382) );
  AOI22_X1 U19523 ( .A1(n28462), .A2(\xmem_data[36][5] ), .B1(n28461), .B2(
        \xmem_data[37][5] ), .ZN(n15381) );
  AOI22_X1 U19524 ( .A1(n14975), .A2(\xmem_data[38][5] ), .B1(n25582), .B2(
        \xmem_data[39][5] ), .ZN(n15380) );
  NAND4_X1 U19525 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15399) );
  AOI22_X1 U19526 ( .A1(n28468), .A2(\xmem_data[40][5] ), .B1(n28467), .B2(
        \xmem_data[41][5] ), .ZN(n15387) );
  AOI22_X1 U19527 ( .A1(n27567), .A2(\xmem_data[42][5] ), .B1(n25408), .B2(
        \xmem_data[43][5] ), .ZN(n15386) );
  AOI22_X1 U19528 ( .A1(n24470), .A2(\xmem_data[44][5] ), .B1(n3413), .B2(
        \xmem_data[45][5] ), .ZN(n15385) );
  AOI22_X1 U19529 ( .A1(n27501), .A2(\xmem_data[46][5] ), .B1(n28470), .B2(
        \xmem_data[47][5] ), .ZN(n15384) );
  NAND4_X1 U19530 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15398) );
  AOI22_X1 U19531 ( .A1(n3222), .A2(\xmem_data[48][5] ), .B1(n29422), .B2(
        \xmem_data[49][5] ), .ZN(n15391) );
  AOI22_X1 U19532 ( .A1(n28476), .A2(\xmem_data[50][5] ), .B1(n28475), .B2(
        \xmem_data[51][5] ), .ZN(n15390) );
  AOI22_X1 U19533 ( .A1(n24633), .A2(\xmem_data[52][5] ), .B1(n30710), .B2(
        \xmem_data[53][5] ), .ZN(n15389) );
  AOI22_X1 U19534 ( .A1(n29306), .A2(\xmem_data[54][5] ), .B1(n28050), .B2(
        \xmem_data[55][5] ), .ZN(n15388) );
  NAND4_X1 U19535 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n15397) );
  AOI22_X1 U19536 ( .A1(n28481), .A2(\xmem_data[56][5] ), .B1(n25424), .B2(
        \xmem_data[57][5] ), .ZN(n15395) );
  AOI22_X1 U19537 ( .A1(n17012), .A2(\xmem_data[58][5] ), .B1(n28334), .B2(
        \xmem_data[59][5] ), .ZN(n15394) );
  AOI22_X1 U19538 ( .A1(n20717), .A2(\xmem_data[60][5] ), .B1(n30303), .B2(
        \xmem_data[61][5] ), .ZN(n15393) );
  AOI22_X1 U19539 ( .A1(n29162), .A2(\xmem_data[62][5] ), .B1(n20800), .B2(
        \xmem_data[63][5] ), .ZN(n15392) );
  NAND4_X1 U19540 ( .A1(n15395), .A2(n15394), .A3(n15393), .A4(n15392), .ZN(
        n15396) );
  OR4_X1 U19541 ( .A1(n15399), .A2(n15398), .A3(n15397), .A4(n15396), .ZN(
        n15400) );
  NAND2_X1 U19542 ( .A1(n15400), .A2(n28490), .ZN(n15401) );
  XOR2_X1 U19543 ( .A(\fmem_data[29][4] ), .B(\fmem_data[29][5] ), .Z(n15404)
         );
  AOI22_X1 U19544 ( .A1(n28058), .A2(\xmem_data[32][6] ), .B1(n29012), .B2(
        \xmem_data[33][6] ), .ZN(n15408) );
  AOI22_X1 U19545 ( .A1(n20941), .A2(\xmem_data[34][6] ), .B1(n24220), .B2(
        \xmem_data[35][6] ), .ZN(n15407) );
  AOI22_X1 U19546 ( .A1(n28462), .A2(\xmem_data[36][6] ), .B1(n28461), .B2(
        \xmem_data[37][6] ), .ZN(n15406) );
  AOI22_X1 U19547 ( .A1(n31362), .A2(\xmem_data[38][6] ), .B1(n29325), .B2(
        \xmem_data[39][6] ), .ZN(n15405) );
  NAND4_X1 U19548 ( .A1(n15408), .A2(n15407), .A3(n15406), .A4(n15405), .ZN(
        n15424) );
  AOI22_X1 U19549 ( .A1(n28468), .A2(\xmem_data[40][6] ), .B1(n28467), .B2(
        \xmem_data[41][6] ), .ZN(n15412) );
  AOI22_X1 U19550 ( .A1(n27567), .A2(\xmem_data[42][6] ), .B1(n30862), .B2(
        \xmem_data[43][6] ), .ZN(n15411) );
  AOI22_X1 U19551 ( .A1(n20709), .A2(\xmem_data[44][6] ), .B1(n3318), .B2(
        \xmem_data[45][6] ), .ZN(n15410) );
  AOI22_X1 U19552 ( .A1(n25485), .A2(\xmem_data[46][6] ), .B1(n28470), .B2(
        \xmem_data[47][6] ), .ZN(n15409) );
  NAND4_X1 U19553 ( .A1(n15412), .A2(n15411), .A3(n15410), .A4(n15409), .ZN(
        n15423) );
  AOI22_X1 U19554 ( .A1(n3221), .A2(\xmem_data[48][6] ), .B1(n30964), .B2(
        \xmem_data[49][6] ), .ZN(n15416) );
  AOI22_X1 U19555 ( .A1(n28476), .A2(\xmem_data[50][6] ), .B1(n28475), .B2(
        \xmem_data[51][6] ), .ZN(n15415) );
  AOI22_X1 U19556 ( .A1(n17061), .A2(\xmem_data[52][6] ), .B1(n3281), .B2(
        \xmem_data[53][6] ), .ZN(n15414) );
  AOI22_X1 U19557 ( .A1(n3231), .A2(\xmem_data[54][6] ), .B1(n25422), .B2(
        \xmem_data[55][6] ), .ZN(n15413) );
  NAND4_X1 U19558 ( .A1(n15416), .A2(n15415), .A3(n15414), .A4(n15413), .ZN(
        n15422) );
  AOI22_X1 U19559 ( .A1(n28481), .A2(\xmem_data[56][6] ), .B1(n20799), .B2(
        \xmem_data[57][6] ), .ZN(n15420) );
  AOI22_X1 U19560 ( .A1(n31326), .A2(\xmem_data[58][6] ), .B1(n3176), .B2(
        \xmem_data[59][6] ), .ZN(n15419) );
  AOI22_X1 U19561 ( .A1(n30513), .A2(\xmem_data[60][6] ), .B1(n28154), .B2(
        \xmem_data[61][6] ), .ZN(n15418) );
  AOI22_X1 U19562 ( .A1(n22677), .A2(\xmem_data[62][6] ), .B1(n24214), .B2(
        \xmem_data[63][6] ), .ZN(n15417) );
  NAND4_X1 U19563 ( .A1(n15420), .A2(n15419), .A3(n15418), .A4(n15417), .ZN(
        n15421) );
  OR4_X1 U19564 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15451) );
  NAND2_X1 U19565 ( .A1(n25450), .A2(\xmem_data[22][6] ), .ZN(n15449) );
  AOI22_X1 U19566 ( .A1(n28500), .A2(\xmem_data[8][6] ), .B1(n29820), .B2(
        \xmem_data[9][6] ), .ZN(n15428) );
  AOI22_X1 U19567 ( .A1(n20579), .A2(\xmem_data[10][6] ), .B1(n30862), .B2(
        \xmem_data[11][6] ), .ZN(n15427) );
  AOI22_X1 U19568 ( .A1(n31346), .A2(\xmem_data[12][6] ), .B1(n29661), .B2(
        \xmem_data[13][6] ), .ZN(n15426) );
  AOI22_X1 U19569 ( .A1(n31347), .A2(\xmem_data[14][6] ), .B1(n27902), .B2(
        \xmem_data[15][6] ), .ZN(n15425) );
  NAND4_X1 U19570 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15447) );
  AOI22_X1 U19571 ( .A1(n25481), .A2(\xmem_data[24][6] ), .B1(n30744), .B2(
        \xmem_data[25][6] ), .ZN(n15432) );
  AOI22_X1 U19572 ( .A1(n28416), .A2(\xmem_data[26][6] ), .B1(n24131), .B2(
        \xmem_data[27][6] ), .ZN(n15431) );
  AOI22_X1 U19573 ( .A1(n22674), .A2(\xmem_data[28][6] ), .B1(n3158), .B2(
        \xmem_data[29][6] ), .ZN(n15430) );
  AOI22_X1 U19574 ( .A1(n27989), .A2(\xmem_data[30][6] ), .B1(n24593), .B2(
        \xmem_data[31][6] ), .ZN(n15429) );
  NAND4_X1 U19575 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15446) );
  AOI22_X1 U19576 ( .A1(n29181), .A2(\xmem_data[20][6] ), .B1(n3345), .B2(
        \xmem_data[21][6] ), .ZN(n15439) );
  AOI22_X1 U19577 ( .A1(n3218), .A2(\xmem_data[16][6] ), .B1(n29288), .B2(
        \xmem_data[17][6] ), .ZN(n15433) );
  INV_X1 U19578 ( .A(n15433), .ZN(n15437) );
  AOI22_X1 U19579 ( .A1(n20500), .A2(\xmem_data[18][6] ), .B1(n14990), .B2(
        \xmem_data[19][6] ), .ZN(n15434) );
  INV_X1 U19580 ( .A(n15434), .ZN(n15436) );
  AND2_X1 U19581 ( .A1(n25422), .A2(\xmem_data[23][6] ), .ZN(n15435) );
  NOR3_X1 U19582 ( .A1(n15437), .A2(n15436), .A3(n15435), .ZN(n15438) );
  NAND2_X1 U19583 ( .A1(n15439), .A2(n15438), .ZN(n15445) );
  AOI22_X1 U19584 ( .A1(n28427), .A2(\xmem_data[0][6] ), .B1(n30872), .B2(
        \xmem_data[1][6] ), .ZN(n15443) );
  AOI22_X1 U19585 ( .A1(n20941), .A2(\xmem_data[2][6] ), .B1(n28428), .B2(
        \xmem_data[3][6] ), .ZN(n15442) );
  AOI22_X1 U19586 ( .A1(n30598), .A2(\xmem_data[4][6] ), .B1(n3302), .B2(
        \xmem_data[5][6] ), .ZN(n15441) );
  AOI22_X1 U19587 ( .A1(n31314), .A2(\xmem_data[6][6] ), .B1(n30525), .B2(
        \xmem_data[7][6] ), .ZN(n15440) );
  NAND4_X1 U19588 ( .A1(n15443), .A2(n15442), .A3(n15441), .A4(n15440), .ZN(
        n15444) );
  NOR4_X1 U19589 ( .A1(n15447), .A2(n15446), .A3(n15445), .A4(n15444), .ZN(
        n15448) );
  AOI21_X1 U19590 ( .B1(n15449), .B2(n15448), .A(n15043), .ZN(n15450) );
  AOI21_X1 U19591 ( .B1(n15451), .B2(n28490), .A(n15450), .ZN(n15496) );
  AOI22_X1 U19592 ( .A1(n28492), .A2(\xmem_data[96][6] ), .B1(n30893), .B2(
        \xmem_data[97][6] ), .ZN(n15455) );
  AOI22_X1 U19593 ( .A1(n27523), .A2(\xmem_data[98][6] ), .B1(n28493), .B2(
        \xmem_data[99][6] ), .ZN(n15454) );
  AOI22_X1 U19594 ( .A1(n28494), .A2(\xmem_data[100][6] ), .B1(n30686), .B2(
        \xmem_data[101][6] ), .ZN(n15453) );
  AOI22_X1 U19595 ( .A1(n28495), .A2(\xmem_data[102][6] ), .B1(n27847), .B2(
        \xmem_data[103][6] ), .ZN(n15452) );
  NAND4_X1 U19596 ( .A1(n15455), .A2(n15454), .A3(n15453), .A4(n15452), .ZN(
        n15471) );
  AOI22_X1 U19597 ( .A1(n28500), .A2(\xmem_data[104][6] ), .B1(n27498), .B2(
        \xmem_data[105][6] ), .ZN(n15459) );
  AOI22_X1 U19598 ( .A1(n25388), .A2(\xmem_data[106][6] ), .B1(n27436), .B2(
        \xmem_data[107][6] ), .ZN(n15458) );
  AOI22_X1 U19599 ( .A1(n29118), .A2(\xmem_data[108][6] ), .B1(n21308), .B2(
        \xmem_data[109][6] ), .ZN(n15457) );
  AOI22_X1 U19600 ( .A1(n28501), .A2(\xmem_data[110][6] ), .B1(n28503), .B2(
        \xmem_data[111][6] ), .ZN(n15456) );
  NAND4_X1 U19601 ( .A1(n15459), .A2(n15458), .A3(n15457), .A4(n15456), .ZN(
        n15470) );
  AOI22_X1 U19602 ( .A1(n3219), .A2(\xmem_data[112][6] ), .B1(n30593), .B2(
        \xmem_data[113][6] ), .ZN(n15463) );
  AOI22_X1 U19603 ( .A1(n28508), .A2(\xmem_data[114][6] ), .B1(n3341), .B2(
        \xmem_data[115][6] ), .ZN(n15462) );
  AOI22_X1 U19604 ( .A1(n28509), .A2(\xmem_data[116][6] ), .B1(n28084), .B2(
        \xmem_data[117][6] ), .ZN(n15461) );
  AOI22_X1 U19605 ( .A1(n3231), .A2(\xmem_data[118][6] ), .B1(n28374), .B2(
        \xmem_data[119][6] ), .ZN(n15460) );
  NAND4_X1 U19606 ( .A1(n15463), .A2(n15462), .A3(n15461), .A4(n15460), .ZN(
        n15469) );
  AOI22_X1 U19607 ( .A1(n28415), .A2(\xmem_data[120][6] ), .B1(n20545), .B2(
        \xmem_data[121][6] ), .ZN(n15467) );
  AOI22_X1 U19608 ( .A1(n28515), .A2(\xmem_data[122][6] ), .B1(n29023), .B2(
        \xmem_data[123][6] ), .ZN(n15466) );
  AOI22_X1 U19609 ( .A1(n28517), .A2(\xmem_data[124][6] ), .B1(n30948), .B2(
        \xmem_data[125][6] ), .ZN(n15465) );
  AOI22_X1 U19610 ( .A1(n30615), .A2(\xmem_data[126][6] ), .B1(n23764), .B2(
        \xmem_data[127][6] ), .ZN(n15464) );
  NAND4_X1 U19611 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15468) );
  OR4_X1 U19612 ( .A1(n15471), .A2(n15470), .A3(n15469), .A4(n15468), .ZN(
        n15494) );
  AOI22_X1 U19613 ( .A1(n25677), .A2(\xmem_data[64][6] ), .B1(n24115), .B2(
        \xmem_data[65][6] ), .ZN(n15475) );
  AOI22_X1 U19614 ( .A1(n30515), .A2(n20682), .B1(n20593), .B2(
        \xmem_data[67][6] ), .ZN(n15474) );
  AOI22_X1 U19615 ( .A1(n28462), .A2(\xmem_data[68][6] ), .B1(n28461), .B2(
        \xmem_data[69][6] ), .ZN(n15473) );
  AOI22_X1 U19616 ( .A1(n24622), .A2(\xmem_data[70][6] ), .B1(n3171), .B2(
        \xmem_data[71][6] ), .ZN(n15472) );
  NAND4_X1 U19617 ( .A1(n15475), .A2(n15474), .A3(n15473), .A4(n15472), .ZN(
        n15492) );
  AOI22_X1 U19618 ( .A1(n28468), .A2(\xmem_data[72][6] ), .B1(n28467), .B2(
        \xmem_data[73][6] ), .ZN(n15480) );
  AOI22_X1 U19619 ( .A1(n20707), .A2(\xmem_data[74][6] ), .B1(n25686), .B2(
        \xmem_data[75][6] ), .ZN(n15479) );
  AOI22_X1 U19620 ( .A1(n27958), .A2(\xmem_data[76][6] ), .B1(n3333), .B2(
        \xmem_data[77][6] ), .ZN(n15478) );
  AND2_X1 U19621 ( .A1(n28501), .A2(\xmem_data[78][6] ), .ZN(n15476) );
  AOI21_X1 U19622 ( .B1(n28470), .B2(\xmem_data[79][6] ), .A(n15476), .ZN(
        n15477) );
  NAND4_X1 U19623 ( .A1(n15480), .A2(n15479), .A3(n15478), .A4(n15477), .ZN(
        n15491) );
  AOI22_X1 U19624 ( .A1(n3218), .A2(\xmem_data[80][6] ), .B1(n25414), .B2(
        \xmem_data[81][6] ), .ZN(n15484) );
  AOI22_X1 U19625 ( .A1(n28476), .A2(\xmem_data[82][6] ), .B1(n28475), .B2(
        \xmem_data[83][6] ), .ZN(n15483) );
  AOI22_X1 U19626 ( .A1(n30882), .A2(\xmem_data[84][6] ), .B1(n24702), .B2(
        \xmem_data[85][6] ), .ZN(n15482) );
  AOI22_X1 U19627 ( .A1(n28045), .A2(\xmem_data[86][6] ), .B1(n23813), .B2(
        \xmem_data[87][6] ), .ZN(n15481) );
  NAND4_X1 U19628 ( .A1(n15484), .A2(n15483), .A3(n15482), .A4(n15481), .ZN(
        n15490) );
  AOI22_X1 U19629 ( .A1(n28481), .A2(\xmem_data[88][6] ), .B1(n29308), .B2(
        \xmem_data[89][6] ), .ZN(n15488) );
  AOI22_X1 U19630 ( .A1(n25605), .A2(\xmem_data[90][6] ), .B1(n28334), .B2(
        \xmem_data[91][6] ), .ZN(n15487) );
  AOI22_X1 U19631 ( .A1(n28090), .A2(\xmem_data[92][6] ), .B1(n23795), .B2(
        \xmem_data[93][6] ), .ZN(n15486) );
  AOI22_X1 U19632 ( .A1(n28993), .A2(\xmem_data[94][6] ), .B1(n24708), .B2(
        \xmem_data[95][6] ), .ZN(n15485) );
  NAND4_X1 U19633 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        n15489) );
  OR4_X1 U19634 ( .A1(n15492), .A2(n15491), .A3(n15490), .A4(n15489), .ZN(
        n15493) );
  AOI22_X1 U19635 ( .A1(n28458), .A2(n15494), .B1(n28526), .B2(n15493), .ZN(
        n15495) );
  XNOR2_X1 U19636 ( .A(n31800), .B(\fmem_data[29][5] ), .ZN(n33131) );
  AOI22_X1 U19637 ( .A1(n29786), .A2(\xmem_data[96][3] ), .B1(n29785), .B2(
        \xmem_data[97][3] ), .ZN(n15500) );
  AOI22_X1 U19638 ( .A1(n29830), .A2(\xmem_data[98][3] ), .B1(n24693), .B2(
        \xmem_data[99][3] ), .ZN(n15499) );
  AOI22_X1 U19639 ( .A1(n27741), .A2(\xmem_data[100][3] ), .B1(n30182), .B2(
        \xmem_data[101][3] ), .ZN(n15498) );
  AOI22_X1 U19640 ( .A1(n29790), .A2(\xmem_data[102][3] ), .B1(n29832), .B2(
        \xmem_data[103][3] ), .ZN(n15497) );
  NAND4_X1 U19641 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15516) );
  AOI22_X1 U19642 ( .A1(n29799), .A2(\xmem_data[104][3] ), .B1(n29629), .B2(
        \xmem_data[105][3] ), .ZN(n15504) );
  AOI22_X1 U19643 ( .A1(n29800), .A2(\xmem_data[106][3] ), .B1(n3375), .B2(
        \xmem_data[107][3] ), .ZN(n15503) );
  AOI22_X1 U19644 ( .A1(n29590), .A2(\xmem_data[108][3] ), .B1(n30662), .B2(
        \xmem_data[109][3] ), .ZN(n15502) );
  AOI22_X1 U19645 ( .A1(n29802), .A2(\xmem_data[110][3] ), .B1(n28233), .B2(
        \xmem_data[111][3] ), .ZN(n15501) );
  NAND4_X1 U19646 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15515) );
  AOI22_X1 U19647 ( .A1(n30745), .A2(\xmem_data[112][3] ), .B1(n30193), .B2(
        \xmem_data[113][3] ), .ZN(n15508) );
  AOI22_X1 U19648 ( .A1(n29771), .A2(\xmem_data[114][3] ), .B1(n29807), .B2(
        \xmem_data[115][3] ), .ZN(n15507) );
  AOI22_X1 U19649 ( .A1(n3165), .A2(\xmem_data[116][3] ), .B1(n3182), .B2(
        \xmem_data[117][3] ), .ZN(n15506) );
  AOI22_X1 U19650 ( .A1(n30715), .A2(\xmem_data[118][3] ), .B1(n24115), .B2(
        \xmem_data[119][3] ), .ZN(n15505) );
  NAND4_X1 U19651 ( .A1(n15508), .A2(n15507), .A3(n15506), .A4(n15505), .ZN(
        n15514) );
  AOI22_X1 U19652 ( .A1(n30198), .A2(\xmem_data[120][3] ), .B1(n29640), .B2(
        \xmem_data[121][3] ), .ZN(n15512) );
  AOI22_X1 U19653 ( .A1(n29817), .A2(\xmem_data[122][3] ), .B1(n29816), .B2(
        \xmem_data[123][3] ), .ZN(n15511) );
  AOI22_X1 U19654 ( .A1(n29819), .A2(\xmem_data[124][3] ), .B1(n29818), .B2(
        \xmem_data[125][3] ), .ZN(n15510) );
  AOI22_X1 U19655 ( .A1(n29821), .A2(\xmem_data[126][3] ), .B1(n29820), .B2(
        \xmem_data[127][3] ), .ZN(n15509) );
  NAND4_X1 U19656 ( .A1(n15512), .A2(n15511), .A3(n15510), .A4(n15509), .ZN(
        n15513) );
  OR4_X1 U19657 ( .A1(n15516), .A2(n15515), .A3(n15514), .A4(n15513), .ZN(
        n15540) );
  AOI22_X1 U19658 ( .A1(n29786), .A2(\xmem_data[64][3] ), .B1(n29785), .B2(
        \xmem_data[65][3] ), .ZN(n15520) );
  AOI22_X1 U19659 ( .A1(n29830), .A2(\xmem_data[66][3] ), .B1(n28677), .B2(
        \xmem_data[67][3] ), .ZN(n15519) );
  AOI22_X1 U19660 ( .A1(n29433), .A2(\xmem_data[68][3] ), .B1(n27013), .B2(
        \xmem_data[69][3] ), .ZN(n15518) );
  AOI22_X1 U19661 ( .A1(n28138), .A2(\xmem_data[70][3] ), .B1(n29832), .B2(
        \xmem_data[71][3] ), .ZN(n15517) );
  NAND4_X1 U19662 ( .A1(n15520), .A2(n15519), .A3(n15518), .A4(n15517), .ZN(
        n15538) );
  AOI22_X1 U19663 ( .A1(n29799), .A2(\xmem_data[72][3] ), .B1(n28208), .B2(
        \xmem_data[73][3] ), .ZN(n15524) );
  AOI22_X1 U19664 ( .A1(n29800), .A2(\xmem_data[74][3] ), .B1(n3375), .B2(
        \xmem_data[75][3] ), .ZN(n15523) );
  AOI22_X1 U19665 ( .A1(n29446), .A2(\xmem_data[76][3] ), .B1(n30662), .B2(
        \xmem_data[77][3] ), .ZN(n15522) );
  AOI22_X1 U19666 ( .A1(n29802), .A2(\xmem_data[78][3] ), .B1(n28089), .B2(
        \xmem_data[79][3] ), .ZN(n15521) );
  NAND4_X1 U19667 ( .A1(n15524), .A2(n15523), .A3(n15522), .A4(n15521), .ZN(
        n15537) );
  AOI22_X1 U19668 ( .A1(n3164), .A2(\xmem_data[84][3] ), .B1(n3188), .B2(
        \xmem_data[85][3] ), .ZN(n15530) );
  BUF_X1 U19669 ( .A(n15525), .Z(n29740) );
  AOI22_X1 U19670 ( .A1(n29740), .A2(\xmem_data[82][3] ), .B1(n29807), .B2(
        \xmem_data[83][3] ), .ZN(n15529) );
  AOI22_X1 U19671 ( .A1(n30302), .A2(\xmem_data[80][3] ), .B1(n30249), .B2(
        \xmem_data[81][3] ), .ZN(n15528) );
  AND2_X1 U19672 ( .A1(n28754), .A2(\xmem_data[87][3] ), .ZN(n15526) );
  AOI21_X1 U19673 ( .B1(n30310), .B2(\xmem_data[86][3] ), .A(n15526), .ZN(
        n15527) );
  NAND4_X1 U19674 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15536) );
  AOI22_X1 U19675 ( .A1(n28173), .A2(\xmem_data[88][3] ), .B1(n29721), .B2(
        \xmem_data[89][3] ), .ZN(n15534) );
  AOI22_X1 U19676 ( .A1(n29817), .A2(\xmem_data[90][3] ), .B1(n29816), .B2(
        \xmem_data[91][3] ), .ZN(n15533) );
  AOI22_X1 U19677 ( .A1(n29819), .A2(\xmem_data[92][3] ), .B1(n29818), .B2(
        \xmem_data[93][3] ), .ZN(n15532) );
  AOI22_X1 U19678 ( .A1(n29821), .A2(\xmem_data[94][3] ), .B1(n29820), .B2(
        \xmem_data[95][3] ), .ZN(n15531) );
  NAND4_X1 U19679 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15535) );
  AOI22_X1 U19680 ( .A1(n29829), .A2(\xmem_data[32][3] ), .B1(n29785), .B2(
        \xmem_data[33][3] ), .ZN(n15544) );
  AOI22_X1 U19681 ( .A1(n29787), .A2(\xmem_data[34][3] ), .B1(n23754), .B2(
        \xmem_data[35][3] ), .ZN(n15543) );
  AOI22_X1 U19682 ( .A1(n29433), .A2(\xmem_data[36][3] ), .B1(n30707), .B2(
        \xmem_data[37][3] ), .ZN(n15542) );
  AOI22_X1 U19683 ( .A1(n3392), .A2(\xmem_data[38][3] ), .B1(n29789), .B2(
        \xmem_data[39][3] ), .ZN(n15541) );
  NAND4_X1 U19684 ( .A1(n15544), .A2(n15543), .A3(n15542), .A4(n15541), .ZN(
        n15561) );
  AOI22_X1 U19685 ( .A1(n27701), .A2(\xmem_data[40][3] ), .B1(n27833), .B2(
        \xmem_data[41][3] ), .ZN(n15548) );
  AOI22_X1 U19686 ( .A1(n29707), .A2(\xmem_data[42][3] ), .B1(n29706), .B2(
        \xmem_data[43][3] ), .ZN(n15547) );
  AOI22_X1 U19687 ( .A1(n30633), .A2(\xmem_data[44][3] ), .B1(n28238), .B2(
        \xmem_data[45][3] ), .ZN(n15546) );
  AOI22_X1 U19688 ( .A1(n29763), .A2(\xmem_data[46][3] ), .B1(n29403), .B2(
        \xmem_data[47][3] ), .ZN(n15545) );
  NAND4_X1 U19689 ( .A1(n15548), .A2(n15547), .A3(n15546), .A4(n15545), .ZN(
        n15560) );
  AOI22_X1 U19690 ( .A1(n29436), .A2(\xmem_data[48][3] ), .B1(n30090), .B2(
        \xmem_data[49][3] ), .ZN(n15553) );
  AOI22_X1 U19691 ( .A1(n29740), .A2(\xmem_data[50][3] ), .B1(n29237), .B2(
        \xmem_data[51][3] ), .ZN(n15552) );
  AOI22_X1 U19692 ( .A1(n3168), .A2(\xmem_data[52][3] ), .B1(n3191), .B2(
        \xmem_data[53][3] ), .ZN(n15551) );
  BUF_X1 U19693 ( .A(n15549), .Z(n29476) );
  AOI22_X1 U19694 ( .A1(n29476), .A2(\xmem_data[54][3] ), .B1(n20730), .B2(
        \xmem_data[55][3] ), .ZN(n15550) );
  NAND4_X1 U19695 ( .A1(n15553), .A2(n15552), .A3(n15551), .A4(n15550), .ZN(
        n15559) );
  AOI22_X1 U19696 ( .A1(n29488), .A2(\xmem_data[56][3] ), .B1(n29721), .B2(
        \xmem_data[57][3] ), .ZN(n15557) );
  AOI22_X1 U19697 ( .A1(n3226), .A2(\xmem_data[58][3] ), .B1(n3151), .B2(
        \xmem_data[59][3] ), .ZN(n15556) );
  AOI22_X1 U19698 ( .A1(n29724), .A2(\xmem_data[60][3] ), .B1(n29723), .B2(
        \xmem_data[61][3] ), .ZN(n15555) );
  AOI22_X1 U19699 ( .A1(n29726), .A2(\xmem_data[62][3] ), .B1(n29725), .B2(
        \xmem_data[63][3] ), .ZN(n15554) );
  NAND4_X1 U19700 ( .A1(n15557), .A2(n15556), .A3(n15555), .A4(n15554), .ZN(
        n15558) );
  OR4_X1 U19701 ( .A1(n15561), .A2(n15560), .A3(n15559), .A4(n15558), .ZN(
        n15583) );
  AOI22_X1 U19702 ( .A1(n29829), .A2(\xmem_data[0][3] ), .B1(n29695), .B2(
        \xmem_data[1][3] ), .ZN(n15565) );
  AOI22_X1 U19703 ( .A1(n29696), .A2(\xmem_data[2][3] ), .B1(n28245), .B2(
        \xmem_data[3][3] ), .ZN(n15564) );
  AOI22_X1 U19704 ( .A1(n29433), .A2(\xmem_data[4][3] ), .B1(n26616), .B2(
        \xmem_data[5][3] ), .ZN(n15563) );
  AOI22_X1 U19705 ( .A1(n28700), .A2(\xmem_data[6][3] ), .B1(n29698), .B2(
        \xmem_data[7][3] ), .ZN(n15562) );
  NAND4_X1 U19706 ( .A1(n15565), .A2(n15564), .A3(n15563), .A4(n15562), .ZN(
        n15581) );
  AOI22_X1 U19707 ( .A1(n30697), .A2(\xmem_data[8][3] ), .B1(n30293), .B2(
        \xmem_data[9][3] ), .ZN(n15569) );
  AOI22_X1 U19708 ( .A1(n29707), .A2(\xmem_data[10][3] ), .B1(n29762), .B2(
        \xmem_data[11][3] ), .ZN(n15568) );
  AOI22_X1 U19709 ( .A1(n30743), .A2(\xmem_data[12][3] ), .B1(n29347), .B2(
        \xmem_data[13][3] ), .ZN(n15567) );
  AOI22_X1 U19710 ( .A1(n29709), .A2(\xmem_data[14][3] ), .B1(n28671), .B2(
        \xmem_data[15][3] ), .ZN(n15566) );
  NAND4_X1 U19711 ( .A1(n15569), .A2(n15568), .A3(n15567), .A4(n15566), .ZN(
        n15580) );
  AOI22_X1 U19712 ( .A1(n28779), .A2(\xmem_data[16][3] ), .B1(n30090), .B2(
        \xmem_data[17][3] ), .ZN(n15573) );
  AOI22_X1 U19713 ( .A1(n29771), .A2(\xmem_data[18][3] ), .B1(n29605), .B2(
        \xmem_data[19][3] ), .ZN(n15572) );
  AOI22_X1 U19714 ( .A1(n3163), .A2(\xmem_data[20][3] ), .B1(n3182), .B2(
        \xmem_data[21][3] ), .ZN(n15571) );
  AOI22_X1 U19715 ( .A1(n30764), .A2(\xmem_data[22][3] ), .B1(n22682), .B2(
        \xmem_data[23][3] ), .ZN(n15570) );
  NAND4_X1 U19716 ( .A1(n15573), .A2(n15572), .A3(n15571), .A4(n15570), .ZN(
        n15579) );
  AOI22_X1 U19717 ( .A1(n29547), .A2(\xmem_data[24][3] ), .B1(n30170), .B2(
        \xmem_data[25][3] ), .ZN(n15577) );
  AOI22_X1 U19718 ( .A1(n3226), .A2(\xmem_data[26][3] ), .B1(n3337), .B2(
        \xmem_data[27][3] ), .ZN(n15576) );
  AOI22_X1 U19719 ( .A1(n29777), .A2(\xmem_data[28][3] ), .B1(n29776), .B2(
        \xmem_data[29][3] ), .ZN(n15575) );
  AOI22_X1 U19720 ( .A1(n28727), .A2(\xmem_data[30][3] ), .B1(n21060), .B2(
        \xmem_data[31][3] ), .ZN(n15574) );
  NAND4_X1 U19721 ( .A1(n15577), .A2(n15576), .A3(n15575), .A4(n15574), .ZN(
        n15578) );
  AOI22_X1 U19722 ( .A1(n29795), .A2(n15583), .B1(n29733), .B2(n15582), .ZN(
        n15584) );
  XNOR2_X1 U19723 ( .A(n3257), .B(\fmem_data[19][7] ), .ZN(n31976) );
  AOI22_X1 U19724 ( .A1(n29786), .A2(\xmem_data[64][2] ), .B1(n29785), .B2(
        \xmem_data[65][2] ), .ZN(n15586) );
  AOI22_X1 U19725 ( .A1(n29602), .A2(\xmem_data[76][2] ), .B1(n3369), .B2(
        \xmem_data[77][2] ), .ZN(n15591) );
  AOI22_X1 U19726 ( .A1(n28779), .A2(\xmem_data[80][2] ), .B1(n30084), .B2(
        \xmem_data[81][2] ), .ZN(n15590) );
  AOI22_X1 U19727 ( .A1(n29830), .A2(\xmem_data[66][2] ), .B1(n24630), .B2(
        \xmem_data[67][2] ), .ZN(n15589) );
  AOI22_X1 U19728 ( .A1(n29802), .A2(\xmem_data[78][2] ), .B1(n28346), .B2(
        \xmem_data[79][2] ), .ZN(n15588) );
  AOI22_X1 U19729 ( .A1(n29800), .A2(\xmem_data[74][2] ), .B1(n3375), .B2(
        \xmem_data[75][2] ), .ZN(n15587) );
  AOI22_X1 U19730 ( .A1(n28138), .A2(\xmem_data[70][2] ), .B1(n29832), .B2(
        \xmem_data[71][2] ), .ZN(n15592) );
  AOI22_X1 U19731 ( .A1(n29363), .A2(\xmem_data[88][2] ), .B1(n30685), .B2(
        \xmem_data[89][2] ), .ZN(n15595) );
  AND2_X1 U19732 ( .A1(n30893), .A2(\xmem_data[87][2] ), .ZN(n15593) );
  AOI21_X1 U19733 ( .B1(n23901), .B2(\xmem_data[86][2] ), .A(n15593), .ZN(
        n15594) );
  NAND3_X1 U19734 ( .A1(n3479), .A2(n15592), .A3(n3552), .ZN(n15607) );
  AOI22_X1 U19735 ( .A1(n29788), .A2(\xmem_data[68][2] ), .B1(n27013), .B2(
        \xmem_data[69][2] ), .ZN(n15605) );
  AOI22_X1 U19736 ( .A1(n3161), .A2(\xmem_data[84][2] ), .B1(n3187), .B2(
        \xmem_data[85][2] ), .ZN(n15596) );
  AOI22_X1 U19737 ( .A1(n29821), .A2(\xmem_data[94][2] ), .B1(n29820), .B2(
        \xmem_data[95][2] ), .ZN(n15599) );
  AOI22_X1 U19738 ( .A1(n29740), .A2(\xmem_data[82][2] ), .B1(n29807), .B2(
        \xmem_data[83][2] ), .ZN(n15598) );
  AOI22_X1 U19739 ( .A1(n29817), .A2(\xmem_data[90][2] ), .B1(n29816), .B2(
        \xmem_data[91][2] ), .ZN(n15597) );
  AOI22_X1 U19740 ( .A1(n29819), .A2(\xmem_data[92][2] ), .B1(n29818), .B2(
        \xmem_data[93][2] ), .ZN(n15600) );
  INV_X1 U19741 ( .A(n15600), .ZN(n15601) );
  NOR2_X1 U19742 ( .A1(n15602), .A2(n15601), .ZN(n15604) );
  AOI22_X1 U19743 ( .A1(n29799), .A2(\xmem_data[72][2] ), .B1(n29708), .B2(
        \xmem_data[73][2] ), .ZN(n15603) );
  NAND4_X1 U19744 ( .A1(n15605), .A2(n15596), .A3(n15604), .A4(n15603), .ZN(
        n15606) );
  OAI21_X1 U19745 ( .B1(n15607), .B2(n15606), .A(n29758), .ZN(n15695) );
  AOI22_X1 U19746 ( .A1(n30248), .A2(\xmem_data[108][2] ), .B1(n29482), .B2(
        \xmem_data[109][2] ), .ZN(n15611) );
  AOI22_X1 U19747 ( .A1(n29800), .A2(\xmem_data[106][2] ), .B1(n29762), .B2(
        \xmem_data[107][2] ), .ZN(n15610) );
  AOI22_X1 U19748 ( .A1(n29799), .A2(\xmem_data[104][2] ), .B1(n28786), .B2(
        \xmem_data[105][2] ), .ZN(n15609) );
  AOI22_X1 U19749 ( .A1(n29802), .A2(\xmem_data[110][2] ), .B1(n27514), .B2(
        \xmem_data[111][2] ), .ZN(n15608) );
  AOI22_X1 U19750 ( .A1(n30766), .A2(\xmem_data[120][2] ), .B1(n30266), .B2(
        \xmem_data[121][2] ), .ZN(n15618) );
  AOI22_X1 U19751 ( .A1(n29777), .A2(\xmem_data[124][2] ), .B1(n29776), .B2(
        \xmem_data[125][2] ), .ZN(n15612) );
  INV_X1 U19752 ( .A(n15612), .ZN(n15616) );
  AOI22_X1 U19753 ( .A1(n29726), .A2(\xmem_data[126][2] ), .B1(n25407), .B2(
        \xmem_data[127][2] ), .ZN(n15614) );
  AOI22_X1 U19754 ( .A1(n29817), .A2(\xmem_data[122][2] ), .B1(n28701), .B2(
        \xmem_data[123][2] ), .ZN(n15613) );
  NAND2_X1 U19755 ( .A1(n15614), .A2(n15613), .ZN(n15615) );
  NOR2_X1 U19756 ( .A1(n15616), .A2(n15615), .ZN(n15617) );
  AOI22_X1 U19757 ( .A1(n28685), .A2(\xmem_data[112][2] ), .B1(n26884), .B2(
        \xmem_data[113][2] ), .ZN(n15619) );
  INV_X1 U19758 ( .A(n15619), .ZN(n15623) );
  AOI22_X1 U19759 ( .A1(n3164), .A2(\xmem_data[116][2] ), .B1(n3182), .B2(
        \xmem_data[117][2] ), .ZN(n15621) );
  AOI22_X1 U19760 ( .A1(n29740), .A2(\xmem_data[114][2] ), .B1(n29807), .B2(
        \xmem_data[115][2] ), .ZN(n15620) );
  NAND2_X1 U19761 ( .A1(n15621), .A2(n15620), .ZN(n15622) );
  NOR2_X1 U19762 ( .A1(n15623), .A2(n15622), .ZN(n15627) );
  NAND2_X1 U19763 ( .A1(n30070), .A2(\xmem_data[118][2] ), .ZN(n15625) );
  NAND2_X1 U19764 ( .A1(n29410), .A2(\xmem_data[119][2] ), .ZN(n15624) );
  NAND4_X1 U19765 ( .A1(n15628), .A2(n3930), .A3(n15627), .A4(n15626), .ZN(
        n15634) );
  AOI22_X1 U19766 ( .A1(n28717), .A2(\xmem_data[96][2] ), .B1(n7691), .B2(
        \xmem_data[97][2] ), .ZN(n15632) );
  AOI22_X1 U19767 ( .A1(n29830), .A2(\xmem_data[98][2] ), .B1(n3414), .B2(
        \xmem_data[99][2] ), .ZN(n15631) );
  AOI22_X1 U19768 ( .A1(n29421), .A2(\xmem_data[100][2] ), .B1(n30654), .B2(
        \xmem_data[101][2] ), .ZN(n15630) );
  AOI22_X1 U19769 ( .A1(n29628), .A2(\xmem_data[102][2] ), .B1(n29832), .B2(
        \xmem_data[103][2] ), .ZN(n15629) );
  NAND4_X1 U19770 ( .A1(n15632), .A2(n15631), .A3(n15630), .A4(n15629), .ZN(
        n15633) );
  OAI21_X1 U19771 ( .B1(n15634), .B2(n15633), .A(n29837), .ZN(n15694) );
  AOI22_X1 U19772 ( .A1(n28739), .A2(\xmem_data[12][2] ), .B1(n29389), .B2(
        \xmem_data[13][2] ), .ZN(n15635) );
  INV_X1 U19773 ( .A(n15635), .ZN(n15651) );
  AOI22_X1 U19774 ( .A1(n29699), .A2(\xmem_data[6][2] ), .B1(n29698), .B2(
        \xmem_data[7][2] ), .ZN(n15637) );
  AOI22_X1 U19775 ( .A1(n27710), .A2(\xmem_data[4][2] ), .B1(n27832), .B2(
        \xmem_data[5][2] ), .ZN(n15636) );
  NAND2_X1 U19776 ( .A1(n15637), .A2(n15636), .ZN(n15650) );
  AOI22_X1 U19777 ( .A1(n30294), .A2(\xmem_data[8][2] ), .B1(n29761), .B2(
        \xmem_data[9][2] ), .ZN(n15648) );
  AOI22_X1 U19778 ( .A1(n28717), .A2(\xmem_data[0][2] ), .B1(n29695), .B2(
        \xmem_data[1][2] ), .ZN(n15638) );
  INV_X1 U19779 ( .A(n15638), .ZN(n15646) );
  NAND2_X1 U19780 ( .A1(n29696), .A2(\xmem_data[2][2] ), .ZN(n15644) );
  NAND2_X1 U19781 ( .A1(n29707), .A2(\xmem_data[10][2] ), .ZN(n15643) );
  NAND2_X1 U19782 ( .A1(n31327), .A2(\xmem_data[15][2] ), .ZN(n15641) );
  NAND2_X1 U19783 ( .A1(n30864), .A2(\xmem_data[3][2] ), .ZN(n15640) );
  NAND2_X1 U19784 ( .A1(n29762), .A2(\xmem_data[11][2] ), .ZN(n15639) );
  NAND2_X1 U19785 ( .A1(n29709), .A2(\xmem_data[14][2] ), .ZN(n15642) );
  NAND4_X1 U19786 ( .A1(n15644), .A2(n15643), .A3(n3935), .A4(n15642), .ZN(
        n15645) );
  NOR2_X1 U19787 ( .A1(n15646), .A2(n15645), .ZN(n15647) );
  NAND2_X1 U19788 ( .A1(n15648), .A2(n15647), .ZN(n15649) );
  AOI22_X1 U19789 ( .A1(n29714), .A2(\xmem_data[16][2] ), .B1(n28778), .B2(
        \xmem_data[17][2] ), .ZN(n15655) );
  AOI22_X1 U19790 ( .A1(n29740), .A2(\xmem_data[18][2] ), .B1(n30543), .B2(
        \xmem_data[19][2] ), .ZN(n15654) );
  AOI22_X1 U19791 ( .A1(n3168), .A2(\xmem_data[20][2] ), .B1(n3191), .B2(
        \xmem_data[21][2] ), .ZN(n15653) );
  AOI22_X1 U19792 ( .A1(n29716), .A2(\xmem_data[22][2] ), .B1(n28232), .B2(
        \xmem_data[23][2] ), .ZN(n15652) );
  AOI22_X1 U19793 ( .A1(n29815), .A2(\xmem_data[24][2] ), .B1(n30685), .B2(
        \xmem_data[25][2] ), .ZN(n15656) );
  INV_X1 U19794 ( .A(n15656), .ZN(n15661) );
  AOI22_X1 U19795 ( .A1(n29724), .A2(\xmem_data[28][2] ), .B1(n29776), .B2(
        \xmem_data[29][2] ), .ZN(n15659) );
  AOI22_X1 U19796 ( .A1(n29726), .A2(\xmem_data[30][2] ), .B1(n17051), .B2(
        \xmem_data[31][2] ), .ZN(n15658) );
  AOI22_X1 U19797 ( .A1(n3226), .A2(\xmem_data[26][2] ), .B1(n30269), .B2(
        \xmem_data[27][2] ), .ZN(n15657) );
  NOR2_X1 U19798 ( .A1(n15661), .A2(n15660), .ZN(n15662) );
  NAND2_X1 U19799 ( .A1(n3816), .A2(n15662), .ZN(n15663) );
  OAI21_X1 U19800 ( .B1(n3919), .B2(n15663), .A(n29733), .ZN(n15693) );
  AOI22_X1 U19801 ( .A1(n29547), .A2(\xmem_data[56][2] ), .B1(n30765), .B2(
        \xmem_data[57][2] ), .ZN(n15670) );
  AOI22_X1 U19802 ( .A1(n29724), .A2(\xmem_data[60][2] ), .B1(n29723), .B2(
        \xmem_data[61][2] ), .ZN(n15664) );
  INV_X1 U19803 ( .A(n15664), .ZN(n15668) );
  AOI22_X1 U19804 ( .A1(n29726), .A2(\xmem_data[62][2] ), .B1(n29725), .B2(
        \xmem_data[63][2] ), .ZN(n15666) );
  AOI22_X1 U19805 ( .A1(n3226), .A2(\xmem_data[58][2] ), .B1(n28701), .B2(
        \xmem_data[59][2] ), .ZN(n15665) );
  NAND2_X1 U19806 ( .A1(n15666), .A2(n15665), .ZN(n15667) );
  NOR2_X1 U19807 ( .A1(n15668), .A2(n15667), .ZN(n15669) );
  AOI22_X1 U19808 ( .A1(n29647), .A2(\xmem_data[44][2] ), .B1(n27761), .B2(
        \xmem_data[45][2] ), .ZN(n15671) );
  INV_X1 U19809 ( .A(n15671), .ZN(n15674) );
  AOI22_X1 U19810 ( .A1(n28685), .A2(\xmem_data[48][2] ), .B1(n29648), .B2(
        \xmem_data[49][2] ), .ZN(n15672) );
  INV_X1 U19811 ( .A(n15672), .ZN(n15673) );
  NOR2_X1 U19812 ( .A1(n15674), .A2(n15673), .ZN(n15685) );
  AOI22_X1 U19813 ( .A1(n27771), .A2(\xmem_data[40][2] ), .B1(n30696), .B2(
        \xmem_data[41][2] ), .ZN(n15684) );
  AOI22_X1 U19814 ( .A1(n29716), .A2(\xmem_data[54][2] ), .B1(n20730), .B2(
        \xmem_data[55][2] ), .ZN(n15675) );
  INV_X1 U19815 ( .A(n15675), .ZN(n15682) );
  AOI22_X1 U19816 ( .A1(n3161), .A2(\xmem_data[52][2] ), .B1(n3184), .B2(
        \xmem_data[53][2] ), .ZN(n15680) );
  AOI22_X1 U19817 ( .A1(n29707), .A2(\xmem_data[42][2] ), .B1(n29706), .B2(
        \xmem_data[43][2] ), .ZN(n15678) );
  AOI22_X1 U19818 ( .A1(n29763), .A2(\xmem_data[46][2] ), .B1(n29591), .B2(
        \xmem_data[47][2] ), .ZN(n15677) );
  AOI22_X1 U19819 ( .A1(n29740), .A2(\xmem_data[50][2] ), .B1(n3121), .B2(
        \xmem_data[51][2] ), .ZN(n15676) );
  NAND2_X1 U19820 ( .A1(n15680), .A2(n15679), .ZN(n15681) );
  NOR2_X1 U19821 ( .A1(n15682), .A2(n15681), .ZN(n15683) );
  NAND4_X1 U19822 ( .A1(n3936), .A2(n15685), .A3(n15684), .A4(n15683), .ZN(
        n15691) );
  AOI22_X1 U19823 ( .A1(n28765), .A2(\xmem_data[32][2] ), .B1(n29785), .B2(
        \xmem_data[33][2] ), .ZN(n15689) );
  AOI22_X1 U19824 ( .A1(n29787), .A2(\xmem_data[34][2] ), .B1(n3142), .B2(
        \xmem_data[35][2] ), .ZN(n15688) );
  AOI22_X1 U19825 ( .A1(n29421), .A2(\xmem_data[36][2] ), .B1(n26616), .B2(
        \xmem_data[37][2] ), .ZN(n15687) );
  AOI22_X1 U19826 ( .A1(n29628), .A2(\xmem_data[38][2] ), .B1(n29789), .B2(
        \xmem_data[39][2] ), .ZN(n15686) );
  NAND4_X1 U19827 ( .A1(n15689), .A2(n15688), .A3(n15687), .A4(n15686), .ZN(
        n15690) );
  OAI21_X1 U19828 ( .B1(n15691), .B2(n15690), .A(n29795), .ZN(n15692) );
  XNOR2_X1 U19829 ( .A(n32936), .B(\fmem_data[19][7] ), .ZN(n30369) );
  XOR2_X1 U19830 ( .A(\fmem_data[19][6] ), .B(\fmem_data[19][7] ), .Z(n15696)
         );
  OAI22_X1 U19831 ( .A1(n31976), .A2(n35656), .B1(n30369), .B2(n35655), .ZN(
        n34257) );
  AOI22_X1 U19832 ( .A1(n28146), .A2(\xmem_data[96][7] ), .B1(n28145), .B2(
        \xmem_data[97][7] ), .ZN(n15700) );
  AOI22_X1 U19833 ( .A1(n3239), .A2(\xmem_data[98][7] ), .B1(n29591), .B2(
        \xmem_data[99][7] ), .ZN(n15699) );
  AOI22_X1 U19834 ( .A1(n28685), .A2(\xmem_data[100][7] ), .B1(n30301), .B2(
        \xmem_data[101][7] ), .ZN(n15698) );
  AOI22_X1 U19835 ( .A1(n29593), .A2(\xmem_data[102][7] ), .B1(n29437), .B2(
        \xmem_data[103][7] ), .ZN(n15697) );
  NAND4_X1 U19836 ( .A1(n15700), .A2(n15699), .A3(n15698), .A4(n15697), .ZN(
        n15716) );
  AOI22_X1 U19837 ( .A1(n3167), .A2(\xmem_data[104][7] ), .B1(n3184), .B2(
        \xmem_data[105][7] ), .ZN(n15704) );
  AOI22_X1 U19838 ( .A1(n30070), .A2(\xmem_data[106][7] ), .B1(n29639), .B2(
        \xmem_data[107][7] ), .ZN(n15703) );
  AOI22_X1 U19839 ( .A1(n28173), .A2(\xmem_data[108][7] ), .B1(n30716), .B2(
        \xmem_data[109][7] ), .ZN(n15702) );
  AOI22_X1 U19840 ( .A1(n29574), .A2(\xmem_data[110][7] ), .B1(n29573), .B2(
        \xmem_data[111][7] ), .ZN(n15701) );
  NAND4_X1 U19841 ( .A1(n15704), .A2(n15703), .A3(n15702), .A4(n15701), .ZN(
        n15715) );
  AOI22_X1 U19842 ( .A1(n29580), .A2(\xmem_data[112][7] ), .B1(n29615), .B2(
        \xmem_data[113][7] ), .ZN(n15708) );
  AOI22_X1 U19843 ( .A1(n29581), .A2(\xmem_data[114][7] ), .B1(n30754), .B2(
        \xmem_data[115][7] ), .ZN(n15707) );
  AOI22_X1 U19844 ( .A1(n29583), .A2(\xmem_data[116][7] ), .B1(n29582), .B2(
        \xmem_data[117][7] ), .ZN(n15706) );
  AOI22_X1 U19845 ( .A1(n29584), .A2(\xmem_data[118][7] ), .B1(n3434), .B2(
        \xmem_data[119][7] ), .ZN(n15705) );
  NAND4_X1 U19846 ( .A1(n15708), .A2(n15707), .A3(n15706), .A4(n15705), .ZN(
        n15714) );
  AOI22_X1 U19847 ( .A1(n30708), .A2(\xmem_data[120][7] ), .B1(n29753), .B2(
        \xmem_data[121][7] ), .ZN(n15712) );
  AOI22_X1 U19848 ( .A1(n29699), .A2(\xmem_data[122][7] ), .B1(n29565), .B2(
        \xmem_data[123][7] ), .ZN(n15711) );
  AOI22_X1 U19849 ( .A1(n29566), .A2(\xmem_data[124][7] ), .B1(n30217), .B2(
        \xmem_data[125][7] ), .ZN(n15710) );
  AOI22_X1 U19850 ( .A1(n29568), .A2(\xmem_data[126][7] ), .B1(n3345), .B2(
        \xmem_data[127][7] ), .ZN(n15709) );
  NAND4_X1 U19851 ( .A1(n15712), .A2(n15711), .A3(n15710), .A4(n15709), .ZN(
        n15713) );
  OR4_X1 U19852 ( .A1(n15716), .A2(n15715), .A3(n15714), .A4(n15713), .ZN(
        n15738) );
  AOI22_X1 U19853 ( .A1(n28146), .A2(\xmem_data[64][7] ), .B1(n29589), .B2(
        \xmem_data[65][7] ), .ZN(n15720) );
  AOI22_X1 U19854 ( .A1(n29603), .A2(\xmem_data[66][7] ), .B1(n30943), .B2(
        \xmem_data[67][7] ), .ZN(n15719) );
  AOI22_X1 U19855 ( .A1(n27811), .A2(\xmem_data[68][7] ), .B1(n29592), .B2(
        \xmem_data[69][7] ), .ZN(n15718) );
  AOI22_X1 U19856 ( .A1(n29649), .A2(\xmem_data[70][7] ), .B1(n25461), .B2(
        \xmem_data[71][7] ), .ZN(n15717) );
  NAND4_X1 U19857 ( .A1(n15720), .A2(n15719), .A3(n15718), .A4(n15717), .ZN(
        n15736) );
  AOI22_X1 U19858 ( .A1(n29616), .A2(\xmem_data[80][7] ), .B1(n29615), .B2(
        \xmem_data[81][7] ), .ZN(n15724) );
  AOI22_X1 U19859 ( .A1(n29617), .A2(\xmem_data[82][7] ), .B1(n28036), .B2(
        \xmem_data[83][7] ), .ZN(n15723) );
  AOI22_X1 U19860 ( .A1(n29619), .A2(\xmem_data[84][7] ), .B1(n29618), .B2(
        \xmem_data[85][7] ), .ZN(n15722) );
  AOI22_X1 U19861 ( .A1(n29621), .A2(\xmem_data[86][7] ), .B1(n3142), .B2(
        \xmem_data[87][7] ), .ZN(n15721) );
  NAND4_X1 U19862 ( .A1(n15724), .A2(n15723), .A3(n15722), .A4(n15721), .ZN(
        n15735) );
  AOI22_X1 U19863 ( .A1(n3166), .A2(\xmem_data[72][7] ), .B1(n3182), .B2(
        \xmem_data[73][7] ), .ZN(n15728) );
  AOI22_X1 U19864 ( .A1(n30310), .A2(\xmem_data[74][7] ), .B1(n29639), .B2(
        \xmem_data[75][7] ), .ZN(n15727) );
  AOI22_X1 U19865 ( .A1(n28173), .A2(\xmem_data[76][7] ), .B1(n29640), .B2(
        \xmem_data[77][7] ), .ZN(n15726) );
  AOI22_X1 U19866 ( .A1(n29641), .A2(\xmem_data[78][7] ), .B1(n3300), .B2(
        \xmem_data[79][7] ), .ZN(n15725) );
  NAND4_X1 U19867 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        n15734) );
  AOI22_X1 U19868 ( .A1(n29630), .A2(\xmem_data[92][7] ), .B1(n30293), .B2(
        \xmem_data[93][7] ), .ZN(n15732) );
  AOI22_X1 U19869 ( .A1(n28734), .A2(\xmem_data[88][7] ), .B1(n26510), .B2(
        \xmem_data[89][7] ), .ZN(n15731) );
  AOI22_X1 U19870 ( .A1(n3392), .A2(\xmem_data[90][7] ), .B1(n29627), .B2(
        \xmem_data[91][7] ), .ZN(n15730) );
  AOI22_X1 U19871 ( .A1(n29667), .A2(\xmem_data[94][7] ), .B1(n3146), .B2(
        \xmem_data[95][7] ), .ZN(n15729) );
  NAND4_X1 U19872 ( .A1(n15732), .A2(n15731), .A3(n15730), .A4(n15729), .ZN(
        n15733) );
  AOI22_X1 U19873 ( .A1(n15738), .A2(n29598), .B1(n15737), .B2(n29600), .ZN(
        n15782) );
  AOI22_X1 U19874 ( .A1(n30743), .A2(\xmem_data[32][7] ), .B1(n28665), .B2(
        \xmem_data[33][7] ), .ZN(n15742) );
  AOI22_X1 U19875 ( .A1(n29603), .A2(\xmem_data[34][7] ), .B1(n28233), .B2(
        \xmem_data[35][7] ), .ZN(n15741) );
  AOI22_X1 U19876 ( .A1(n28751), .A2(\xmem_data[36][7] ), .B1(n29739), .B2(
        \xmem_data[37][7] ), .ZN(n15740) );
  AOI22_X1 U19877 ( .A1(n29649), .A2(\xmem_data[38][7] ), .B1(n30303), .B2(
        \xmem_data[39][7] ), .ZN(n15739) );
  NAND4_X1 U19878 ( .A1(n15742), .A2(n15741), .A3(n15740), .A4(n15739), .ZN(
        n15758) );
  AOI22_X1 U19879 ( .A1(n3167), .A2(\xmem_data[40][7] ), .B1(n3183), .B2(
        \xmem_data[41][7] ), .ZN(n15746) );
  AOI22_X1 U19880 ( .A1(n27031), .A2(\xmem_data[42][7] ), .B1(n29319), .B2(
        \xmem_data[43][7] ), .ZN(n15745) );
  AOI22_X1 U19881 ( .A1(n28680), .A2(\xmem_data[44][7] ), .B1(n30765), .B2(
        \xmem_data[45][7] ), .ZN(n15744) );
  AOI22_X1 U19882 ( .A1(n29641), .A2(\xmem_data[46][7] ), .B1(n3269), .B2(
        \xmem_data[47][7] ), .ZN(n15743) );
  NAND4_X1 U19883 ( .A1(n15746), .A2(n15745), .A3(n15744), .A4(n15743), .ZN(
        n15757) );
  AOI22_X1 U19884 ( .A1(n29616), .A2(\xmem_data[48][7] ), .B1(n29579), .B2(
        \xmem_data[49][7] ), .ZN(n15750) );
  AOI22_X1 U19885 ( .A1(n29617), .A2(\xmem_data[50][7] ), .B1(n29383), .B2(
        \xmem_data[51][7] ), .ZN(n15749) );
  AOI22_X1 U19886 ( .A1(n29619), .A2(\xmem_data[52][7] ), .B1(n29618), .B2(
        \xmem_data[53][7] ), .ZN(n15748) );
  AOI22_X1 U19887 ( .A1(n29621), .A2(\xmem_data[54][7] ), .B1(n3142), .B2(
        \xmem_data[55][7] ), .ZN(n15747) );
  NAND4_X1 U19888 ( .A1(n15750), .A2(n15749), .A3(n15748), .A4(n15747), .ZN(
        n15756) );
  AOI22_X1 U19889 ( .A1(n28136), .A2(\xmem_data[56][7] ), .B1(n29697), .B2(
        \xmem_data[57][7] ), .ZN(n15754) );
  AOI22_X1 U19890 ( .A1(n28138), .A2(\xmem_data[58][7] ), .B1(n29627), .B2(
        \xmem_data[59][7] ), .ZN(n15753) );
  AOI22_X1 U19891 ( .A1(n29630), .A2(\xmem_data[60][7] ), .B1(n3198), .B2(
        \xmem_data[61][7] ), .ZN(n15752) );
  AOI22_X1 U19892 ( .A1(n29667), .A2(\xmem_data[62][7] ), .B1(n28308), .B2(
        \xmem_data[63][7] ), .ZN(n15751) );
  NAND4_X1 U19893 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        n15755) );
  OR4_X1 U19894 ( .A1(n15758), .A2(n15757), .A3(n15756), .A4(n15755), .ZN(
        n15780) );
  AOI22_X1 U19895 ( .A1(n29421), .A2(\xmem_data[24][7] ), .B1(n26510), .B2(
        \xmem_data[25][7] ), .ZN(n15762) );
  AOI22_X1 U19896 ( .A1(n30215), .A2(\xmem_data[26][7] ), .B1(n28218), .B2(
        \xmem_data[27][7] ), .ZN(n15761) );
  AOI22_X1 U19897 ( .A1(n29674), .A2(\xmem_data[28][7] ), .B1(n28786), .B2(
        \xmem_data[29][7] ), .ZN(n15760) );
  AOI22_X1 U19898 ( .A1(n29667), .A2(\xmem_data[30][7] ), .B1(n30698), .B2(
        \xmem_data[31][7] ), .ZN(n15759) );
  NAND4_X1 U19899 ( .A1(n15762), .A2(n15761), .A3(n15760), .A4(n15759), .ZN(
        n15778) );
  AOI22_X1 U19900 ( .A1(n3165), .A2(\xmem_data[8][7] ), .B1(n3190), .B2(
        \xmem_data[9][7] ), .ZN(n15766) );
  AOI22_X1 U19901 ( .A1(n30310), .A2(\xmem_data[10][7] ), .B1(n29639), .B2(
        \xmem_data[11][7] ), .ZN(n15765) );
  AOI22_X1 U19902 ( .A1(n30063), .A2(\xmem_data[12][7] ), .B1(n30765), .B2(
        \xmem_data[13][7] ), .ZN(n15764) );
  AOI22_X1 U19903 ( .A1(n29641), .A2(\xmem_data[14][7] ), .B1(n3328), .B2(
        \xmem_data[15][7] ), .ZN(n15763) );
  NAND4_X1 U19904 ( .A1(n15766), .A2(n15765), .A3(n15764), .A4(n15763), .ZN(
        n15777) );
  AOI22_X1 U19905 ( .A1(n28180), .A2(\xmem_data[0][7] ), .B1(n29704), .B2(
        \xmem_data[1][7] ), .ZN(n15770) );
  AOI22_X1 U19906 ( .A1(n3239), .A2(\xmem_data[2][7] ), .B1(n29591), .B2(
        \xmem_data[3][7] ), .ZN(n15769) );
  AOI22_X1 U19907 ( .A1(n3174), .A2(\xmem_data[4][7] ), .B1(n29739), .B2(
        \xmem_data[5][7] ), .ZN(n15768) );
  AOI22_X1 U19908 ( .A1(n29649), .A2(\xmem_data[6][7] ), .B1(n30746), .B2(
        \xmem_data[7][7] ), .ZN(n15767) );
  NAND4_X1 U19909 ( .A1(n15770), .A2(n15769), .A3(n15768), .A4(n15767), .ZN(
        n15776) );
  AOI22_X1 U19910 ( .A1(n29656), .A2(\xmem_data[16][7] ), .B1(n29615), .B2(
        \xmem_data[17][7] ), .ZN(n15774) );
  AOI22_X1 U19911 ( .A1(n29658), .A2(\xmem_data[18][7] ), .B1(n29657), .B2(
        \xmem_data[19][7] ), .ZN(n15773) );
  AOI22_X1 U19912 ( .A1(n29660), .A2(\xmem_data[20][7] ), .B1(n29659), .B2(
        \xmem_data[21][7] ), .ZN(n15772) );
  AOI22_X1 U19913 ( .A1(n29662), .A2(\xmem_data[22][7] ), .B1(n29661), .B2(
        \xmem_data[23][7] ), .ZN(n15771) );
  NAND4_X1 U19914 ( .A1(n15774), .A2(n15773), .A3(n15772), .A4(n15771), .ZN(
        n15775) );
  OR4_X1 U19915 ( .A1(n15778), .A2(n15777), .A3(n15776), .A4(n15775), .ZN(
        n15779) );
  AOI22_X1 U19916 ( .A1(n15780), .A2(n29683), .B1(n29681), .B2(n15779), .ZN(
        n15781) );
  NAND2_X1 U19917 ( .A1(n15782), .A2(n15781), .ZN(n35359) );
  XNOR2_X1 U19918 ( .A(n35359), .B(\fmem_data[7][3] ), .ZN(n30347) );
  AOI22_X1 U19919 ( .A1(n28734), .A2(\xmem_data[120][6] ), .B1(n29697), .B2(
        \xmem_data[121][6] ), .ZN(n15784) );
  AOI22_X1 U19920 ( .A1(n29674), .A2(\xmem_data[124][6] ), .B1(n28208), .B2(
        \xmem_data[125][6] ), .ZN(n15783) );
  NAND2_X1 U19921 ( .A1(n15784), .A2(n15783), .ZN(n15790) );
  AOI22_X1 U19922 ( .A1(n3161), .A2(\xmem_data[104][6] ), .B1(n3184), .B2(
        \xmem_data[105][6] ), .ZN(n15788) );
  AOI22_X1 U19923 ( .A1(n30062), .A2(\xmem_data[106][6] ), .B1(n27825), .B2(
        \xmem_data[107][6] ), .ZN(n15787) );
  AOI22_X1 U19924 ( .A1(n29815), .A2(\xmem_data[108][6] ), .B1(n30644), .B2(
        \xmem_data[109][6] ), .ZN(n15786) );
  AOI22_X1 U19925 ( .A1(n29574), .A2(\xmem_data[110][6] ), .B1(n29573), .B2(
        \xmem_data[111][6] ), .ZN(n15785) );
  NAND4_X1 U19926 ( .A1(n15788), .A2(n15787), .A3(n15786), .A4(n15785), .ZN(
        n15789) );
  OR2_X1 U19927 ( .A1(n15790), .A2(n15789), .ZN(n15806) );
  AOI22_X1 U19928 ( .A1(n3392), .A2(\xmem_data[122][6] ), .B1(n29565), .B2(
        \xmem_data[123][6] ), .ZN(n15804) );
  AOI22_X1 U19929 ( .A1(n28180), .A2(\xmem_data[96][6] ), .B1(n3368), .B2(
        \xmem_data[97][6] ), .ZN(n15803) );
  AOI22_X1 U19930 ( .A1(n28685), .A2(\xmem_data[100][6] ), .B1(n29648), .B2(
        \xmem_data[101][6] ), .ZN(n15791) );
  INV_X1 U19931 ( .A(n15791), .ZN(n15801) );
  AOI22_X1 U19932 ( .A1(n29656), .A2(\xmem_data[112][6] ), .B1(n29615), .B2(
        \xmem_data[113][6] ), .ZN(n15795) );
  AOI22_X1 U19933 ( .A1(n29658), .A2(\xmem_data[114][6] ), .B1(n31345), .B2(
        \xmem_data[115][6] ), .ZN(n15794) );
  AOI22_X1 U19934 ( .A1(n29583), .A2(\xmem_data[116][6] ), .B1(n29582), .B2(
        \xmem_data[117][6] ), .ZN(n15793) );
  AOI22_X1 U19935 ( .A1(n29584), .A2(\xmem_data[118][6] ), .B1(n24630), .B2(
        \xmem_data[119][6] ), .ZN(n15792) );
  NAND4_X1 U19936 ( .A1(n15795), .A2(n15794), .A3(n15793), .A4(n15792), .ZN(
        n15800) );
  AOI22_X1 U19937 ( .A1(n29593), .A2(\xmem_data[102][6] ), .B1(n28516), .B2(
        \xmem_data[103][6] ), .ZN(n15798) );
  AOI22_X1 U19938 ( .A1(n3239), .A2(\xmem_data[98][6] ), .B1(n29591), .B2(
        \xmem_data[99][6] ), .ZN(n15797) );
  AOI22_X1 U19939 ( .A1(n29568), .A2(\xmem_data[126][6] ), .B1(n3345), .B2(
        \xmem_data[127][6] ), .ZN(n15796) );
  NOR3_X1 U19940 ( .A1(n15801), .A2(n15800), .A3(n15799), .ZN(n15802) );
  OAI21_X1 U19941 ( .B1(n15806), .B2(n15805), .A(n29598), .ZN(n15884) );
  AOI22_X1 U19942 ( .A1(n3161), .A2(\xmem_data[72][6] ), .B1(n3183), .B2(
        \xmem_data[73][6] ), .ZN(n15810) );
  AOI22_X1 U19943 ( .A1(n29810), .A2(\xmem_data[74][6] ), .B1(n22682), .B2(
        \xmem_data[75][6] ), .ZN(n15809) );
  AOI22_X1 U19944 ( .A1(n30766), .A2(\xmem_data[76][6] ), .B1(n29640), .B2(
        \xmem_data[77][6] ), .ZN(n15808) );
  AOI22_X1 U19945 ( .A1(n29641), .A2(\xmem_data[78][6] ), .B1(n3302), .B2(
        \xmem_data[79][6] ), .ZN(n15807) );
  AOI22_X1 U19946 ( .A1(n27754), .A2(\xmem_data[68][6] ), .B1(n30237), .B2(
        \xmem_data[69][6] ), .ZN(n15811) );
  INV_X1 U19947 ( .A(n15811), .ZN(n15818) );
  AOI22_X1 U19948 ( .A1(n29566), .A2(\xmem_data[92][6] ), .B1(n27833), .B2(
        \xmem_data[93][6] ), .ZN(n15814) );
  AOI22_X1 U19949 ( .A1(n29649), .A2(\xmem_data[70][6] ), .B1(n28516), .B2(
        \xmem_data[71][6] ), .ZN(n15813) );
  AOI22_X1 U19950 ( .A1(n29603), .A2(n20682), .B1(n28346), .B2(
        \xmem_data[67][6] ), .ZN(n15812) );
  NAND2_X1 U19951 ( .A1(n15814), .A2(n3921), .ZN(n15817) );
  AOI22_X1 U19952 ( .A1(n3249), .A2(\xmem_data[64][6] ), .B1(n3368), .B2(
        \xmem_data[65][6] ), .ZN(n15815) );
  INV_X1 U19953 ( .A(n15815), .ZN(n15816) );
  NOR3_X1 U19954 ( .A1(n15818), .A2(n15817), .A3(n15816), .ZN(n15819) );
  NAND2_X1 U19955 ( .A1(n3778), .A2(n15819), .ZN(n15832) );
  AOI22_X1 U19956 ( .A1(n29580), .A2(\xmem_data[80][6] ), .B1(n29579), .B2(
        \xmem_data[81][6] ), .ZN(n15823) );
  AOI22_X1 U19957 ( .A1(n29581), .A2(\xmem_data[82][6] ), .B1(n23730), .B2(
        \xmem_data[83][6] ), .ZN(n15822) );
  AOI22_X1 U19958 ( .A1(n29619), .A2(\xmem_data[84][6] ), .B1(n29618), .B2(
        \xmem_data[85][6] ), .ZN(n15821) );
  AOI22_X1 U19959 ( .A1(n29621), .A2(\xmem_data[86][6] ), .B1(n3142), .B2(
        \xmem_data[87][6] ), .ZN(n15820) );
  NAND4_X1 U19960 ( .A1(n15823), .A2(n15822), .A3(n15821), .A4(n15820), .ZN(
        n15826) );
  AOI22_X1 U19961 ( .A1(n29667), .A2(\xmem_data[94][6] ), .B1(n30710), .B2(
        \xmem_data[95][6] ), .ZN(n15824) );
  INV_X1 U19962 ( .A(n15824), .ZN(n15825) );
  NOR2_X1 U19963 ( .A1(n15826), .A2(n15825), .ZN(n15830) );
  AND2_X1 U19964 ( .A1(n29627), .A2(\xmem_data[91][6] ), .ZN(n15827) );
  AOI21_X1 U19965 ( .B1(n28207), .B2(\xmem_data[90][6] ), .A(n15827), .ZN(
        n15829) );
  AOI22_X1 U19966 ( .A1(n28136), .A2(\xmem_data[88][6] ), .B1(n30654), .B2(
        \xmem_data[89][6] ), .ZN(n15828) );
  OAI21_X1 U19967 ( .B1(n15832), .B2(n15831), .A(n29600), .ZN(n15883) );
  AOI22_X1 U19968 ( .A1(n27703), .A2(\xmem_data[0][6] ), .B1(n29646), .B2(
        \xmem_data[1][6] ), .ZN(n15837) );
  AOI22_X1 U19969 ( .A1(n3239), .A2(\xmem_data[2][6] ), .B1(n29591), .B2(
        \xmem_data[3][6] ), .ZN(n15836) );
  AOI22_X1 U19970 ( .A1(n28751), .A2(\xmem_data[4][6] ), .B1(n30237), .B2(
        \xmem_data[5][6] ), .ZN(n15835) );
  AOI22_X1 U19971 ( .A1(n15833), .A2(\xmem_data[6][6] ), .B1(n24213), .B2(
        \xmem_data[7][6] ), .ZN(n15834) );
  AOI22_X1 U19972 ( .A1(n29674), .A2(\xmem_data[28][6] ), .B1(n3170), .B2(
        \xmem_data[29][6] ), .ZN(n15839) );
  AOI22_X1 U19973 ( .A1(n29788), .A2(\xmem_data[24][6] ), .B1(n30182), .B2(
        \xmem_data[25][6] ), .ZN(n15838) );
  AOI22_X1 U19974 ( .A1(n3165), .A2(\xmem_data[8][6] ), .B1(n3189), .B2(
        \xmem_data[9][6] ), .ZN(n15850) );
  AOI22_X1 U19975 ( .A1(n29667), .A2(\xmem_data[30][6] ), .B1(n3132), .B2(
        \xmem_data[31][6] ), .ZN(n15849) );
  AOI22_X1 U19976 ( .A1(n29656), .A2(\xmem_data[16][6] ), .B1(n29655), .B2(
        \xmem_data[17][6] ), .ZN(n15843) );
  AOI22_X1 U19977 ( .A1(n29658), .A2(\xmem_data[18][6] ), .B1(n29657), .B2(
        \xmem_data[19][6] ), .ZN(n15842) );
  AOI22_X1 U19978 ( .A1(n29660), .A2(\xmem_data[20][6] ), .B1(n29659), .B2(
        \xmem_data[21][6] ), .ZN(n15841) );
  AOI22_X1 U19979 ( .A1(n29662), .A2(\xmem_data[22][6] ), .B1(n29661), .B2(
        \xmem_data[23][6] ), .ZN(n15840) );
  NAND4_X1 U19980 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        n15847) );
  AOI22_X1 U19981 ( .A1(n15844), .A2(\xmem_data[14][6] ), .B1(n3302), .B2(
        \xmem_data[15][6] ), .ZN(n15845) );
  INV_X1 U19982 ( .A(n15845), .ZN(n15846) );
  NAND3_X1 U19983 ( .A1(n15850), .A2(n15849), .A3(n15848), .ZN(n15853) );
  AOI22_X1 U19984 ( .A1(n29628), .A2(\xmem_data[26][6] ), .B1(n29789), .B2(
        \xmem_data[27][6] ), .ZN(n15851) );
  INV_X1 U19985 ( .A(n15851), .ZN(n15852) );
  NOR2_X1 U19986 ( .A1(n15853), .A2(n15852), .ZN(n15856) );
  AOI22_X1 U19987 ( .A1(n30715), .A2(\xmem_data[10][6] ), .B1(n23777), .B2(
        \xmem_data[11][6] ), .ZN(n15855) );
  AOI22_X1 U19988 ( .A1(n30063), .A2(\xmem_data[12][6] ), .B1(n30170), .B2(
        \xmem_data[13][6] ), .ZN(n15854) );
  NAND4_X1 U19989 ( .A1(n3546), .A2(n15857), .A3(n15856), .A4(n3922), .ZN(
        n15858) );
  NAND2_X1 U19990 ( .A1(n15858), .A2(n29681), .ZN(n15882) );
  AOI22_X1 U19991 ( .A1(n29590), .A2(\xmem_data[32][6] ), .B1(n28238), .B2(
        \xmem_data[33][6] ), .ZN(n15861) );
  AOI22_X1 U19992 ( .A1(n29790), .A2(\xmem_data[58][6] ), .B1(n29627), .B2(
        \xmem_data[59][6] ), .ZN(n15860) );
  AOI22_X1 U19993 ( .A1(n29566), .A2(\xmem_data[60][6] ), .B1(n27833), .B2(
        \xmem_data[61][6] ), .ZN(n15859) );
  NAND3_X1 U19994 ( .A1(n15861), .A2(n15860), .A3(n15859), .ZN(n15867) );
  AOI22_X1 U19995 ( .A1(n3164), .A2(\xmem_data[40][6] ), .B1(n3183), .B2(
        \xmem_data[41][6] ), .ZN(n15865) );
  AOI22_X1 U19996 ( .A1(n29716), .A2(\xmem_data[42][6] ), .B1(n31255), .B2(
        \xmem_data[43][6] ), .ZN(n15864) );
  AOI22_X1 U19997 ( .A1(n29815), .A2(\xmem_data[44][6] ), .B1(n30685), .B2(
        \xmem_data[45][6] ), .ZN(n15863) );
  AOI22_X1 U19998 ( .A1(n29641), .A2(\xmem_data[46][6] ), .B1(n29054), .B2(
        \xmem_data[47][6] ), .ZN(n15862) );
  NAND4_X1 U19999 ( .A1(n15865), .A2(n15864), .A3(n15863), .A4(n15862), .ZN(
        n15866) );
  AOI22_X1 U20000 ( .A1(n29433), .A2(\xmem_data[56][6] ), .B1(n27013), .B2(
        \xmem_data[57][6] ), .ZN(n15868) );
  INV_X1 U20001 ( .A(n15868), .ZN(n15878) );
  AOI22_X1 U20002 ( .A1(n29714), .A2(\xmem_data[36][6] ), .B1(n30249), .B2(
        \xmem_data[37][6] ), .ZN(n15876) );
  AOI22_X1 U20003 ( .A1(n29649), .A2(\xmem_data[38][6] ), .B1(n31354), .B2(
        \xmem_data[39][6] ), .ZN(n15870) );
  AOI22_X1 U20004 ( .A1(n29603), .A2(\xmem_data[34][6] ), .B1(n29403), .B2(
        \xmem_data[35][6] ), .ZN(n15869) );
  AOI22_X1 U20005 ( .A1(n29667), .A2(\xmem_data[62][6] ), .B1(n28084), .B2(
        \xmem_data[63][6] ), .ZN(n15875) );
  AOI22_X1 U20006 ( .A1(n29580), .A2(\xmem_data[48][6] ), .B1(n29579), .B2(
        \xmem_data[49][6] ), .ZN(n15874) );
  AOI22_X1 U20007 ( .A1(n29581), .A2(\xmem_data[50][6] ), .B1(n28192), .B2(
        \xmem_data[51][6] ), .ZN(n15873) );
  AOI22_X1 U20008 ( .A1(n29619), .A2(\xmem_data[52][6] ), .B1(n29618), .B2(
        \xmem_data[53][6] ), .ZN(n15872) );
  AOI22_X1 U20009 ( .A1(n29621), .A2(\xmem_data[54][6] ), .B1(n3142), .B2(
        \xmem_data[55][6] ), .ZN(n15871) );
  NAND4_X1 U20010 ( .A1(n15876), .A2(n3933), .A3(n15875), .A4(n3503), .ZN(
        n15877) );
  NAND4_X1 U20011 ( .A1(n15884), .A2(n15883), .A3(n15882), .A4(n15881), .ZN(
        n35140) );
  XNOR2_X1 U20012 ( .A(n35140), .B(\fmem_data[7][3] ), .ZN(n29542) );
  XOR2_X1 U20013 ( .A(\fmem_data[7][2] ), .B(\fmem_data[7][3] ), .Z(n15885) );
  AOI22_X1 U20014 ( .A1(n28462), .A2(\xmem_data[96][5] ), .B1(n28226), .B2(
        \xmem_data[97][5] ), .ZN(n15889) );
  AOI22_X1 U20015 ( .A1(n31314), .A2(\xmem_data[98][5] ), .B1(n27542), .B2(
        \xmem_data[99][5] ), .ZN(n15888) );
  AOI22_X1 U20016 ( .A1(n28468), .A2(\xmem_data[100][5] ), .B1(n29657), .B2(
        \xmem_data[101][5] ), .ZN(n15887) );
  AOI22_X1 U20017 ( .A1(n29248), .A2(\xmem_data[102][5] ), .B1(n28354), .B2(
        \xmem_data[103][5] ), .ZN(n15886) );
  NAND4_X1 U20018 ( .A1(n15889), .A2(n15888), .A3(n15887), .A4(n15886), .ZN(
        n15905) );
  AOI22_X1 U20019 ( .A1(n29173), .A2(\xmem_data[106][5] ), .B1(n28044), .B2(
        \xmem_data[107][5] ), .ZN(n15893) );
  AOI22_X1 U20020 ( .A1(n21309), .A2(\xmem_data[104][5] ), .B1(n23754), .B2(
        \xmem_data[105][5] ), .ZN(n15892) );
  AOI22_X1 U20021 ( .A1(n3222), .A2(\xmem_data[108][5] ), .B1(n29494), .B2(
        \xmem_data[109][5] ), .ZN(n15891) );
  AOI22_X1 U20022 ( .A1(n25562), .A2(\xmem_data[110][5] ), .B1(n29174), .B2(
        \xmem_data[111][5] ), .ZN(n15890) );
  NAND4_X1 U20023 ( .A1(n15893), .A2(n15892), .A3(n15891), .A4(n15890), .ZN(
        n15904) );
  AOI22_X1 U20024 ( .A1(n29181), .A2(\xmem_data[112][5] ), .B1(n29157), .B2(
        \xmem_data[113][5] ), .ZN(n15897) );
  AOI22_X1 U20025 ( .A1(n25514), .A2(\xmem_data[114][5] ), .B1(n27447), .B2(
        \xmem_data[115][5] ), .ZN(n15896) );
  AOI22_X1 U20026 ( .A1(n29180), .A2(\xmem_data[116][5] ), .B1(n29179), .B2(
        \xmem_data[117][5] ), .ZN(n15895) );
  AOI22_X1 U20027 ( .A1(n28345), .A2(\xmem_data[118][5] ), .B1(n28334), .B2(
        \xmem_data[119][5] ), .ZN(n15894) );
  NAND4_X1 U20028 ( .A1(n15897), .A2(n15896), .A3(n15895), .A4(n15894), .ZN(
        n15903) );
  AOI22_X1 U20029 ( .A1(n23793), .A2(\xmem_data[120][5] ), .B1(n29187), .B2(
        \xmem_data[121][5] ), .ZN(n15901) );
  AOI22_X1 U20030 ( .A1(n23716), .A2(\xmem_data[122][5] ), .B1(n23717), .B2(
        \xmem_data[123][5] ), .ZN(n15900) );
  AOI22_X1 U20031 ( .A1(n27918), .A2(\xmem_data[124][5] ), .B1(n23777), .B2(
        \xmem_data[125][5] ), .ZN(n15899) );
  AOI22_X1 U20032 ( .A1(n29190), .A2(\xmem_data[126][5] ), .B1(n3206), .B2(
        \xmem_data[127][5] ), .ZN(n15898) );
  NAND4_X1 U20033 ( .A1(n15901), .A2(n15900), .A3(n15899), .A4(n15898), .ZN(
        n15902) );
  OR4_X1 U20034 ( .A1(n15905), .A2(n15904), .A3(n15903), .A4(n15902), .ZN(
        n15928) );
  AOI22_X1 U20035 ( .A1(n29089), .A2(\xmem_data[64][5] ), .B1(n30645), .B2(
        \xmem_data[65][5] ), .ZN(n15909) );
  AOI22_X1 U20036 ( .A1(n27365), .A2(\xmem_data[66][5] ), .B1(n24685), .B2(
        \xmem_data[67][5] ), .ZN(n15908) );
  AOI22_X1 U20037 ( .A1(n29086), .A2(\xmem_data[68][5] ), .B1(n27568), .B2(
        \xmem_data[69][5] ), .ZN(n15907) );
  AOI22_X1 U20038 ( .A1(n30601), .A2(\xmem_data[70][5] ), .B1(n25408), .B2(
        \xmem_data[71][5] ), .ZN(n15906) );
  NAND4_X1 U20039 ( .A1(n15909), .A2(n15908), .A3(n15907), .A4(n15906), .ZN(
        n15926) );
  AND2_X1 U20040 ( .A1(n28501), .A2(\xmem_data[74][5] ), .ZN(n15910) );
  AOI21_X1 U20041 ( .B1(n20991), .B2(\xmem_data[75][5] ), .A(n15910), .ZN(
        n15914) );
  AOI22_X1 U20042 ( .A1(n27563), .A2(\xmem_data[72][5] ), .B1(n3305), .B2(
        \xmem_data[73][5] ), .ZN(n15913) );
  AOI22_X1 U20043 ( .A1(n3222), .A2(\xmem_data[76][5] ), .B1(n23740), .B2(
        \xmem_data[77][5] ), .ZN(n15912) );
  AOI22_X1 U20044 ( .A1(n29095), .A2(\xmem_data[78][5] ), .B1(n17010), .B2(
        \xmem_data[79][5] ), .ZN(n15911) );
  NAND4_X1 U20045 ( .A1(n15914), .A2(n15913), .A3(n15912), .A4(n15911), .ZN(
        n15925) );
  AOI22_X1 U20046 ( .A1(n29104), .A2(\xmem_data[80][5] ), .B1(n29762), .B2(
        \xmem_data[81][5] ), .ZN(n15918) );
  AOI22_X1 U20047 ( .A1(n29103), .A2(\xmem_data[82][5] ), .B1(n22712), .B2(
        \xmem_data[83][5] ), .ZN(n15917) );
  AOI22_X1 U20048 ( .A1(n27943), .A2(\xmem_data[84][5] ), .B1(n27514), .B2(
        \xmem_data[85][5] ), .ZN(n15916) );
  AOI22_X1 U20049 ( .A1(n24212), .A2(\xmem_data[86][5] ), .B1(n29109), .B2(
        \xmem_data[87][5] ), .ZN(n15915) );
  NAND4_X1 U20050 ( .A1(n15918), .A2(n15917), .A3(n15916), .A4(n15915), .ZN(
        n15924) );
  AOI22_X1 U20051 ( .A1(n28090), .A2(\xmem_data[88][5] ), .B1(n29187), .B2(
        \xmem_data[89][5] ), .ZN(n15922) );
  AOI22_X1 U20052 ( .A1(n29162), .A2(\xmem_data[90][5] ), .B1(n25573), .B2(
        \xmem_data[91][5] ), .ZN(n15921) );
  AOI22_X1 U20053 ( .A1(n25398), .A2(\xmem_data[92][5] ), .B1(n22682), .B2(
        \xmem_data[93][5] ), .ZN(n15920) );
  AOI22_X1 U20054 ( .A1(n29101), .A2(\xmem_data[94][5] ), .B1(n3326), .B2(
        \xmem_data[95][5] ), .ZN(n15919) );
  NAND4_X1 U20055 ( .A1(n15922), .A2(n15921), .A3(n15920), .A4(n15919), .ZN(
        n15923) );
  OR4_X1 U20056 ( .A1(n15926), .A2(n15925), .A3(n15924), .A4(n15923), .ZN(
        n15927) );
  AOI22_X1 U20057 ( .A1(n15928), .A2(n29171), .B1(n15927), .B2(n29201), .ZN(
        n15975) );
  AOI22_X1 U20058 ( .A1(n30598), .A2(\xmem_data[0][5] ), .B1(n28226), .B2(
        \xmem_data[1][5] ), .ZN(n15932) );
  AOI22_X1 U20059 ( .A1(n27365), .A2(\xmem_data[2][5] ), .B1(n20818), .B2(
        \xmem_data[3][5] ), .ZN(n15931) );
  AOI22_X1 U20060 ( .A1(n29136), .A2(\xmem_data[4][5] ), .B1(n29657), .B2(
        \xmem_data[5][5] ), .ZN(n15930) );
  AOI22_X1 U20061 ( .A1(n29125), .A2(\xmem_data[6][5] ), .B1(n29124), .B2(
        \xmem_data[7][5] ), .ZN(n15929) );
  NAND4_X1 U20062 ( .A1(n15932), .A2(n15931), .A3(n15930), .A4(n15929), .ZN(
        n15949) );
  AOI22_X1 U20063 ( .A1(n29118), .A2(\xmem_data[8][5] ), .B1(n3332), .B2(
        \xmem_data[9][5] ), .ZN(n15937) );
  AND2_X1 U20064 ( .A1(n30589), .A2(\xmem_data[10][5] ), .ZN(n15933) );
  AOI21_X1 U20065 ( .B1(n25354), .B2(\xmem_data[11][5] ), .A(n15933), .ZN(
        n15936) );
  AOI22_X1 U20066 ( .A1(n3221), .A2(\xmem_data[12][5] ), .B1(n29494), .B2(
        \xmem_data[13][5] ), .ZN(n15935) );
  AOI22_X1 U20067 ( .A1(n25562), .A2(\xmem_data[14][5] ), .B1(n30883), .B2(
        \xmem_data[15][5] ), .ZN(n15934) );
  NAND4_X1 U20068 ( .A1(n15937), .A2(n15936), .A3(n15935), .A4(n15934), .ZN(
        n15948) );
  AOI22_X1 U20069 ( .A1(n28509), .A2(\xmem_data[16][5] ), .B1(n27396), .B2(
        \xmem_data[17][5] ), .ZN(n15941) );
  AOI22_X1 U20070 ( .A1(n3231), .A2(\xmem_data[18][5] ), .B1(n27447), .B2(
        \xmem_data[19][5] ), .ZN(n15940) );
  AOI22_X1 U20071 ( .A1(n28415), .A2(\xmem_data[20][5] ), .B1(n28051), .B2(
        \xmem_data[21][5] ), .ZN(n15939) );
  AOI22_X1 U20072 ( .A1(n24212), .A2(\xmem_data[22][5] ), .B1(n28334), .B2(
        \xmem_data[23][5] ), .ZN(n15938) );
  NAND4_X1 U20073 ( .A1(n15941), .A2(n15940), .A3(n15939), .A4(n15938), .ZN(
        n15947) );
  AOI22_X1 U20074 ( .A1(n23793), .A2(\xmem_data[24][5] ), .B1(n3464), .B2(
        \xmem_data[25][5] ), .ZN(n15945) );
  AOI22_X1 U20075 ( .A1(n3208), .A2(\xmem_data[26][5] ), .B1(n25573), .B2(
        \xmem_data[27][5] ), .ZN(n15944) );
  AOI22_X1 U20076 ( .A1(n25520), .A2(\xmem_data[28][5] ), .B1(n17044), .B2(
        \xmem_data[29][5] ), .ZN(n15943) );
  AOI22_X1 U20077 ( .A1(n20814), .A2(\xmem_data[30][5] ), .B1(n28428), .B2(
        \xmem_data[31][5] ), .ZN(n15942) );
  NAND4_X1 U20078 ( .A1(n15945), .A2(n15944), .A3(n15943), .A4(n15942), .ZN(
        n15946) );
  OR4_X1 U20079 ( .A1(n15949), .A2(n15948), .A3(n15947), .A4(n15946), .ZN(
        n15973) );
  AND2_X1 U20080 ( .A1(n24439), .A2(\xmem_data[42][5] ), .ZN(n15950) );
  AOI21_X1 U20081 ( .B1(n20991), .B2(\xmem_data[43][5] ), .A(n15950), .ZN(
        n15954) );
  AOI22_X1 U20082 ( .A1(n24470), .A2(\xmem_data[40][5] ), .B1(n27813), .B2(
        \xmem_data[41][5] ), .ZN(n15953) );
  AOI22_X1 U20083 ( .A1(n3222), .A2(\xmem_data[44][5] ), .B1(n24696), .B2(
        \xmem_data[45][5] ), .ZN(n15952) );
  AOI22_X1 U20084 ( .A1(n29095), .A2(\xmem_data[46][5] ), .B1(n27938), .B2(
        \xmem_data[47][5] ), .ZN(n15951) );
  NAND4_X1 U20085 ( .A1(n15954), .A2(n15953), .A3(n15952), .A4(n15951), .ZN(
        n15971) );
  AOI22_X1 U20086 ( .A1(n29089), .A2(\xmem_data[32][5] ), .B1(n23724), .B2(
        \xmem_data[33][5] ), .ZN(n15959) );
  AOI22_X1 U20087 ( .A1(n27365), .A2(\xmem_data[34][5] ), .B1(n29151), .B2(
        \xmem_data[35][5] ), .ZN(n15958) );
  AND2_X1 U20088 ( .A1(n29086), .A2(\xmem_data[36][5] ), .ZN(n15955) );
  AOI21_X1 U20089 ( .B1(n31345), .B2(\xmem_data[37][5] ), .A(n15955), .ZN(
        n15957) );
  AOI22_X1 U20090 ( .A1(n22727), .A2(\xmem_data[38][5] ), .B1(n25724), .B2(
        \xmem_data[39][5] ), .ZN(n15956) );
  NAND4_X1 U20091 ( .A1(n15959), .A2(n15958), .A3(n15957), .A4(n15956), .ZN(
        n15970) );
  AOI22_X1 U20092 ( .A1(n29104), .A2(\xmem_data[48][5] ), .B1(n29157), .B2(
        \xmem_data[49][5] ), .ZN(n15963) );
  AOI22_X1 U20093 ( .A1(n29103), .A2(\xmem_data[50][5] ), .B1(n30607), .B2(
        \xmem_data[51][5] ), .ZN(n15962) );
  AOI22_X1 U20094 ( .A1(n25456), .A2(\xmem_data[52][5] ), .B1(n28346), .B2(
        \xmem_data[53][5] ), .ZN(n15961) );
  AOI22_X1 U20095 ( .A1(n22740), .A2(\xmem_data[54][5] ), .B1(n29109), .B2(
        \xmem_data[55][5] ), .ZN(n15960) );
  NAND4_X1 U20096 ( .A1(n15963), .A2(n15962), .A3(n15961), .A4(n15960), .ZN(
        n15969) );
  AOI22_X1 U20097 ( .A1(n22703), .A2(\xmem_data[56][5] ), .B1(n3464), .B2(
        \xmem_data[57][5] ), .ZN(n15967) );
  AOI22_X1 U20098 ( .A1(n29162), .A2(\xmem_data[58][5] ), .B1(n25573), .B2(
        \xmem_data[59][5] ), .ZN(n15966) );
  AOI22_X1 U20099 ( .A1(n31270), .A2(\xmem_data[60][5] ), .B1(n22717), .B2(
        \xmem_data[61][5] ), .ZN(n15965) );
  AOI22_X1 U20100 ( .A1(n29101), .A2(\xmem_data[62][5] ), .B1(n30899), .B2(
        \xmem_data[63][5] ), .ZN(n15964) );
  NAND4_X1 U20101 ( .A1(n15967), .A2(n15966), .A3(n15965), .A4(n15964), .ZN(
        n15968) );
  OR4_X1 U20102 ( .A1(n15971), .A2(n15970), .A3(n15969), .A4(n15968), .ZN(
        n15972) );
  AOI22_X1 U20103 ( .A1(n15973), .A2(n29143), .B1(n15972), .B2(n29145), .ZN(
        n15974) );
  NAND2_X1 U20104 ( .A1(n15975), .A2(n15974), .ZN(n34859) );
  XNOR2_X1 U20105 ( .A(n34859), .B(\fmem_data[25][3] ), .ZN(n29208) );
  AOI22_X1 U20106 ( .A1(n29089), .A2(\xmem_data[32][6] ), .B1(n30600), .B2(
        \xmem_data[33][6] ), .ZN(n15979) );
  AOI22_X1 U20107 ( .A1(n20553), .A2(\xmem_data[34][6] ), .B1(n24685), .B2(
        \xmem_data[35][6] ), .ZN(n15978) );
  AOI22_X1 U20108 ( .A1(n29086), .A2(\xmem_data[36][6] ), .B1(n28467), .B2(
        \xmem_data[37][6] ), .ZN(n15977) );
  AOI22_X1 U20109 ( .A1(n17050), .A2(\xmem_data[38][6] ), .B1(n25441), .B2(
        \xmem_data[39][6] ), .ZN(n15976) );
  NAND4_X1 U20110 ( .A1(n15979), .A2(n15978), .A3(n15977), .A4(n15976), .ZN(
        n15995) );
  AOI22_X1 U20111 ( .A1(n30861), .A2(\xmem_data[40][6] ), .B1(n3412), .B2(
        \xmem_data[41][6] ), .ZN(n15983) );
  AOI22_X1 U20112 ( .A1(n30589), .A2(\xmem_data[42][6] ), .B1(n20576), .B2(
        \xmem_data[43][6] ), .ZN(n15982) );
  AOI22_X1 U20113 ( .A1(n3220), .A2(\xmem_data[44][6] ), .B1(n25414), .B2(
        \xmem_data[45][6] ), .ZN(n15981) );
  AOI22_X1 U20114 ( .A1(n29095), .A2(\xmem_data[46][6] ), .B1(n25490), .B2(
        \xmem_data[47][6] ), .ZN(n15980) );
  NAND4_X1 U20115 ( .A1(n15983), .A2(n15982), .A3(n15981), .A4(n15980), .ZN(
        n15994) );
  AOI22_X1 U20116 ( .A1(n29104), .A2(\xmem_data[48][6] ), .B1(n29157), .B2(
        \xmem_data[49][6] ), .ZN(n15987) );
  AOI22_X1 U20117 ( .A1(n29103), .A2(\xmem_data[50][6] ), .B1(n27447), .B2(
        \xmem_data[51][6] ), .ZN(n15986) );
  AOI22_X1 U20118 ( .A1(n27943), .A2(\xmem_data[52][6] ), .B1(n29308), .B2(
        \xmem_data[53][6] ), .ZN(n15985) );
  AOI22_X1 U20119 ( .A1(n25423), .A2(\xmem_data[54][6] ), .B1(n29109), .B2(
        \xmem_data[55][6] ), .ZN(n15984) );
  NAND4_X1 U20120 ( .A1(n15987), .A2(n15986), .A3(n15985), .A4(n15984), .ZN(
        n15993) );
  AOI22_X1 U20121 ( .A1(n25382), .A2(\xmem_data[56][6] ), .B1(n30303), .B2(
        \xmem_data[57][6] ), .ZN(n15991) );
  AOI22_X1 U20122 ( .A1(n3213), .A2(\xmem_data[58][6] ), .B1(n24509), .B2(
        \xmem_data[59][6] ), .ZN(n15990) );
  AOI22_X1 U20123 ( .A1(n25398), .A2(\xmem_data[60][6] ), .B1(n20942), .B2(
        \xmem_data[61][6] ), .ZN(n15989) );
  AOI22_X1 U20124 ( .A1(n29101), .A2(\xmem_data[62][6] ), .B1(n17002), .B2(
        \xmem_data[63][6] ), .ZN(n15988) );
  NAND4_X1 U20125 ( .A1(n15991), .A2(n15990), .A3(n15989), .A4(n15988), .ZN(
        n15992) );
  OR4_X1 U20126 ( .A1(n15995), .A2(n15994), .A3(n15993), .A4(n15992), .ZN(
        n16018) );
  AND2_X1 U20127 ( .A1(n30589), .A2(\xmem_data[10][6] ), .ZN(n15996) );
  AOI21_X1 U20128 ( .B1(n27502), .B2(\xmem_data[11][6] ), .A(n15996), .ZN(
        n16000) );
  AOI22_X1 U20129 ( .A1(n29118), .A2(\xmem_data[8][6] ), .B1(n28039), .B2(
        \xmem_data[9][6] ), .ZN(n15999) );
  AOI22_X1 U20130 ( .A1(n3221), .A2(\xmem_data[12][6] ), .B1(n31368), .B2(
        \xmem_data[13][6] ), .ZN(n15998) );
  AOI22_X1 U20131 ( .A1(n25562), .A2(\xmem_data[14][6] ), .B1(n3340), .B2(
        \xmem_data[15][6] ), .ZN(n15997) );
  NAND4_X1 U20132 ( .A1(n16000), .A2(n15999), .A3(n15998), .A4(n15997), .ZN(
        n16016) );
  AOI22_X1 U20133 ( .A1(n31361), .A2(\xmem_data[0][6] ), .B1(n28202), .B2(
        \xmem_data[1][6] ), .ZN(n16004) );
  AOI22_X1 U20134 ( .A1(n27365), .A2(\xmem_data[2][6] ), .B1(n29151), .B2(
        \xmem_data[3][6] ), .ZN(n16003) );
  AOI22_X1 U20135 ( .A1(n29136), .A2(\xmem_data[4][6] ), .B1(n14982), .B2(
        \xmem_data[5][6] ), .ZN(n16002) );
  AOI22_X1 U20136 ( .A1(n29125), .A2(\xmem_data[6][6] ), .B1(n29124), .B2(
        \xmem_data[7][6] ), .ZN(n16001) );
  NAND4_X1 U20137 ( .A1(n16004), .A2(n16003), .A3(n16002), .A4(n16001), .ZN(
        n16015) );
  AOI22_X1 U20138 ( .A1(n24633), .A2(\xmem_data[16][6] ), .B1(n29157), .B2(
        \xmem_data[17][6] ), .ZN(n16008) );
  AOI22_X1 U20139 ( .A1(n3231), .A2(\xmem_data[18][6] ), .B1(n27447), .B2(
        \xmem_data[19][6] ), .ZN(n16007) );
  AOI22_X1 U20140 ( .A1(n20588), .A2(\xmem_data[20][6] ), .B1(n17013), .B2(
        \xmem_data[21][6] ), .ZN(n16006) );
  AOI22_X1 U20141 ( .A1(n22740), .A2(\xmem_data[22][6] ), .B1(n20541), .B2(
        \xmem_data[23][6] ), .ZN(n16005) );
  NAND4_X1 U20142 ( .A1(n16008), .A2(n16007), .A3(n16006), .A4(n16005), .ZN(
        n16014) );
  AOI22_X1 U20143 ( .A1(n22703), .A2(\xmem_data[24][6] ), .B1(n27455), .B2(
        \xmem_data[25][6] ), .ZN(n16012) );
  AOI22_X1 U20144 ( .A1(n27516), .A2(\xmem_data[26][6] ), .B1(n28059), .B2(
        \xmem_data[27][6] ), .ZN(n16011) );
  AOI22_X1 U20145 ( .A1(n27518), .A2(\xmem_data[28][6] ), .B1(n23802), .B2(
        \xmem_data[29][6] ), .ZN(n16010) );
  AOI22_X1 U20146 ( .A1(n29280), .A2(\xmem_data[30][6] ), .B1(n24615), .B2(
        \xmem_data[31][6] ), .ZN(n16009) );
  NAND4_X1 U20147 ( .A1(n16012), .A2(n16011), .A3(n16010), .A4(n16009), .ZN(
        n16013) );
  OR4_X1 U20148 ( .A1(n16016), .A2(n16015), .A3(n16014), .A4(n16013), .ZN(
        n16017) );
  AOI22_X1 U20149 ( .A1(n16018), .A2(n29145), .B1(n16017), .B2(n29143), .ZN(
        n16064) );
  AOI22_X1 U20150 ( .A1(n28494), .A2(\xmem_data[96][6] ), .B1(n25401), .B2(
        \xmem_data[97][6] ), .ZN(n16022) );
  AOI22_X1 U20151 ( .A1(n29126), .A2(\xmem_data[98][6] ), .B1(n29151), .B2(
        \xmem_data[99][6] ), .ZN(n16021) );
  AOI22_X1 U20152 ( .A1(n17003), .A2(\xmem_data[100][6] ), .B1(n25628), .B2(
        \xmem_data[101][6] ), .ZN(n16020) );
  AOI22_X1 U20153 ( .A1(n20579), .A2(\xmem_data[102][6] ), .B1(n25408), .B2(
        \xmem_data[103][6] ), .ZN(n16019) );
  NAND4_X1 U20154 ( .A1(n16022), .A2(n16021), .A3(n16020), .A4(n16019), .ZN(
        n16038) );
  AOI22_X1 U20155 ( .A1(n28317), .A2(\xmem_data[104][6] ), .B1(n3332), .B2(
        \xmem_data[105][6] ), .ZN(n16026) );
  AOI22_X1 U20156 ( .A1(n29173), .A2(\xmem_data[106][6] ), .B1(n29254), .B2(
        \xmem_data[107][6] ), .ZN(n16025) );
  AOI22_X1 U20157 ( .A1(n3219), .A2(\xmem_data[108][6] ), .B1(n20805), .B2(
        \xmem_data[109][6] ), .ZN(n16024) );
  AOI22_X1 U20158 ( .A1(n24207), .A2(\xmem_data[110][6] ), .B1(n29174), .B2(
        \xmem_data[111][6] ), .ZN(n16023) );
  NAND4_X1 U20159 ( .A1(n16026), .A2(n16025), .A3(n16024), .A4(n16023), .ZN(
        n16037) );
  AOI22_X1 U20160 ( .A1(n29181), .A2(\xmem_data[112][6] ), .B1(n27396), .B2(
        \xmem_data[113][6] ), .ZN(n16030) );
  AOI22_X1 U20161 ( .A1(n30877), .A2(\xmem_data[114][6] ), .B1(n23813), .B2(
        \xmem_data[115][6] ), .ZN(n16029) );
  AOI22_X1 U20162 ( .A1(n29180), .A2(\xmem_data[116][6] ), .B1(n29179), .B2(
        \xmem_data[117][6] ), .ZN(n16028) );
  AOI22_X1 U20163 ( .A1(n24639), .A2(\xmem_data[118][6] ), .B1(n20959), .B2(
        \xmem_data[119][6] ), .ZN(n16027) );
  NAND4_X1 U20164 ( .A1(n16030), .A2(n16029), .A3(n16028), .A4(n16027), .ZN(
        n16036) );
  AOI22_X1 U20165 ( .A1(n22741), .A2(\xmem_data[120][6] ), .B1(n21005), .B2(
        \xmem_data[121][6] ), .ZN(n16034) );
  AOI22_X1 U20166 ( .A1(n29188), .A2(\xmem_data[122][6] ), .B1(n24509), .B2(
        \xmem_data[123][6] ), .ZN(n16033) );
  AOI22_X1 U20167 ( .A1(n24707), .A2(\xmem_data[124][6] ), .B1(n29047), .B2(
        \xmem_data[125][6] ), .ZN(n16032) );
  AOI22_X1 U20168 ( .A1(n29190), .A2(\xmem_data[126][6] ), .B1(n3206), .B2(
        \xmem_data[127][6] ), .ZN(n16031) );
  NAND4_X1 U20169 ( .A1(n16034), .A2(n16033), .A3(n16032), .A4(n16031), .ZN(
        n16035) );
  OR4_X1 U20170 ( .A1(n16038), .A2(n16037), .A3(n16036), .A4(n16035), .ZN(
        n16062) );
  AOI22_X1 U20171 ( .A1(n29089), .A2(\xmem_data[64][6] ), .B1(n28202), .B2(
        \xmem_data[65][6] ), .ZN(n16043) );
  AOI22_X1 U20172 ( .A1(n27365), .A2(n20682), .B1(n22684), .B2(
        \xmem_data[67][6] ), .ZN(n16042) );
  AND2_X1 U20173 ( .A1(n29086), .A2(\xmem_data[68][6] ), .ZN(n16039) );
  AOI21_X1 U20174 ( .B1(n20952), .B2(\xmem_data[69][6] ), .A(n16039), .ZN(
        n16041) );
  AOI22_X1 U20175 ( .A1(n29125), .A2(\xmem_data[70][6] ), .B1(n20710), .B2(
        \xmem_data[71][6] ), .ZN(n16040) );
  NAND4_X1 U20176 ( .A1(n16043), .A2(n16042), .A3(n16041), .A4(n16040), .ZN(
        n16060) );
  AOI22_X1 U20177 ( .A1(n29104), .A2(\xmem_data[80][6] ), .B1(n27396), .B2(
        \xmem_data[81][6] ), .ZN(n16047) );
  AOI22_X1 U20178 ( .A1(n29103), .A2(\xmem_data[82][6] ), .B1(n25604), .B2(
        \xmem_data[83][6] ), .ZN(n16046) );
  AOI22_X1 U20179 ( .A1(n20546), .A2(\xmem_data[84][6] ), .B1(n25708), .B2(
        \xmem_data[85][6] ), .ZN(n16045) );
  AOI22_X1 U20180 ( .A1(n27452), .A2(\xmem_data[86][6] ), .B1(n29109), .B2(
        \xmem_data[87][6] ), .ZN(n16044) );
  NAND4_X1 U20181 ( .A1(n16047), .A2(n16046), .A3(n16045), .A4(n16044), .ZN(
        n16059) );
  AOI22_X1 U20182 ( .A1(n25606), .A2(\xmem_data[88][6] ), .B1(n28091), .B2(
        \xmem_data[89][6] ), .ZN(n16051) );
  AOI22_X1 U20183 ( .A1(n25383), .A2(\xmem_data[90][6] ), .B1(n24593), .B2(
        \xmem_data[91][6] ), .ZN(n16050) );
  AOI22_X1 U20184 ( .A1(n20505), .A2(\xmem_data[92][6] ), .B1(n22682), .B2(
        \xmem_data[93][6] ), .ZN(n16049) );
  AOI22_X1 U20185 ( .A1(n29101), .A2(\xmem_data[94][6] ), .B1(n24220), .B2(
        \xmem_data[95][6] ), .ZN(n16048) );
  NAND4_X1 U20186 ( .A1(n16051), .A2(n16050), .A3(n16049), .A4(n16048), .ZN(
        n16058) );
  AND2_X1 U20187 ( .A1(n14875), .A2(\xmem_data[74][6] ), .ZN(n16052) );
  AOI21_X1 U20188 ( .B1(n25692), .B2(\xmem_data[75][6] ), .A(n16052), .ZN(
        n16056) );
  AOI22_X1 U20189 ( .A1(n24573), .A2(\xmem_data[72][6] ), .B1(n3382), .B2(
        \xmem_data[73][6] ), .ZN(n16055) );
  AOI22_X1 U20190 ( .A1(n3218), .A2(\xmem_data[76][6] ), .B1(n29065), .B2(
        \xmem_data[77][6] ), .ZN(n16054) );
  AOI22_X1 U20191 ( .A1(n29095), .A2(\xmem_data[78][6] ), .B1(n25490), .B2(
        \xmem_data[79][6] ), .ZN(n16053) );
  NAND4_X1 U20192 ( .A1(n16056), .A2(n16055), .A3(n16054), .A4(n16053), .ZN(
        n16057) );
  OR4_X1 U20193 ( .A1(n16060), .A2(n16059), .A3(n16058), .A4(n16057), .ZN(
        n16061) );
  AOI22_X1 U20194 ( .A1(n16062), .A2(n29171), .B1(n16061), .B2(n29201), .ZN(
        n16063) );
  XNOR2_X1 U20195 ( .A(n34982), .B(\fmem_data[25][3] ), .ZN(n33058) );
  AOI22_X1 U20196 ( .A1(n28428), .A2(\xmem_data[32][3] ), .B1(n30495), .B2(
        \xmem_data[33][3] ), .ZN(n16068) );
  AOI22_X1 U20197 ( .A1(n14974), .A2(\xmem_data[34][3] ), .B1(n23779), .B2(
        \xmem_data[35][3] ), .ZN(n16067) );
  AOI22_X1 U20198 ( .A1(n30497), .A2(\xmem_data[36][3] ), .B1(n30496), .B2(
        \xmem_data[37][3] ), .ZN(n16066) );
  AOI22_X1 U20199 ( .A1(n28036), .A2(\xmem_data[38][3] ), .B1(n30498), .B2(
        \xmem_data[39][3] ), .ZN(n16065) );
  AOI22_X1 U20200 ( .A1(n30503), .A2(\xmem_data[44][3] ), .B1(n3220), .B2(
        \xmem_data[45][3] ), .ZN(n16083) );
  AOI22_X1 U20201 ( .A1(n20994), .A2(\xmem_data[48][3] ), .B1(n3256), .B2(
        \xmem_data[49][3] ), .ZN(n16072) );
  AOI22_X1 U20202 ( .A1(n3375), .A2(\xmem_data[50][3] ), .B1(n25514), .B2(
        \xmem_data[51][3] ), .ZN(n16071) );
  AOI22_X1 U20203 ( .A1(n25422), .A2(\xmem_data[52][3] ), .B1(n20588), .B2(
        \xmem_data[53][3] ), .ZN(n16070) );
  AOI22_X1 U20204 ( .A1(n30508), .A2(\xmem_data[54][3] ), .B1(n22740), .B2(
        \xmem_data[55][3] ), .ZN(n16069) );
  NAND4_X1 U20205 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        n16077) );
  AOI22_X1 U20206 ( .A1(n27925), .A2(\xmem_data[40][3] ), .B1(n24573), .B2(
        \xmem_data[41][3] ), .ZN(n16075) );
  AOI22_X1 U20207 ( .A1(n24563), .A2(\xmem_data[46][3] ), .B1(n23739), .B2(
        \xmem_data[47][3] ), .ZN(n16074) );
  AOI22_X1 U20208 ( .A1(n22728), .A2(\xmem_data[42][3] ), .B1(n31347), .B2(
        \xmem_data[43][3] ), .ZN(n16073) );
  NOR2_X1 U20209 ( .A1(n16077), .A2(n16076), .ZN(n16082) );
  AOI22_X1 U20210 ( .A1(n30514), .A2(\xmem_data[56][3] ), .B1(n30513), .B2(
        \xmem_data[57][3] ), .ZN(n16081) );
  AOI22_X1 U20211 ( .A1(n27755), .A2(\xmem_data[58][3] ), .B1(n22742), .B2(
        \xmem_data[59][3] ), .ZN(n16080) );
  AOI22_X1 U20212 ( .A1(n31330), .A2(\xmem_data[60][3] ), .B1(n24645), .B2(
        \xmem_data[61][3] ), .ZN(n16079) );
  AOI22_X1 U20213 ( .A1(n30872), .A2(\xmem_data[62][3] ), .B1(n30515), .B2(
        \xmem_data[63][3] ), .ZN(n16078) );
  NAND4_X1 U20214 ( .A1(n3865), .A2(n16083), .A3(n16082), .A4(n3528), .ZN(
        n16084) );
  NAND2_X1 U20215 ( .A1(n16084), .A2(n30565), .ZN(n16155) );
  AOI22_X1 U20216 ( .A1(n30592), .A2(\xmem_data[108][3] ), .B1(n3218), .B2(
        \xmem_data[109][3] ), .ZN(n16088) );
  AOI22_X1 U20217 ( .A1(n3348), .A2(\xmem_data[106][3] ), .B1(n30589), .B2(
        \xmem_data[107][3] ), .ZN(n16087) );
  AOI22_X1 U20218 ( .A1(n30588), .A2(\xmem_data[104][3] ), .B1(n30571), .B2(
        \xmem_data[105][3] ), .ZN(n16086) );
  AOI22_X1 U20219 ( .A1(n30593), .A2(\xmem_data[110][3] ), .B1(n28356), .B2(
        \xmem_data[111][3] ), .ZN(n16085) );
  NAND4_X1 U20220 ( .A1(n16088), .A2(n16087), .A3(n16086), .A4(n16085), .ZN(
        n16106) );
  AOI22_X1 U20221 ( .A1(n3326), .A2(\xmem_data[96][3] ), .B1(n21051), .B2(
        \xmem_data[97][3] ), .ZN(n16092) );
  AOI22_X1 U20222 ( .A1(n30600), .A2(\xmem_data[98][3] ), .B1(n30599), .B2(
        \xmem_data[99][3] ), .ZN(n16091) );
  AOI22_X1 U20223 ( .A1(n20734), .A2(\xmem_data[100][3] ), .B1(n27526), .B2(
        \xmem_data[101][3] ), .ZN(n16090) );
  AOI22_X1 U20224 ( .A1(n29383), .A2(\xmem_data[102][3] ), .B1(n30601), .B2(
        \xmem_data[103][3] ), .ZN(n16089) );
  NAND4_X1 U20225 ( .A1(n16092), .A2(n16091), .A3(n16090), .A4(n16089), .ZN(
        n16104) );
  AOI22_X1 U20226 ( .A1(n30606), .A2(\xmem_data[112][3] ), .B1(n30882), .B2(
        \xmem_data[113][3] ), .ZN(n16096) );
  AOI22_X1 U20227 ( .A1(n3280), .A2(\xmem_data[114][3] ), .B1(n28045), .B2(
        \xmem_data[115][3] ), .ZN(n16095) );
  AOI22_X1 U20228 ( .A1(n30607), .A2(\xmem_data[116][3] ), .B1(n29180), .B2(
        \xmem_data[117][3] ), .ZN(n16094) );
  AOI22_X1 U20229 ( .A1(n30608), .A2(\xmem_data[118][3] ), .B1(n21015), .B2(
        \xmem_data[119][3] ), .ZN(n16093) );
  NAND4_X1 U20230 ( .A1(n16096), .A2(n16095), .A3(n16094), .A4(n16093), .ZN(
        n16102) );
  AOI22_X1 U20231 ( .A1(n30614), .A2(\xmem_data[120][3] ), .B1(n30613), .B2(
        \xmem_data[121][3] ), .ZN(n16100) );
  AOI22_X1 U20232 ( .A1(n21005), .A2(\xmem_data[122][3] ), .B1(n30615), .B2(
        \xmem_data[123][3] ), .ZN(n16099) );
  AOI22_X1 U20233 ( .A1(n24509), .A2(\xmem_data[124][3] ), .B1(n16989), .B2(
        \xmem_data[125][3] ), .ZN(n16098) );
  AOI22_X1 U20234 ( .A1(n30617), .A2(\xmem_data[126][3] ), .B1(n30616), .B2(
        \xmem_data[127][3] ), .ZN(n16097) );
  NAND4_X1 U20235 ( .A1(n16100), .A2(n16099), .A3(n16098), .A4(n16097), .ZN(
        n16101) );
  OR2_X1 U20236 ( .A1(n16102), .A2(n16101), .ZN(n16103) );
  OR2_X1 U20237 ( .A1(n16104), .A2(n16103), .ZN(n16105) );
  OAI21_X1 U20238 ( .B1(n16106), .B2(n16105), .A(n30626), .ZN(n16154) );
  AOI22_X1 U20239 ( .A1(n3178), .A2(\xmem_data[64][3] ), .B1(n27856), .B2(
        \xmem_data[65][3] ), .ZN(n16111) );
  AOI22_X1 U20240 ( .A1(n30600), .A2(\xmem_data[66][3] ), .B1(n30599), .B2(
        \xmem_data[67][3] ), .ZN(n16110) );
  AOI22_X1 U20241 ( .A1(n28293), .A2(\xmem_data[68][3] ), .B1(n28468), .B2(
        \xmem_data[69][3] ), .ZN(n16109) );
  AND2_X1 U20242 ( .A1(n30601), .A2(\xmem_data[71][3] ), .ZN(n16107) );
  AOI21_X1 U20243 ( .B1(n30754), .B2(\xmem_data[70][3] ), .A(n16107), .ZN(
        n16108) );
  AOI22_X1 U20244 ( .A1(n30588), .A2(\xmem_data[72][3] ), .B1(n30861), .B2(
        \xmem_data[73][3] ), .ZN(n16112) );
  INV_X1 U20245 ( .A(n16112), .ZN(n16116) );
  AOI22_X1 U20246 ( .A1(n30593), .A2(\xmem_data[78][3] ), .B1(n20558), .B2(
        \xmem_data[79][3] ), .ZN(n16114) );
  AOI22_X1 U20247 ( .A1(n3348), .A2(\xmem_data[74][3] ), .B1(n30589), .B2(
        \xmem_data[75][3] ), .ZN(n16113) );
  NAND2_X1 U20248 ( .A1(n16114), .A2(n16113), .ZN(n16115) );
  NOR2_X1 U20249 ( .A1(n16116), .A2(n16115), .ZN(n16129) );
  AOI22_X1 U20250 ( .A1(n30614), .A2(\xmem_data[88][3] ), .B1(n30613), .B2(
        \xmem_data[89][3] ), .ZN(n16120) );
  AOI22_X1 U20251 ( .A1(n23795), .A2(\xmem_data[90][3] ), .B1(n30615), .B2(
        \xmem_data[91][3] ), .ZN(n16119) );
  AOI22_X1 U20252 ( .A1(n23717), .A2(\xmem_data[92][3] ), .B1(n28492), .B2(
        \xmem_data[93][3] ), .ZN(n16118) );
  AOI22_X1 U20253 ( .A1(n30617), .A2(\xmem_data[94][3] ), .B1(n30616), .B2(
        \xmem_data[95][3] ), .ZN(n16117) );
  NAND4_X1 U20254 ( .A1(n16120), .A2(n16119), .A3(n16118), .A4(n16117), .ZN(
        n16126) );
  AOI22_X1 U20255 ( .A1(n30606), .A2(\xmem_data[80][3] ), .B1(n30882), .B2(
        \xmem_data[81][3] ), .ZN(n16124) );
  AOI22_X1 U20256 ( .A1(n24702), .A2(\xmem_data[82][3] ), .B1(n25450), .B2(
        \xmem_data[83][3] ), .ZN(n16123) );
  AOI22_X1 U20257 ( .A1(n30607), .A2(\xmem_data[84][3] ), .B1(n20982), .B2(
        \xmem_data[85][3] ), .ZN(n16122) );
  AOI22_X1 U20258 ( .A1(n30608), .A2(\xmem_data[86][3] ), .B1(n20958), .B2(
        \xmem_data[87][3] ), .ZN(n16121) );
  NAND4_X1 U20259 ( .A1(n16124), .A2(n16123), .A3(n16122), .A4(n16121), .ZN(
        n16125) );
  NOR2_X1 U20260 ( .A1(n16126), .A2(n16125), .ZN(n16128) );
  AOI22_X1 U20261 ( .A1(n30592), .A2(\xmem_data[76][3] ), .B1(n3220), .B2(
        \xmem_data[77][3] ), .ZN(n16127) );
  NAND4_X1 U20262 ( .A1(n3866), .A2(n16129), .A3(n16128), .A4(n16127), .ZN(
        n16130) );
  NAND2_X1 U20263 ( .A1(n16130), .A2(n30628), .ZN(n16153) );
  AOI22_X1 U20264 ( .A1(n30557), .A2(\xmem_data[0][3] ), .B1(n28494), .B2(
        \xmem_data[1][3] ), .ZN(n16134) );
  AOI22_X1 U20265 ( .A1(n28226), .A2(\xmem_data[2][3] ), .B1(n27975), .B2(
        \xmem_data[3][3] ), .ZN(n16133) );
  AOI22_X1 U20266 ( .A1(n3172), .A2(\xmem_data[4][3] ), .B1(n28292), .B2(
        \xmem_data[5][3] ), .ZN(n16132) );
  AOI22_X1 U20267 ( .A1(n27498), .A2(\xmem_data[6][3] ), .B1(n30524), .B2(
        \xmem_data[7][3] ), .ZN(n16131) );
  NAND4_X1 U20268 ( .A1(n16134), .A2(n16133), .A3(n16132), .A4(n16131), .ZN(
        n16150) );
  AOI22_X1 U20269 ( .A1(n24607), .A2(\xmem_data[8][3] ), .B1(n29118), .B2(
        \xmem_data[9][3] ), .ZN(n16138) );
  AOI22_X1 U20270 ( .A1(n3412), .A2(\xmem_data[10][3] ), .B1(n28501), .B2(
        \xmem_data[11][3] ), .ZN(n16137) );
  AOI22_X1 U20271 ( .A1(n25413), .A2(\xmem_data[12][3] ), .B1(n3222), .B2(
        \xmem_data[13][3] ), .ZN(n16136) );
  AOI22_X1 U20272 ( .A1(n20724), .A2(\xmem_data[14][3] ), .B1(n30534), .B2(
        \xmem_data[15][3] ), .ZN(n16135) );
  NAND4_X1 U20273 ( .A1(n16138), .A2(n16137), .A3(n16136), .A4(n16135), .ZN(
        n16149) );
  AOI22_X1 U20274 ( .A1(n25416), .A2(\xmem_data[16][3] ), .B1(n30550), .B2(
        \xmem_data[17][3] ), .ZN(n16142) );
  AOI22_X1 U20275 ( .A1(n24702), .A2(\xmem_data[18][3] ), .B1(n29045), .B2(
        \xmem_data[19][3] ), .ZN(n16141) );
  AOI22_X1 U20276 ( .A1(n30551), .A2(\xmem_data[20][3] ), .B1(n27943), .B2(
        \xmem_data[21][3] ), .ZN(n16140) );
  AOI22_X1 U20277 ( .A1(n20716), .A2(\xmem_data[22][3] ), .B1(n30552), .B2(
        \xmem_data[23][3] ), .ZN(n16139) );
  NAND4_X1 U20278 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        n16148) );
  AOI22_X1 U20279 ( .A1(n27537), .A2(\xmem_data[24][3] ), .B1(n30541), .B2(
        \xmem_data[25][3] ), .ZN(n16146) );
  AOI22_X1 U20280 ( .A1(n3119), .A2(\xmem_data[26][3] ), .B1(n30542), .B2(
        \xmem_data[27][3] ), .ZN(n16145) );
  AOI22_X1 U20281 ( .A1(n28337), .A2(\xmem_data[28][3] ), .B1(n30544), .B2(
        \xmem_data[29][3] ), .ZN(n16144) );
  AOI22_X1 U20282 ( .A1(n21008), .A2(\xmem_data[30][3] ), .B1(n30545), .B2(
        \xmem_data[31][3] ), .ZN(n16143) );
  NAND4_X1 U20283 ( .A1(n16146), .A2(n16145), .A3(n16144), .A4(n16143), .ZN(
        n16147) );
  OR4_X1 U20284 ( .A1(n16150), .A2(n16149), .A3(n16148), .A4(n16147), .ZN(
        n16151) );
  NAND2_X1 U20285 ( .A1(n16151), .A2(n30563), .ZN(n16152) );
  XNOR2_X1 U20286 ( .A(n31219), .B(\fmem_data[26][5] ), .ZN(n30387) );
  XNOR2_X1 U20287 ( .A(n3276), .B(\fmem_data[26][5] ), .ZN(n33045) );
  OAI22_X1 U20288 ( .A1(n30387), .A2(n35033), .B1(n33045), .B2(n35034), .ZN(
        n34076) );
  AOI22_X1 U20289 ( .A1(n16986), .A2(\xmem_data[96][1] ), .B1(n20798), .B2(
        \xmem_data[97][1] ), .ZN(n16159) );
  AOI22_X1 U20290 ( .A1(n16988), .A2(\xmem_data[98][1] ), .B1(n17019), .B2(
        \xmem_data[99][1] ), .ZN(n16158) );
  AOI22_X1 U20291 ( .A1(n21007), .A2(\xmem_data[100][1] ), .B1(n16989), .B2(
        \xmem_data[101][1] ), .ZN(n16157) );
  AOI22_X1 U20292 ( .A1(n16990), .A2(\xmem_data[102][1] ), .B1(n31360), .B2(
        \xmem_data[103][1] ), .ZN(n16156) );
  NAND4_X1 U20293 ( .A1(n16159), .A2(n16158), .A3(n16157), .A4(n16156), .ZN(
        n16176) );
  AOI22_X1 U20294 ( .A1(n30557), .A2(\xmem_data[104][1] ), .B1(n20943), .B2(
        \xmem_data[105][1] ), .ZN(n16163) );
  AOI22_X1 U20295 ( .A1(n3270), .A2(\xmem_data[106][1] ), .B1(n3201), .B2(
        \xmem_data[107][1] ), .ZN(n16162) );
  AOI22_X1 U20296 ( .A1(n25582), .A2(\xmem_data[108][1] ), .B1(n25723), .B2(
        \xmem_data[109][1] ), .ZN(n16161) );
  AOI22_X1 U20297 ( .A1(n25584), .A2(\xmem_data[110][1] ), .B1(n27567), .B2(
        \xmem_data[111][1] ), .ZN(n16160) );
  NAND4_X1 U20298 ( .A1(n16163), .A2(n16162), .A3(n16161), .A4(n16160), .ZN(
        n16175) );
  AOI22_X1 U20299 ( .A1(n28082), .A2(\xmem_data[116][1] ), .B1(n3217), .B2(
        \xmem_data[117][1] ), .ZN(n16168) );
  AOI22_X1 U20300 ( .A1(n30909), .A2(\xmem_data[112][1] ), .B1(n27499), .B2(
        \xmem_data[113][1] ), .ZN(n16167) );
  AOI22_X1 U20301 ( .A1(n21067), .A2(\xmem_data[118][1] ), .B1(n20723), .B2(
        \xmem_data[119][1] ), .ZN(n16165) );
  AOI22_X1 U20302 ( .A1(n16980), .A2(\xmem_data[114][1] ), .B1(n16979), .B2(
        \xmem_data[115][1] ), .ZN(n16164) );
  NAND3_X1 U20303 ( .A1(n16168), .A2(n16167), .A3(n16166), .ZN(n16174) );
  AOI22_X1 U20304 ( .A1(n28083), .A2(\xmem_data[120][1] ), .B1(n30550), .B2(
        \xmem_data[121][1] ), .ZN(n16172) );
  AOI22_X1 U20305 ( .A1(n16973), .A2(\xmem_data[122][1] ), .B1(n16972), .B2(
        \xmem_data[123][1] ), .ZN(n16171) );
  AOI22_X1 U20306 ( .A1(n16974), .A2(\xmem_data[124][1] ), .B1(n29180), .B2(
        \xmem_data[125][1] ), .ZN(n16170) );
  AOI22_X1 U20307 ( .A1(n31327), .A2(\xmem_data[126][1] ), .B1(n20958), .B2(
        \xmem_data[127][1] ), .ZN(n16169) );
  NAND4_X1 U20308 ( .A1(n16172), .A2(n16171), .A3(n16170), .A4(n16169), .ZN(
        n16173) );
  OR4_X1 U20309 ( .A1(n16176), .A2(n16175), .A3(n16174), .A4(n16173), .ZN(
        n16198) );
  AOI22_X1 U20310 ( .A1(n16986), .A2(\xmem_data[64][1] ), .B1(n21076), .B2(
        \xmem_data[65][1] ), .ZN(n16180) );
  AOI22_X1 U20311 ( .A1(n16988), .A2(\xmem_data[66][1] ), .B1(n17019), .B2(
        \xmem_data[67][1] ), .ZN(n16179) );
  AOI22_X1 U20312 ( .A1(n23717), .A2(\xmem_data[68][1] ), .B1(n16989), .B2(
        \xmem_data[69][1] ), .ZN(n16178) );
  AOI22_X1 U20313 ( .A1(n16990), .A2(\xmem_data[70][1] ), .B1(n25399), .B2(
        \xmem_data[71][1] ), .ZN(n16177) );
  NAND4_X1 U20314 ( .A1(n16180), .A2(n16179), .A3(n16178), .A4(n16177), .ZN(
        n16196) );
  AOI22_X1 U20315 ( .A1(n29240), .A2(\xmem_data[72][1] ), .B1(n30495), .B2(
        \xmem_data[73][1] ), .ZN(n16184) );
  AOI22_X1 U20316 ( .A1(n3271), .A2(\xmem_data[74][1] ), .B1(n3199), .B2(
        \xmem_data[75][1] ), .ZN(n16183) );
  AOI22_X1 U20317 ( .A1(n24685), .A2(\xmem_data[76][1] ), .B1(n29247), .B2(
        \xmem_data[77][1] ), .ZN(n16182) );
  AOI22_X1 U20318 ( .A1(n25628), .A2(\xmem_data[78][1] ), .B1(n30601), .B2(
        \xmem_data[79][1] ), .ZN(n16181) );
  NAND4_X1 U20319 ( .A1(n16184), .A2(n16183), .A3(n16182), .A4(n16181), .ZN(
        n16195) );
  AOI22_X1 U20320 ( .A1(n28082), .A2(\xmem_data[84][1] ), .B1(n3222), .B2(
        \xmem_data[85][1] ), .ZN(n16188) );
  AOI22_X1 U20321 ( .A1(n16980), .A2(\xmem_data[82][1] ), .B1(n16979), .B2(
        \xmem_data[83][1] ), .ZN(n16187) );
  AOI22_X1 U20322 ( .A1(n24526), .A2(\xmem_data[80][1] ), .B1(n31262), .B2(
        \xmem_data[81][1] ), .ZN(n16186) );
  AOI22_X1 U20323 ( .A1(n31368), .A2(\xmem_data[86][1] ), .B1(n20500), .B2(
        \xmem_data[87][1] ), .ZN(n16185) );
  NAND4_X1 U20324 ( .A1(n16188), .A2(n16187), .A3(n16186), .A4(n16185), .ZN(
        n16194) );
  AOI22_X1 U20325 ( .A1(n3342), .A2(\xmem_data[88][1] ), .B1(n22711), .B2(
        \xmem_data[89][1] ), .ZN(n16192) );
  AOI22_X1 U20326 ( .A1(n16973), .A2(\xmem_data[90][1] ), .B1(n16972), .B2(
        \xmem_data[91][1] ), .ZN(n16191) );
  AOI22_X1 U20327 ( .A1(n16974), .A2(\xmem_data[92][1] ), .B1(n29180), .B2(
        \xmem_data[93][1] ), .ZN(n16190) );
  AOI22_X1 U20328 ( .A1(n30886), .A2(\xmem_data[94][1] ), .B1(n24516), .B2(
        \xmem_data[95][1] ), .ZN(n16189) );
  NAND4_X1 U20329 ( .A1(n16192), .A2(n16191), .A3(n16190), .A4(n16189), .ZN(
        n16193) );
  OR4_X1 U20330 ( .A1(n16196), .A2(n16195), .A3(n16194), .A4(n16193), .ZN(
        n16197) );
  AOI22_X1 U20331 ( .A1(n16997), .A2(n16198), .B1(n16966), .B2(n16197), .ZN(
        n16247) );
  AOI22_X1 U20332 ( .A1(n16986), .A2(\xmem_data[32][1] ), .B1(n22741), .B2(
        \xmem_data[33][1] ), .ZN(n16202) );
  AOI22_X1 U20333 ( .A1(n27945), .A2(\xmem_data[34][1] ), .B1(n16987), .B2(
        \xmem_data[35][1] ), .ZN(n16201) );
  AOI22_X1 U20334 ( .A1(n17020), .A2(\xmem_data[36][1] ), .B1(n31355), .B2(
        \xmem_data[37][1] ), .ZN(n16200) );
  AOI22_X1 U20335 ( .A1(n17021), .A2(\xmem_data[38][1] ), .B1(n24592), .B2(
        \xmem_data[39][1] ), .ZN(n16199) );
  NAND4_X1 U20336 ( .A1(n16202), .A2(n16201), .A3(n16200), .A4(n16199), .ZN(
        n16218) );
  AOI22_X1 U20337 ( .A1(n24220), .A2(\xmem_data[40][1] ), .B1(n17001), .B2(
        \xmem_data[41][1] ), .ZN(n16206) );
  AOI22_X1 U20338 ( .A1(n17004), .A2(\xmem_data[42][1] ), .B1(n3199), .B2(
        \xmem_data[43][1] ), .ZN(n16205) );
  AOI22_X1 U20339 ( .A1(n22719), .A2(\xmem_data[44][1] ), .B1(n17003), .B2(
        \xmem_data[45][1] ), .ZN(n16204) );
  AOI22_X1 U20340 ( .A1(n30754), .A2(\xmem_data[46][1] ), .B1(n16999), .B2(
        \xmem_data[47][1] ), .ZN(n16203) );
  NAND4_X1 U20341 ( .A1(n16206), .A2(n16205), .A3(n16204), .A4(n16203), .ZN(
        n16217) );
  AOI22_X1 U20342 ( .A1(n17030), .A2(\xmem_data[48][1] ), .B1(n28317), .B2(
        \xmem_data[49][1] ), .ZN(n16210) );
  AOI22_X1 U20343 ( .A1(n3388), .A2(\xmem_data[50][1] ), .B1(n17031), .B2(
        \xmem_data[51][1] ), .ZN(n16209) );
  AOI22_X1 U20344 ( .A1(n28044), .A2(\xmem_data[52][1] ), .B1(n3220), .B2(
        \xmem_data[53][1] ), .ZN(n16208) );
  AOI22_X1 U20345 ( .A1(n17033), .A2(\xmem_data[54][1] ), .B1(n24207), .B2(
        \xmem_data[55][1] ), .ZN(n16207) );
  NAND4_X1 U20346 ( .A1(n16210), .A2(n16209), .A3(n16208), .A4(n16207), .ZN(
        n16216) );
  AOI22_X1 U20347 ( .A1(n17010), .A2(\xmem_data[56][1] ), .B1(n25486), .B2(
        \xmem_data[57][1] ), .ZN(n16214) );
  AOI22_X1 U20348 ( .A1(n21074), .A2(\xmem_data[58][1] ), .B1(n17011), .B2(
        \xmem_data[59][1] ), .ZN(n16213) );
  AOI22_X1 U20349 ( .A1(n25670), .A2(\xmem_data[60][1] ), .B1(n29180), .B2(
        \xmem_data[61][1] ), .ZN(n16212) );
  AOI22_X1 U20350 ( .A1(n17013), .A2(\xmem_data[62][1] ), .B1(n17012), .B2(
        \xmem_data[63][1] ), .ZN(n16211) );
  NAND4_X1 U20351 ( .A1(n16214), .A2(n16213), .A3(n16212), .A4(n16211), .ZN(
        n16215) );
  OR4_X1 U20352 ( .A1(n16218), .A2(n16217), .A3(n16216), .A4(n16215), .ZN(
        n16245) );
  AOI22_X1 U20353 ( .A1(n3177), .A2(\xmem_data[8][1] ), .B1(n25716), .B2(
        \xmem_data[9][1] ), .ZN(n16222) );
  AOI22_X1 U20354 ( .A1(n24623), .A2(\xmem_data[10][1] ), .B1(n3199), .B2(
        \xmem_data[11][1] ), .ZN(n16221) );
  AOI22_X1 U20355 ( .A1(n21058), .A2(\xmem_data[12][1] ), .B1(n17049), .B2(
        \xmem_data[13][1] ), .ZN(n16220) );
  AOI22_X1 U20356 ( .A1(n17051), .A2(\xmem_data[14][1] ), .B1(n17050), .B2(
        \xmem_data[15][1] ), .ZN(n16219) );
  AND4_X1 U20357 ( .A1(n16222), .A2(n16221), .A3(n16220), .A4(n16219), .ZN(
        n16243) );
  NAND2_X1 U20358 ( .A1(n17041), .A2(\xmem_data[0][1] ), .ZN(n16242) );
  AOI22_X1 U20359 ( .A1(n25694), .A2(\xmem_data[24][1] ), .B1(n17061), .B2(
        \xmem_data[25][1] ), .ZN(n16226) );
  AOI22_X1 U20360 ( .A1(n17063), .A2(\xmem_data[26][1] ), .B1(n17062), .B2(
        \xmem_data[27][1] ), .ZN(n16225) );
  AOI22_X1 U20361 ( .A1(n24554), .A2(\xmem_data[28][1] ), .B1(n22701), .B2(
        \xmem_data[29][1] ), .ZN(n16224) );
  AOI22_X1 U20362 ( .A1(n17064), .A2(\xmem_data[30][1] ), .B1(n24132), .B2(
        \xmem_data[31][1] ), .ZN(n16223) );
  NAND4_X1 U20363 ( .A1(n16226), .A2(n16225), .A3(n16224), .A4(n16223), .ZN(
        n16235) );
  AOI22_X1 U20364 ( .A1(n17044), .A2(\xmem_data[6][1] ), .B1(n29280), .B2(
        \xmem_data[7][1] ), .ZN(n16233) );
  AOI22_X1 U20365 ( .A1(n28059), .A2(\xmem_data[4][1] ), .B1(n17043), .B2(
        \xmem_data[5][1] ), .ZN(n16227) );
  INV_X1 U20366 ( .A(n16227), .ZN(n16231) );
  NAND2_X1 U20367 ( .A1(n25382), .A2(\xmem_data[1][1] ), .ZN(n16229) );
  AOI22_X1 U20368 ( .A1(n21005), .A2(\xmem_data[2][1] ), .B1(n3202), .B2(
        \xmem_data[3][1] ), .ZN(n16228) );
  NAND2_X1 U20369 ( .A1(n16229), .A2(n16228), .ZN(n16230) );
  NOR2_X1 U20370 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  NAND2_X1 U20371 ( .A1(n16233), .A2(n16232), .ZN(n16234) );
  NOR2_X1 U20372 ( .A1(n16235), .A2(n16234), .ZN(n16241) );
  AOI22_X1 U20373 ( .A1(n28470), .A2(\xmem_data[20][1] ), .B1(n3222), .B2(
        \xmem_data[21][1] ), .ZN(n16239) );
  AOI22_X1 U20374 ( .A1(n3434), .A2(\xmem_data[18][1] ), .B1(n16979), .B2(
        \xmem_data[19][1] ), .ZN(n16238) );
  AOI22_X1 U20375 ( .A1(n17056), .A2(\xmem_data[16][1] ), .B1(n28317), .B2(
        \xmem_data[17][1] ), .ZN(n16237) );
  AOI22_X1 U20376 ( .A1(n25612), .A2(\xmem_data[22][1] ), .B1(n27444), .B2(
        \xmem_data[23][1] ), .ZN(n16236) );
  AND4_X1 U20377 ( .A1(n16239), .A2(n16238), .A3(n16237), .A4(n16236), .ZN(
        n16240) );
  NAND4_X1 U20378 ( .A1(n16243), .A2(n16242), .A3(n16241), .A4(n16240), .ZN(
        n16244) );
  AOI22_X1 U20379 ( .A1(n16245), .A2(n17038), .B1(n17073), .B2(n16244), .ZN(
        n16246) );
  AOI22_X1 U20380 ( .A1(n31268), .A2(\xmem_data[32][2] ), .B1(n24160), .B2(
        \xmem_data[33][2] ), .ZN(n16251) );
  AOI22_X1 U20381 ( .A1(n27755), .A2(\xmem_data[34][2] ), .B1(n17019), .B2(
        \xmem_data[35][2] ), .ZN(n16250) );
  AOI22_X1 U20382 ( .A1(n17021), .A2(\xmem_data[38][2] ), .B1(n29238), .B2(
        \xmem_data[39][2] ), .ZN(n16249) );
  AOI22_X1 U20383 ( .A1(n17020), .A2(\xmem_data[36][2] ), .B1(n24546), .B2(
        \xmem_data[37][2] ), .ZN(n16248) );
  NAND4_X1 U20384 ( .A1(n16251), .A2(n16250), .A3(n16249), .A4(n16248), .ZN(
        n16257) );
  AOI22_X1 U20385 ( .A1(n17010), .A2(\xmem_data[56][2] ), .B1(n28372), .B2(
        \xmem_data[57][2] ), .ZN(n16255) );
  AOI22_X1 U20386 ( .A1(n25732), .A2(\xmem_data[58][2] ), .B1(n17011), .B2(
        \xmem_data[59][2] ), .ZN(n16254) );
  AOI22_X1 U20387 ( .A1(n23813), .A2(\xmem_data[60][2] ), .B1(n28481), .B2(
        \xmem_data[61][2] ), .ZN(n16253) );
  AOI22_X1 U20388 ( .A1(n17013), .A2(\xmem_data[62][2] ), .B1(n17012), .B2(
        \xmem_data[63][2] ), .ZN(n16252) );
  NAND4_X1 U20389 ( .A1(n16255), .A2(n16254), .A3(n16253), .A4(n16252), .ZN(
        n16256) );
  OR2_X1 U20390 ( .A1(n16257), .A2(n16256), .ZN(n16264) );
  AOI22_X1 U20391 ( .A1(n20593), .A2(\xmem_data[40][2] ), .B1(n17001), .B2(
        \xmem_data[41][2] ), .ZN(n16262) );
  AOI22_X1 U20392 ( .A1(n17004), .A2(\xmem_data[42][2] ), .B1(n3201), .B2(
        \xmem_data[43][2] ), .ZN(n16261) );
  AOI22_X1 U20393 ( .A1(n27847), .A2(\xmem_data[44][2] ), .B1(n17003), .B2(
        \xmem_data[45][2] ), .ZN(n16260) );
  AND2_X1 U20394 ( .A1(n16999), .A2(\xmem_data[47][2] ), .ZN(n16258) );
  AOI21_X1 U20395 ( .B1(n27498), .B2(\xmem_data[46][2] ), .A(n16258), .ZN(
        n16259) );
  NAND4_X1 U20396 ( .A1(n16262), .A2(n16261), .A3(n16260), .A4(n16259), .ZN(
        n16263) );
  OR2_X1 U20397 ( .A1(n16264), .A2(n16263), .ZN(n16273) );
  AOI22_X1 U20398 ( .A1(n27439), .A2(\xmem_data[52][2] ), .B1(n3220), .B2(
        \xmem_data[53][2] ), .ZN(n16271) );
  AOI22_X1 U20399 ( .A1(n17030), .A2(\xmem_data[48][2] ), .B1(n25561), .B2(
        \xmem_data[49][2] ), .ZN(n16270) );
  AOI22_X1 U20400 ( .A1(n17033), .A2(\xmem_data[54][2] ), .B1(n25562), .B2(
        \xmem_data[55][2] ), .ZN(n16265) );
  INV_X1 U20401 ( .A(n16265), .ZN(n16268) );
  AOI22_X1 U20402 ( .A1(n3387), .A2(\xmem_data[50][2] ), .B1(n17031), .B2(
        \xmem_data[51][2] ), .ZN(n16266) );
  INV_X1 U20403 ( .A(n16266), .ZN(n16267) );
  NOR2_X1 U20404 ( .A1(n16268), .A2(n16267), .ZN(n16269) );
  OAI21_X1 U20405 ( .B1(n16273), .B2(n16272), .A(n17038), .ZN(n16351) );
  AOI22_X1 U20406 ( .A1(n30956), .A2(\xmem_data[104][2] ), .B1(n14882), .B2(
        \xmem_data[105][2] ), .ZN(n16277) );
  AOI22_X1 U20407 ( .A1(n3270), .A2(\xmem_data[106][2] ), .B1(n3199), .B2(
        \xmem_data[107][2] ), .ZN(n16276) );
  AOI22_X1 U20408 ( .A1(n24166), .A2(\xmem_data[108][2] ), .B1(n25723), .B2(
        \xmem_data[109][2] ), .ZN(n16275) );
  AOI22_X1 U20409 ( .A1(n23730), .A2(\xmem_data[110][2] ), .B1(n31344), .B2(
        \xmem_data[111][2] ), .ZN(n16274) );
  NAND4_X1 U20410 ( .A1(n16277), .A2(n16276), .A3(n16275), .A4(n16274), .ZN(
        n16280) );
  AOI22_X1 U20411 ( .A1(n25686), .A2(\xmem_data[112][2] ), .B1(n30908), .B2(
        \xmem_data[113][2] ), .ZN(n16278) );
  INV_X1 U20412 ( .A(n16278), .ZN(n16279) );
  NOR2_X1 U20413 ( .A1(n16280), .A2(n16279), .ZN(n16295) );
  AOI22_X1 U20414 ( .A1(n16986), .A2(\xmem_data[96][2] ), .B1(n29046), .B2(
        \xmem_data[97][2] ), .ZN(n16284) );
  AOI22_X1 U20415 ( .A1(n16988), .A2(\xmem_data[98][2] ), .B1(n3202), .B2(
        \xmem_data[99][2] ), .ZN(n16283) );
  AOI22_X1 U20416 ( .A1(n22676), .A2(\xmem_data[100][2] ), .B1(n16989), .B2(
        \xmem_data[101][2] ), .ZN(n16282) );
  AOI22_X1 U20417 ( .A1(n16990), .A2(\xmem_data[102][2] ), .B1(n23801), .B2(
        \xmem_data[103][2] ), .ZN(n16281) );
  NAND4_X1 U20418 ( .A1(n16284), .A2(n16283), .A3(n16282), .A4(n16281), .ZN(
        n16288) );
  AOI22_X1 U20419 ( .A1(n28367), .A2(\xmem_data[118][2] ), .B1(n27507), .B2(
        \xmem_data[119][2] ), .ZN(n16286) );
  AOI22_X1 U20420 ( .A1(n16980), .A2(\xmem_data[114][2] ), .B1(n16979), .B2(
        \xmem_data[115][2] ), .ZN(n16285) );
  NAND2_X1 U20421 ( .A1(n16286), .A2(n16285), .ZN(n16287) );
  NOR2_X1 U20422 ( .A1(n16288), .A2(n16287), .ZN(n16294) );
  AOI22_X1 U20423 ( .A1(n20576), .A2(\xmem_data[116][2] ), .B1(n3222), .B2(
        \xmem_data[117][2] ), .ZN(n16293) );
  AOI22_X1 U20424 ( .A1(n22666), .A2(\xmem_data[120][2] ), .B1(n28372), .B2(
        \xmem_data[121][2] ), .ZN(n16292) );
  AOI22_X1 U20425 ( .A1(n16973), .A2(\xmem_data[122][2] ), .B1(n16972), .B2(
        \xmem_data[123][2] ), .ZN(n16291) );
  AOI22_X1 U20426 ( .A1(n16974), .A2(\xmem_data[124][2] ), .B1(n24590), .B2(
        \xmem_data[125][2] ), .ZN(n16290) );
  AOI22_X1 U20427 ( .A1(n31327), .A2(\xmem_data[126][2] ), .B1(n28345), .B2(
        \xmem_data[127][2] ), .ZN(n16289) );
  NAND4_X1 U20428 ( .A1(n16295), .A2(n16294), .A3(n16293), .A4(n3760), .ZN(
        n16296) );
  NAND2_X1 U20429 ( .A1(n16296), .A2(n16997), .ZN(n16350) );
  AOI22_X1 U20430 ( .A1(n17056), .A2(\xmem_data[16][2] ), .B1(n12471), .B2(
        \xmem_data[17][2] ), .ZN(n16300) );
  AOI22_X1 U20431 ( .A1(n3388), .A2(\xmem_data[18][2] ), .B1(n16979), .B2(
        \xmem_data[19][2] ), .ZN(n16299) );
  AOI22_X1 U20432 ( .A1(n28355), .A2(\xmem_data[20][2] ), .B1(n3218), .B2(
        \xmem_data[21][2] ), .ZN(n16298) );
  AOI22_X1 U20433 ( .A1(n24563), .A2(\xmem_data[22][2] ), .B1(n28508), .B2(
        \xmem_data[23][2] ), .ZN(n16297) );
  NAND4_X1 U20434 ( .A1(n16300), .A2(n16299), .A3(n16298), .A4(n16297), .ZN(
        n16322) );
  AOI22_X1 U20435 ( .A1(n20818), .A2(\xmem_data[12][2] ), .B1(n17049), .B2(
        \xmem_data[13][2] ), .ZN(n16302) );
  NAND2_X1 U20436 ( .A1(n17051), .A2(\xmem_data[14][2] ), .ZN(n16301) );
  AOI22_X1 U20437 ( .A1(n31328), .A2(\xmem_data[2][2] ), .B1(n17019), .B2(
        \xmem_data[3][2] ), .ZN(n16304) );
  AOI22_X1 U20438 ( .A1(n24511), .A2(\xmem_data[8][2] ), .B1(n28327), .B2(
        \xmem_data[9][2] ), .ZN(n16303) );
  NAND2_X1 U20439 ( .A1(n16304), .A2(n16303), .ZN(n16308) );
  AOI22_X1 U20440 ( .A1(n30645), .A2(\xmem_data[10][2] ), .B1(n3199), .B2(
        \xmem_data[11][2] ), .ZN(n16306) );
  NAND2_X1 U20441 ( .A1(n17050), .A2(\xmem_data[15][2] ), .ZN(n16305) );
  NAND2_X1 U20442 ( .A1(n16306), .A2(n16305), .ZN(n16307) );
  AOI22_X1 U20443 ( .A1(n27938), .A2(\xmem_data[24][2] ), .B1(n17061), .B2(
        \xmem_data[25][2] ), .ZN(n16312) );
  AOI22_X1 U20444 ( .A1(n17063), .A2(\xmem_data[26][2] ), .B1(n17062), .B2(
        \xmem_data[27][2] ), .ZN(n16311) );
  AOI22_X1 U20445 ( .A1(n25422), .A2(\xmem_data[28][2] ), .B1(n20982), .B2(
        \xmem_data[29][2] ), .ZN(n16310) );
  AOI22_X1 U20446 ( .A1(n17064), .A2(\xmem_data[30][2] ), .B1(n31326), .B2(
        \xmem_data[31][2] ), .ZN(n16309) );
  AOI22_X1 U20447 ( .A1(n17041), .A2(\xmem_data[0][2] ), .B1(n30541), .B2(
        \xmem_data[1][2] ), .ZN(n16313) );
  INV_X1 U20448 ( .A(n16313), .ZN(n16317) );
  AOI22_X1 U20449 ( .A1(n28096), .A2(\xmem_data[4][2] ), .B1(n17043), .B2(
        \xmem_data[5][2] ), .ZN(n16315) );
  AOI22_X1 U20450 ( .A1(n17044), .A2(\xmem_data[6][2] ), .B1(n29190), .B2(
        \xmem_data[7][2] ), .ZN(n16314) );
  NAND2_X1 U20451 ( .A1(n16315), .A2(n16314), .ZN(n16316) );
  NOR2_X1 U20452 ( .A1(n16317), .A2(n16316), .ZN(n16318) );
  OAI21_X1 U20453 ( .B1(n16322), .B2(n16321), .A(n17073), .ZN(n16349) );
  AND2_X1 U20454 ( .A1(n28354), .A2(\xmem_data[80][2] ), .ZN(n16323) );
  AOI21_X1 U20455 ( .B1(n20709), .B2(\xmem_data[81][2] ), .A(n16323), .ZN(
        n16324) );
  INV_X1 U20456 ( .A(n16324), .ZN(n16331) );
  AOI22_X1 U20457 ( .A1(n28493), .A2(\xmem_data[72][2] ), .B1(n28494), .B2(
        \xmem_data[73][2] ), .ZN(n16329) );
  AOI22_X1 U20458 ( .A1(n3270), .A2(\xmem_data[74][2] ), .B1(n3201), .B2(
        \xmem_data[75][2] ), .ZN(n16328) );
  AOI22_X1 U20459 ( .A1(n3172), .A2(\xmem_data[76][2] ), .B1(n28468), .B2(
        \xmem_data[77][2] ), .ZN(n16327) );
  AND2_X1 U20460 ( .A1(n31261), .A2(\xmem_data[79][2] ), .ZN(n16325) );
  AOI21_X1 U20461 ( .B1(n29383), .B2(\xmem_data[78][2] ), .A(n16325), .ZN(
        n16326) );
  NAND4_X1 U20462 ( .A1(n16329), .A2(n16328), .A3(n16327), .A4(n16326), .ZN(
        n16330) );
  AOI22_X1 U20463 ( .A1(n16986), .A2(\xmem_data[64][2] ), .B1(n27912), .B2(
        \xmem_data[65][2] ), .ZN(n16335) );
  AOI22_X1 U20464 ( .A1(n16988), .A2(\xmem_data[66][2] ), .B1(n16987), .B2(
        \xmem_data[67][2] ), .ZN(n16334) );
  AOI22_X1 U20465 ( .A1(n23764), .A2(\xmem_data[68][2] ), .B1(n16989), .B2(
        \xmem_data[69][2] ), .ZN(n16333) );
  AOI22_X1 U20466 ( .A1(n16990), .A2(\xmem_data[70][2] ), .B1(n24460), .B2(
        \xmem_data[71][2] ), .ZN(n16332) );
  NAND4_X1 U20467 ( .A1(n16335), .A2(n16334), .A3(n16333), .A4(n16332), .ZN(
        n16339) );
  AOI22_X1 U20468 ( .A1(n30964), .A2(\xmem_data[86][2] ), .B1(n20598), .B2(
        \xmem_data[87][2] ), .ZN(n16337) );
  AOI22_X1 U20469 ( .A1(n16980), .A2(\xmem_data[82][2] ), .B1(n16979), .B2(
        \xmem_data[83][2] ), .ZN(n16336) );
  NAND2_X1 U20470 ( .A1(n16337), .A2(n16336), .ZN(n16338) );
  NOR2_X1 U20471 ( .A1(n16339), .A2(n16338), .ZN(n16345) );
  AOI22_X1 U20472 ( .A1(n25449), .A2(\xmem_data[88][2] ), .B1(n31275), .B2(
        \xmem_data[89][2] ), .ZN(n16343) );
  AOI22_X1 U20473 ( .A1(n16973), .A2(\xmem_data[90][2] ), .B1(n16972), .B2(
        \xmem_data[91][2] ), .ZN(n16342) );
  AOI22_X1 U20474 ( .A1(n16974), .A2(\xmem_data[92][2] ), .B1(n29180), .B2(
        \xmem_data[93][2] ), .ZN(n16341) );
  AOI22_X1 U20475 ( .A1(n24157), .A2(\xmem_data[94][2] ), .B1(n31326), .B2(
        \xmem_data[95][2] ), .ZN(n16340) );
  AOI22_X1 U20476 ( .A1(n23756), .A2(\xmem_data[84][2] ), .B1(n3222), .B2(
        \xmem_data[85][2] ), .ZN(n16344) );
  NAND3_X1 U20477 ( .A1(n16345), .A2(n3801), .A3(n16344), .ZN(n16346) );
  OAI21_X1 U20478 ( .B1(n16347), .B2(n16346), .A(n16966), .ZN(n16348) );
  XNOR2_X1 U20479 ( .A(n32787), .B(\fmem_data[2][7] ), .ZN(n32018) );
  OAI22_X1 U20480 ( .A1(n22777), .A2(n35721), .B1(n35722), .B2(n32018), .ZN(
        n34075) );
  OAI21_X1 U20481 ( .B1(n3259), .B2(n18725), .A(n18727), .ZN(n16353) );
  NAND2_X1 U20482 ( .A1(n3259), .A2(n18725), .ZN(n16352) );
  NAND2_X1 U20483 ( .A1(n16353), .A2(n16352), .ZN(n31843) );
  FA_X1 U20484 ( .A(n16356), .B(n16355), .CI(n16354), .CO(n31845), .S(n26263)
         );
  XNOR2_X1 U20485 ( .A(n35256), .B(\fmem_data[31][1] ), .ZN(n32178) );
  AOI22_X1 U20486 ( .A1(n22719), .A2(\xmem_data[104][3] ), .B1(n25406), .B2(
        \xmem_data[105][3] ), .ZN(n16363) );
  AOI22_X1 U20487 ( .A1(n25407), .A2(\xmem_data[106][3] ), .B1(n24468), .B2(
        \xmem_data[107][3] ), .ZN(n16362) );
  AND2_X1 U20488 ( .A1(n25408), .A2(\xmem_data[108][3] ), .ZN(n16359) );
  AOI21_X1 U20489 ( .B1(n31309), .B2(\xmem_data[109][3] ), .A(n16359), .ZN(
        n16361) );
  AOI22_X1 U20490 ( .A1(n3318), .A2(\xmem_data[110][3] ), .B1(n24172), .B2(
        \xmem_data[111][3] ), .ZN(n16360) );
  AND4_X1 U20491 ( .A1(n16363), .A2(n16362), .A3(n16361), .A4(n16360), .ZN(
        n16377) );
  AOI22_X1 U20492 ( .A1(n25422), .A2(\xmem_data[120][3] ), .B1(n22701), .B2(
        \xmem_data[121][3] ), .ZN(n16367) );
  AOI22_X1 U20493 ( .A1(n25424), .A2(\xmem_data[122][3] ), .B1(n25423), .B2(
        \xmem_data[123][3] ), .ZN(n16366) );
  AOI22_X1 U20494 ( .A1(n25425), .A2(\xmem_data[124][3] ), .B1(n25606), .B2(
        \xmem_data[125][3] ), .ZN(n16365) );
  AOI22_X1 U20495 ( .A1(n29396), .A2(\xmem_data[126][3] ), .B1(n20586), .B2(
        \xmem_data[127][3] ), .ZN(n16364) );
  NAND4_X1 U20496 ( .A1(n16367), .A2(n16366), .A3(n16365), .A4(n16364), .ZN(
        n16375) );
  AOI22_X1 U20497 ( .A1(n25413), .A2(\xmem_data[112][3] ), .B1(n3221), .B2(
        \xmem_data[113][3] ), .ZN(n16368) );
  INV_X1 U20498 ( .A(n16368), .ZN(n16374) );
  AOI22_X1 U20499 ( .A1(n25416), .A2(\xmem_data[116][3] ), .B1(n25415), .B2(
        \xmem_data[117][3] ), .ZN(n16369) );
  INV_X1 U20500 ( .A(n16369), .ZN(n16373) );
  AOI22_X1 U20501 ( .A1(n25414), .A2(\xmem_data[114][3] ), .B1(n20558), .B2(
        \xmem_data[115][3] ), .ZN(n16371) );
  NAND2_X1 U20502 ( .A1(n25417), .A2(\xmem_data[118][3] ), .ZN(n16370) );
  NAND2_X1 U20503 ( .A1(n16371), .A2(n16370), .ZN(n16372) );
  NOR3_X1 U20504 ( .A1(n16375), .A2(n16374), .A3(n3996), .ZN(n16376) );
  NAND2_X1 U20505 ( .A1(n16377), .A2(n16376), .ZN(n16383) );
  AOI22_X1 U20506 ( .A1(n31330), .A2(\xmem_data[96][3] ), .B1(n25398), .B2(
        \xmem_data[97][3] ), .ZN(n16381) );
  AOI22_X1 U20507 ( .A1(n25400), .A2(\xmem_data[98][3] ), .B1(n25399), .B2(
        \xmem_data[99][3] ), .ZN(n16380) );
  AOI22_X1 U20508 ( .A1(n24190), .A2(\xmem_data[100][3] ), .B1(n28060), .B2(
        \xmem_data[101][3] ), .ZN(n16379) );
  AOI22_X1 U20509 ( .A1(n25401), .A2(\xmem_data[102][3] ), .B1(n14975), .B2(
        \xmem_data[103][3] ), .ZN(n16378) );
  NAND4_X1 U20510 ( .A1(n16381), .A2(n16380), .A3(n16379), .A4(n16378), .ZN(
        n16382) );
  OAI21_X1 U20511 ( .B1(n3963), .B2(n3498), .A(n25473), .ZN(n16412) );
  NAND2_X1 U20512 ( .A1(n3231), .A2(\xmem_data[87][3] ), .ZN(n16409) );
  AOI22_X1 U20513 ( .A1(n31316), .A2(\xmem_data[72][3] ), .B1(n25406), .B2(
        \xmem_data[73][3] ), .ZN(n16387) );
  AOI22_X1 U20514 ( .A1(n25407), .A2(\xmem_data[74][3] ), .B1(n24122), .B2(
        \xmem_data[75][3] ), .ZN(n16386) );
  AOI22_X1 U20515 ( .A1(n25408), .A2(\xmem_data[76][3] ), .B1(n25561), .B2(
        \xmem_data[77][3] ), .ZN(n16385) );
  AOI22_X1 U20516 ( .A1(n3318), .A2(\xmem_data[78][3] ), .B1(n27501), .B2(
        \xmem_data[79][3] ), .ZN(n16384) );
  AND4_X1 U20517 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        n16395) );
  AOI22_X1 U20518 ( .A1(n25413), .A2(\xmem_data[80][3] ), .B1(n3221), .B2(
        \xmem_data[81][3] ), .ZN(n16394) );
  AOI22_X1 U20519 ( .A1(n25416), .A2(\xmem_data[84][3] ), .B1(n25415), .B2(
        \xmem_data[85][3] ), .ZN(n16388) );
  INV_X1 U20520 ( .A(n16388), .ZN(n16392) );
  AOI22_X1 U20521 ( .A1(n25414), .A2(\xmem_data[82][3] ), .B1(n20500), .B2(
        \xmem_data[83][3] ), .ZN(n16390) );
  NAND2_X1 U20522 ( .A1(n25417), .A2(\xmem_data[86][3] ), .ZN(n16389) );
  NAND2_X1 U20523 ( .A1(n16390), .A2(n16389), .ZN(n16391) );
  NOR2_X1 U20524 ( .A1(n16392), .A2(n16391), .ZN(n16393) );
  NAND3_X1 U20525 ( .A1(n16395), .A2(n16394), .A3(n16393), .ZN(n16407) );
  AOI22_X1 U20526 ( .A1(n25422), .A2(\xmem_data[88][3] ), .B1(n20546), .B2(
        \xmem_data[89][3] ), .ZN(n16399) );
  AOI22_X1 U20527 ( .A1(n25424), .A2(\xmem_data[90][3] ), .B1(n25423), .B2(
        \xmem_data[91][3] ), .ZN(n16398) );
  AOI22_X1 U20528 ( .A1(n25425), .A2(\xmem_data[92][3] ), .B1(n28090), .B2(
        \xmem_data[93][3] ), .ZN(n16397) );
  AOI22_X1 U20529 ( .A1(n24458), .A2(\xmem_data[94][3] ), .B1(n31269), .B2(
        \xmem_data[95][3] ), .ZN(n16396) );
  NAND4_X1 U20530 ( .A1(n16399), .A2(n16398), .A3(n16397), .A4(n16396), .ZN(
        n16405) );
  AOI22_X1 U20531 ( .A1(n21007), .A2(\xmem_data[64][3] ), .B1(n25398), .B2(
        \xmem_data[65][3] ), .ZN(n16403) );
  AOI22_X1 U20532 ( .A1(n25400), .A2(\xmem_data[66][3] ), .B1(n25399), .B2(
        \xmem_data[67][3] ), .ZN(n16402) );
  AOI22_X1 U20533 ( .A1(n3178), .A2(\xmem_data[68][3] ), .B1(n21051), .B2(
        \xmem_data[69][3] ), .ZN(n16401) );
  AOI22_X1 U20534 ( .A1(n25401), .A2(\xmem_data[70][3] ), .B1(n14975), .B2(
        \xmem_data[71][3] ), .ZN(n16400) );
  NAND4_X1 U20535 ( .A1(n16403), .A2(n16402), .A3(n16401), .A4(n16400), .ZN(
        n16404) );
  NAND2_X1 U20536 ( .A1(n16409), .A2(n16408), .ZN(n16410) );
  NAND2_X1 U20537 ( .A1(n16410), .A2(n25471), .ZN(n16411) );
  NAND2_X1 U20538 ( .A1(n16412), .A2(n16411), .ZN(n16468) );
  NAND2_X1 U20539 ( .A1(n25450), .A2(\xmem_data[23][3] ), .ZN(n16442) );
  AOI22_X1 U20540 ( .A1(n17041), .A2(\xmem_data[28][3] ), .B1(n25382), .B2(
        \xmem_data[29][3] ), .ZN(n16431) );
  AOI22_X1 U20541 ( .A1(n17002), .A2(\xmem_data[4][3] ), .B1(n25364), .B2(
        \xmem_data[5][3] ), .ZN(n16430) );
  AOI22_X1 U20542 ( .A1(n3171), .A2(\xmem_data[8][3] ), .B1(n25359), .B2(
        \xmem_data[9][3] ), .ZN(n16416) );
  AOI22_X1 U20543 ( .A1(n27498), .A2(\xmem_data[10][3] ), .B1(n25388), .B2(
        \xmem_data[11][3] ), .ZN(n16415) );
  AOI22_X1 U20544 ( .A1(n25358), .A2(\xmem_data[12][3] ), .B1(n25357), .B2(
        \xmem_data[13][3] ), .ZN(n16414) );
  AOI22_X1 U20545 ( .A1(n3386), .A2(\xmem_data[14][3] ), .B1(n25360), .B2(
        \xmem_data[15][3] ), .ZN(n16413) );
  NAND4_X1 U20546 ( .A1(n16416), .A2(n16415), .A3(n16414), .A4(n16413), .ZN(
        n16428) );
  AOI22_X1 U20547 ( .A1(n30309), .A2(\xmem_data[2][3] ), .B1(n25367), .B2(
        \xmem_data[3][3] ), .ZN(n16426) );
  AOI22_X1 U20548 ( .A1(n30663), .A2(\xmem_data[26][3] ), .B1(n24132), .B2(
        \xmem_data[27][3] ), .ZN(n16425) );
  AOI22_X1 U20549 ( .A1(n27919), .A2(\xmem_data[0][3] ), .B1(n21006), .B2(
        \xmem_data[1][3] ), .ZN(n16417) );
  INV_X1 U20550 ( .A(n16417), .ZN(n16423) );
  AOI22_X1 U20551 ( .A1(n31315), .A2(\xmem_data[6][3] ), .B1(n28098), .B2(
        \xmem_data[7][3] ), .ZN(n16419) );
  AOI22_X1 U20552 ( .A1(n27755), .A2(\xmem_data[30][3] ), .B1(n25383), .B2(
        \xmem_data[31][3] ), .ZN(n16418) );
  NAND2_X1 U20553 ( .A1(n16419), .A2(n16418), .ZN(n16422) );
  AOI22_X1 U20554 ( .A1(n28374), .A2(\xmem_data[24][3] ), .B1(n3358), .B2(
        \xmem_data[25][3] ), .ZN(n16420) );
  INV_X1 U20555 ( .A(n16420), .ZN(n16421) );
  NOR3_X1 U20556 ( .A1(n16423), .A2(n16422), .A3(n16421), .ZN(n16424) );
  NAND3_X1 U20557 ( .A1(n16426), .A2(n16425), .A3(n16424), .ZN(n16427) );
  NOR2_X1 U20558 ( .A1(n16428), .A2(n16427), .ZN(n16429) );
  NAND3_X1 U20559 ( .A1(n16431), .A2(n16430), .A3(n16429), .ZN(n16440) );
  AOI22_X1 U20560 ( .A1(n25354), .A2(\xmem_data[16][3] ), .B1(n3222), .B2(
        \xmem_data[17][3] ), .ZN(n16438) );
  AOI22_X1 U20561 ( .A1(n29289), .A2(\xmem_data[20][3] ), .B1(n27550), .B2(
        \xmem_data[21][3] ), .ZN(n16432) );
  INV_X1 U20562 ( .A(n16432), .ZN(n16436) );
  AOI22_X1 U20563 ( .A1(n30292), .A2(\xmem_data[18][3] ), .B1(n22667), .B2(
        \xmem_data[19][3] ), .ZN(n16434) );
  NAND2_X1 U20564 ( .A1(n25377), .A2(\xmem_data[22][3] ), .ZN(n16433) );
  NAND2_X1 U20565 ( .A1(n16434), .A2(n16433), .ZN(n16435) );
  NOR2_X1 U20566 ( .A1(n16436), .A2(n16435), .ZN(n16437) );
  NAND2_X1 U20567 ( .A1(n16438), .A2(n16437), .ZN(n16439) );
  NOR2_X1 U20568 ( .A1(n16440), .A2(n16439), .ZN(n16441) );
  NAND2_X1 U20569 ( .A1(n16442), .A2(n16441), .ZN(n16444) );
  NAND2_X1 U20570 ( .A1(n16444), .A2(n16443), .ZN(n16466) );
  AOI22_X1 U20571 ( .A1(n25434), .A2(\xmem_data[32][3] ), .B1(n23796), .B2(
        \xmem_data[33][3] ), .ZN(n16448) );
  AOI22_X1 U20572 ( .A1(n23802), .A2(\xmem_data[34][3] ), .B1(n25435), .B2(
        \xmem_data[35][3] ), .ZN(n16447) );
  AOI22_X1 U20573 ( .A1(n28493), .A2(\xmem_data[36][3] ), .B1(n20551), .B2(
        \xmem_data[37][3] ), .ZN(n16446) );
  AOI22_X1 U20574 ( .A1(n3308), .A2(\xmem_data[38][3] ), .B1(n28098), .B2(
        \xmem_data[39][3] ), .ZN(n16445) );
  NAND4_X1 U20575 ( .A1(n16448), .A2(n16447), .A3(n16446), .A4(n16445), .ZN(
        n16464) );
  AOI22_X1 U20576 ( .A1(n3171), .A2(\xmem_data[40][3] ), .B1(n28468), .B2(
        \xmem_data[41][3] ), .ZN(n16452) );
  AOI22_X1 U20577 ( .A1(n29820), .A2(\xmem_data[42][3] ), .B1(n25440), .B2(
        \xmem_data[43][3] ), .ZN(n16451) );
  AOI22_X1 U20578 ( .A1(n25441), .A2(\xmem_data[44][3] ), .B1(n31346), .B2(
        \xmem_data[45][3] ), .ZN(n16450) );
  AOI22_X1 U20579 ( .A1(n25443), .A2(\xmem_data[46][3] ), .B1(n25442), .B2(
        \xmem_data[47][3] ), .ZN(n16449) );
  NAND4_X1 U20580 ( .A1(n16452), .A2(n16451), .A3(n16450), .A4(n16449), .ZN(
        n16463) );
  AOI22_X1 U20581 ( .A1(n28082), .A2(\xmem_data[48][3] ), .B1(n3221), .B2(
        \xmem_data[49][3] ), .ZN(n16456) );
  AOI22_X1 U20582 ( .A1(n25448), .A2(\xmem_data[50][3] ), .B1(n20598), .B2(
        \xmem_data[51][3] ), .ZN(n16455) );
  AOI22_X1 U20583 ( .A1(n25449), .A2(\xmem_data[52][3] ), .B1(n24564), .B2(
        \xmem_data[53][3] ), .ZN(n16454) );
  AOI22_X1 U20584 ( .A1(n25451), .A2(\xmem_data[54][3] ), .B1(n31252), .B2(
        \xmem_data[55][3] ), .ZN(n16453) );
  NAND4_X1 U20585 ( .A1(n16456), .A2(n16455), .A3(n16454), .A4(n16453), .ZN(
        n16462) );
  AOI22_X1 U20586 ( .A1(n16974), .A2(\xmem_data[56][3] ), .B1(n28415), .B2(
        \xmem_data[57][3] ), .ZN(n16460) );
  AOI22_X1 U20587 ( .A1(n25457), .A2(\xmem_data[58][3] ), .B1(n13168), .B2(
        \xmem_data[59][3] ), .ZN(n16459) );
  AOI22_X1 U20588 ( .A1(n25459), .A2(\xmem_data[60][3] ), .B1(n25458), .B2(
        \xmem_data[61][3] ), .ZN(n16458) );
  AOI22_X1 U20589 ( .A1(n30666), .A2(\xmem_data[62][3] ), .B1(n25460), .B2(
        \xmem_data[63][3] ), .ZN(n16457) );
  NAND4_X1 U20590 ( .A1(n16460), .A2(n16459), .A3(n16458), .A4(n16457), .ZN(
        n16461) );
  OR4_X1 U20591 ( .A1(n16464), .A2(n16463), .A3(n16462), .A4(n16461), .ZN(
        n16465) );
  XNOR2_X1 U20592 ( .A(n32612), .B(\fmem_data[30][5] ), .ZN(n30998) );
  AOI22_X1 U20593 ( .A1(n25358), .A2(\xmem_data[12][4] ), .B1(n25357), .B2(
        \xmem_data[13][4] ), .ZN(n16469) );
  AOI22_X1 U20594 ( .A1(n24467), .A2(\xmem_data[8][4] ), .B1(n25359), .B2(
        \xmem_data[9][4] ), .ZN(n16472) );
  NAND2_X1 U20595 ( .A1(n3219), .A2(\xmem_data[17][4] ), .ZN(n16471) );
  NAND2_X1 U20596 ( .A1(n25388), .A2(\xmem_data[11][4] ), .ZN(n16470) );
  AOI22_X1 U20597 ( .A1(n29698), .A2(\xmem_data[18][4] ), .B1(n24695), .B2(
        \xmem_data[19][4] ), .ZN(n16473) );
  NOR2_X1 U20598 ( .A1(n16475), .A2(n16474), .ZN(n16483) );
  NAND2_X1 U20599 ( .A1(n25354), .A2(\xmem_data[16][4] ), .ZN(n16482) );
  AOI22_X1 U20600 ( .A1(n30666), .A2(\xmem_data[30][4] ), .B1(n25383), .B2(
        \xmem_data[31][4] ), .ZN(n16476) );
  INV_X1 U20601 ( .A(n16476), .ZN(n16480) );
  AOI22_X1 U20602 ( .A1(n28374), .A2(\xmem_data[24][4] ), .B1(n22739), .B2(
        \xmem_data[25][4] ), .ZN(n16478) );
  AOI22_X1 U20603 ( .A1(n17041), .A2(\xmem_data[28][4] ), .B1(n25382), .B2(
        \xmem_data[29][4] ), .ZN(n16477) );
  NAND2_X1 U20604 ( .A1(n16478), .A2(n16477), .ZN(n16479) );
  NOR2_X1 U20605 ( .A1(n16480), .A2(n16479), .ZN(n16481) );
  NAND4_X1 U20606 ( .A1(n16469), .A2(n16483), .A3(n16482), .A4(n16481), .ZN(
        n16495) );
  AOI22_X1 U20607 ( .A1(n27919), .A2(\xmem_data[0][4] ), .B1(n24645), .B2(
        \xmem_data[1][4] ), .ZN(n16487) );
  AOI22_X1 U20608 ( .A1(n23722), .A2(\xmem_data[2][4] ), .B1(n25367), .B2(
        \xmem_data[3][4] ), .ZN(n16486) );
  AOI22_X1 U20609 ( .A1(n22683), .A2(\xmem_data[4][4] ), .B1(n25364), .B2(
        \xmem_data[5][4] ), .ZN(n16485) );
  AOI22_X1 U20610 ( .A1(n29246), .A2(\xmem_data[6][4] ), .B1(n28098), .B2(
        \xmem_data[7][4] ), .ZN(n16484) );
  AOI22_X1 U20611 ( .A1(n3229), .A2(\xmem_data[14][4] ), .B1(n25360), .B2(
        \xmem_data[15][4] ), .ZN(n16488) );
  INV_X1 U20612 ( .A(n16488), .ZN(n16489) );
  AOI21_X1 U20613 ( .B1(\xmem_data[10][4] ), .B2(n27717), .A(n16489), .ZN(
        n16493) );
  AOI22_X1 U20614 ( .A1(n27763), .A2(\xmem_data[26][4] ), .B1(n21015), .B2(
        \xmem_data[27][4] ), .ZN(n16492) );
  AOI22_X1 U20615 ( .A1(n28083), .A2(\xmem_data[20][4] ), .B1(n3256), .B2(
        \xmem_data[21][4] ), .ZN(n16491) );
  NAND2_X1 U20616 ( .A1(n25377), .A2(\xmem_data[22][4] ), .ZN(n16490) );
  NAND4_X1 U20617 ( .A1(n3542), .A2(n16493), .A3(n16492), .A4(n3923), .ZN(
        n16494) );
  NOR2_X1 U20618 ( .A1(n16495), .A2(n16494), .ZN(n16497) );
  NAND2_X1 U20619 ( .A1(n23771), .A2(\xmem_data[23][4] ), .ZN(n16496) );
  AOI21_X1 U20620 ( .B1(n16497), .B2(n16496), .A(n25392), .ZN(n16521) );
  AND2_X1 U20621 ( .A1(n3219), .A2(\xmem_data[49][4] ), .ZN(n16498) );
  AOI21_X1 U20622 ( .B1(n24443), .B2(\xmem_data[48][4] ), .A(n16498), .ZN(
        n16502) );
  AOI22_X1 U20623 ( .A1(n25448), .A2(\xmem_data[50][4] ), .B1(n24695), .B2(
        \xmem_data[51][4] ), .ZN(n16501) );
  AOI22_X1 U20624 ( .A1(n25449), .A2(\xmem_data[52][4] ), .B1(n22669), .B2(
        \xmem_data[53][4] ), .ZN(n16500) );
  AOI22_X1 U20625 ( .A1(n25451), .A2(\xmem_data[54][4] ), .B1(n3231), .B2(
        \xmem_data[55][4] ), .ZN(n16499) );
  NAND4_X1 U20626 ( .A1(n16502), .A2(n16501), .A3(n16500), .A4(n16499), .ZN(
        n16518) );
  AOI22_X1 U20627 ( .A1(n3171), .A2(\xmem_data[40][4] ), .B1(n25406), .B2(
        \xmem_data[41][4] ), .ZN(n16506) );
  AOI22_X1 U20628 ( .A1(n28192), .A2(\xmem_data[42][4] ), .B1(n25440), .B2(
        \xmem_data[43][4] ), .ZN(n16505) );
  AOI22_X1 U20629 ( .A1(n25441), .A2(\xmem_data[44][4] ), .B1(n25629), .B2(
        \xmem_data[45][4] ), .ZN(n16504) );
  AOI22_X1 U20630 ( .A1(n25443), .A2(\xmem_data[46][4] ), .B1(n25442), .B2(
        \xmem_data[47][4] ), .ZN(n16503) );
  NAND4_X1 U20631 ( .A1(n16506), .A2(n16505), .A3(n16504), .A4(n16503), .ZN(
        n16517) );
  AOI22_X1 U20632 ( .A1(n24450), .A2(\xmem_data[56][4] ), .B1(n28415), .B2(
        \xmem_data[57][4] ), .ZN(n16510) );
  AOI22_X1 U20633 ( .A1(n25457), .A2(\xmem_data[58][4] ), .B1(n25423), .B2(
        \xmem_data[59][4] ), .ZN(n16509) );
  AOI22_X1 U20634 ( .A1(n25459), .A2(\xmem_data[60][4] ), .B1(n25458), .B2(
        \xmem_data[61][4] ), .ZN(n16508) );
  AOI22_X1 U20635 ( .A1(n28053), .A2(\xmem_data[62][4] ), .B1(n25460), .B2(
        \xmem_data[63][4] ), .ZN(n16507) );
  NAND4_X1 U20636 ( .A1(n16510), .A2(n16509), .A3(n16508), .A4(n16507), .ZN(
        n16516) );
  AOI22_X1 U20637 ( .A1(n25434), .A2(\xmem_data[32][4] ), .B1(n23796), .B2(
        \xmem_data[33][4] ), .ZN(n16514) );
  AOI22_X1 U20638 ( .A1(n29319), .A2(\xmem_data[34][4] ), .B1(n25435), .B2(
        \xmem_data[35][4] ), .ZN(n16513) );
  AOI22_X1 U20639 ( .A1(n3178), .A2(\xmem_data[36][4] ), .B1(n20943), .B2(
        \xmem_data[37][4] ), .ZN(n16512) );
  AOI22_X1 U20640 ( .A1(n3308), .A2(\xmem_data[38][4] ), .B1(n24223), .B2(
        \xmem_data[39][4] ), .ZN(n16511) );
  NAND4_X1 U20641 ( .A1(n16514), .A2(n16513), .A3(n16512), .A4(n16511), .ZN(
        n16515) );
  OR4_X1 U20642 ( .A1(n16518), .A2(n16517), .A3(n16516), .A4(n16515), .ZN(
        n16519) );
  AND2_X1 U20643 ( .A1(n16519), .A2(n25396), .ZN(n16520) );
  NOR2_X1 U20644 ( .A1(n16521), .A2(n16520), .ZN(n16565) );
  AOI22_X1 U20645 ( .A1(n28059), .A2(\xmem_data[96][4] ), .B1(n25398), .B2(
        \xmem_data[97][4] ), .ZN(n16525) );
  AOI22_X1 U20646 ( .A1(n25400), .A2(\xmem_data[98][4] ), .B1(n25399), .B2(
        \xmem_data[99][4] ), .ZN(n16524) );
  AOI22_X1 U20647 ( .A1(n27974), .A2(\xmem_data[100][4] ), .B1(n24222), .B2(
        \xmem_data[101][4] ), .ZN(n16523) );
  AOI22_X1 U20648 ( .A1(n25401), .A2(\xmem_data[102][4] ), .B1(n14975), .B2(
        \xmem_data[103][4] ), .ZN(n16522) );
  NAND4_X1 U20649 ( .A1(n16525), .A2(n16524), .A3(n16523), .A4(n16522), .ZN(
        n16541) );
  AOI22_X1 U20650 ( .A1(n3179), .A2(\xmem_data[104][4] ), .B1(n25406), .B2(
        \xmem_data[105][4] ), .ZN(n16529) );
  AOI22_X1 U20651 ( .A1(n25407), .A2(\xmem_data[106][4] ), .B1(n24686), .B2(
        \xmem_data[107][4] ), .ZN(n16528) );
  AOI22_X1 U20652 ( .A1(n25408), .A2(\xmem_data[108][4] ), .B1(n20489), .B2(
        \xmem_data[109][4] ), .ZN(n16527) );
  AOI22_X1 U20653 ( .A1(n3318), .A2(\xmem_data[110][4] ), .B1(n27501), .B2(
        \xmem_data[111][4] ), .ZN(n16526) );
  NAND4_X1 U20654 ( .A1(n16529), .A2(n16528), .A3(n16527), .A4(n16526), .ZN(
        n16540) );
  AOI22_X1 U20655 ( .A1(n25413), .A2(\xmem_data[112][4] ), .B1(n3221), .B2(
        \xmem_data[113][4] ), .ZN(n16533) );
  AOI22_X1 U20656 ( .A1(n25414), .A2(\xmem_data[114][4] ), .B1(n24695), .B2(
        \xmem_data[115][4] ), .ZN(n16532) );
  AOI22_X1 U20657 ( .A1(n25416), .A2(\xmem_data[116][4] ), .B1(n25415), .B2(
        \xmem_data[117][4] ), .ZN(n16531) );
  AOI22_X1 U20658 ( .A1(n25417), .A2(\xmem_data[118][4] ), .B1(n24657), .B2(
        \xmem_data[119][4] ), .ZN(n16530) );
  NAND4_X1 U20659 ( .A1(n16533), .A2(n16532), .A3(n16531), .A4(n16530), .ZN(
        n16539) );
  AOI22_X1 U20660 ( .A1(n25422), .A2(\xmem_data[120][4] ), .B1(n29307), .B2(
        \xmem_data[121][4] ), .ZN(n16537) );
  AOI22_X1 U20661 ( .A1(n25424), .A2(\xmem_data[122][4] ), .B1(n25423), .B2(
        \xmem_data[123][4] ), .ZN(n16536) );
  AOI22_X1 U20662 ( .A1(n25425), .A2(\xmem_data[124][4] ), .B1(n14898), .B2(
        \xmem_data[125][4] ), .ZN(n16535) );
  AOI22_X1 U20663 ( .A1(n28336), .A2(\xmem_data[126][4] ), .B1(n3207), .B2(
        \xmem_data[127][4] ), .ZN(n16534) );
  NAND4_X1 U20664 ( .A1(n16537), .A2(n16536), .A3(n16535), .A4(n16534), .ZN(
        n16538) );
  OR4_X1 U20665 ( .A1(n16541), .A2(n16540), .A3(n16539), .A4(n16538), .ZN(
        n16563) );
  AOI22_X1 U20666 ( .A1(n25434), .A2(\xmem_data[64][4] ), .B1(n28427), .B2(
        \xmem_data[65][4] ), .ZN(n16545) );
  AOI22_X1 U20667 ( .A1(n27855), .A2(\xmem_data[66][4] ), .B1(n25435), .B2(
        \xmem_data[67][4] ), .ZN(n16544) );
  AOI22_X1 U20668 ( .A1(n27974), .A2(\xmem_data[68][4] ), .B1(n31361), .B2(
        \xmem_data[69][4] ), .ZN(n16543) );
  AOI22_X1 U20669 ( .A1(n3308), .A2(\xmem_data[70][4] ), .B1(n22685), .B2(
        \xmem_data[71][4] ), .ZN(n16542) );
  NAND4_X1 U20670 ( .A1(n16545), .A2(n16544), .A3(n16543), .A4(n16542), .ZN(
        n16561) );
  AOI22_X1 U20671 ( .A1(n3171), .A2(\xmem_data[72][4] ), .B1(n28468), .B2(
        \xmem_data[73][4] ), .ZN(n16549) );
  AOI22_X1 U20672 ( .A1(n29383), .A2(\xmem_data[74][4] ), .B1(n25440), .B2(
        \xmem_data[75][4] ), .ZN(n16548) );
  AOI22_X1 U20673 ( .A1(n25441), .A2(\xmem_data[76][4] ), .B1(n20489), .B2(
        \xmem_data[77][4] ), .ZN(n16547) );
  AOI22_X1 U20674 ( .A1(n25443), .A2(\xmem_data[78][4] ), .B1(n25442), .B2(
        \xmem_data[79][4] ), .ZN(n16546) );
  NAND4_X1 U20675 ( .A1(n16549), .A2(n16548), .A3(n16547), .A4(n16546), .ZN(
        n16560) );
  AOI22_X1 U20676 ( .A1(n23734), .A2(\xmem_data[80][4] ), .B1(n3218), .B2(
        \xmem_data[81][4] ), .ZN(n16553) );
  AOI22_X1 U20677 ( .A1(n25448), .A2(\xmem_data[82][4] ), .B1(n31367), .B2(
        \xmem_data[83][4] ), .ZN(n16552) );
  AOI22_X1 U20678 ( .A1(n25449), .A2(\xmem_data[84][4] ), .B1(n25486), .B2(
        \xmem_data[85][4] ), .ZN(n16551) );
  AOI22_X1 U20679 ( .A1(n25451), .A2(\xmem_data[86][4] ), .B1(n31252), .B2(
        \xmem_data[87][4] ), .ZN(n16550) );
  NAND4_X1 U20680 ( .A1(n16553), .A2(n16552), .A3(n16551), .A4(n16550), .ZN(
        n16559) );
  AOI22_X1 U20681 ( .A1(n30885), .A2(\xmem_data[88][4] ), .B1(n27988), .B2(
        \xmem_data[89][4] ), .ZN(n16557) );
  AOI22_X1 U20682 ( .A1(n25457), .A2(\xmem_data[90][4] ), .B1(n24159), .B2(
        \xmem_data[91][4] ), .ZN(n16556) );
  AOI22_X1 U20683 ( .A1(n25459), .A2(\xmem_data[92][4] ), .B1(n25458), .B2(
        \xmem_data[93][4] ), .ZN(n16555) );
  AOI22_X1 U20684 ( .A1(n29605), .A2(\xmem_data[94][4] ), .B1(n25460), .B2(
        \xmem_data[95][4] ), .ZN(n16554) );
  NAND4_X1 U20685 ( .A1(n16557), .A2(n16556), .A3(n16555), .A4(n16554), .ZN(
        n16558) );
  OR4_X1 U20686 ( .A1(n16561), .A2(n16560), .A3(n16559), .A4(n16558), .ZN(
        n16562) );
  AOI22_X1 U20687 ( .A1(n25473), .A2(n16563), .B1(n25471), .B2(n16562), .ZN(
        n16564) );
  XNOR2_X1 U20688 ( .A(n31655), .B(\fmem_data[30][5] ), .ZN(n30419) );
  OAI22_X1 U20689 ( .A1(n30998), .A2(n33103), .B1(n30419), .B2(n33105), .ZN(
        n26798) );
  OAI21_X1 U20690 ( .B1(n16566), .B2(n3586), .A(n26798), .ZN(n16568) );
  NAND2_X1 U20691 ( .A1(n16568), .A2(n16567), .ZN(n26794) );
  AOI22_X1 U20692 ( .A1(n24697), .A2(\xmem_data[96][7] ), .B1(n27994), .B2(
        \xmem_data[97][7] ), .ZN(n16572) );
  AOI22_X1 U20693 ( .A1(n3129), .A2(\xmem_data[98][7] ), .B1(n27547), .B2(
        \xmem_data[99][7] ), .ZN(n16571) );
  AOI22_X1 U20694 ( .A1(n27551), .A2(\xmem_data[100][7] ), .B1(n24158), .B2(
        \xmem_data[101][7] ), .ZN(n16570) );
  AOI22_X1 U20695 ( .A1(n30943), .A2(\xmem_data[102][7] ), .B1(n28515), .B2(
        \xmem_data[103][7] ), .ZN(n16569) );
  NAND4_X1 U20696 ( .A1(n16572), .A2(n16571), .A3(n16570), .A4(n16569), .ZN(
        n16588) );
  AOI22_X1 U20697 ( .A1(n16986), .A2(\xmem_data[104][7] ), .B1(n25671), .B2(
        \xmem_data[105][7] ), .ZN(n16576) );
  AOI22_X1 U20698 ( .A1(n3465), .A2(\xmem_data[106][7] ), .B1(n13188), .B2(
        \xmem_data[107][7] ), .ZN(n16575) );
  AOI22_X1 U20699 ( .A1(n30949), .A2(\xmem_data[108][7] ), .B1(n17043), .B2(
        \xmem_data[109][7] ), .ZN(n16574) );
  AOI22_X1 U20700 ( .A1(n30950), .A2(\xmem_data[110][7] ), .B1(n30616), .B2(
        \xmem_data[111][7] ), .ZN(n16573) );
  NAND4_X1 U20701 ( .A1(n16576), .A2(n16575), .A3(n16574), .A4(n16573), .ZN(
        n16587) );
  AOI22_X1 U20702 ( .A1(n30956), .A2(\xmem_data[112][7] ), .B1(n30955), .B2(
        \xmem_data[113][7] ), .ZN(n16580) );
  AOI22_X1 U20703 ( .A1(n28461), .A2(\xmem_data[114][7] ), .B1(n27365), .B2(
        \xmem_data[115][7] ), .ZN(n16579) );
  AOI22_X1 U20704 ( .A1(n3171), .A2(\xmem_data[116][7] ), .B1(n28500), .B2(
        \xmem_data[117][7] ), .ZN(n16578) );
  AOI22_X1 U20705 ( .A1(n29383), .A2(\xmem_data[118][7] ), .B1(n25440), .B2(
        \xmem_data[119][7] ), .ZN(n16577) );
  NAND4_X1 U20706 ( .A1(n16580), .A2(n16579), .A3(n16578), .A4(n16577), .ZN(
        n16586) );
  AOI22_X1 U20707 ( .A1(n3380), .A2(\xmem_data[120][7] ), .B1(n20489), .B2(
        \xmem_data[121][7] ), .ZN(n16584) );
  AOI22_X1 U20708 ( .A1(n3333), .A2(\xmem_data[122][7] ), .B1(n3247), .B2(
        \xmem_data[123][7] ), .ZN(n16583) );
  AOI22_X1 U20709 ( .A1(n30962), .A2(\xmem_data[124][7] ), .B1(n3217), .B2(
        \xmem_data[125][7] ), .ZN(n16582) );
  AOI22_X1 U20710 ( .A1(n30964), .A2(\xmem_data[126][7] ), .B1(n30963), .B2(
        \xmem_data[127][7] ), .ZN(n16581) );
  NAND4_X1 U20711 ( .A1(n16584), .A2(n16583), .A3(n16582), .A4(n16581), .ZN(
        n16585) );
  OR4_X1 U20712 ( .A1(n16588), .A2(n16587), .A3(n16586), .A4(n16585), .ZN(
        n16610) );
  AOI22_X1 U20713 ( .A1(n30883), .A2(\xmem_data[64][7] ), .B1(n30882), .B2(
        \xmem_data[65][7] ), .ZN(n16592) );
  AOI22_X1 U20714 ( .A1(n28344), .A2(\xmem_data[66][7] ), .B1(n28007), .B2(
        \xmem_data[67][7] ), .ZN(n16591) );
  AOI22_X1 U20715 ( .A1(n30885), .A2(\xmem_data[68][7] ), .B1(n30884), .B2(
        \xmem_data[69][7] ), .ZN(n16590) );
  AOI22_X1 U20716 ( .A1(n30886), .A2(\xmem_data[70][7] ), .B1(n24132), .B2(
        \xmem_data[71][7] ), .ZN(n16589) );
  NAND4_X1 U20717 ( .A1(n16592), .A2(n16591), .A3(n16590), .A4(n16589), .ZN(
        n16608) );
  AOI22_X1 U20718 ( .A1(n24131), .A2(\xmem_data[72][7] ), .B1(n30513), .B2(
        \xmem_data[73][7] ), .ZN(n16596) );
  AOI22_X1 U20719 ( .A1(n20776), .A2(\xmem_data[74][7] ), .B1(n27989), .B2(
        \xmem_data[75][7] ), .ZN(n16595) );
  AOI22_X1 U20720 ( .A1(n20542), .A2(\xmem_data[76][7] ), .B1(n25677), .B2(
        \xmem_data[77][7] ), .ZN(n16594) );
  AOI22_X1 U20721 ( .A1(n30893), .A2(\xmem_data[78][7] ), .B1(n24592), .B2(
        \xmem_data[79][7] ), .ZN(n16593) );
  NAND4_X1 U20722 ( .A1(n16596), .A2(n16595), .A3(n16594), .A4(n16593), .ZN(
        n16607) );
  AOI22_X1 U20723 ( .A1(n3325), .A2(\xmem_data[80][7] ), .B1(n30898), .B2(
        \xmem_data[81][7] ), .ZN(n16600) );
  AOI22_X1 U20724 ( .A1(n3301), .A2(\xmem_data[82][7] ), .B1(n31314), .B2(
        \xmem_data[83][7] ), .ZN(n16599) );
  AOI22_X1 U20725 ( .A1(n25582), .A2(\xmem_data[84][7] ), .B1(n27526), .B2(
        \xmem_data[85][7] ), .ZN(n16598) );
  AOI22_X1 U20726 ( .A1(n30901), .A2(\xmem_data[86][7] ), .B1(n30900), .B2(
        \xmem_data[87][7] ), .ZN(n16597) );
  NAND4_X1 U20727 ( .A1(n16600), .A2(n16599), .A3(n16598), .A4(n16597), .ZN(
        n16606) );
  AOI22_X1 U20728 ( .A1(n30909), .A2(\xmem_data[88][7] ), .B1(n30908), .B2(
        \xmem_data[89][7] ), .ZN(n16604) );
  AOI22_X1 U20729 ( .A1(n3351), .A2(\xmem_data[90][7] ), .B1(n23731), .B2(
        \xmem_data[91][7] ), .ZN(n16603) );
  AOI22_X1 U20730 ( .A1(n30906), .A2(\xmem_data[92][7] ), .B1(n3217), .B2(
        \xmem_data[93][7] ), .ZN(n16602) );
  AOI22_X1 U20731 ( .A1(n20724), .A2(\xmem_data[94][7] ), .B1(n27507), .B2(
        \xmem_data[95][7] ), .ZN(n16601) );
  NAND4_X1 U20732 ( .A1(n16604), .A2(n16603), .A3(n16602), .A4(n16601), .ZN(
        n16605) );
  OR4_X1 U20733 ( .A1(n16608), .A2(n16607), .A3(n16606), .A4(n16605), .ZN(
        n16609) );
  AOI22_X1 U20734 ( .A1(n30976), .A2(n16610), .B1(n30974), .B2(n16609), .ZN(
        n16661) );
  AOI22_X1 U20735 ( .A1(n30883), .A2(\xmem_data[32][7] ), .B1(n30882), .B2(
        \xmem_data[33][7] ), .ZN(n16614) );
  AOI22_X1 U20736 ( .A1(n27905), .A2(\xmem_data[34][7] ), .B1(n25514), .B2(
        \xmem_data[35][7] ), .ZN(n16613) );
  AOI22_X1 U20737 ( .A1(n30885), .A2(\xmem_data[36][7] ), .B1(n30884), .B2(
        \xmem_data[37][7] ), .ZN(n16612) );
  AOI22_X1 U20738 ( .A1(n30886), .A2(\xmem_data[38][7] ), .B1(n24516), .B2(
        \xmem_data[39][7] ), .ZN(n16611) );
  NAND4_X1 U20739 ( .A1(n16614), .A2(n16613), .A3(n16612), .A4(n16611), .ZN(
        n16630) );
  AOI22_X1 U20740 ( .A1(n27537), .A2(\xmem_data[40][7] ), .B1(n14898), .B2(
        \xmem_data[41][7] ), .ZN(n16618) );
  AOI22_X1 U20741 ( .A1(n28752), .A2(\xmem_data[42][7] ), .B1(n29188), .B2(
        \xmem_data[43][7] ), .ZN(n16617) );
  AOI22_X1 U20742 ( .A1(n25573), .A2(\xmem_data[44][7] ), .B1(n25520), .B2(
        \xmem_data[45][7] ), .ZN(n16616) );
  AOI22_X1 U20743 ( .A1(n30893), .A2(\xmem_data[46][7] ), .B1(n23776), .B2(
        \xmem_data[47][7] ), .ZN(n16615) );
  NAND4_X1 U20744 ( .A1(n16618), .A2(n16617), .A3(n16616), .A4(n16615), .ZN(
        n16629) );
  AOI22_X1 U20745 ( .A1(n25717), .A2(\xmem_data[48][7] ), .B1(n30898), .B2(
        \xmem_data[49][7] ), .ZN(n16622) );
  AOI22_X1 U20746 ( .A1(n3302), .A2(\xmem_data[50][7] ), .B1(n28098), .B2(
        \xmem_data[51][7] ), .ZN(n16621) );
  AOI22_X1 U20747 ( .A1(n3179), .A2(\xmem_data[52][7] ), .B1(n17049), .B2(
        \xmem_data[53][7] ), .ZN(n16620) );
  AOI22_X1 U20748 ( .A1(n30901), .A2(\xmem_data[54][7] ), .B1(n30900), .B2(
        \xmem_data[55][7] ), .ZN(n16619) );
  NAND4_X1 U20749 ( .A1(n16622), .A2(n16621), .A3(n16620), .A4(n16619), .ZN(
        n16628) );
  AOI22_X1 U20750 ( .A1(n30909), .A2(\xmem_data[56][7] ), .B1(n30908), .B2(
        \xmem_data[57][7] ), .ZN(n16626) );
  AOI22_X1 U20751 ( .A1(n3352), .A2(\xmem_data[58][7] ), .B1(n25687), .B2(
        \xmem_data[59][7] ), .ZN(n16625) );
  AOI22_X1 U20752 ( .A1(n30906), .A2(\xmem_data[60][7] ), .B1(n3217), .B2(
        \xmem_data[61][7] ), .ZN(n16624) );
  AOI22_X1 U20753 ( .A1(n23740), .A2(\xmem_data[62][7] ), .B1(n20500), .B2(
        \xmem_data[63][7] ), .ZN(n16623) );
  NAND4_X1 U20754 ( .A1(n16626), .A2(n16625), .A3(n16624), .A4(n16623), .ZN(
        n16627) );
  OR4_X1 U20755 ( .A1(n16630), .A2(n16629), .A3(n16628), .A4(n16627), .ZN(
        n16659) );
  AOI22_X1 U20756 ( .A1(n24640), .A2(\xmem_data[6][7] ), .B1(n24212), .B2(
        \xmem_data[7][7] ), .ZN(n16642) );
  AOI22_X1 U20757 ( .A1(n25449), .A2(\xmem_data[0][7] ), .B1(n25415), .B2(
        \xmem_data[1][7] ), .ZN(n16633) );
  AOI22_X1 U20758 ( .A1(n23813), .A2(\xmem_data[4][7] ), .B1(n30854), .B2(
        \xmem_data[5][7] ), .ZN(n16632) );
  NAND2_X1 U20759 ( .A1(n3129), .A2(\xmem_data[2][7] ), .ZN(n16631) );
  NAND3_X1 U20760 ( .A1(n16633), .A2(n16632), .A3(n16631), .ZN(n16640) );
  AOI22_X1 U20761 ( .A1(n30674), .A2(\xmem_data[22][7] ), .B1(n27435), .B2(
        \xmem_data[23][7] ), .ZN(n16634) );
  INV_X1 U20762 ( .A(n16634), .ZN(n16639) );
  AOI22_X1 U20763 ( .A1(n30849), .A2(\xmem_data[16][7] ), .B1(n25716), .B2(
        \xmem_data[17][7] ), .ZN(n16637) );
  AOI22_X1 U20764 ( .A1(n25582), .A2(\xmem_data[20][7] ), .B1(n21057), .B2(
        \xmem_data[21][7] ), .ZN(n16636) );
  AOI22_X1 U20765 ( .A1(n23724), .A2(\xmem_data[18][7] ), .B1(n14975), .B2(
        \xmem_data[19][7] ), .ZN(n16635) );
  NOR3_X1 U20766 ( .A1(n16640), .A2(n16639), .A3(n16638), .ZN(n16641) );
  NAND2_X1 U20767 ( .A1(n16642), .A2(n16641), .ZN(n16655) );
  AOI22_X1 U20768 ( .A1(n30614), .A2(\xmem_data[8][7] ), .B1(n24160), .B2(
        \xmem_data[9][7] ), .ZN(n16646) );
  AOI22_X1 U20769 ( .A1(n21048), .A2(\xmem_data[10][7] ), .B1(n23716), .B2(
        \xmem_data[11][7] ), .ZN(n16645) );
  AOI22_X1 U20770 ( .A1(n24214), .A2(\xmem_data[12][7] ), .B1(n22718), .B2(
        \xmem_data[13][7] ), .ZN(n16644) );
  AOI22_X1 U20771 ( .A1(n30872), .A2(\xmem_data[14][7] ), .B1(n30871), .B2(
        \xmem_data[15][7] ), .ZN(n16643) );
  AOI22_X1 U20772 ( .A1(n24563), .A2(\xmem_data[30][7] ), .B1(n30963), .B2(
        \xmem_data[31][7] ), .ZN(n16647) );
  INV_X1 U20773 ( .A(n16647), .ZN(n16650) );
  AOI22_X1 U20774 ( .A1(n30864), .A2(\xmem_data[26][7] ), .B1(n30863), .B2(
        \xmem_data[27][7] ), .ZN(n16648) );
  INV_X1 U20775 ( .A(n16648), .ZN(n16649) );
  NOR2_X1 U20776 ( .A1(n16650), .A2(n16649), .ZN(n16653) );
  AOI22_X1 U20777 ( .A1(n30862), .A2(\xmem_data[24][7] ), .B1(n30861), .B2(
        \xmem_data[25][7] ), .ZN(n16652) );
  AOI22_X1 U20778 ( .A1(n28470), .A2(\xmem_data[28][7] ), .B1(n3217), .B2(
        \xmem_data[29][7] ), .ZN(n16651) );
  NAND4_X1 U20779 ( .A1(n3851), .A2(n16653), .A3(n16652), .A4(n16651), .ZN(
        n16654) );
  NOR2_X1 U20780 ( .A1(n16655), .A2(n16654), .ZN(n16657) );
  NAND2_X1 U20781 ( .A1(n25450), .A2(\xmem_data[3][7] ), .ZN(n16656) );
  AOI21_X1 U20782 ( .B1(n16657), .B2(n16656), .A(n30879), .ZN(n16658) );
  AOI21_X1 U20783 ( .B1(n16659), .B2(n30918), .A(n16658), .ZN(n16660) );
  XNOR2_X1 U20784 ( .A(n35355), .B(\fmem_data[10][3] ), .ZN(n33031) );
  XNOR2_X1 U20785 ( .A(n31674), .B(\fmem_data[10][3] ), .ZN(n31948) );
  XOR2_X1 U20786 ( .A(\fmem_data[10][3] ), .B(\fmem_data[10][2] ), .Z(n16662)
         );
  OAI22_X1 U20787 ( .A1(n33031), .A2(n34736), .B1(n31948), .B2(n33690), .ZN(
        n23830) );
  AOI22_X1 U20788 ( .A1(n28492), .A2(\xmem_data[96][7] ), .B1(n21008), .B2(
        \xmem_data[97][7] ), .ZN(n16666) );
  AOI22_X1 U20789 ( .A1(n24460), .A2(\xmem_data[98][7] ), .B1(n28493), .B2(
        \xmem_data[99][7] ), .ZN(n16665) );
  AOI22_X1 U20790 ( .A1(n28494), .A2(\xmem_data[100][7] ), .B1(n31315), .B2(
        \xmem_data[101][7] ), .ZN(n16664) );
  AOI22_X1 U20791 ( .A1(n28495), .A2(\xmem_data[102][7] ), .B1(n30497), .B2(
        \xmem_data[103][7] ), .ZN(n16663) );
  NAND4_X1 U20792 ( .A1(n16666), .A2(n16665), .A3(n16664), .A4(n16663), .ZN(
        n16682) );
  AOI22_X1 U20793 ( .A1(n28500), .A2(\xmem_data[104][7] ), .B1(n28241), .B2(
        \xmem_data[105][7] ), .ZN(n16670) );
  AOI22_X1 U20794 ( .A1(n20707), .A2(\xmem_data[106][7] ), .B1(n29057), .B2(
        \xmem_data[107][7] ), .ZN(n16669) );
  AOI22_X1 U20795 ( .A1(n29118), .A2(\xmem_data[108][7] ), .B1(n28677), .B2(
        \xmem_data[109][7] ), .ZN(n16668) );
  AOI22_X1 U20796 ( .A1(n28501), .A2(\xmem_data[110][7] ), .B1(n28503), .B2(
        \xmem_data[111][7] ), .ZN(n16667) );
  NAND4_X1 U20797 ( .A1(n16670), .A2(n16669), .A3(n16668), .A4(n16667), .ZN(
        n16681) );
  AOI22_X1 U20798 ( .A1(n3221), .A2(\xmem_data[112][7] ), .B1(n29627), .B2(
        \xmem_data[113][7] ), .ZN(n16674) );
  AOI22_X1 U20799 ( .A1(n28508), .A2(\xmem_data[114][7] ), .B1(n24534), .B2(
        \xmem_data[115][7] ), .ZN(n16673) );
  AOI22_X1 U20800 ( .A1(n28509), .A2(\xmem_data[116][7] ), .B1(n3126), .B2(
        \xmem_data[117][7] ), .ZN(n16672) );
  AOI22_X1 U20801 ( .A1(n25450), .A2(\xmem_data[118][7] ), .B1(n28374), .B2(
        \xmem_data[119][7] ), .ZN(n16671) );
  NAND4_X1 U20802 ( .A1(n16674), .A2(n16673), .A3(n16672), .A4(n16671), .ZN(
        n16680) );
  AOI22_X1 U20803 ( .A1(n27943), .A2(\xmem_data[120][7] ), .B1(n25708), .B2(
        \xmem_data[121][7] ), .ZN(n16678) );
  AOI22_X1 U20804 ( .A1(n28515), .A2(\xmem_data[122][7] ), .B1(n25425), .B2(
        \xmem_data[123][7] ), .ZN(n16677) );
  AOI22_X1 U20805 ( .A1(n28517), .A2(\xmem_data[124][7] ), .B1(n3465), .B2(
        \xmem_data[125][7] ), .ZN(n16676) );
  AOI22_X1 U20806 ( .A1(n22742), .A2(\xmem_data[126][7] ), .B1(n28337), .B2(
        \xmem_data[127][7] ), .ZN(n16675) );
  NAND4_X1 U20807 ( .A1(n16678), .A2(n16677), .A3(n16676), .A4(n16675), .ZN(
        n16679) );
  OR4_X1 U20808 ( .A1(n16682), .A2(n16681), .A3(n16680), .A4(n16679), .ZN(
        n16704) );
  AOI22_X1 U20809 ( .A1(n20940), .A2(\xmem_data[64][7] ), .B1(n21050), .B2(
        \xmem_data[65][7] ), .ZN(n16686) );
  AOI22_X1 U20810 ( .A1(n25399), .A2(\xmem_data[66][7] ), .B1(n30899), .B2(
        \xmem_data[67][7] ), .ZN(n16685) );
  AOI22_X1 U20811 ( .A1(n28462), .A2(\xmem_data[68][7] ), .B1(n28461), .B2(
        \xmem_data[69][7] ), .ZN(n16684) );
  AOI22_X1 U20812 ( .A1(n24521), .A2(\xmem_data[70][7] ), .B1(n24685), .B2(
        \xmem_data[71][7] ), .ZN(n16683) );
  NAND4_X1 U20813 ( .A1(n16686), .A2(n16685), .A3(n16684), .A4(n16683), .ZN(
        n16702) );
  AOI22_X1 U20814 ( .A1(n28468), .A2(\xmem_data[72][7] ), .B1(n28467), .B2(
        \xmem_data[73][7] ), .ZN(n16690) );
  AOI22_X1 U20815 ( .A1(n31261), .A2(\xmem_data[74][7] ), .B1(n25441), .B2(
        \xmem_data[75][7] ), .ZN(n16689) );
  AOI22_X1 U20816 ( .A1(n28317), .A2(\xmem_data[76][7] ), .B1(n3318), .B2(
        \xmem_data[77][7] ), .ZN(n16688) );
  AOI22_X1 U20817 ( .A1(n20568), .A2(\xmem_data[78][7] ), .B1(n28470), .B2(
        \xmem_data[79][7] ), .ZN(n16687) );
  NAND4_X1 U20818 ( .A1(n16690), .A2(n16689), .A3(n16688), .A4(n16687), .ZN(
        n16701) );
  AOI22_X1 U20819 ( .A1(n3221), .A2(\xmem_data[80][7] ), .B1(n27831), .B2(
        \xmem_data[81][7] ), .ZN(n16694) );
  AOI22_X1 U20820 ( .A1(n28476), .A2(\xmem_data[82][7] ), .B1(n28475), .B2(
        \xmem_data[83][7] ), .ZN(n16693) );
  AOI22_X1 U20821 ( .A1(n27994), .A2(\xmem_data[84][7] ), .B1(n29231), .B2(
        \xmem_data[85][7] ), .ZN(n16692) );
  AOI22_X1 U20822 ( .A1(n29045), .A2(\xmem_data[86][7] ), .B1(n23813), .B2(
        \xmem_data[87][7] ), .ZN(n16691) );
  NAND4_X1 U20823 ( .A1(n16694), .A2(n16693), .A3(n16692), .A4(n16691), .ZN(
        n16700) );
  AOI22_X1 U20824 ( .A1(n25458), .A2(\xmem_data[92][7] ), .B1(n25672), .B2(
        \xmem_data[93][7] ), .ZN(n16698) );
  AOI22_X1 U20825 ( .A1(n28375), .A2(\xmem_data[90][7] ), .B1(n31268), .B2(
        \xmem_data[91][7] ), .ZN(n16697) );
  AOI22_X1 U20826 ( .A1(n28481), .A2(\xmem_data[88][7] ), .B1(n25424), .B2(
        \xmem_data[89][7] ), .ZN(n16696) );
  AOI22_X1 U20827 ( .A1(n31269), .A2(\xmem_data[94][7] ), .B1(n25573), .B2(
        \xmem_data[95][7] ), .ZN(n16695) );
  NAND4_X1 U20828 ( .A1(n16698), .A2(n16697), .A3(n16696), .A4(n16695), .ZN(
        n16699) );
  OR4_X1 U20829 ( .A1(n16702), .A2(n16701), .A3(n16700), .A4(n16699), .ZN(
        n16703) );
  AOI22_X1 U20830 ( .A1(n28458), .A2(n16704), .B1(n28526), .B2(n16703), .ZN(
        n16752) );
  AOI22_X1 U20831 ( .A1(n25450), .A2(\xmem_data[22][7] ), .B1(n25422), .B2(
        \xmem_data[23][7] ), .ZN(n16727) );
  AOI22_X1 U20832 ( .A1(n28500), .A2(\xmem_data[8][7] ), .B1(n24687), .B2(
        \xmem_data[9][7] ), .ZN(n16709) );
  AOI22_X1 U20833 ( .A1(n27567), .A2(\xmem_data[10][7] ), .B1(n20953), .B2(
        \xmem_data[11][7] ), .ZN(n16708) );
  AOI22_X1 U20834 ( .A1(n20709), .A2(\xmem_data[12][7] ), .B1(n28718), .B2(
        \xmem_data[13][7] ), .ZN(n16707) );
  AND2_X1 U20835 ( .A1(n25485), .A2(\xmem_data[14][7] ), .ZN(n16705) );
  AOI21_X1 U20836 ( .B1(n28470), .B2(\xmem_data[15][7] ), .A(n16705), .ZN(
        n16706) );
  NAND4_X1 U20837 ( .A1(n16709), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16725) );
  AOI22_X1 U20838 ( .A1(n28427), .A2(\xmem_data[0][7] ), .B1(n29319), .B2(
        \xmem_data[1][7] ), .ZN(n16713) );
  AOI22_X1 U20839 ( .A1(n24592), .A2(\xmem_data[2][7] ), .B1(n28428), .B2(
        \xmem_data[3][7] ), .ZN(n16712) );
  AOI22_X1 U20840 ( .A1(n25679), .A2(\xmem_data[4][7] ), .B1(n28461), .B2(
        \xmem_data[5][7] ), .ZN(n16711) );
  AOI22_X1 U20841 ( .A1(n29126), .A2(\xmem_data[6][7] ), .B1(n24606), .B2(
        \xmem_data[7][7] ), .ZN(n16710) );
  NAND4_X1 U20842 ( .A1(n16713), .A2(n16712), .A3(n16711), .A4(n16710), .ZN(
        n16723) );
  AOI22_X1 U20843 ( .A1(n3358), .A2(\xmem_data[24][7] ), .B1(n28671), .B2(
        \xmem_data[25][7] ), .ZN(n16717) );
  AOI22_X1 U20844 ( .A1(n28416), .A2(\xmem_data[26][7] ), .B1(n31268), .B2(
        \xmem_data[27][7] ), .ZN(n16716) );
  AOI22_X1 U20845 ( .A1(n29009), .A2(\xmem_data[28][7] ), .B1(n27755), .B2(
        \xmem_data[29][7] ), .ZN(n16715) );
  AOI22_X1 U20846 ( .A1(n27989), .A2(\xmem_data[30][7] ), .B1(n25635), .B2(
        \xmem_data[31][7] ), .ZN(n16714) );
  NAND4_X1 U20847 ( .A1(n16717), .A2(n16716), .A3(n16715), .A4(n16714), .ZN(
        n16722) );
  AOI22_X1 U20848 ( .A1(n24564), .A2(\xmem_data[20][7] ), .B1(n27905), .B2(
        \xmem_data[21][7] ), .ZN(n16720) );
  AOI22_X1 U20849 ( .A1(n20723), .A2(\xmem_data[18][7] ), .B1(n25416), .B2(
        \xmem_data[19][7] ), .ZN(n16719) );
  AOI22_X1 U20850 ( .A1(n3219), .A2(\xmem_data[16][7] ), .B1(n29431), .B2(
        \xmem_data[17][7] ), .ZN(n16718) );
  NAND3_X1 U20851 ( .A1(n16720), .A2(n16719), .A3(n16718), .ZN(n16721) );
  OR3_X1 U20852 ( .A1(n16723), .A2(n16722), .A3(n16721), .ZN(n16724) );
  NOR2_X1 U20853 ( .A1(n16725), .A2(n16724), .ZN(n16726) );
  AOI21_X1 U20854 ( .B1(n16727), .B2(n16726), .A(n15043), .ZN(n16728) );
  AOI22_X1 U20855 ( .A1(n25520), .A2(\xmem_data[32][7] ), .B1(n30872), .B2(
        \xmem_data[33][7] ), .ZN(n16732) );
  AOI22_X1 U20856 ( .A1(n25399), .A2(\xmem_data[34][7] ), .B1(n24615), .B2(
        \xmem_data[35][7] ), .ZN(n16731) );
  AOI22_X1 U20857 ( .A1(n28462), .A2(\xmem_data[36][7] ), .B1(n28461), .B2(
        \xmem_data[37][7] ), .ZN(n16730) );
  AOI22_X1 U20858 ( .A1(n24570), .A2(\xmem_data[38][7] ), .B1(n27847), .B2(
        \xmem_data[39][7] ), .ZN(n16729) );
  NAND4_X1 U20859 ( .A1(n16732), .A2(n16731), .A3(n16730), .A4(n16729), .ZN(
        n16748) );
  AOI22_X1 U20860 ( .A1(n28468), .A2(\xmem_data[40][7] ), .B1(n28467), .B2(
        \xmem_data[41][7] ), .ZN(n16736) );
  AOI22_X1 U20861 ( .A1(n27435), .A2(\xmem_data[42][7] ), .B1(n20827), .B2(
        \xmem_data[43][7] ), .ZN(n16735) );
  AOI22_X1 U20862 ( .A1(n30861), .A2(\xmem_data[44][7] ), .B1(n3348), .B2(
        \xmem_data[45][7] ), .ZN(n16734) );
  AOI22_X1 U20863 ( .A1(n24439), .A2(\xmem_data[46][7] ), .B1(n28470), .B2(
        \xmem_data[47][7] ), .ZN(n16733) );
  NAND4_X1 U20864 ( .A1(n16736), .A2(n16735), .A3(n16734), .A4(n16733), .ZN(
        n16747) );
  AOI22_X1 U20865 ( .A1(n3217), .A2(\xmem_data[48][7] ), .B1(n28137), .B2(
        \xmem_data[49][7] ), .ZN(n16740) );
  AOI22_X1 U20866 ( .A1(n28476), .A2(\xmem_data[50][7] ), .B1(n28475), .B2(
        \xmem_data[51][7] ), .ZN(n16739) );
  AOI22_X1 U20867 ( .A1(n27903), .A2(\xmem_data[52][7] ), .B1(n29231), .B2(
        \xmem_data[53][7] ), .ZN(n16738) );
  AOI22_X1 U20868 ( .A1(n25514), .A2(\xmem_data[54][7] ), .B1(n23813), .B2(
        \xmem_data[55][7] ), .ZN(n16737) );
  NAND4_X1 U20869 ( .A1(n16740), .A2(n16739), .A3(n16738), .A4(n16737), .ZN(
        n16746) );
  AOI22_X1 U20870 ( .A1(n28481), .A2(\xmem_data[56][7] ), .B1(n23792), .B2(
        \xmem_data[57][7] ), .ZN(n16744) );
  AOI22_X1 U20871 ( .A1(n30552), .A2(\xmem_data[58][7] ), .B1(n29272), .B2(
        \xmem_data[59][7] ), .ZN(n16743) );
  AOI22_X1 U20872 ( .A1(n23793), .A2(\xmem_data[60][7] ), .B1(n29315), .B2(
        \xmem_data[61][7] ), .ZN(n16742) );
  AOI22_X1 U20873 ( .A1(n23716), .A2(\xmem_data[62][7] ), .B1(n25434), .B2(
        \xmem_data[63][7] ), .ZN(n16741) );
  NAND4_X1 U20874 ( .A1(n16744), .A2(n16743), .A3(n16742), .A4(n16741), .ZN(
        n16745) );
  OR4_X1 U20875 ( .A1(n16748), .A2(n16747), .A3(n16746), .A4(n16745), .ZN(
        n16749) );
  XOR2_X1 U20876 ( .A(\fmem_data[29][2] ), .B(\fmem_data[29][3] ), .Z(n16753)
         );
  AOI22_X1 U20877 ( .A1(n27902), .A2(\xmem_data[96][3] ), .B1(n3217), .B2(
        \xmem_data[97][3] ), .ZN(n16757) );
  AOI22_X1 U20878 ( .A1(n28367), .A2(\xmem_data[98][3] ), .B1(n29255), .B2(
        \xmem_data[99][3] ), .ZN(n16756) );
  AOI22_X1 U20879 ( .A1(n27904), .A2(\xmem_data[100][3] ), .B1(n27903), .B2(
        \xmem_data[101][3] ), .ZN(n16755) );
  AOI22_X1 U20880 ( .A1(n27905), .A2(\xmem_data[102][3] ), .B1(n25514), .B2(
        \xmem_data[103][3] ), .ZN(n16754) );
  NAND4_X1 U20881 ( .A1(n16757), .A2(n16756), .A3(n16755), .A4(n16754), .ZN(
        n16773) );
  AOI22_X1 U20882 ( .A1(n27910), .A2(\xmem_data[104][3] ), .B1(n29180), .B2(
        \xmem_data[105][3] ), .ZN(n16761) );
  AOI22_X1 U20883 ( .A1(n27911), .A2(\xmem_data[106][3] ), .B1(n25605), .B2(
        \xmem_data[107][3] ), .ZN(n16760) );
  AOI22_X1 U20884 ( .A1(n3176), .A2(\xmem_data[108][3] ), .B1(n27912), .B2(
        \xmem_data[109][3] ), .ZN(n16759) );
  AOI22_X1 U20885 ( .A1(n20718), .A2(\xmem_data[110][3] ), .B1(n22742), .B2(
        \xmem_data[111][3] ), .ZN(n16758) );
  NAND4_X1 U20886 ( .A1(n16761), .A2(n16760), .A3(n16759), .A4(n16758), .ZN(
        n16772) );
  AOI22_X1 U20887 ( .A1(n27919), .A2(\xmem_data[112][3] ), .B1(n27918), .B2(
        \xmem_data[113][3] ), .ZN(n16765) );
  AOI22_X1 U20888 ( .A1(n29319), .A2(\xmem_data[114][3] ), .B1(n27920), .B2(
        \xmem_data[115][3] ), .ZN(n16764) );
  AOI22_X1 U20889 ( .A1(n22683), .A2(\xmem_data[116][3] ), .B1(n28429), .B2(
        \xmem_data[117][3] ), .ZN(n16763) );
  AOI22_X1 U20890 ( .A1(n3330), .A2(\xmem_data[118][3] ), .B1(n29126), .B2(
        \xmem_data[119][3] ), .ZN(n16762) );
  NAND4_X1 U20891 ( .A1(n16765), .A2(n16764), .A3(n16763), .A4(n16762), .ZN(
        n16771) );
  AOI22_X1 U20892 ( .A1(n20782), .A2(\xmem_data[120][3] ), .B1(n29136), .B2(
        \xmem_data[121][3] ), .ZN(n16769) );
  AOI22_X1 U20893 ( .A1(n31345), .A2(\xmem_data[122][3] ), .B1(n20769), .B2(
        \xmem_data[123][3] ), .ZN(n16768) );
  AOI22_X1 U20894 ( .A1(n27925), .A2(\xmem_data[124][3] ), .B1(n27563), .B2(
        \xmem_data[125][3] ), .ZN(n16767) );
  AOI22_X1 U20895 ( .A1(n24630), .A2(\xmem_data[126][3] ), .B1(n3247), .B2(
        \xmem_data[127][3] ), .ZN(n16766) );
  NAND4_X1 U20896 ( .A1(n16769), .A2(n16768), .A3(n16767), .A4(n16766), .ZN(
        n16770) );
  OR4_X1 U20897 ( .A1(n16773), .A2(n16772), .A3(n16771), .A4(n16770), .ZN(
        n16795) );
  AOI22_X1 U20898 ( .A1(n27902), .A2(\xmem_data[64][3] ), .B1(n3218), .B2(
        \xmem_data[65][3] ), .ZN(n16777) );
  AOI22_X1 U20899 ( .A1(n23770), .A2(\xmem_data[66][3] ), .B1(n25562), .B2(
        \xmem_data[67][3] ), .ZN(n16776) );
  AOI22_X1 U20900 ( .A1(n27904), .A2(\xmem_data[68][3] ), .B1(n27903), .B2(
        \xmem_data[69][3] ), .ZN(n16775) );
  AOI22_X1 U20901 ( .A1(n27905), .A2(\xmem_data[70][3] ), .B1(n30877), .B2(
        \xmem_data[71][3] ), .ZN(n16774) );
  NAND4_X1 U20902 ( .A1(n16777), .A2(n16776), .A3(n16775), .A4(n16774), .ZN(
        n16793) );
  AOI22_X1 U20903 ( .A1(n27910), .A2(\xmem_data[72][3] ), .B1(n29180), .B2(
        \xmem_data[73][3] ), .ZN(n16781) );
  AOI22_X1 U20904 ( .A1(n27911), .A2(\xmem_data[74][3] ), .B1(n29232), .B2(
        \xmem_data[75][3] ), .ZN(n16780) );
  AOI22_X1 U20905 ( .A1(n3176), .A2(\xmem_data[76][3] ), .B1(n27912), .B2(
        \xmem_data[77][3] ), .ZN(n16779) );
  AOI22_X1 U20906 ( .A1(n23795), .A2(\xmem_data[78][3] ), .B1(n3208), .B2(
        \xmem_data[79][3] ), .ZN(n16778) );
  NAND4_X1 U20907 ( .A1(n16781), .A2(n16780), .A3(n16779), .A4(n16778), .ZN(
        n16792) );
  AOI22_X1 U20908 ( .A1(n27919), .A2(\xmem_data[80][3] ), .B1(n27918), .B2(
        \xmem_data[81][3] ), .ZN(n16785) );
  AOI22_X1 U20909 ( .A1(n29012), .A2(\xmem_data[82][3] ), .B1(n27920), .B2(
        \xmem_data[83][3] ), .ZN(n16784) );
  AOI22_X1 U20910 ( .A1(n27952), .A2(\xmem_data[84][3] ), .B1(n20506), .B2(
        \xmem_data[85][3] ), .ZN(n16783) );
  AOI22_X1 U20911 ( .A1(n3308), .A2(\xmem_data[86][3] ), .B1(n24570), .B2(
        \xmem_data[87][3] ), .ZN(n16782) );
  NAND4_X1 U20912 ( .A1(n16785), .A2(n16784), .A3(n16783), .A4(n16782), .ZN(
        n16791) );
  AOI22_X1 U20913 ( .A1(n29325), .A2(\xmem_data[88][3] ), .B1(n29247), .B2(
        \xmem_data[89][3] ), .ZN(n16789) );
  AOI22_X1 U20914 ( .A1(n20985), .A2(\xmem_data[90][3] ), .B1(n20579), .B2(
        \xmem_data[91][3] ), .ZN(n16788) );
  AOI22_X1 U20915 ( .A1(n27925), .A2(\xmem_data[92][3] ), .B1(n25357), .B2(
        \xmem_data[93][3] ), .ZN(n16787) );
  AOI22_X1 U20916 ( .A1(n3333), .A2(\xmem_data[94][3] ), .B1(n25687), .B2(
        \xmem_data[95][3] ), .ZN(n16786) );
  NAND4_X1 U20917 ( .A1(n16789), .A2(n16788), .A3(n16787), .A4(n16786), .ZN(
        n16790) );
  OR4_X1 U20918 ( .A1(n16793), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        n16794) );
  AOI22_X1 U20919 ( .A1(n27937), .A2(n16795), .B1(n27935), .B2(n16794), .ZN(
        n16849) );
  NOR2_X1 U20920 ( .A1(n27877), .A2(n39017), .ZN(n16796) );
  NAND2_X1 U20921 ( .A1(n28007), .A2(n16796), .ZN(n16848) );
  AOI22_X1 U20922 ( .A1(n28337), .A2(\xmem_data[16][3] ), .B1(n24546), .B2(
        \xmem_data[17][3] ), .ZN(n16800) );
  AOI22_X1 U20923 ( .A1(n27855), .A2(\xmem_data[18][3] ), .B1(n25399), .B2(
        \xmem_data[19][3] ), .ZN(n16799) );
  AOI22_X1 U20924 ( .A1(n30849), .A2(\xmem_data[20][3] ), .B1(n20816), .B2(
        \xmem_data[21][3] ), .ZN(n16798) );
  AOI22_X1 U20925 ( .A1(n3301), .A2(\xmem_data[22][3] ), .B1(n28495), .B2(
        \xmem_data[23][3] ), .ZN(n16797) );
  NAND4_X1 U20926 ( .A1(n16800), .A2(n16799), .A3(n16798), .A4(n16797), .ZN(
        n16806) );
  AOI22_X1 U20927 ( .A1(n27847), .A2(\xmem_data[24][3] ), .B1(n28468), .B2(
        \xmem_data[25][3] ), .ZN(n16804) );
  AOI22_X1 U20928 ( .A1(n27852), .A2(\xmem_data[26][3] ), .B1(n20951), .B2(
        \xmem_data[27][3] ), .ZN(n16803) );
  AOI22_X1 U20929 ( .A1(n25408), .A2(\xmem_data[28][3] ), .B1(n29118), .B2(
        \xmem_data[29][3] ), .ZN(n16802) );
  AOI22_X1 U20930 ( .A1(n3414), .A2(\xmem_data[30][3] ), .B1(n29286), .B2(
        \xmem_data[31][3] ), .ZN(n16801) );
  NAND4_X1 U20931 ( .A1(n16804), .A2(n16803), .A3(n16802), .A4(n16801), .ZN(
        n16805) );
  OR2_X1 U20932 ( .A1(n16806), .A2(n16805), .ZN(n16822) );
  AOI22_X1 U20933 ( .A1(n20991), .A2(\xmem_data[0][3] ), .B1(n3218), .B2(
        \xmem_data[1][3] ), .ZN(n16807) );
  INV_X1 U20934 ( .A(n16807), .ZN(n16811) );
  AOI22_X1 U20935 ( .A1(n23812), .A2(\xmem_data[4][3] ), .B1(n30550), .B2(
        \xmem_data[5][3] ), .ZN(n16809) );
  NAND2_X1 U20936 ( .A1(n3137), .A2(\xmem_data[6][3] ), .ZN(n16808) );
  NAND2_X1 U20937 ( .A1(n16809), .A2(n16808), .ZN(n16810) );
  NOR2_X1 U20938 ( .A1(n16811), .A2(n16810), .ZN(n16820) );
  AOI22_X1 U20939 ( .A1(n30551), .A2(\xmem_data[8][3] ), .B1(n27863), .B2(
        \xmem_data[9][3] ), .ZN(n16815) );
  AOI22_X1 U20940 ( .A1(n28671), .A2(\xmem_data[10][3] ), .B1(n24516), .B2(
        \xmem_data[11][3] ), .ZN(n16814) );
  AOI22_X1 U20941 ( .A1(n30514), .A2(\xmem_data[12][3] ), .B1(n29046), .B2(
        \xmem_data[13][3] ), .ZN(n16813) );
  AOI22_X1 U20942 ( .A1(n30666), .A2(\xmem_data[14][3] ), .B1(n27864), .B2(
        \xmem_data[15][3] ), .ZN(n16812) );
  NAND4_X1 U20943 ( .A1(n16815), .A2(n16814), .A3(n16813), .A4(n16812), .ZN(
        n16818) );
  AOI22_X1 U20944 ( .A1(n29627), .A2(\xmem_data[2][3] ), .B1(n27869), .B2(
        \xmem_data[3][3] ), .ZN(n16816) );
  NOR2_X1 U20945 ( .A1(n16818), .A2(n16817), .ZN(n16819) );
  NAND2_X1 U20946 ( .A1(n16820), .A2(n16819), .ZN(n16821) );
  NOR2_X1 U20947 ( .A1(n16822), .A2(n16821), .ZN(n16823) );
  NOR2_X1 U20948 ( .A1(n16823), .A2(n27877), .ZN(n16846) );
  AOI22_X1 U20949 ( .A1(n30962), .A2(\xmem_data[32][3] ), .B1(n3222), .B2(
        \xmem_data[33][3] ), .ZN(n16827) );
  AOI22_X1 U20950 ( .A1(n29494), .A2(\xmem_data[34][3] ), .B1(n28508), .B2(
        \xmem_data[35][3] ), .ZN(n16826) );
  AOI22_X1 U20951 ( .A1(n27938), .A2(\xmem_data[36][3] ), .B1(n25616), .B2(
        \xmem_data[37][3] ), .ZN(n16825) );
  AOI22_X1 U20952 ( .A1(n20962), .A2(\xmem_data[38][3] ), .B1(n28307), .B2(
        \xmem_data[39][3] ), .ZN(n16824) );
  NAND4_X1 U20953 ( .A1(n16827), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        n16843) );
  AOI22_X1 U20954 ( .A1(n25422), .A2(\xmem_data[40][3] ), .B1(n27943), .B2(
        \xmem_data[41][3] ), .ZN(n16831) );
  AOI22_X1 U20955 ( .A1(n27944), .A2(\xmem_data[42][3] ), .B1(n17012), .B2(
        \xmem_data[43][3] ), .ZN(n16830) );
  AOI22_X1 U20956 ( .A1(n31268), .A2(\xmem_data[44][3] ), .B1(n29009), .B2(
        \xmem_data[45][3] ), .ZN(n16829) );
  AOI22_X1 U20957 ( .A1(n27945), .A2(\xmem_data[46][3] ), .B1(n27516), .B2(
        \xmem_data[47][3] ), .ZN(n16828) );
  NAND4_X1 U20958 ( .A1(n16831), .A2(n16830), .A3(n16829), .A4(n16828), .ZN(
        n16842) );
  AOI22_X1 U20959 ( .A1(n29317), .A2(\xmem_data[48][3] ), .B1(n14970), .B2(
        \xmem_data[49][3] ), .ZN(n16835) );
  AOI22_X1 U20960 ( .A1(n23722), .A2(\xmem_data[50][3] ), .B1(n27950), .B2(
        \xmem_data[51][3] ), .ZN(n16834) );
  AOI22_X1 U20961 ( .A1(n27952), .A2(\xmem_data[52][3] ), .B1(n27951), .B2(
        \xmem_data[53][3] ), .ZN(n16833) );
  AOI22_X1 U20962 ( .A1(n3270), .A2(\xmem_data[54][3] ), .B1(n20507), .B2(
        \xmem_data[55][3] ), .ZN(n16832) );
  NAND4_X1 U20963 ( .A1(n16835), .A2(n16834), .A3(n16833), .A4(n16832), .ZN(
        n16841) );
  AOI22_X1 U20964 ( .A1(n24685), .A2(\xmem_data[56][3] ), .B1(n28292), .B2(
        \xmem_data[57][3] ), .ZN(n16839) );
  AOI22_X1 U20965 ( .A1(n31308), .A2(\xmem_data[58][3] ), .B1(n27957), .B2(
        \xmem_data[59][3] ), .ZN(n16838) );
  AOI22_X1 U20966 ( .A1(n27959), .A2(\xmem_data[60][3] ), .B1(n27958), .B2(
        \xmem_data[61][3] ), .ZN(n16837) );
  AOI22_X1 U20967 ( .A1(n22728), .A2(\xmem_data[62][3] ), .B1(n20711), .B2(
        \xmem_data[63][3] ), .ZN(n16836) );
  NAND4_X1 U20968 ( .A1(n16839), .A2(n16838), .A3(n16837), .A4(n16836), .ZN(
        n16840) );
  OR4_X1 U20969 ( .A1(n16843), .A2(n16842), .A3(n16841), .A4(n16840), .ZN(
        n16844) );
  AND2_X1 U20970 ( .A1(n16844), .A2(n27968), .ZN(n16845) );
  NOR2_X1 U20971 ( .A1(n16846), .A2(n16845), .ZN(n16847) );
  AOI22_X1 U20972 ( .A1(n20518), .A2(\xmem_data[32][2] ), .B1(n3221), .B2(
        \xmem_data[33][2] ), .ZN(n16853) );
  AOI22_X1 U20973 ( .A1(n30964), .A2(\xmem_data[34][2] ), .B1(n28319), .B2(
        \xmem_data[35][2] ), .ZN(n16852) );
  AOI22_X1 U20974 ( .A1(n27938), .A2(\xmem_data[36][2] ), .B1(n30550), .B2(
        \xmem_data[37][2] ), .ZN(n16851) );
  AOI22_X1 U20975 ( .A1(n30698), .A2(\xmem_data[38][2] ), .B1(n29103), .B2(
        \xmem_data[39][2] ), .ZN(n16850) );
  NAND4_X1 U20976 ( .A1(n16853), .A2(n16852), .A3(n16851), .A4(n16850), .ZN(
        n16869) );
  AOI22_X1 U20977 ( .A1(n25422), .A2(\xmem_data[40][2] ), .B1(n25456), .B2(
        \xmem_data[41][2] ), .ZN(n16857) );
  AOI22_X1 U20978 ( .A1(n27944), .A2(\xmem_data[42][2] ), .B1(n29232), .B2(
        \xmem_data[43][2] ), .ZN(n16856) );
  AOI22_X1 U20979 ( .A1(n28334), .A2(\xmem_data[44][2] ), .B1(n28517), .B2(
        \xmem_data[45][2] ), .ZN(n16855) );
  AOI22_X1 U20980 ( .A1(n30746), .A2(\xmem_data[46][2] ), .B1(n25383), .B2(
        \xmem_data[47][2] ), .ZN(n16854) );
  NAND4_X1 U20981 ( .A1(n16857), .A2(n16856), .A3(n16855), .A4(n16854), .ZN(
        n16868) );
  AOI22_X1 U20982 ( .A1(n13149), .A2(\xmem_data[48][2] ), .B1(n27518), .B2(
        \xmem_data[49][2] ), .ZN(n16861) );
  AOI22_X1 U20983 ( .A1(n28687), .A2(\xmem_data[50][2] ), .B1(n27950), .B2(
        \xmem_data[51][2] ), .ZN(n16860) );
  AOI22_X1 U20984 ( .A1(n27952), .A2(\xmem_data[52][2] ), .B1(n27951), .B2(
        \xmem_data[53][2] ), .ZN(n16859) );
  AOI22_X1 U20985 ( .A1(n20984), .A2(\xmem_data[54][2] ), .B1(n14975), .B2(
        \xmem_data[55][2] ), .ZN(n16858) );
  NAND4_X1 U20986 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        n16867) );
  AOI22_X1 U20987 ( .A1(n3209), .A2(\xmem_data[56][2] ), .B1(n28500), .B2(
        \xmem_data[57][2] ), .ZN(n16865) );
  AOI22_X1 U20988 ( .A1(n30674), .A2(\xmem_data[58][2] ), .B1(n27957), .B2(
        \xmem_data[59][2] ), .ZN(n16864) );
  AOI22_X1 U20989 ( .A1(n27959), .A2(\xmem_data[60][2] ), .B1(n27958), .B2(
        \xmem_data[61][2] ), .ZN(n16863) );
  AOI22_X1 U20990 ( .A1(n3350), .A2(\xmem_data[62][2] ), .B1(n3247), .B2(
        \xmem_data[63][2] ), .ZN(n16862) );
  NAND4_X1 U20991 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        n16866) );
  OR4_X1 U20992 ( .A1(n16869), .A2(n16868), .A3(n16867), .A4(n16866), .ZN(
        n16899) );
  AOI22_X1 U20993 ( .A1(n20800), .A2(\xmem_data[16][2] ), .B1(n27918), .B2(
        \xmem_data[17][2] ), .ZN(n16873) );
  AOI22_X1 U20994 ( .A1(n27855), .A2(\xmem_data[18][2] ), .B1(n24165), .B2(
        \xmem_data[19][2] ), .ZN(n16872) );
  AOI22_X1 U20995 ( .A1(n28493), .A2(\xmem_data[20][2] ), .B1(n28327), .B2(
        \xmem_data[21][2] ), .ZN(n16871) );
  AOI22_X1 U20996 ( .A1(n25718), .A2(\xmem_data[22][2] ), .B1(n28098), .B2(
        \xmem_data[23][2] ), .ZN(n16870) );
  AOI22_X1 U20997 ( .A1(n27852), .A2(\xmem_data[26][2] ), .B1(n24468), .B2(
        \xmem_data[27][2] ), .ZN(n16880) );
  AOI22_X1 U20998 ( .A1(n27847), .A2(\xmem_data[24][2] ), .B1(n17003), .B2(
        \xmem_data[25][2] ), .ZN(n16874) );
  INV_X1 U20999 ( .A(n16874), .ZN(n16877) );
  AOI22_X1 U21000 ( .A1(n3317), .A2(\xmem_data[30][2] ), .B1(n31347), .B2(
        \xmem_data[31][2] ), .ZN(n16875) );
  INV_X1 U21001 ( .A(n16875), .ZN(n16876) );
  NOR2_X1 U21002 ( .A1(n16877), .A2(n16876), .ZN(n16879) );
  AOI22_X1 U21003 ( .A1(n25630), .A2(\xmem_data[28][2] ), .B1(n3203), .B2(
        \xmem_data[29][2] ), .ZN(n16878) );
  NAND4_X1 U21004 ( .A1(n3852), .A2(n16880), .A3(n16879), .A4(n16878), .ZN(
        n16895) );
  AOI22_X1 U21005 ( .A1(n27447), .A2(\xmem_data[8][2] ), .B1(n27863), .B2(
        \xmem_data[9][2] ), .ZN(n16884) );
  AOI22_X1 U21006 ( .A1(n29451), .A2(\xmem_data[10][2] ), .B1(n28416), .B2(
        \xmem_data[11][2] ), .ZN(n16883) );
  AOI22_X1 U21007 ( .A1(n3176), .A2(\xmem_data[12][2] ), .B1(n24160), .B2(
        \xmem_data[13][2] ), .ZN(n16882) );
  AOI22_X1 U21008 ( .A1(n24545), .A2(\xmem_data[14][2] ), .B1(n27864), .B2(
        \xmem_data[15][2] ), .ZN(n16881) );
  NAND4_X1 U21009 ( .A1(n16884), .A2(n16883), .A3(n16882), .A4(n16881), .ZN(
        n16893) );
  AOI22_X1 U21010 ( .A1(n27902), .A2(\xmem_data[0][2] ), .B1(n3222), .B2(
        \xmem_data[1][2] ), .ZN(n16891) );
  AOI22_X1 U21011 ( .A1(n27938), .A2(\xmem_data[4][2] ), .B1(n13444), .B2(
        \xmem_data[5][2] ), .ZN(n16885) );
  INV_X1 U21012 ( .A(n16885), .ZN(n16889) );
  AOI22_X1 U21013 ( .A1(n29698), .A2(\xmem_data[2][2] ), .B1(n27869), .B2(
        \xmem_data[3][2] ), .ZN(n16887) );
  NAND2_X1 U21014 ( .A1(n3282), .A2(\xmem_data[6][2] ), .ZN(n16886) );
  NAND2_X1 U21015 ( .A1(n16887), .A2(n16886), .ZN(n16888) );
  NOR2_X1 U21016 ( .A1(n16889), .A2(n16888), .ZN(n16890) );
  NAND2_X1 U21017 ( .A1(n16891), .A2(n16890), .ZN(n16892) );
  OR2_X1 U21018 ( .A1(n16893), .A2(n16892), .ZN(n16894) );
  NOR2_X1 U21019 ( .A1(n16895), .A2(n16894), .ZN(n16897) );
  NAND2_X1 U21020 ( .A1(n25450), .A2(\xmem_data[7][2] ), .ZN(n16896) );
  AOI21_X1 U21021 ( .B1(n16897), .B2(n16896), .A(n27877), .ZN(n16898) );
  AOI21_X1 U21022 ( .B1(n16899), .B2(n27968), .A(n16898), .ZN(n16943) );
  AOI22_X1 U21023 ( .A1(n27902), .A2(\xmem_data[96][2] ), .B1(n3218), .B2(
        \xmem_data[97][2] ), .ZN(n16903) );
  AOI22_X1 U21024 ( .A1(n23740), .A2(\xmem_data[98][2] ), .B1(n27444), .B2(
        \xmem_data[99][2] ), .ZN(n16902) );
  AOI22_X1 U21025 ( .A1(n27904), .A2(\xmem_data[100][2] ), .B1(n27903), .B2(
        \xmem_data[101][2] ), .ZN(n16901) );
  AOI22_X1 U21026 ( .A1(n27905), .A2(\xmem_data[102][2] ), .B1(n28510), .B2(
        \xmem_data[103][2] ), .ZN(n16900) );
  NAND4_X1 U21027 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16919) );
  AOI22_X1 U21028 ( .A1(n27910), .A2(\xmem_data[104][2] ), .B1(n30854), .B2(
        \xmem_data[105][2] ), .ZN(n16907) );
  AOI22_X1 U21029 ( .A1(n27911), .A2(\xmem_data[106][2] ), .B1(n23761), .B2(
        \xmem_data[107][2] ), .ZN(n16906) );
  AOI22_X1 U21030 ( .A1(n3176), .A2(\xmem_data[108][2] ), .B1(n27912), .B2(
        \xmem_data[109][2] ), .ZN(n16905) );
  AOI22_X1 U21031 ( .A1(n28154), .A2(\xmem_data[110][2] ), .B1(n29188), .B2(
        \xmem_data[111][2] ), .ZN(n16904) );
  NAND4_X1 U21032 ( .A1(n16907), .A2(n16906), .A3(n16905), .A4(n16904), .ZN(
        n16918) );
  AOI22_X1 U21033 ( .A1(n27919), .A2(\xmem_data[112][2] ), .B1(n27918), .B2(
        \xmem_data[113][2] ), .ZN(n16911) );
  AOI22_X1 U21034 ( .A1(n23777), .A2(\xmem_data[114][2] ), .B1(n27920), .B2(
        \xmem_data[115][2] ), .ZN(n16910) );
  AOI22_X1 U21035 ( .A1(n27974), .A2(\xmem_data[116][2] ), .B1(n20816), .B2(
        \xmem_data[117][2] ), .ZN(n16909) );
  AOI22_X1 U21036 ( .A1(n29324), .A2(\xmem_data[118][2] ), .B1(n28983), .B2(
        \xmem_data[119][2] ), .ZN(n16908) );
  NAND4_X1 U21037 ( .A1(n16911), .A2(n16910), .A3(n16909), .A4(n16908), .ZN(
        n16917) );
  AOI22_X1 U21038 ( .A1(n24685), .A2(\xmem_data[120][2] ), .B1(n28468), .B2(
        \xmem_data[121][2] ), .ZN(n16915) );
  AOI22_X1 U21039 ( .A1(n28772), .A2(\xmem_data[122][2] ), .B1(n25440), .B2(
        \xmem_data[123][2] ), .ZN(n16914) );
  AOI22_X1 U21040 ( .A1(n27925), .A2(\xmem_data[124][2] ), .B1(n28075), .B2(
        \xmem_data[125][2] ), .ZN(n16913) );
  AOI22_X1 U21041 ( .A1(n20828), .A2(\xmem_data[126][2] ), .B1(n22753), .B2(
        \xmem_data[127][2] ), .ZN(n16912) );
  NAND4_X1 U21042 ( .A1(n16915), .A2(n16914), .A3(n16913), .A4(n16912), .ZN(
        n16916) );
  OR4_X1 U21043 ( .A1(n16919), .A2(n16918), .A3(n16917), .A4(n16916), .ZN(
        n16941) );
  AOI22_X1 U21044 ( .A1(n27902), .A2(\xmem_data[64][2] ), .B1(n3221), .B2(
        \xmem_data[65][2] ), .ZN(n16923) );
  AOI22_X1 U21045 ( .A1(n24696), .A2(\xmem_data[66][2] ), .B1(n13469), .B2(
        \xmem_data[67][2] ), .ZN(n16922) );
  AOI22_X1 U21046 ( .A1(n27904), .A2(\xmem_data[68][2] ), .B1(n27903), .B2(
        \xmem_data[69][2] ), .ZN(n16921) );
  AOI22_X1 U21047 ( .A1(n27905), .A2(\xmem_data[70][2] ), .B1(n25514), .B2(
        \xmem_data[71][2] ), .ZN(n16920) );
  NAND4_X1 U21048 ( .A1(n16923), .A2(n16922), .A3(n16921), .A4(n16920), .ZN(
        n16939) );
  AOI22_X1 U21049 ( .A1(n27910), .A2(\xmem_data[72][2] ), .B1(n24130), .B2(
        \xmem_data[73][2] ), .ZN(n16927) );
  AOI22_X1 U21050 ( .A1(n27911), .A2(\xmem_data[74][2] ), .B1(n28416), .B2(
        \xmem_data[75][2] ), .ZN(n16926) );
  AOI22_X1 U21051 ( .A1(n3176), .A2(\xmem_data[76][2] ), .B1(n27912), .B2(
        \xmem_data[77][2] ), .ZN(n16925) );
  AOI22_X1 U21052 ( .A1(n3466), .A2(\xmem_data[78][2] ), .B1(n3213), .B2(
        \xmem_data[79][2] ), .ZN(n16924) );
  NAND4_X1 U21053 ( .A1(n16927), .A2(n16926), .A3(n16925), .A4(n16924), .ZN(
        n16938) );
  AOI22_X1 U21054 ( .A1(n27919), .A2(\xmem_data[80][2] ), .B1(n27918), .B2(
        \xmem_data[81][2] ), .ZN(n16931) );
  AOI22_X1 U21055 ( .A1(n20942), .A2(\xmem_data[82][2] ), .B1(n27920), .B2(
        \xmem_data[83][2] ), .ZN(n16930) );
  AOI22_X1 U21056 ( .A1(n21010), .A2(\xmem_data[84][2] ), .B1(n25679), .B2(
        \xmem_data[85][2] ), .ZN(n16929) );
  AOI22_X1 U21057 ( .A1(n29297), .A2(\xmem_data[86][2] ), .B1(n28062), .B2(
        \xmem_data[87][2] ), .ZN(n16928) );
  NAND4_X1 U21058 ( .A1(n16931), .A2(n16930), .A3(n16929), .A4(n16928), .ZN(
        n16937) );
  AOI22_X1 U21059 ( .A1(n20782), .A2(\xmem_data[88][2] ), .B1(n11008), .B2(
        \xmem_data[89][2] ), .ZN(n16935) );
  AOI22_X1 U21060 ( .A1(n29327), .A2(\xmem_data[90][2] ), .B1(n20769), .B2(
        \xmem_data[91][2] ), .ZN(n16934) );
  AOI22_X1 U21061 ( .A1(n27925), .A2(\xmem_data[92][2] ), .B1(n25357), .B2(
        \xmem_data[93][2] ), .ZN(n16933) );
  AOI22_X1 U21062 ( .A1(n3305), .A2(\xmem_data[94][2] ), .B1(n29253), .B2(
        \xmem_data[95][2] ), .ZN(n16932) );
  NAND4_X1 U21063 ( .A1(n16935), .A2(n16934), .A3(n16933), .A4(n16932), .ZN(
        n16936) );
  OR4_X1 U21064 ( .A1(n16939), .A2(n16938), .A3(n16937), .A4(n16936), .ZN(
        n16940) );
  AOI22_X1 U21065 ( .A1(n27937), .A2(n16941), .B1(n27935), .B2(n16940), .ZN(
        n16942) );
  XOR2_X1 U21066 ( .A(\fmem_data[14][6] ), .B(\fmem_data[14][7] ), .Z(n16944)
         );
  OAI22_X1 U21067 ( .A1(n33228), .A2(n35577), .B1(n31952), .B2(n35576), .ZN(
        n23828) );
  NOR2_X1 U21068 ( .A1(n26794), .A2(n26795), .ZN(n17748) );
  XNOR2_X1 U21069 ( .A(n31895), .B(\fmem_data[4][3] ), .ZN(n33177) );
  XNOR2_X1 U21070 ( .A(n32584), .B(\fmem_data[4][3] ), .ZN(n28265) );
  XOR2_X1 U21071 ( .A(\fmem_data[4][3] ), .B(\fmem_data[4][2] ), .Z(n16945) );
  OAI22_X1 U21072 ( .A1(n33177), .A2(n33174), .B1(n28265), .B2(n33176), .ZN(
        n23585) );
  AOI22_X1 U21073 ( .A1(n16986), .A2(\xmem_data[64][0] ), .B1(n24160), .B2(
        \xmem_data[65][0] ), .ZN(n16949) );
  AOI22_X1 U21074 ( .A1(n16988), .A2(\xmem_data[66][0] ), .B1(n16987), .B2(
        \xmem_data[67][0] ), .ZN(n16948) );
  AOI22_X1 U21075 ( .A1(n20585), .A2(\xmem_data[68][0] ), .B1(n16989), .B2(
        \xmem_data[69][0] ), .ZN(n16947) );
  AOI22_X1 U21076 ( .A1(n16990), .A2(\xmem_data[70][0] ), .B1(n31254), .B2(
        \xmem_data[71][0] ), .ZN(n16946) );
  NAND4_X1 U21077 ( .A1(n16949), .A2(n16948), .A3(n16947), .A4(n16946), .ZN(
        n16965) );
  AOI22_X1 U21078 ( .A1(n25575), .A2(\xmem_data[72][0] ), .B1(n21051), .B2(
        \xmem_data[73][0] ), .ZN(n16953) );
  AOI22_X1 U21079 ( .A1(n3271), .A2(\xmem_data[74][0] ), .B1(n3201), .B2(
        \xmem_data[75][0] ), .ZN(n16952) );
  AOI22_X1 U21080 ( .A1(n3179), .A2(\xmem_data[76][0] ), .B1(n28328), .B2(
        \xmem_data[77][0] ), .ZN(n16951) );
  AOI22_X1 U21081 ( .A1(n24687), .A2(\xmem_data[78][0] ), .B1(n29248), .B2(
        \xmem_data[79][0] ), .ZN(n16950) );
  NAND4_X1 U21082 ( .A1(n16953), .A2(n16952), .A3(n16951), .A4(n16950), .ZN(
        n16964) );
  AOI22_X1 U21083 ( .A1(n30906), .A2(\xmem_data[84][0] ), .B1(n3221), .B2(
        \xmem_data[85][0] ), .ZN(n16957) );
  AOI22_X1 U21084 ( .A1(n16980), .A2(\xmem_data[82][0] ), .B1(n16979), .B2(
        \xmem_data[83][0] ), .ZN(n16956) );
  AOI22_X1 U21085 ( .A1(n24688), .A2(\xmem_data[80][0] ), .B1(n27958), .B2(
        \xmem_data[81][0] ), .ZN(n16955) );
  AOI22_X1 U21086 ( .A1(n23770), .A2(\xmem_data[86][0] ), .B1(n24695), .B2(
        \xmem_data[87][0] ), .ZN(n16954) );
  NAND4_X1 U21087 ( .A1(n16957), .A2(n16956), .A3(n16955), .A4(n16954), .ZN(
        n16963) );
  AOI22_X1 U21088 ( .A1(n20807), .A2(\xmem_data[88][0] ), .B1(n25616), .B2(
        \xmem_data[89][0] ), .ZN(n16961) );
  AOI22_X1 U21089 ( .A1(n16973), .A2(\xmem_data[90][0] ), .B1(n16972), .B2(
        \xmem_data[91][0] ), .ZN(n16960) );
  AOI22_X1 U21090 ( .A1(n16974), .A2(\xmem_data[92][0] ), .B1(n29180), .B2(
        \xmem_data[93][0] ), .ZN(n16959) );
  AOI22_X1 U21091 ( .A1(n31353), .A2(\xmem_data[94][0] ), .B1(n28515), .B2(
        \xmem_data[95][0] ), .ZN(n16958) );
  NAND4_X1 U21092 ( .A1(n16961), .A2(n16960), .A3(n16959), .A4(n16958), .ZN(
        n16962) );
  OR4_X1 U21093 ( .A1(n16965), .A2(n16964), .A3(n16963), .A4(n16962), .ZN(
        n16967) );
  NAND2_X1 U21094 ( .A1(n16967), .A2(n16966), .ZN(n17078) );
  AOI22_X1 U21095 ( .A1(n22683), .A2(\xmem_data[104][0] ), .B1(n20506), .B2(
        \xmem_data[105][0] ), .ZN(n16971) );
  AOI22_X1 U21096 ( .A1(n3270), .A2(\xmem_data[106][0] ), .B1(n3199), .B2(
        \xmem_data[107][0] ), .ZN(n16970) );
  AOI22_X1 U21097 ( .A1(n14976), .A2(\xmem_data[108][0] ), .B1(n29136), .B2(
        \xmem_data[109][0] ), .ZN(n16969) );
  AOI22_X1 U21098 ( .A1(n21060), .A2(\xmem_data[110][0] ), .B1(n17050), .B2(
        \xmem_data[111][0] ), .ZN(n16968) );
  AOI22_X1 U21099 ( .A1(n29254), .A2(\xmem_data[116][0] ), .B1(n3221), .B2(
        \xmem_data[117][0] ), .ZN(n16996) );
  AOI22_X1 U21100 ( .A1(n29257), .A2(\xmem_data[120][0] ), .B1(n30882), .B2(
        \xmem_data[121][0] ), .ZN(n16978) );
  AOI22_X1 U21101 ( .A1(n16973), .A2(\xmem_data[122][0] ), .B1(n16972), .B2(
        \xmem_data[123][0] ), .ZN(n16977) );
  AOI22_X1 U21102 ( .A1(n16974), .A2(\xmem_data[124][0] ), .B1(n3357), .B2(
        \xmem_data[125][0] ), .ZN(n16976) );
  AOI22_X1 U21103 ( .A1(n28671), .A2(\xmem_data[126][0] ), .B1(n27535), .B2(
        \xmem_data[127][0] ), .ZN(n16975) );
  NAND4_X1 U21104 ( .A1(n16978), .A2(n16977), .A3(n16976), .A4(n16975), .ZN(
        n16985) );
  AOI22_X1 U21105 ( .A1(n25630), .A2(\xmem_data[112][0] ), .B1(n31262), .B2(
        \xmem_data[113][0] ), .ZN(n16983) );
  AOI22_X1 U21106 ( .A1(n29288), .A2(\xmem_data[118][0] ), .B1(n20787), .B2(
        \xmem_data[119][0] ), .ZN(n16982) );
  AOI22_X1 U21107 ( .A1(n16980), .A2(\xmem_data[114][0] ), .B1(n16979), .B2(
        \xmem_data[115][0] ), .ZN(n16981) );
  NAND3_X1 U21108 ( .A1(n16983), .A2(n16982), .A3(n16981), .ZN(n16984) );
  NOR2_X1 U21109 ( .A1(n16985), .A2(n16984), .ZN(n16995) );
  AOI22_X1 U21110 ( .A1(n16986), .A2(\xmem_data[96][0] ), .B1(n20798), .B2(
        \xmem_data[97][0] ), .ZN(n16994) );
  AOI22_X1 U21111 ( .A1(n16988), .A2(\xmem_data[98][0] ), .B1(n17019), .B2(
        \xmem_data[99][0] ), .ZN(n16993) );
  AOI22_X1 U21112 ( .A1(n29010), .A2(\xmem_data[100][0] ), .B1(n16989), .B2(
        \xmem_data[101][0] ), .ZN(n16992) );
  AOI22_X1 U21113 ( .A1(n16990), .A2(\xmem_data[102][0] ), .B1(n23801), .B2(
        \xmem_data[103][0] ), .ZN(n16991) );
  NAND4_X1 U21114 ( .A1(n3836), .A2(n16996), .A3(n16995), .A4(n3505), .ZN(
        n16998) );
  NAND2_X1 U21115 ( .A1(n16998), .A2(n16997), .ZN(n17077) );
  AOI22_X1 U21116 ( .A1(n30257), .A2(\xmem_data[46][0] ), .B1(n16999), .B2(
        \xmem_data[47][0] ), .ZN(n17000) );
  INV_X1 U21117 ( .A(n17000), .ZN(n17009) );
  AOI22_X1 U21118 ( .A1(n24615), .A2(\xmem_data[40][0] ), .B1(n17001), .B2(
        \xmem_data[41][0] ), .ZN(n17007) );
  AOI22_X1 U21119 ( .A1(n28293), .A2(\xmem_data[44][0] ), .B1(n17003), .B2(
        \xmem_data[45][0] ), .ZN(n17006) );
  AOI22_X1 U21120 ( .A1(n17004), .A2(\xmem_data[42][0] ), .B1(n3200), .B2(
        \xmem_data[43][0] ), .ZN(n17005) );
  NOR2_X1 U21121 ( .A1(n17009), .A2(n17008), .ZN(n17029) );
  AOI22_X1 U21122 ( .A1(n17010), .A2(\xmem_data[56][0] ), .B1(n25616), .B2(
        \xmem_data[57][0] ), .ZN(n17017) );
  AOI22_X1 U21123 ( .A1(n17063), .A2(\xmem_data[58][0] ), .B1(n17011), .B2(
        \xmem_data[59][0] ), .ZN(n17016) );
  AOI22_X1 U21124 ( .A1(n28374), .A2(\xmem_data[60][0] ), .B1(n28481), .B2(
        \xmem_data[61][0] ), .ZN(n17015) );
  AOI22_X1 U21125 ( .A1(n17013), .A2(\xmem_data[62][0] ), .B1(n17012), .B2(
        \xmem_data[63][0] ), .ZN(n17014) );
  NAND4_X1 U21126 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n17014), .ZN(
        n17027) );
  AOI22_X1 U21127 ( .A1(n17019), .A2(\xmem_data[35][0] ), .B1(n31354), .B2(
        \xmem_data[34][0] ), .ZN(n17025) );
  AOI22_X1 U21128 ( .A1(n31268), .A2(\xmem_data[32][0] ), .B1(n27912), .B2(
        \xmem_data[33][0] ), .ZN(n17024) );
  AOI22_X1 U21129 ( .A1(n17020), .A2(\xmem_data[36][0] ), .B1(n27518), .B2(
        \xmem_data[37][0] ), .ZN(n17023) );
  AOI22_X1 U21130 ( .A1(n17021), .A2(\xmem_data[38][0] ), .B1(n29190), .B2(
        \xmem_data[39][0] ), .ZN(n17022) );
  NAND4_X1 U21131 ( .A1(n17025), .A2(n17024), .A3(n17023), .A4(n17022), .ZN(
        n17026) );
  NOR2_X1 U21132 ( .A1(n17027), .A2(n17026), .ZN(n17028) );
  NAND2_X1 U21133 ( .A1(n17029), .A2(n17028), .ZN(n17040) );
  AOI22_X1 U21134 ( .A1(n17030), .A2(\xmem_data[48][0] ), .B1(n27499), .B2(
        \xmem_data[49][0] ), .ZN(n17037) );
  AOI22_X1 U21135 ( .A1(n3388), .A2(\xmem_data[50][0] ), .B1(n17031), .B2(
        \xmem_data[51][0] ), .ZN(n17036) );
  AOI22_X1 U21136 ( .A1(n30592), .A2(\xmem_data[52][0] ), .B1(n3219), .B2(
        \xmem_data[53][0] ), .ZN(n17035) );
  AOI22_X1 U21137 ( .A1(n17033), .A2(\xmem_data[54][0] ), .B1(n30963), .B2(
        \xmem_data[55][0] ), .ZN(n17034) );
  NAND4_X1 U21138 ( .A1(n17037), .A2(n17036), .A3(n17035), .A4(n17034), .ZN(
        n17039) );
  AOI22_X1 U21139 ( .A1(n17041), .A2(\xmem_data[0][0] ), .B1(n29046), .B2(
        \xmem_data[1][0] ), .ZN(n17048) );
  AOI22_X1 U21140 ( .A1(n29008), .A2(\xmem_data[2][0] ), .B1(n17019), .B2(
        \xmem_data[3][0] ), .ZN(n17047) );
  AOI22_X1 U21141 ( .A1(n31330), .A2(\xmem_data[4][0] ), .B1(n17043), .B2(
        \xmem_data[5][0] ), .ZN(n17046) );
  AOI22_X1 U21142 ( .A1(n17044), .A2(\xmem_data[6][0] ), .B1(n28097), .B2(
        \xmem_data[7][0] ), .ZN(n17045) );
  NAND4_X1 U21143 ( .A1(n17048), .A2(n17047), .A3(n17046), .A4(n17045), .ZN(
        n17072) );
  AOI22_X1 U21144 ( .A1(n28061), .A2(\xmem_data[8][0] ), .B1(n3372), .B2(
        \xmem_data[9][0] ), .ZN(n17055) );
  AOI22_X1 U21145 ( .A1(n24522), .A2(\xmem_data[10][0] ), .B1(n3199), .B2(
        \xmem_data[11][0] ), .ZN(n17054) );
  AOI22_X1 U21146 ( .A1(n22719), .A2(\xmem_data[12][0] ), .B1(n17049), .B2(
        \xmem_data[13][0] ), .ZN(n17053) );
  AOI22_X1 U21147 ( .A1(n17051), .A2(\xmem_data[14][0] ), .B1(n17050), .B2(
        \xmem_data[15][0] ), .ZN(n17052) );
  NAND4_X1 U21148 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17071) );
  AOI22_X1 U21149 ( .A1(n17056), .A2(\xmem_data[16][0] ), .B1(n24525), .B2(
        \xmem_data[17][0] ), .ZN(n17060) );
  AOI22_X1 U21150 ( .A1(n3305), .A2(\xmem_data[18][0] ), .B1(n16979), .B2(
        \xmem_data[19][0] ), .ZN(n17059) );
  AOI22_X1 U21151 ( .A1(n29064), .A2(\xmem_data[20][0] ), .B1(n3218), .B2(
        \xmem_data[21][0] ), .ZN(n17058) );
  AOI22_X1 U21152 ( .A1(n24533), .A2(\xmem_data[22][0] ), .B1(n23739), .B2(
        \xmem_data[23][0] ), .ZN(n17057) );
  NAND4_X1 U21153 ( .A1(n17060), .A2(n17059), .A3(n17058), .A4(n17057), .ZN(
        n17070) );
  AOI22_X1 U21154 ( .A1(n17010), .A2(\xmem_data[24][0] ), .B1(n17061), .B2(
        \xmem_data[25][0] ), .ZN(n17068) );
  AOI22_X1 U21155 ( .A1(n17063), .A2(\xmem_data[26][0] ), .B1(n17062), .B2(
        \xmem_data[27][0] ), .ZN(n17067) );
  AOI22_X1 U21156 ( .A1(n25422), .A2(\xmem_data[28][0] ), .B1(n25481), .B2(
        \xmem_data[29][0] ), .ZN(n17066) );
  AOI22_X1 U21157 ( .A1(n17064), .A2(\xmem_data[30][0] ), .B1(n24516), .B2(
        \xmem_data[31][0] ), .ZN(n17065) );
  NAND4_X1 U21158 ( .A1(n17068), .A2(n17067), .A3(n17066), .A4(n17065), .ZN(
        n17069) );
  OR4_X1 U21159 ( .A1(n17072), .A2(n17071), .A3(n17070), .A4(n17069), .ZN(
        n17074) );
  NAND2_X1 U21160 ( .A1(n17074), .A2(n17073), .ZN(n17075) );
  INV_X1 U21161 ( .A(n35722), .ZN(n17079) );
  NAND2_X1 U21162 ( .A1(n20952), .A2(\xmem_data[44][0] ), .ZN(n17081) );
  NAND2_X1 U21163 ( .A1(n20951), .A2(\xmem_data[45][0] ), .ZN(n17080) );
  NAND2_X1 U21164 ( .A1(n17081), .A2(n17080), .ZN(n17089) );
  AOI22_X1 U21165 ( .A1(n20959), .A2(\xmem_data[62][0] ), .B1(n29009), .B2(
        \xmem_data[63][0] ), .ZN(n17083) );
  AOI22_X1 U21166 ( .A1(n20961), .A2(\xmem_data[58][0] ), .B1(n27988), .B2(
        \xmem_data[59][0] ), .ZN(n17082) );
  NAND2_X1 U21167 ( .A1(n17083), .A2(n17082), .ZN(n17087) );
  AOI22_X1 U21168 ( .A1(n20969), .A2(\xmem_data[54][0] ), .B1(n28372), .B2(
        \xmem_data[55][0] ), .ZN(n17085) );
  AOI22_X1 U21169 ( .A1(n17033), .A2(\xmem_data[52][0] ), .B1(n23739), .B2(
        \xmem_data[53][0] ), .ZN(n17084) );
  NAND2_X1 U21170 ( .A1(n17085), .A2(n17084), .ZN(n17086) );
  OR2_X1 U21171 ( .A1(n17087), .A2(n17086), .ZN(n17088) );
  AOI22_X1 U21172 ( .A1(n20939), .A2(\xmem_data[32][0] ), .B1(n20938), .B2(
        \xmem_data[33][0] ), .ZN(n17093) );
  AOI22_X1 U21173 ( .A1(n21007), .A2(\xmem_data[34][0] ), .B1(n20940), .B2(
        \xmem_data[35][0] ), .ZN(n17092) );
  AOI22_X1 U21174 ( .A1(n20942), .A2(\xmem_data[36][0] ), .B1(n20941), .B2(
        \xmem_data[37][0] ), .ZN(n17091) );
  AOI22_X1 U21175 ( .A1(n20593), .A2(\xmem_data[38][0] ), .B1(n20943), .B2(
        \xmem_data[39][0] ), .ZN(n17090) );
  NAND4_X1 U21176 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17101) );
  AOI22_X1 U21177 ( .A1(n29403), .A2(\xmem_data[60][0] ), .B1(n20958), .B2(
        \xmem_data[61][0] ), .ZN(n17099) );
  AOI22_X1 U21178 ( .A1(n20962), .A2(\xmem_data[56][0] ), .B1(n23771), .B2(
        \xmem_data[57][0] ), .ZN(n17098) );
  AOI22_X1 U21179 ( .A1(n29325), .A2(\xmem_data[42][0] ), .B1(n23781), .B2(
        \xmem_data[43][0] ), .ZN(n17097) );
  AOI22_X1 U21180 ( .A1(n21308), .A2(\xmem_data[48][0] ), .B1(n24172), .B2(
        \xmem_data[49][0] ), .ZN(n17095) );
  AOI22_X1 U21181 ( .A1(n20950), .A2(\xmem_data[40][0] ), .B1(n20949), .B2(
        \xmem_data[41][0] ), .ZN(n17094) );
  NAND4_X1 U21182 ( .A1(n17099), .A2(n17098), .A3(n17097), .A4(n17096), .ZN(
        n17100) );
  NOR2_X1 U21183 ( .A1(n17101), .A2(n17100), .ZN(n17104) );
  AOI22_X1 U21184 ( .A1(n28355), .A2(\xmem_data[50][0] ), .B1(n3217), .B2(
        \xmem_data[51][0] ), .ZN(n17103) );
  AOI22_X1 U21185 ( .A1(n20953), .A2(\xmem_data[46][0] ), .B1(n27563), .B2(
        \xmem_data[47][0] ), .ZN(n17102) );
  NAND3_X1 U21186 ( .A1(n17104), .A2(n17103), .A3(n17102), .ZN(n17105) );
  AOI22_X1 U21187 ( .A1(n21005), .A2(\xmem_data[0][0] ), .B1(n22742), .B2(
        \xmem_data[1][0] ), .ZN(n17109) );
  AOI22_X1 U21188 ( .A1(n21007), .A2(\xmem_data[2][0] ), .B1(n21006), .B2(
        \xmem_data[3][0] ), .ZN(n17108) );
  AOI22_X1 U21189 ( .A1(n21008), .A2(\xmem_data[4][0] ), .B1(n24592), .B2(
        \xmem_data[5][0] ), .ZN(n17107) );
  AOI22_X1 U21190 ( .A1(n21010), .A2(\xmem_data[6][0] ), .B1(n25581), .B2(
        \xmem_data[7][0] ), .ZN(n17106) );
  NAND4_X1 U21191 ( .A1(n17109), .A2(n17108), .A3(n17107), .A4(n17106), .ZN(
        n17115) );
  AOI22_X1 U21192 ( .A1(n24638), .A2(\xmem_data[26][0] ), .B1(n20982), .B2(
        \xmem_data[27][0] ), .ZN(n17113) );
  AOI22_X1 U21193 ( .A1(n24157), .A2(\xmem_data[28][0] ), .B1(n21015), .B2(
        \xmem_data[29][0] ), .ZN(n17112) );
  AOI22_X1 U21194 ( .A1(n25425), .A2(\xmem_data[30][0] ), .B1(n27536), .B2(
        \xmem_data[31][0] ), .ZN(n17111) );
  AOI22_X1 U21195 ( .A1(n20808), .A2(\xmem_data[24][0] ), .B1(n28343), .B2(
        \xmem_data[25][0] ), .ZN(n17110) );
  AOI22_X1 U21196 ( .A1(n30907), .A2(\xmem_data[16][0] ), .B1(n14875), .B2(
        \xmem_data[17][0] ), .ZN(n17116) );
  INV_X1 U21197 ( .A(n17116), .ZN(n17117) );
  AOI21_X1 U21198 ( .B1(\xmem_data[12][0] ), .B2(n20985), .A(n17117), .ZN(
        n17123) );
  AOI22_X1 U21199 ( .A1(n20984), .A2(\xmem_data[8][0] ), .B1(n20983), .B2(
        \xmem_data[9][0] ), .ZN(n17119) );
  AOI22_X1 U21200 ( .A1(\xmem_data[13][0] ), .A2(n30601), .B1(n3218), .B2(
        \xmem_data[19][0] ), .ZN(n17118) );
  AND2_X1 U21201 ( .A1(n17119), .A2(n17118), .ZN(n17122) );
  AOI22_X1 U21202 ( .A1(n3209), .A2(\xmem_data[10][0] ), .B1(n28292), .B2(
        \xmem_data[11][0] ), .ZN(n17121) );
  NAND2_X1 U21203 ( .A1(n20991), .A2(\xmem_data[18][0] ), .ZN(n17120) );
  NAND4_X1 U21204 ( .A1(n17123), .A2(n17122), .A3(n17121), .A4(n17120), .ZN(
        n17127) );
  AOI22_X1 U21205 ( .A1(n20994), .A2(\xmem_data[22][0] ), .B1(n20993), .B2(
        \xmem_data[23][0] ), .ZN(n17125) );
  AOI22_X1 U21206 ( .A1(n27831), .A2(\xmem_data[20][0] ), .B1(n20992), .B2(
        \xmem_data[21][0] ), .ZN(n17124) );
  NAND2_X1 U21207 ( .A1(n17125), .A2(n17124), .ZN(n17126) );
  NOR2_X1 U21208 ( .A1(n17127), .A2(n17126), .ZN(n17129) );
  AOI22_X1 U21209 ( .A1(n20986), .A2(\xmem_data[14][0] ), .B1(n25357), .B2(
        \xmem_data[15][0] ), .ZN(n17128) );
  NAND2_X1 U21210 ( .A1(n17129), .A2(n17128), .ZN(n17130) );
  OAI21_X1 U21211 ( .B1(n3987), .B2(n17130), .A(n20980), .ZN(n17178) );
  AOI22_X1 U21212 ( .A1(n30514), .A2(\xmem_data[126][0] ), .B1(n21076), .B2(
        \xmem_data[127][0] ), .ZN(n17132) );
  AOI22_X1 U21213 ( .A1(n20961), .A2(\xmem_data[122][0] ), .B1(n28373), .B2(
        \xmem_data[123][0] ), .ZN(n17131) );
  NAND2_X1 U21214 ( .A1(n17132), .A2(n17131), .ZN(n17138) );
  AOI22_X1 U21215 ( .A1(n21060), .A2(\xmem_data[108][0] ), .B1(n21059), .B2(
        \xmem_data[109][0] ), .ZN(n17133) );
  INV_X1 U21216 ( .A(n17133), .ZN(n17137) );
  AOI22_X1 U21217 ( .A1(n21069), .A2(\xmem_data[118][0] ), .B1(n21068), .B2(
        \xmem_data[119][0] ), .ZN(n17135) );
  AOI22_X1 U21218 ( .A1(n21067), .A2(\xmem_data[116][0] ), .B1(n25491), .B2(
        \xmem_data[117][0] ), .ZN(n17134) );
  NAND2_X1 U21219 ( .A1(n17135), .A2(n17134), .ZN(n17136) );
  AOI22_X1 U21220 ( .A1(n21048), .A2(\xmem_data[96][0] ), .B1(n30615), .B2(
        \xmem_data[97][0] ), .ZN(n17142) );
  AOI22_X1 U21221 ( .A1(n24509), .A2(\xmem_data[98][0] ), .B1(n27918), .B2(
        \xmem_data[99][0] ), .ZN(n17141) );
  AOI22_X1 U21222 ( .A1(n21050), .A2(\xmem_data[100][0] ), .B1(n21049), .B2(
        \xmem_data[101][0] ), .ZN(n17140) );
  AOI22_X1 U21223 ( .A1(n28428), .A2(\xmem_data[102][0] ), .B1(n23778), .B2(
        \xmem_data[103][0] ), .ZN(n17139) );
  NAND4_X1 U21224 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17150) );
  AOI22_X1 U21225 ( .A1(n23792), .A2(\xmem_data[124][0] ), .B1(n21075), .B2(
        \xmem_data[125][0] ), .ZN(n17148) );
  AOI22_X1 U21226 ( .A1(n21074), .A2(\xmem_data[120][0] ), .B1(n25450), .B2(
        \xmem_data[121][0] ), .ZN(n17147) );
  AOI22_X1 U21227 ( .A1(n21058), .A2(\xmem_data[106][0] ), .B1(n21057), .B2(
        \xmem_data[107][0] ), .ZN(n17146) );
  AOI22_X1 U21228 ( .A1(n30590), .A2(\xmem_data[112][0] ), .B1(n3247), .B2(
        \xmem_data[113][0] ), .ZN(n17144) );
  AOI22_X1 U21229 ( .A1(n21056), .A2(\xmem_data[104][0] ), .B1(n20983), .B2(
        \xmem_data[105][0] ), .ZN(n17143) );
  NAND4_X1 U21230 ( .A1(n17148), .A2(n17147), .A3(n17146), .A4(n17145), .ZN(
        n17149) );
  NOR2_X1 U21231 ( .A1(n17150), .A2(n17149), .ZN(n17153) );
  AOI22_X1 U21232 ( .A1(n21066), .A2(\xmem_data[114][0] ), .B1(n3220), .B2(
        \xmem_data[115][0] ), .ZN(n17152) );
  AOI22_X1 U21233 ( .A1(n21061), .A2(\xmem_data[110][0] ), .B1(n22729), .B2(
        \xmem_data[111][0] ), .ZN(n17151) );
  NAND3_X1 U21234 ( .A1(n17153), .A2(n17152), .A3(n17151), .ZN(n17154) );
  AOI22_X1 U21235 ( .A1(n22728), .A2(\xmem_data[80][0] ), .B1(n28501), .B2(
        \xmem_data[81][0] ), .ZN(n17158) );
  AOI22_X1 U21236 ( .A1(n21066), .A2(\xmem_data[82][0] ), .B1(n3222), .B2(
        \xmem_data[83][0] ), .ZN(n17157) );
  AOI22_X1 U21237 ( .A1(n21067), .A2(\xmem_data[84][0] ), .B1(n20992), .B2(
        \xmem_data[85][0] ), .ZN(n17156) );
  AOI22_X1 U21238 ( .A1(n21069), .A2(\xmem_data[86][0] ), .B1(n21068), .B2(
        \xmem_data[87][0] ), .ZN(n17155) );
  NAND4_X1 U21239 ( .A1(n17158), .A2(n17157), .A3(n17156), .A4(n17155), .ZN(
        n17175) );
  AOI22_X1 U21240 ( .A1(n21048), .A2(\xmem_data[64][0] ), .B1(n22677), .B2(
        \xmem_data[65][0] ), .ZN(n17162) );
  AOI22_X1 U21241 ( .A1(n24509), .A2(\xmem_data[66][0] ), .B1(n25677), .B2(
        \xmem_data[67][0] ), .ZN(n17161) );
  AOI22_X1 U21242 ( .A1(n21050), .A2(\xmem_data[68][0] ), .B1(n21049), .B2(
        \xmem_data[69][0] ), .ZN(n17160) );
  AOI22_X1 U21243 ( .A1(n30849), .A2(\xmem_data[70][0] ), .B1(n21051), .B2(
        \xmem_data[71][0] ), .ZN(n17159) );
  NAND4_X1 U21244 ( .A1(n17162), .A2(n17161), .A3(n17160), .A4(n17159), .ZN(
        n17167) );
  AOI22_X1 U21245 ( .A1(n21060), .A2(\xmem_data[76][0] ), .B1(n21059), .B2(
        \xmem_data[77][0] ), .ZN(n17165) );
  AOI22_X1 U21246 ( .A1(n21056), .A2(\xmem_data[72][0] ), .B1(n28098), .B2(
        \xmem_data[73][0] ), .ZN(n17164) );
  AOI22_X1 U21247 ( .A1(n21058), .A2(\xmem_data[74][0] ), .B1(n21057), .B2(
        \xmem_data[75][0] ), .ZN(n17163) );
  NAND3_X1 U21248 ( .A1(n17165), .A2(n17164), .A3(n17163), .ZN(n17166) );
  NOR2_X1 U21249 ( .A1(n17167), .A2(n17166), .ZN(n17173) );
  AOI22_X1 U21250 ( .A1(n21074), .A2(\xmem_data[88][0] ), .B1(n29103), .B2(
        \xmem_data[89][0] ), .ZN(n17171) );
  AOI22_X1 U21251 ( .A1(n28374), .A2(\xmem_data[90][0] ), .B1(n25481), .B2(
        \xmem_data[91][0] ), .ZN(n17170) );
  AOI22_X1 U21252 ( .A1(n28089), .A2(\xmem_data[92][0] ), .B1(n21075), .B2(
        \xmem_data[93][0] ), .ZN(n17169) );
  AOI22_X1 U21253 ( .A1(n28298), .A2(\xmem_data[94][0] ), .B1(n21076), .B2(
        \xmem_data[95][0] ), .ZN(n17168) );
  AOI22_X1 U21254 ( .A1(n21061), .A2(\xmem_data[78][0] ), .B1(n31346), .B2(
        \xmem_data[79][0] ), .ZN(n17172) );
  NAND3_X1 U21255 ( .A1(n17173), .A2(n3787), .A3(n17172), .ZN(n17174) );
  OAI21_X1 U21256 ( .B1(n17175), .B2(n17174), .A(n21086), .ZN(n17176) );
  INV_X1 U21257 ( .A(n35494), .ZN(n17180) );
  AOI22_X1 U21258 ( .A1(n21050), .A2(\xmem_data[24][0] ), .B1(n13452), .B2(
        \xmem_data[25][0] ), .ZN(n17184) );
  AOI22_X1 U21259 ( .A1(n30899), .A2(\xmem_data[26][0] ), .B1(n28462), .B2(
        \xmem_data[27][0] ), .ZN(n17183) );
  AOI22_X1 U21260 ( .A1(n28226), .A2(\xmem_data[28][0] ), .B1(n24622), .B2(
        \xmem_data[29][0] ), .ZN(n17182) );
  AOI22_X1 U21261 ( .A1(n27542), .A2(\xmem_data[30][0] ), .B1(n29017), .B2(
        \xmem_data[31][0] ), .ZN(n17181) );
  NAND4_X1 U21262 ( .A1(n17184), .A2(n17183), .A3(n17182), .A4(n17181), .ZN(
        n17202) );
  AOI22_X1 U21263 ( .A1(n27568), .A2(\xmem_data[0][0] ), .B1(n27567), .B2(
        \xmem_data[1][0] ), .ZN(n17189) );
  AOI22_X1 U21264 ( .A1(n27564), .A2(\xmem_data[2][0] ), .B1(n27563), .B2(
        \xmem_data[3][0] ), .ZN(n17188) );
  AOI22_X1 U21265 ( .A1(n24693), .A2(\xmem_data[4][0] ), .B1(n25360), .B2(
        \xmem_data[5][0] ), .ZN(n17187) );
  AND2_X1 U21266 ( .A1(n3218), .A2(\xmem_data[7][0] ), .ZN(n17185) );
  AOI21_X1 U21267 ( .B1(n20518), .B2(\xmem_data[6][0] ), .A(n17185), .ZN(
        n17186) );
  NAND4_X1 U21268 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17201) );
  AOI22_X1 U21269 ( .A1(n30608), .A2(\xmem_data[16][0] ), .B1(n27535), .B2(
        \xmem_data[17][0] ), .ZN(n17193) );
  AOI22_X1 U21270 ( .A1(n25710), .A2(\xmem_data[18][0] ), .B1(n27536), .B2(
        \xmem_data[19][0] ), .ZN(n17192) );
  AOI22_X1 U21271 ( .A1(n30303), .A2(\xmem_data[20][0] ), .B1(n29188), .B2(
        \xmem_data[21][0] ), .ZN(n17191) );
  AOI22_X1 U21272 ( .A1(n28059), .A2(\xmem_data[22][0] ), .B1(n28058), .B2(
        \xmem_data[23][0] ), .ZN(n17190) );
  NAND4_X1 U21273 ( .A1(n17193), .A2(n17192), .A3(n17191), .A4(n17190), .ZN(
        n17200) );
  AND2_X1 U21274 ( .A1(n28952), .A2(\xmem_data[12][0] ), .ZN(n17196) );
  AND2_X1 U21275 ( .A1(n29288), .A2(\xmem_data[8][0] ), .ZN(n17195) );
  NOR3_X1 U21276 ( .A1(n17196), .A2(n17195), .A3(n17194), .ZN(n17198) );
  AOI22_X1 U21277 ( .A1(n20725), .A2(\xmem_data[10][0] ), .B1(n27550), .B2(
        \xmem_data[11][0] ), .ZN(n17197) );
  NAND4_X1 U21278 ( .A1(n3997), .A2(n3555), .A3(n17198), .A4(n17197), .ZN(
        n17199) );
  NOR4_X1 U21279 ( .A1(n17202), .A2(n17201), .A3(n17200), .A4(n17199), .ZN(
        n17204) );
  NAND2_X1 U21280 ( .A1(n3231), .A2(\xmem_data[13][0] ), .ZN(n17203) );
  AOI21_X1 U21281 ( .B1(n17204), .B2(n17203), .A(n27573), .ZN(n17205) );
  INV_X1 U21282 ( .A(n17205), .ZN(n17274) );
  AOI22_X1 U21283 ( .A1(n27445), .A2(\xmem_data[72][0] ), .B1(n27444), .B2(
        \xmem_data[73][0] ), .ZN(n17209) );
  AOI22_X1 U21284 ( .A1(n23741), .A2(\xmem_data[74][0] ), .B1(n13444), .B2(
        \xmem_data[75][0] ), .ZN(n17208) );
  AOI22_X1 U21285 ( .A1(n29706), .A2(\xmem_data[76][0] ), .B1(n27446), .B2(
        \xmem_data[77][0] ), .ZN(n17207) );
  AOI22_X1 U21286 ( .A1(n27447), .A2(\xmem_data[78][0] ), .B1(n20546), .B2(
        \xmem_data[79][0] ), .ZN(n17206) );
  NAND4_X1 U21287 ( .A1(n17209), .A2(n17208), .A3(n17207), .A4(n17206), .ZN(
        n17220) );
  AOI22_X1 U21288 ( .A1(n27453), .A2(\xmem_data[80][0] ), .B1(n27452), .B2(
        \xmem_data[81][0] ), .ZN(n17213) );
  AOI22_X1 U21289 ( .A1(n23763), .A2(\xmem_data[82][0] ), .B1(n22674), .B2(
        \xmem_data[83][0] ), .ZN(n17212) );
  AOI22_X1 U21290 ( .A1(n28231), .A2(\xmem_data[84][0] ), .B1(n27454), .B2(
        \xmem_data[85][0] ), .ZN(n17211) );
  AOI22_X1 U21291 ( .A1(n20800), .A2(\xmem_data[86][0] ), .B1(n28492), .B2(
        \xmem_data[87][0] ), .ZN(n17210) );
  NAND4_X1 U21292 ( .A1(n17213), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17219) );
  AOI22_X1 U21293 ( .A1(n17021), .A2(\xmem_data[88][0] ), .B1(n27460), .B2(
        \xmem_data[89][0] ), .ZN(n17217) );
  AOI22_X1 U21294 ( .A1(n27462), .A2(\xmem_data[90][0] ), .B1(n27461), .B2(
        \xmem_data[91][0] ), .ZN(n17216) );
  AOI22_X1 U21295 ( .A1(n24623), .A2(\xmem_data[92][0] ), .B1(n23723), .B2(
        \xmem_data[93][0] ), .ZN(n17215) );
  AOI22_X1 U21296 ( .A1(n25582), .A2(\xmem_data[94][0] ), .B1(n27463), .B2(
        \xmem_data[95][0] ), .ZN(n17214) );
  NAND4_X1 U21297 ( .A1(n17217), .A2(n17216), .A3(n17215), .A4(n17214), .ZN(
        n17218) );
  OR3_X1 U21298 ( .A1(n17220), .A2(n17219), .A3(n17218), .ZN(n17226) );
  AOI22_X1 U21299 ( .A1(n25584), .A2(\xmem_data[64][0] ), .B1(n27435), .B2(
        \xmem_data[65][0] ), .ZN(n17224) );
  AOI22_X1 U21300 ( .A1(n27436), .A2(\xmem_data[66][0] ), .B1(n24573), .B2(
        \xmem_data[67][0] ), .ZN(n17223) );
  AOI22_X1 U21301 ( .A1(n3424), .A2(\xmem_data[68][0] ), .B1(n27437), .B2(
        \xmem_data[69][0] ), .ZN(n17222) );
  AOI22_X1 U21302 ( .A1(n27439), .A2(\xmem_data[70][0] ), .B1(n3217), .B2(
        \xmem_data[71][0] ), .ZN(n17221) );
  NAND4_X1 U21303 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17225) );
  OAI21_X1 U21304 ( .B1(n17226), .B2(n17225), .A(n27494), .ZN(n17273) );
  AOI22_X1 U21305 ( .A1(n27498), .A2(\xmem_data[32][0] ), .B1(n20951), .B2(
        \xmem_data[33][0] ), .ZN(n17231) );
  AOI22_X1 U21306 ( .A1(n27500), .A2(\xmem_data[34][0] ), .B1(n27499), .B2(
        \xmem_data[35][0] ), .ZN(n17230) );
  AOI22_X1 U21307 ( .A1(n3424), .A2(\xmem_data[36][0] ), .B1(n27501), .B2(
        \xmem_data[37][0] ), .ZN(n17229) );
  AND2_X1 U21308 ( .A1(n3222), .A2(\xmem_data[39][0] ), .ZN(n17227) );
  AOI21_X1 U21309 ( .B1(n27502), .B2(\xmem_data[38][0] ), .A(n17227), .ZN(
        n17228) );
  NAND4_X1 U21310 ( .A1(n17231), .A2(n17230), .A3(n17229), .A4(n17228), .ZN(
        n17247) );
  AOI22_X1 U21311 ( .A1(n24563), .A2(\xmem_data[40][0] ), .B1(n27507), .B2(
        \xmem_data[41][0] ), .ZN(n17235) );
  AOI22_X1 U21312 ( .A1(n17010), .A2(\xmem_data[42][0] ), .B1(n13444), .B2(
        \xmem_data[43][0] ), .ZN(n17234) );
  AOI22_X1 U21313 ( .A1(n30710), .A2(\xmem_data[44][0] ), .B1(n28007), .B2(
        \xmem_data[45][0] ), .ZN(n17233) );
  AOI22_X1 U21314 ( .A1(n27508), .A2(\xmem_data[46][0] ), .B1(n25456), .B2(
        \xmem_data[47][0] ), .ZN(n17232) );
  NAND4_X1 U21315 ( .A1(n17235), .A2(n17234), .A3(n17233), .A4(n17232), .ZN(
        n17246) );
  AOI22_X1 U21316 ( .A1(n27514), .A2(\xmem_data[48][0] ), .B1(n27513), .B2(
        \xmem_data[49][0] ), .ZN(n17239) );
  AOI22_X1 U21317 ( .A1(n27515), .A2(\xmem_data[50][0] ), .B1(n25572), .B2(
        \xmem_data[51][0] ), .ZN(n17238) );
  AOI22_X1 U21318 ( .A1(n24213), .A2(\xmem_data[52][0] ), .B1(n27516), .B2(
        \xmem_data[53][0] ), .ZN(n17237) );
  AOI22_X1 U21319 ( .A1(n23764), .A2(\xmem_data[54][0] ), .B1(n27518), .B2(
        \xmem_data[55][0] ), .ZN(n17236) );
  NAND4_X1 U21320 ( .A1(n17239), .A2(n17238), .A3(n17237), .A4(n17236), .ZN(
        n17245) );
  AOI22_X1 U21321 ( .A1(n21008), .A2(\xmem_data[56][0] ), .B1(n27523), .B2(
        \xmem_data[57][0] ), .ZN(n17243) );
  AOI22_X1 U21322 ( .A1(n27524), .A2(\xmem_data[58][0] ), .B1(n25364), .B2(
        \xmem_data[59][0] ), .ZN(n17242) );
  AOI22_X1 U21323 ( .A1(n29246), .A2(\xmem_data[60][0] ), .B1(n27525), .B2(
        \xmem_data[61][0] ), .ZN(n17241) );
  AOI22_X1 U21324 ( .A1(n24606), .A2(\xmem_data[62][0] ), .B1(n27526), .B2(
        \xmem_data[63][0] ), .ZN(n17240) );
  NAND4_X1 U21325 ( .A1(n17243), .A2(n17242), .A3(n17241), .A4(n17240), .ZN(
        n17244) );
  OR4_X1 U21326 ( .A1(n17247), .A2(n17246), .A3(n17245), .A4(n17244), .ZN(
        n17248) );
  NAND2_X1 U21327 ( .A1(n17248), .A2(n27577), .ZN(n17272) );
  AOI22_X1 U21328 ( .A1(n20577), .A2(\xmem_data[96][0] ), .B1(n27435), .B2(
        \xmem_data[97][0] ), .ZN(n17253) );
  AOI22_X1 U21329 ( .A1(n27436), .A2(\xmem_data[98][0] ), .B1(n29118), .B2(
        \xmem_data[99][0] ), .ZN(n17252) );
  AOI22_X1 U21330 ( .A1(n29661), .A2(\xmem_data[100][0] ), .B1(n27437), .B2(
        \xmem_data[101][0] ), .ZN(n17251) );
  AND2_X1 U21331 ( .A1(n3217), .A2(\xmem_data[103][0] ), .ZN(n17249) );
  AOI21_X1 U21332 ( .B1(n27439), .B2(\xmem_data[102][0] ), .A(n17249), .ZN(
        n17250) );
  NAND4_X1 U21333 ( .A1(n17253), .A2(n17252), .A3(n17251), .A4(n17250), .ZN(
        n17269) );
  AOI22_X1 U21334 ( .A1(n27445), .A2(\xmem_data[104][0] ), .B1(n27444), .B2(
        \xmem_data[105][0] ), .ZN(n17257) );
  AOI22_X1 U21335 ( .A1(n22709), .A2(\xmem_data[106][0] ), .B1(n30550), .B2(
        \xmem_data[107][0] ), .ZN(n17256) );
  AOI22_X1 U21336 ( .A1(n25417), .A2(\xmem_data[108][0] ), .B1(n27446), .B2(
        \xmem_data[109][0] ), .ZN(n17255) );
  AOI22_X1 U21337 ( .A1(n27447), .A2(\xmem_data[110][0] ), .B1(n20546), .B2(
        \xmem_data[111][0] ), .ZN(n17254) );
  NAND4_X1 U21338 ( .A1(n17257), .A2(n17256), .A3(n17255), .A4(n17254), .ZN(
        n17268) );
  AOI22_X1 U21339 ( .A1(n27453), .A2(\xmem_data[112][0] ), .B1(n27452), .B2(
        \xmem_data[113][0] ), .ZN(n17261) );
  AOI22_X1 U21340 ( .A1(n30614), .A2(\xmem_data[114][0] ), .B1(n30541), .B2(
        \xmem_data[115][0] ), .ZN(n17260) );
  AOI22_X1 U21341 ( .A1(n28053), .A2(\xmem_data[116][0] ), .B1(n27454), .B2(
        \xmem_data[117][0] ), .ZN(n17259) );
  AOI22_X1 U21342 ( .A1(n31330), .A2(\xmem_data[118][0] ), .B1(n20505), .B2(
        \xmem_data[119][0] ), .ZN(n17258) );
  NAND4_X1 U21343 ( .A1(n17261), .A2(n17260), .A3(n17259), .A4(n17258), .ZN(
        n17267) );
  AOI22_X1 U21344 ( .A1(n23777), .A2(\xmem_data[120][0] ), .B1(n27460), .B2(
        \xmem_data[121][0] ), .ZN(n17265) );
  AOI22_X1 U21345 ( .A1(n27462), .A2(\xmem_data[122][0] ), .B1(n27461), .B2(
        \xmem_data[123][0] ), .ZN(n17264) );
  AOI22_X1 U21346 ( .A1(n30600), .A2(\xmem_data[124][0] ), .B1(n29245), .B2(
        \xmem_data[125][0] ), .ZN(n17263) );
  AOI22_X1 U21347 ( .A1(n25582), .A2(\xmem_data[126][0] ), .B1(n27463), .B2(
        \xmem_data[127][0] ), .ZN(n17262) );
  NAND4_X1 U21348 ( .A1(n17265), .A2(n17264), .A3(n17263), .A4(n17262), .ZN(
        n17266) );
  OR4_X1 U21349 ( .A1(n17269), .A2(n17268), .A3(n17267), .A4(n17266), .ZN(
        n17270) );
  NAND2_X1 U21350 ( .A1(n17270), .A2(n27496), .ZN(n17271) );
  AOI22_X1 U21351 ( .A1(n3218), .A2(\xmem_data[32][1] ), .B1(n28733), .B2(
        \xmem_data[33][1] ), .ZN(n17278) );
  AOI22_X1 U21352 ( .A1(n24207), .A2(\xmem_data[34][1] ), .B1(n30883), .B2(
        \xmem_data[35][1] ), .ZN(n17277) );
  AOI22_X1 U21353 ( .A1(n24140), .A2(\xmem_data[36][1] ), .B1(n3134), .B2(
        \xmem_data[37][1] ), .ZN(n17276) );
  AOI22_X1 U21354 ( .A1(n28007), .A2(\xmem_data[38][1] ), .B1(n25604), .B2(
        \xmem_data[39][1] ), .ZN(n17275) );
  NAND4_X1 U21355 ( .A1(n17278), .A2(n17277), .A3(n17276), .A4(n17275), .ZN(
        n17295) );
  AOI22_X1 U21356 ( .A1(n27943), .A2(\xmem_data[40][1] ), .B1(n23762), .B2(
        \xmem_data[41][1] ), .ZN(n17282) );
  AOI22_X1 U21357 ( .A1(n24212), .A2(\xmem_data[42][1] ), .B1(n17041), .B2(
        \xmem_data[43][1] ), .ZN(n17281) );
  AOI22_X1 U21358 ( .A1(n28090), .A2(\xmem_data[44][1] ), .B1(n20718), .B2(
        \xmem_data[45][1] ), .ZN(n17280) );
  AOI22_X1 U21359 ( .A1(n23716), .A2(\xmem_data[46][1] ), .B1(n24214), .B2(
        \xmem_data[47][1] ), .ZN(n17279) );
  NAND4_X1 U21360 ( .A1(n17282), .A2(n17281), .A3(n17280), .A4(n17279), .ZN(
        n17294) );
  AOI22_X1 U21361 ( .A1(n24219), .A2(\xmem_data[48][1] ), .B1(n24710), .B2(
        \xmem_data[49][1] ), .ZN(n17286) );
  AOI22_X1 U21362 ( .A1(n24221), .A2(\xmem_data[50][1] ), .B1(n27524), .B2(
        \xmem_data[51][1] ), .ZN(n17285) );
  AOI22_X1 U21363 ( .A1(n24222), .A2(\xmem_data[52][1] ), .B1(n25401), .B2(
        \xmem_data[53][1] ), .ZN(n17284) );
  AOI22_X1 U21364 ( .A1(n24223), .A2(\xmem_data[54][1] ), .B1(n25582), .B2(
        \xmem_data[55][1] ), .ZN(n17283) );
  NAND4_X1 U21365 ( .A1(n17286), .A2(n17285), .A3(n17284), .A4(n17283), .ZN(
        n17293) );
  AOI22_X1 U21366 ( .A1(n25527), .A2(\xmem_data[56][1] ), .B1(n29298), .B2(
        \xmem_data[57][1] ), .ZN(n17291) );
  AOI22_X1 U21367 ( .A1(n20579), .A2(\xmem_data[58][1] ), .B1(n24526), .B2(
        \xmem_data[59][1] ), .ZN(n17290) );
  AOI22_X1 U21368 ( .A1(n27499), .A2(\xmem_data[60][1] ), .B1(n16980), .B2(
        \xmem_data[61][1] ), .ZN(n17289) );
  AND2_X1 U21369 ( .A1(n25360), .A2(\xmem_data[62][1] ), .ZN(n17287) );
  AOI21_X1 U21370 ( .B1(n20576), .B2(\xmem_data[63][1] ), .A(n17287), .ZN(
        n17288) );
  NAND4_X1 U21371 ( .A1(n17291), .A2(n17290), .A3(n17289), .A4(n17288), .ZN(
        n17292) );
  OR4_X1 U21372 ( .A1(n17295), .A2(n17294), .A3(n17293), .A4(n17292), .ZN(
        n17296) );
  AOI22_X1 U21373 ( .A1(n25458), .A2(\xmem_data[12][1] ), .B1(n31354), .B2(
        \xmem_data[13][1] ), .ZN(n17300) );
  AOI22_X1 U21374 ( .A1(n24132), .A2(\xmem_data[10][1] ), .B1(n24131), .B2(
        \xmem_data[11][1] ), .ZN(n17299) );
  AOI22_X1 U21375 ( .A1(n24130), .A2(\xmem_data[8][1] ), .B1(n22738), .B2(
        \xmem_data[9][1] ), .ZN(n17298) );
  AOI22_X1 U21376 ( .A1(n24134), .A2(\xmem_data[14][1] ), .B1(n24133), .B2(
        \xmem_data[15][1] ), .ZN(n17297) );
  AOI22_X1 U21377 ( .A1(n23781), .A2(\xmem_data[24][1] ), .B1(n29298), .B2(
        \xmem_data[25][1] ), .ZN(n17305) );
  AOI22_X1 U21378 ( .A1(n24122), .A2(\xmem_data[26][1] ), .B1(n29124), .B2(
        \xmem_data[27][1] ), .ZN(n17304) );
  AOI22_X1 U21379 ( .A1(n24525), .A2(\xmem_data[28][1] ), .B1(n3335), .B2(
        \xmem_data[29][1] ), .ZN(n17303) );
  AND2_X1 U21380 ( .A1(n3247), .A2(\xmem_data[30][1] ), .ZN(n17301) );
  AOI21_X1 U21381 ( .B1(n21066), .B2(\xmem_data[31][1] ), .A(n17301), .ZN(
        n17302) );
  NAND4_X1 U21382 ( .A1(n17305), .A2(n17304), .A3(n17303), .A4(n17302), .ZN(
        n17316) );
  AOI22_X1 U21383 ( .A1(n20787), .A2(\xmem_data[2][1] ), .B1(n24141), .B2(
        \xmem_data[3][1] ), .ZN(n17309) );
  AOI22_X1 U21384 ( .A1(n24140), .A2(\xmem_data[4][1] ), .B1(n14991), .B2(
        \xmem_data[5][1] ), .ZN(n17308) );
  AOI22_X1 U21385 ( .A1(n3217), .A2(\xmem_data[0][1] ), .B1(n24139), .B2(
        \xmem_data[1][1] ), .ZN(n17307) );
  NAND2_X1 U21386 ( .A1(n23813), .A2(\xmem_data[7][1] ), .ZN(n17306) );
  AOI22_X1 U21387 ( .A1(n16989), .A2(\xmem_data[16][1] ), .B1(n24115), .B2(
        \xmem_data[17][1] ), .ZN(n17313) );
  AOI22_X1 U21388 ( .A1(n24116), .A2(\xmem_data[18][1] ), .B1(n28460), .B2(
        \xmem_data[19][1] ), .ZN(n17312) );
  AOI22_X1 U21389 ( .A1(n24117), .A2(\xmem_data[20][1] ), .B1(n21056), .B2(
        \xmem_data[21][1] ), .ZN(n17311) );
  AOI22_X1 U21390 ( .A1(n29126), .A2(\xmem_data[22][1] ), .B1(n20734), .B2(
        \xmem_data[23][1] ), .ZN(n17310) );
  NAND4_X1 U21391 ( .A1(n17313), .A2(n17312), .A3(n17311), .A4(n17310), .ZN(
        n17314) );
  OR4_X1 U21392 ( .A1(n17317), .A2(n17316), .A3(n17315), .A4(n17314), .ZN(
        n17318) );
  INV_X1 U21393 ( .A(n17389), .ZN(n24151) );
  NOR2_X1 U21394 ( .A1(n24151), .A2(n39025), .ZN(n17319) );
  NOR2_X1 U21395 ( .A1(n17320), .A2(n3962), .ZN(n17367) );
  AOI22_X1 U21396 ( .A1(n3217), .A2(\xmem_data[96][1] ), .B1(n24696), .B2(
        \xmem_data[97][1] ), .ZN(n17324) );
  AOI22_X1 U21397 ( .A1(n24695), .A2(\xmem_data[98][1] ), .B1(n29257), .B2(
        \xmem_data[99][1] ), .ZN(n17323) );
  AOI22_X1 U21398 ( .A1(n20559), .A2(\xmem_data[100][1] ), .B1(n30710), .B2(
        \xmem_data[101][1] ), .ZN(n17322) );
  AOI22_X1 U21399 ( .A1(n23771), .A2(\xmem_data[102][1] ), .B1(n28374), .B2(
        \xmem_data[103][1] ), .ZN(n17321) );
  NAND4_X1 U21400 ( .A1(n17324), .A2(n17323), .A3(n17322), .A4(n17321), .ZN(
        n17341) );
  AOI22_X1 U21401 ( .A1(n24158), .A2(\xmem_data[104][1] ), .B1(n24157), .B2(
        \xmem_data[105][1] ), .ZN(n17328) );
  AOI22_X1 U21402 ( .A1(n24159), .A2(\xmem_data[106][1] ), .B1(n17041), .B2(
        \xmem_data[107][1] ), .ZN(n17327) );
  AOI22_X1 U21403 ( .A1(n24160), .A2(\xmem_data[108][1] ), .B1(n20718), .B2(
        \xmem_data[109][1] ), .ZN(n17326) );
  AOI22_X1 U21404 ( .A1(n23716), .A2(\xmem_data[110][1] ), .B1(n31330), .B2(
        \xmem_data[111][1] ), .ZN(n17325) );
  NAND4_X1 U21405 ( .A1(n17328), .A2(n17327), .A3(n17326), .A4(n17325), .ZN(
        n17340) );
  AOI22_X1 U21406 ( .A1(n25520), .A2(\xmem_data[112][1] ), .B1(n20815), .B2(
        \xmem_data[113][1] ), .ZN(n17332) );
  AOI22_X1 U21407 ( .A1(n24165), .A2(\xmem_data[114][1] ), .B1(n25575), .B2(
        \xmem_data[115][1] ), .ZN(n17331) );
  AOI22_X1 U21408 ( .A1(n30898), .A2(\xmem_data[116][1] ), .B1(n3330), .B2(
        \xmem_data[117][1] ), .ZN(n17330) );
  AOI22_X1 U21409 ( .A1(n24167), .A2(\xmem_data[118][1] ), .B1(n24166), .B2(
        \xmem_data[119][1] ), .ZN(n17329) );
  NAND4_X1 U21410 ( .A1(n17332), .A2(n17331), .A3(n17330), .A4(n17329), .ZN(
        n17339) );
  AOI22_X1 U21411 ( .A1(n11008), .A2(\xmem_data[120][1] ), .B1(n20985), .B2(
        \xmem_data[121][1] ), .ZN(n17337) );
  AOI22_X1 U21412 ( .A1(n20707), .A2(\xmem_data[122][1] ), .B1(n20710), .B2(
        \xmem_data[123][1] ), .ZN(n17336) );
  AOI22_X1 U21413 ( .A1(n30571), .A2(\xmem_data[124][1] ), .B1(n3317), .B2(
        \xmem_data[125][1] ), .ZN(n17335) );
  AND2_X1 U21414 ( .A1(n24172), .A2(\xmem_data[126][1] ), .ZN(n17333) );
  AOI21_X1 U21415 ( .B1(n25354), .B2(\xmem_data[127][1] ), .A(n17333), .ZN(
        n17334) );
  NAND4_X1 U21416 ( .A1(n17337), .A2(n17336), .A3(n17335), .A4(n17334), .ZN(
        n17338) );
  OR4_X1 U21417 ( .A1(n17341), .A2(n17340), .A3(n17339), .A4(n17338), .ZN(
        n17342) );
  NAND2_X1 U21418 ( .A1(n17342), .A2(n24205), .ZN(n17366) );
  AOI22_X1 U21419 ( .A1(n3219), .A2(\xmem_data[64][1] ), .B1(n23740), .B2(
        \xmem_data[65][1] ), .ZN(n17346) );
  AOI22_X1 U21420 ( .A1(n27507), .A2(\xmem_data[66][1] ), .B1(n29257), .B2(
        \xmem_data[67][1] ), .ZN(n17345) );
  AOI22_X1 U21421 ( .A1(n20806), .A2(\xmem_data[68][1] ), .B1(n23742), .B2(
        \xmem_data[69][1] ), .ZN(n17344) );
  AOI22_X1 U21422 ( .A1(n28045), .A2(\xmem_data[70][1] ), .B1(n28374), .B2(
        \xmem_data[71][1] ), .ZN(n17343) );
  NAND4_X1 U21423 ( .A1(n17346), .A2(n17345), .A3(n17344), .A4(n17343), .ZN(
        n17363) );
  AOI22_X1 U21424 ( .A1(n24158), .A2(\xmem_data[72][1] ), .B1(n24157), .B2(
        \xmem_data[73][1] ), .ZN(n17350) );
  AOI22_X1 U21425 ( .A1(n24159), .A2(\xmem_data[74][1] ), .B1(n17041), .B2(
        \xmem_data[75][1] ), .ZN(n17349) );
  AOI22_X1 U21426 ( .A1(n24160), .A2(\xmem_data[76][1] ), .B1(n25461), .B2(
        \xmem_data[77][1] ), .ZN(n17348) );
  AOI22_X1 U21427 ( .A1(n29279), .A2(\xmem_data[78][1] ), .B1(n22676), .B2(
        \xmem_data[79][1] ), .ZN(n17347) );
  NAND4_X1 U21428 ( .A1(n17350), .A2(n17349), .A3(n17348), .A4(n17347), .ZN(
        n17362) );
  AOI22_X1 U21429 ( .A1(n24219), .A2(\xmem_data[80][1] ), .B1(n28687), .B2(
        \xmem_data[81][1] ), .ZN(n17354) );
  AOI22_X1 U21430 ( .A1(n24165), .A2(\xmem_data[82][1] ), .B1(n24548), .B2(
        \xmem_data[83][1] ), .ZN(n17353) );
  AOI22_X1 U21431 ( .A1(n30495), .A2(\xmem_data[84][1] ), .B1(n30269), .B2(
        \xmem_data[85][1] ), .ZN(n17352) );
  AOI22_X1 U21432 ( .A1(n24167), .A2(\xmem_data[86][1] ), .B1(n24166), .B2(
        \xmem_data[87][1] ), .ZN(n17351) );
  NAND4_X1 U21433 ( .A1(n17354), .A2(n17353), .A3(n17352), .A4(n17351), .ZN(
        n17361) );
  AOI22_X1 U21434 ( .A1(n25723), .A2(\xmem_data[88][1] ), .B1(n20770), .B2(
        \xmem_data[89][1] ), .ZN(n17359) );
  AOI22_X1 U21435 ( .A1(n24686), .A2(\xmem_data[90][1] ), .B1(n30909), .B2(
        \xmem_data[91][1] ), .ZN(n17358) );
  AOI22_X1 U21436 ( .A1(n30571), .A2(\xmem_data[92][1] ), .B1(n3449), .B2(
        \xmem_data[93][1] ), .ZN(n17357) );
  AND2_X1 U21437 ( .A1(n24172), .A2(\xmem_data[94][1] ), .ZN(n17355) );
  AOI21_X1 U21438 ( .B1(n20991), .B2(\xmem_data[95][1] ), .A(n17355), .ZN(
        n17356) );
  NAND4_X1 U21439 ( .A1(n17359), .A2(n17358), .A3(n17357), .A4(n17356), .ZN(
        n17360) );
  OR4_X1 U21440 ( .A1(n17363), .A2(n17362), .A3(n17361), .A4(n17360), .ZN(
        n17364) );
  NAND2_X1 U21441 ( .A1(n17364), .A2(n24204), .ZN(n17365) );
  AOI22_X1 U21442 ( .A1(n3220), .A2(\xmem_data[0][0] ), .B1(n24139), .B2(
        \xmem_data[1][0] ), .ZN(n17372) );
  AOI22_X1 U21443 ( .A1(n28476), .A2(\xmem_data[2][0] ), .B1(n24141), .B2(
        \xmem_data[3][0] ), .ZN(n17371) );
  AOI22_X1 U21444 ( .A1(n24140), .A2(\xmem_data[4][0] ), .B1(n3128), .B2(
        \xmem_data[5][0] ), .ZN(n17370) );
  AOI22_X1 U21445 ( .A1(n30877), .A2(\xmem_data[6][0] ), .B1(n23813), .B2(
        \xmem_data[7][0] ), .ZN(n17369) );
  NAND4_X1 U21446 ( .A1(n17372), .A2(n17371), .A3(n17370), .A4(n17369), .ZN(
        n17388) );
  AOI22_X1 U21447 ( .A1(n24130), .A2(\xmem_data[8][0] ), .B1(n23762), .B2(
        \xmem_data[9][0] ), .ZN(n17376) );
  AOI22_X1 U21448 ( .A1(n24132), .A2(\xmem_data[10][0] ), .B1(n27537), .B2(
        \xmem_data[11][0] ), .ZN(n17375) );
  AOI22_X1 U21449 ( .A1(n22674), .A2(\xmem_data[12][0] ), .B1(n28336), .B2(
        \xmem_data[13][0] ), .ZN(n17374) );
  AOI22_X1 U21450 ( .A1(n24134), .A2(\xmem_data[14][0] ), .B1(n24133), .B2(
        \xmem_data[15][0] ), .ZN(n17373) );
  NAND4_X1 U21451 ( .A1(n17376), .A2(n17375), .A3(n17374), .A4(n17373), .ZN(
        n17387) );
  AOI22_X1 U21452 ( .A1(n16989), .A2(\xmem_data[16][0] ), .B1(n24115), .B2(
        \xmem_data[17][0] ), .ZN(n17380) );
  AOI22_X1 U21453 ( .A1(n24116), .A2(\xmem_data[18][0] ), .B1(n24615), .B2(
        \xmem_data[19][0] ), .ZN(n17379) );
  AOI22_X1 U21454 ( .A1(n24117), .A2(\xmem_data[20][0] ), .B1(n28202), .B2(
        \xmem_data[21][0] ), .ZN(n17378) );
  AOI22_X1 U21455 ( .A1(n24622), .A2(\xmem_data[22][0] ), .B1(n20782), .B2(
        \xmem_data[23][0] ), .ZN(n17377) );
  NAND4_X1 U21456 ( .A1(n17380), .A2(n17379), .A3(n17378), .A4(n17377), .ZN(
        n17386) );
  AOI22_X1 U21457 ( .A1(n25527), .A2(\xmem_data[24][0] ), .B1(n13420), .B2(
        \xmem_data[25][0] ), .ZN(n17384) );
  AOI22_X1 U21458 ( .A1(n24122), .A2(\xmem_data[26][0] ), .B1(n21061), .B2(
        \xmem_data[27][0] ), .ZN(n17383) );
  AOI22_X1 U21459 ( .A1(n29118), .A2(\xmem_data[28][0] ), .B1(n3433), .B2(
        \xmem_data[29][0] ), .ZN(n17382) );
  AOI22_X1 U21460 ( .A1(n30589), .A2(\xmem_data[30][0] ), .B1(n25730), .B2(
        \xmem_data[31][0] ), .ZN(n17381) );
  NAND4_X1 U21461 ( .A1(n17384), .A2(n17383), .A3(n17382), .A4(n17381), .ZN(
        n17385) );
  OR4_X1 U21462 ( .A1(n17388), .A2(n17387), .A3(n17386), .A4(n17385), .ZN(
        n17390) );
  AOI22_X1 U21463 ( .A1(n23781), .A2(\xmem_data[56][0] ), .B1(n27568), .B2(
        \xmem_data[57][0] ), .ZN(n17395) );
  AOI22_X1 U21464 ( .A1(n13487), .A2(\xmem_data[58][0] ), .B1(n28354), .B2(
        \xmem_data[59][0] ), .ZN(n17394) );
  AOI22_X1 U21465 ( .A1(n29328), .A2(\xmem_data[60][0] ), .B1(n3348), .B2(
        \xmem_data[61][0] ), .ZN(n17393) );
  AND2_X1 U21466 ( .A1(n27437), .A2(\xmem_data[62][0] ), .ZN(n17391) );
  AOI21_X1 U21467 ( .B1(n25413), .B2(\xmem_data[63][0] ), .A(n17391), .ZN(
        n17392) );
  NAND4_X1 U21468 ( .A1(n17395), .A2(n17394), .A3(n17393), .A4(n17392), .ZN(
        n17412) );
  AOI22_X1 U21469 ( .A1(n27943), .A2(\xmem_data[40][0] ), .B1(n28671), .B2(
        \xmem_data[41][0] ), .ZN(n17399) );
  AOI22_X1 U21470 ( .A1(n24212), .A2(\xmem_data[42][0] ), .B1(n16986), .B2(
        \xmem_data[43][0] ), .ZN(n17398) );
  AOI22_X1 U21471 ( .A1(n25606), .A2(\xmem_data[44][0] ), .B1(n30948), .B2(
        \xmem_data[45][0] ), .ZN(n17397) );
  AOI22_X1 U21472 ( .A1(n31269), .A2(\xmem_data[46][0] ), .B1(n24214), .B2(
        \xmem_data[47][0] ), .ZN(n17396) );
  NAND4_X1 U21473 ( .A1(n17399), .A2(n17398), .A3(n17397), .A4(n17396), .ZN(
        n17410) );
  AOI22_X1 U21474 ( .A1(n24219), .A2(\xmem_data[48][0] ), .B1(n28302), .B2(
        \xmem_data[49][0] ), .ZN(n17403) );
  AOI22_X1 U21475 ( .A1(n24221), .A2(\xmem_data[50][0] ), .B1(n30899), .B2(
        \xmem_data[51][0] ), .ZN(n17402) );
  AOI22_X1 U21476 ( .A1(n24222), .A2(\xmem_data[52][0] ), .B1(n20817), .B2(
        \xmem_data[53][0] ), .ZN(n17401) );
  AOI22_X1 U21477 ( .A1(n24223), .A2(\xmem_data[54][0] ), .B1(n20782), .B2(
        \xmem_data[55][0] ), .ZN(n17400) );
  NAND4_X1 U21478 ( .A1(n17403), .A2(n17402), .A3(n17401), .A4(n17400), .ZN(
        n17409) );
  AOI22_X1 U21479 ( .A1(n3222), .A2(\xmem_data[32][0] ), .B1(n17033), .B2(
        \xmem_data[33][0] ), .ZN(n17407) );
  AOI22_X1 U21480 ( .A1(n24207), .A2(\xmem_data[34][0] ), .B1(n22758), .B2(
        \xmem_data[35][0] ), .ZN(n17406) );
  AOI22_X1 U21481 ( .A1(n20559), .A2(\xmem_data[36][0] ), .B1(n3282), .B2(
        \xmem_data[37][0] ), .ZN(n17405) );
  AOI22_X1 U21482 ( .A1(n25450), .A2(\xmem_data[38][0] ), .B1(n25604), .B2(
        \xmem_data[39][0] ), .ZN(n17404) );
  NAND4_X1 U21483 ( .A1(n17407), .A2(n17406), .A3(n17405), .A4(n17404), .ZN(
        n17408) );
  AOI22_X1 U21484 ( .A1(n25359), .A2(\xmem_data[88][0] ), .B1(n28241), .B2(
        \xmem_data[89][0] ), .ZN(n17417) );
  AOI22_X1 U21485 ( .A1(n30498), .A2(\xmem_data[90][0] ), .B1(n25408), .B2(
        \xmem_data[91][0] ), .ZN(n17416) );
  AOI22_X1 U21486 ( .A1(n12471), .A2(\xmem_data[92][0] ), .B1(n3388), .B2(
        \xmem_data[93][0] ), .ZN(n17415) );
  AND2_X1 U21487 ( .A1(n24172), .A2(\xmem_data[94][0] ), .ZN(n17413) );
  AOI21_X1 U21488 ( .B1(n20576), .B2(\xmem_data[95][0] ), .A(n17413), .ZN(
        n17414) );
  NAND4_X1 U21489 ( .A1(n17417), .A2(n17416), .A3(n17415), .A4(n17414), .ZN(
        n17435) );
  AOI22_X1 U21490 ( .A1(n24158), .A2(\xmem_data[72][0] ), .B1(n24157), .B2(
        \xmem_data[73][0] ), .ZN(n17421) );
  AOI22_X1 U21491 ( .A1(n24159), .A2(\xmem_data[74][0] ), .B1(n17041), .B2(
        \xmem_data[75][0] ), .ZN(n17420) );
  AOI22_X1 U21492 ( .A1(n24160), .A2(\xmem_data[76][0] ), .B1(n3466), .B2(
        \xmem_data[77][0] ), .ZN(n17419) );
  AOI22_X1 U21493 ( .A1(n28993), .A2(\xmem_data[78][0] ), .B1(n20585), .B2(
        \xmem_data[79][0] ), .ZN(n17418) );
  NAND4_X1 U21494 ( .A1(n17421), .A2(n17420), .A3(n17419), .A4(n17418), .ZN(
        n17433) );
  AOI22_X1 U21495 ( .A1(n3220), .A2(\xmem_data[64][0] ), .B1(n22708), .B2(
        \xmem_data[65][0] ), .ZN(n17425) );
  AOI22_X1 U21496 ( .A1(n20500), .A2(\xmem_data[66][0] ), .B1(n23812), .B2(
        \xmem_data[67][0] ), .ZN(n17424) );
  AOI22_X1 U21497 ( .A1(n13444), .A2(\xmem_data[68][0] ), .B1(n17063), .B2(
        \xmem_data[69][0] ), .ZN(n17423) );
  AOI22_X1 U21498 ( .A1(n28045), .A2(\xmem_data[70][0] ), .B1(n28374), .B2(
        \xmem_data[71][0] ), .ZN(n17422) );
  NAND4_X1 U21499 ( .A1(n17425), .A2(n17424), .A3(n17423), .A4(n17422), .ZN(
        n17431) );
  AOI22_X1 U21500 ( .A1(n20505), .A2(\xmem_data[80][0] ), .B1(n28994), .B2(
        \xmem_data[81][0] ), .ZN(n17429) );
  AOI22_X1 U21501 ( .A1(n24165), .A2(\xmem_data[82][0] ), .B1(n24548), .B2(
        \xmem_data[83][0] ), .ZN(n17428) );
  AOI22_X1 U21502 ( .A1(n24117), .A2(\xmem_data[84][0] ), .B1(n25636), .B2(
        \xmem_data[85][0] ), .ZN(n17427) );
  AOI22_X1 U21503 ( .A1(n24167), .A2(\xmem_data[86][0] ), .B1(n24166), .B2(
        \xmem_data[87][0] ), .ZN(n17426) );
  NAND4_X1 U21504 ( .A1(n17429), .A2(n17428), .A3(n17427), .A4(n17426), .ZN(
        n17430) );
  AOI22_X1 U21505 ( .A1(n28500), .A2(\xmem_data[120][0] ), .B1(n29820), .B2(
        \xmem_data[121][0] ), .ZN(n17440) );
  AOI22_X1 U21506 ( .A1(n24624), .A2(\xmem_data[122][0] ), .B1(n30862), .B2(
        \xmem_data[123][0] ), .ZN(n17439) );
  AOI22_X1 U21507 ( .A1(n29118), .A2(\xmem_data[124][0] ), .B1(n3351), .B2(
        \xmem_data[125][0] ), .ZN(n17438) );
  AND2_X1 U21508 ( .A1(n24172), .A2(\xmem_data[126][0] ), .ZN(n17436) );
  AOI21_X1 U21509 ( .B1(n24694), .B2(\xmem_data[127][0] ), .A(n17436), .ZN(
        n17437) );
  NAND4_X1 U21510 ( .A1(n17440), .A2(n17439), .A3(n17438), .A4(n17437), .ZN(
        n17458) );
  AOI22_X1 U21511 ( .A1(n3220), .A2(\xmem_data[96][0] ), .B1(n24139), .B2(
        \xmem_data[97][0] ), .ZN(n17444) );
  AOI22_X1 U21512 ( .A1(n20787), .A2(\xmem_data[98][0] ), .B1(n23812), .B2(
        \xmem_data[99][0] ), .ZN(n17443) );
  AOI22_X1 U21513 ( .A1(n24140), .A2(\xmem_data[100][0] ), .B1(n17063), .B2(
        \xmem_data[101][0] ), .ZN(n17442) );
  AOI22_X1 U21514 ( .A1(n29103), .A2(\xmem_data[102][0] ), .B1(n28374), .B2(
        \xmem_data[103][0] ), .ZN(n17441) );
  NAND4_X1 U21515 ( .A1(n17444), .A2(n17443), .A3(n17442), .A4(n17441), .ZN(
        n17450) );
  AOI22_X1 U21516 ( .A1(n23796), .A2(\xmem_data[112][0] ), .B1(n24115), .B2(
        \xmem_data[113][0] ), .ZN(n17448) );
  AOI22_X1 U21517 ( .A1(n24165), .A2(\xmem_data[114][0] ), .B1(n25717), .B2(
        \xmem_data[115][0] ), .ZN(n17447) );
  AOI22_X1 U21518 ( .A1(n20943), .A2(\xmem_data[116][0] ), .B1(n3300), .B2(
        \xmem_data[117][0] ), .ZN(n17446) );
  AOI22_X1 U21519 ( .A1(n24167), .A2(\xmem_data[118][0] ), .B1(n24166), .B2(
        \xmem_data[119][0] ), .ZN(n17445) );
  NAND4_X1 U21520 ( .A1(n17448), .A2(n17447), .A3(n17446), .A4(n17445), .ZN(
        n17449) );
  AOI22_X1 U21521 ( .A1(n24158), .A2(\xmem_data[104][0] ), .B1(n24157), .B2(
        \xmem_data[105][0] ), .ZN(n17454) );
  AOI22_X1 U21522 ( .A1(n24159), .A2(\xmem_data[106][0] ), .B1(n23763), .B2(
        \xmem_data[107][0] ), .ZN(n17453) );
  AOI22_X1 U21523 ( .A1(n24160), .A2(\xmem_data[108][0] ), .B1(n3121), .B2(
        \xmem_data[109][0] ), .ZN(n17452) );
  AOI22_X1 U21524 ( .A1(n25383), .A2(\xmem_data[110][0] ), .B1(n20585), .B2(
        \xmem_data[111][0] ), .ZN(n17451) );
  NAND4_X1 U21525 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17455) );
  XOR2_X1 U21526 ( .A(\fmem_data[13][6] ), .B(\fmem_data[13][7] ), .Z(n17463)
         );
  AOI22_X1 U21527 ( .A1(n3334), .A2(\xmem_data[96][0] ), .B1(n29173), .B2(
        \xmem_data[97][0] ), .ZN(n17468) );
  AOI22_X1 U21528 ( .A1(n24532), .A2(\xmem_data[98][0] ), .B1(n3219), .B2(
        \xmem_data[99][0] ), .ZN(n17467) );
  AOI22_X1 U21529 ( .A1(n24533), .A2(\xmem_data[100][0] ), .B1(n20598), .B2(
        \xmem_data[101][0] ), .ZN(n17466) );
  AOI22_X1 U21530 ( .A1(n24534), .A2(\xmem_data[102][0] ), .B1(n28372), .B2(
        \xmem_data[103][0] ), .ZN(n17465) );
  NAND4_X1 U21531 ( .A1(n17468), .A2(n17467), .A3(n17466), .A4(n17465), .ZN(
        n17484) );
  AOI22_X1 U21532 ( .A1(n3375), .A2(\xmem_data[104][0] ), .B1(n28045), .B2(
        \xmem_data[105][0] ), .ZN(n17472) );
  AOI22_X1 U21533 ( .A1(n27551), .A2(\xmem_data[106][0] ), .B1(n28481), .B2(
        \xmem_data[107][0] ), .ZN(n17471) );
  AOI22_X1 U21534 ( .A1(n27911), .A2(\xmem_data[108][0] ), .B1(n24516), .B2(
        \xmem_data[109][0] ), .ZN(n17470) );
  AOI22_X1 U21535 ( .A1(n3175), .A2(\xmem_data[110][0] ), .B1(n20544), .B2(
        \xmem_data[111][0] ), .ZN(n17469) );
  NAND4_X1 U21536 ( .A1(n17472), .A2(n17471), .A3(n17470), .A4(n17469), .ZN(
        n17483) );
  AOI22_X1 U21537 ( .A1(n25461), .A2(\xmem_data[112][0] ), .B1(n27454), .B2(
        \xmem_data[113][0] ), .ZN(n17476) );
  AOI22_X1 U21538 ( .A1(n24509), .A2(\xmem_data[114][0] ), .B1(n24459), .B2(
        \xmem_data[115][0] ), .ZN(n17475) );
  AOI22_X1 U21539 ( .A1(n20815), .A2(\xmem_data[116][0] ), .B1(n24510), .B2(
        \xmem_data[117][0] ), .ZN(n17474) );
  AOI22_X1 U21540 ( .A1(n24511), .A2(\xmem_data[118][0] ), .B1(n25364), .B2(
        \xmem_data[119][0] ), .ZN(n17473) );
  NAND4_X1 U21541 ( .A1(n17476), .A2(n17475), .A3(n17474), .A4(n17473), .ZN(
        n17482) );
  AOI22_X1 U21542 ( .A1(n24522), .A2(\xmem_data[120][0] ), .B1(n24521), .B2(
        \xmem_data[121][0] ), .ZN(n17480) );
  AOI22_X1 U21543 ( .A1(n3209), .A2(\xmem_data[122][0] ), .B1(n17049), .B2(
        \xmem_data[123][0] ), .ZN(n17479) );
  AOI22_X1 U21544 ( .A1(n29327), .A2(\xmem_data[124][0] ), .B1(n24524), .B2(
        \xmem_data[125][0] ), .ZN(n17478) );
  AOI22_X1 U21545 ( .A1(n24526), .A2(\xmem_data[126][0] ), .B1(n24525), .B2(
        \xmem_data[127][0] ), .ZN(n17477) );
  NAND4_X1 U21546 ( .A1(n17480), .A2(n17479), .A3(n17478), .A4(n17477), .ZN(
        n17481) );
  OR4_X1 U21547 ( .A1(n17484), .A2(n17483), .A3(n17482), .A4(n17481), .ZN(
        n17506) );
  AOI22_X1 U21548 ( .A1(n22728), .A2(\xmem_data[64][0] ), .B1(n24439), .B2(
        \xmem_data[65][0] ), .ZN(n17488) );
  AOI22_X1 U21549 ( .A1(n24532), .A2(\xmem_data[66][0] ), .B1(n3218), .B2(
        \xmem_data[67][0] ), .ZN(n17487) );
  AOI22_X1 U21550 ( .A1(n24533), .A2(\xmem_data[68][0] ), .B1(n25509), .B2(
        \xmem_data[69][0] ), .ZN(n17486) );
  AOI22_X1 U21551 ( .A1(n24534), .A2(\xmem_data[70][0] ), .B1(n20559), .B2(
        \xmem_data[71][0] ), .ZN(n17485) );
  NAND4_X1 U21552 ( .A1(n17488), .A2(n17487), .A3(n17486), .A4(n17485), .ZN(
        n17504) );
  AOI22_X1 U21553 ( .A1(n25451), .A2(\xmem_data[72][0] ), .B1(n25514), .B2(
        \xmem_data[73][0] ), .ZN(n17492) );
  AOI22_X1 U21554 ( .A1(n27551), .A2(\xmem_data[74][0] ), .B1(n3358), .B2(
        \xmem_data[75][0] ), .ZN(n17491) );
  AOI22_X1 U21555 ( .A1(n28233), .A2(\xmem_data[76][0] ), .B1(n24516), .B2(
        \xmem_data[77][0] ), .ZN(n17490) );
  AOI22_X1 U21556 ( .A1(n3175), .A2(\xmem_data[78][0] ), .B1(n24160), .B2(
        \xmem_data[79][0] ), .ZN(n17489) );
  NAND4_X1 U21557 ( .A1(n17492), .A2(n17491), .A3(n17490), .A4(n17489), .ZN(
        n17503) );
  AOI22_X1 U21558 ( .A1(n27517), .A2(\xmem_data[80][0] ), .B1(n25460), .B2(
        \xmem_data[81][0] ), .ZN(n17496) );
  AOI22_X1 U21559 ( .A1(n24509), .A2(\xmem_data[82][0] ), .B1(n20940), .B2(
        \xmem_data[83][0] ), .ZN(n17495) );
  AOI22_X1 U21560 ( .A1(n20942), .A2(\xmem_data[84][0] ), .B1(n24510), .B2(
        \xmem_data[85][0] ), .ZN(n17494) );
  AOI22_X1 U21561 ( .A1(n24511), .A2(\xmem_data[86][0] ), .B1(n24222), .B2(
        \xmem_data[87][0] ), .ZN(n17493) );
  NAND4_X1 U21562 ( .A1(n17496), .A2(n17495), .A3(n17494), .A4(n17493), .ZN(
        n17502) );
  AOI22_X1 U21563 ( .A1(n24522), .A2(\xmem_data[88][0] ), .B1(n24521), .B2(
        \xmem_data[89][0] ), .ZN(n17500) );
  AOI22_X1 U21564 ( .A1(n3209), .A2(\xmem_data[90][0] ), .B1(n28468), .B2(
        \xmem_data[91][0] ), .ZN(n17499) );
  AOI22_X1 U21565 ( .A1(n30674), .A2(\xmem_data[92][0] ), .B1(n24524), .B2(
        \xmem_data[93][0] ), .ZN(n17498) );
  AOI22_X1 U21566 ( .A1(n24526), .A2(\xmem_data[94][0] ), .B1(n24525), .B2(
        \xmem_data[95][0] ), .ZN(n17497) );
  NAND4_X1 U21567 ( .A1(n17500), .A2(n17499), .A3(n17498), .A4(n17497), .ZN(
        n17501) );
  AOI22_X1 U21568 ( .A1(n24542), .A2(n17506), .B1(n24581), .B2(n17505), .ZN(
        n17554) );
  AOI22_X1 U21569 ( .A1(n3149), .A2(\xmem_data[32][0] ), .B1(n3247), .B2(
        \xmem_data[33][0] ), .ZN(n17510) );
  AOI22_X1 U21570 ( .A1(n24562), .A2(\xmem_data[34][0] ), .B1(n3222), .B2(
        \xmem_data[35][0] ), .ZN(n17509) );
  AOI22_X1 U21571 ( .A1(n24563), .A2(\xmem_data[36][0] ), .B1(n22667), .B2(
        \xmem_data[37][0] ), .ZN(n17508) );
  AOI22_X1 U21572 ( .A1(n24565), .A2(\xmem_data[38][0] ), .B1(n24564), .B2(
        \xmem_data[39][0] ), .ZN(n17507) );
  NAND4_X1 U21573 ( .A1(n17510), .A2(n17509), .A3(n17508), .A4(n17507), .ZN(
        n17526) );
  AOI22_X1 U21574 ( .A1(n30295), .A2(\xmem_data[40][0] ), .B1(n24553), .B2(
        \xmem_data[41][0] ), .ZN(n17514) );
  AOI22_X1 U21575 ( .A1(n24554), .A2(\xmem_data[42][0] ), .B1(n25481), .B2(
        \xmem_data[43][0] ), .ZN(n17513) );
  AOI22_X1 U21576 ( .A1(n24556), .A2(\xmem_data[44][0] ), .B1(n24555), .B2(
        \xmem_data[45][0] ), .ZN(n17512) );
  AOI22_X1 U21577 ( .A1(n17041), .A2(\xmem_data[46][0] ), .B1(n30541), .B2(
        \xmem_data[47][0] ), .ZN(n17511) );
  NAND4_X1 U21578 ( .A1(n17514), .A2(n17513), .A3(n17512), .A4(n17511), .ZN(
        n17525) );
  AOI22_X1 U21579 ( .A1(n24545), .A2(\xmem_data[48][0] ), .B1(n28993), .B2(
        \xmem_data[49][0] ), .ZN(n17518) );
  AOI22_X1 U21580 ( .A1(n24547), .A2(\xmem_data[50][0] ), .B1(n24546), .B2(
        \xmem_data[51][0] ), .ZN(n17517) );
  AOI22_X1 U21581 ( .A1(n29047), .A2(\xmem_data[52][0] ), .B1(n28097), .B2(
        \xmem_data[53][0] ), .ZN(n17516) );
  AOI22_X1 U21582 ( .A1(n24548), .A2(\xmem_data[54][0] ), .B1(n25716), .B2(
        \xmem_data[55][0] ), .ZN(n17515) );
  NAND4_X1 U21583 ( .A1(n17518), .A2(n17517), .A3(n17516), .A4(n17515), .ZN(
        n17524) );
  AOI22_X1 U21584 ( .A1(n24571), .A2(\xmem_data[56][0] ), .B1(n24570), .B2(
        \xmem_data[57][0] ), .ZN(n17522) );
  AOI22_X1 U21585 ( .A1(n24572), .A2(\xmem_data[58][0] ), .B1(n25723), .B2(
        \xmem_data[59][0] ), .ZN(n17521) );
  AOI22_X1 U21586 ( .A1(n21060), .A2(\xmem_data[60][0] ), .B1(n22727), .B2(
        \xmem_data[61][0] ), .ZN(n17520) );
  AOI22_X1 U21587 ( .A1(n28038), .A2(\xmem_data[62][0] ), .B1(n24573), .B2(
        \xmem_data[63][0] ), .ZN(n17519) );
  NAND4_X1 U21588 ( .A1(n17522), .A2(n17521), .A3(n17520), .A4(n17519), .ZN(
        n17523) );
  OR4_X1 U21589 ( .A1(n17526), .A2(n17525), .A3(n17524), .A4(n17523), .ZN(
        n17527) );
  AOI22_X1 U21590 ( .A1(n3144), .A2(\xmem_data[0][0] ), .B1(n24439), .B2(
        \xmem_data[1][0] ), .ZN(n17531) );
  AOI22_X1 U21591 ( .A1(n24443), .A2(\xmem_data[2][0] ), .B1(n3221), .B2(
        \xmem_data[3][0] ), .ZN(n17530) );
  AOI22_X1 U21592 ( .A1(n30278), .A2(\xmem_data[4][0] ), .B1(n29095), .B2(
        \xmem_data[5][0] ), .ZN(n17529) );
  AOI22_X1 U21593 ( .A1(n24438), .A2(\xmem_data[6][0] ), .B1(n30882), .B2(
        \xmem_data[7][0] ), .ZN(n17528) );
  AND4_X1 U21594 ( .A1(n17531), .A2(n17530), .A3(n17529), .A4(n17528), .ZN(
        n17544) );
  AOI22_X1 U21595 ( .A1(n3338), .A2(\xmem_data[24][0] ), .B1(n20781), .B2(
        \xmem_data[25][0] ), .ZN(n17535) );
  AOI22_X1 U21596 ( .A1(n24467), .A2(\xmem_data[26][0] ), .B1(n27526), .B2(
        \xmem_data[27][0] ), .ZN(n17534) );
  AOI22_X1 U21597 ( .A1(n29820), .A2(\xmem_data[28][0] ), .B1(n24468), .B2(
        \xmem_data[29][0] ), .ZN(n17533) );
  AOI22_X1 U21598 ( .A1(n30862), .A2(\xmem_data[30][0] ), .B1(n24470), .B2(
        \xmem_data[31][0] ), .ZN(n17532) );
  NAND4_X1 U21599 ( .A1(n17535), .A2(n17534), .A3(n17533), .A4(n17532), .ZN(
        n17542) );
  AOI22_X1 U21600 ( .A1(n29451), .A2(\xmem_data[12][0] ), .B1(n24448), .B2(
        \xmem_data[13][0] ), .ZN(n17536) );
  INV_X1 U21601 ( .A(n17536), .ZN(n17541) );
  AOI22_X1 U21602 ( .A1(n16986), .A2(\xmem_data[14][0] ), .B1(n24160), .B2(
        \xmem_data[15][0] ), .ZN(n17539) );
  AOI22_X1 U21603 ( .A1(n24450), .A2(\xmem_data[10][0] ), .B1(n30884), .B2(
        \xmem_data[11][0] ), .ZN(n17538) );
  NAND2_X1 U21604 ( .A1(n3132), .A2(\xmem_data[8][0] ), .ZN(n17537) );
  NAND3_X1 U21605 ( .A1(n17539), .A2(n17538), .A3(n17537), .ZN(n17540) );
  NOR3_X1 U21606 ( .A1(n17542), .A2(n17541), .A3(n17540), .ZN(n17543) );
  NAND2_X1 U21607 ( .A1(n17544), .A2(n17543), .ZN(n17551) );
  AOI22_X1 U21608 ( .A1(n24458), .A2(\xmem_data[16][0] ), .B1(n24457), .B2(
        \xmem_data[17][0] ), .ZN(n17548) );
  AOI22_X1 U21609 ( .A1(n23717), .A2(\xmem_data[18][0] ), .B1(n24459), .B2(
        \xmem_data[19][0] ), .ZN(n17547) );
  AOI22_X1 U21610 ( .A1(n28994), .A2(\xmem_data[20][0] ), .B1(n24460), .B2(
        \xmem_data[21][0] ), .ZN(n17546) );
  AOI22_X1 U21611 ( .A1(n3178), .A2(\xmem_data[22][0] ), .B1(n20551), .B2(
        \xmem_data[23][0] ), .ZN(n17545) );
  NAND4_X1 U21612 ( .A1(n17548), .A2(n17547), .A3(n17546), .A4(n17545), .ZN(
        n17549) );
  XNOR2_X1 U21613 ( .A(n31704), .B(\fmem_data[17][3] ), .ZN(n32646) );
  XNOR2_X1 U21614 ( .A(n32543), .B(\fmem_data[17][3] ), .ZN(n30791) );
  OAI22_X1 U21615 ( .A1(n32646), .A2(n33250), .B1(n33249), .B2(n30791), .ZN(
        n26383) );
  AOI22_X1 U21616 ( .A1(n29231), .A2(\xmem_data[96][1] ), .B1(n28510), .B2(
        \xmem_data[97][1] ), .ZN(n17560) );
  AOI22_X1 U21617 ( .A1(n27447), .A2(\xmem_data[98][1] ), .B1(n13475), .B2(
        \xmem_data[99][1] ), .ZN(n17559) );
  AOI22_X1 U21618 ( .A1(n20716), .A2(\xmem_data[100][1] ), .B1(n29232), .B2(
        \xmem_data[101][1] ), .ZN(n17558) );
  AOI22_X1 U21619 ( .A1(n31268), .A2(\xmem_data[102][1] ), .B1(n23793), .B2(
        \xmem_data[103][1] ), .ZN(n17557) );
  NAND4_X1 U21620 ( .A1(n17560), .A2(n17559), .A3(n17558), .A4(n17557), .ZN(
        n17576) );
  AOI22_X1 U21621 ( .A1(n24213), .A2(\xmem_data[104][1] ), .B1(n3208), .B2(
        \xmem_data[105][1] ), .ZN(n17564) );
  AOI22_X1 U21622 ( .A1(n24509), .A2(\xmem_data[106][1] ), .B1(n24459), .B2(
        \xmem_data[107][1] ), .ZN(n17563) );
  AOI22_X1 U21623 ( .A1(n29239), .A2(\xmem_data[108][1] ), .B1(n29238), .B2(
        \xmem_data[109][1] ), .ZN(n17562) );
  AOI22_X1 U21624 ( .A1(n29240), .A2(\xmem_data[110][1] ), .B1(n20506), .B2(
        \xmem_data[111][1] ), .ZN(n17561) );
  NAND4_X1 U21625 ( .A1(n17564), .A2(n17563), .A3(n17562), .A4(n17561), .ZN(
        n17575) );
  AOI22_X1 U21626 ( .A1(n29246), .A2(\xmem_data[112][1] ), .B1(n29245), .B2(
        \xmem_data[113][1] ), .ZN(n17568) );
  AOI22_X1 U21627 ( .A1(n3172), .A2(\xmem_data[114][1] ), .B1(n29247), .B2(
        \xmem_data[115][1] ), .ZN(n17567) );
  AOI22_X1 U21628 ( .A1(n29657), .A2(\xmem_data[116][1] ), .B1(n29248), .B2(
        \xmem_data[117][1] ), .ZN(n17566) );
  AOI22_X1 U21629 ( .A1(n30909), .A2(\xmem_data[118][1] ), .B1(n27499), .B2(
        \xmem_data[119][1] ), .ZN(n17565) );
  NAND4_X1 U21630 ( .A1(n17568), .A2(n17567), .A3(n17566), .A4(n17565), .ZN(
        n17574) );
  AOI22_X1 U21631 ( .A1(n20828), .A2(\xmem_data[120][1] ), .B1(n29253), .B2(
        \xmem_data[121][1] ), .ZN(n17572) );
  AOI22_X1 U21632 ( .A1(n29254), .A2(\xmem_data[122][1] ), .B1(n3220), .B2(
        \xmem_data[123][1] ), .ZN(n17571) );
  AOI22_X1 U21633 ( .A1(n29256), .A2(\xmem_data[124][1] ), .B1(n29255), .B2(
        \xmem_data[125][1] ), .ZN(n17570) );
  AOI22_X1 U21634 ( .A1(n29257), .A2(\xmem_data[126][1] ), .B1(n29181), .B2(
        \xmem_data[127][1] ), .ZN(n17569) );
  NAND4_X1 U21635 ( .A1(n17572), .A2(n17571), .A3(n17570), .A4(n17569), .ZN(
        n17573) );
  OR4_X1 U21636 ( .A1(n17576), .A2(n17575), .A3(n17574), .A4(n17573), .ZN(
        n17598) );
  AOI22_X1 U21637 ( .A1(n29231), .A2(\xmem_data[64][1] ), .B1(n28045), .B2(
        \xmem_data[65][1] ), .ZN(n17580) );
  AOI22_X1 U21638 ( .A1(n27447), .A2(\xmem_data[66][1] ), .B1(n20982), .B2(
        \xmem_data[67][1] ), .ZN(n17579) );
  AOI22_X1 U21639 ( .A1(n28051), .A2(\xmem_data[68][1] ), .B1(n29232), .B2(
        \xmem_data[69][1] ), .ZN(n17578) );
  AOI22_X1 U21640 ( .A1(n3176), .A2(\xmem_data[70][1] ), .B1(n22741), .B2(
        \xmem_data[71][1] ), .ZN(n17577) );
  NAND4_X1 U21641 ( .A1(n17580), .A2(n17579), .A3(n17578), .A4(n17577), .ZN(
        n17596) );
  AOI22_X1 U21642 ( .A1(n24213), .A2(\xmem_data[72][1] ), .B1(n28335), .B2(
        \xmem_data[73][1] ), .ZN(n17584) );
  AOI22_X1 U21643 ( .A1(n24509), .A2(\xmem_data[74][1] ), .B1(n31329), .B2(
        \xmem_data[75][1] ), .ZN(n17583) );
  AOI22_X1 U21644 ( .A1(n29239), .A2(\xmem_data[76][1] ), .B1(n29238), .B2(
        \xmem_data[77][1] ), .ZN(n17582) );
  AOI22_X1 U21645 ( .A1(n29240), .A2(\xmem_data[78][1] ), .B1(n30598), .B2(
        \xmem_data[79][1] ), .ZN(n17581) );
  NAND4_X1 U21646 ( .A1(n17584), .A2(n17583), .A3(n17582), .A4(n17581), .ZN(
        n17595) );
  AOI22_X1 U21647 ( .A1(n29246), .A2(\xmem_data[80][1] ), .B1(n29245), .B2(
        \xmem_data[81][1] ), .ZN(n17588) );
  AOI22_X1 U21648 ( .A1(n21058), .A2(\xmem_data[82][1] ), .B1(n29247), .B2(
        \xmem_data[83][1] ), .ZN(n17587) );
  AOI22_X1 U21649 ( .A1(n14982), .A2(\xmem_data[84][1] ), .B1(n29248), .B2(
        \xmem_data[85][1] ), .ZN(n17586) );
  AOI22_X1 U21650 ( .A1(n17056), .A2(\xmem_data[86][1] ), .B1(n31346), .B2(
        \xmem_data[87][1] ), .ZN(n17585) );
  NAND4_X1 U21651 ( .A1(n17588), .A2(n17587), .A3(n17586), .A4(n17585), .ZN(
        n17594) );
  AOI22_X1 U21652 ( .A1(n29661), .A2(\xmem_data[88][1] ), .B1(n29253), .B2(
        \xmem_data[89][1] ), .ZN(n17592) );
  AOI22_X1 U21653 ( .A1(n29254), .A2(\xmem_data[90][1] ), .B1(n3217), .B2(
        \xmem_data[91][1] ), .ZN(n17591) );
  AOI22_X1 U21654 ( .A1(n29256), .A2(\xmem_data[92][1] ), .B1(n29255), .B2(
        \xmem_data[93][1] ), .ZN(n17590) );
  AOI22_X1 U21655 ( .A1(n29257), .A2(\xmem_data[94][1] ), .B1(n28509), .B2(
        \xmem_data[95][1] ), .ZN(n17589) );
  NAND4_X1 U21656 ( .A1(n17592), .A2(n17591), .A3(n17590), .A4(n17589), .ZN(
        n17593) );
  OR4_X1 U21657 ( .A1(n17596), .A2(n17595), .A3(n17594), .A4(n17593), .ZN(
        n17597) );
  AOI22_X1 U21658 ( .A1(n29269), .A2(n17598), .B1(n29267), .B2(n17597), .ZN(
        n17649) );
  AOI22_X1 U21659 ( .A1(n3126), .A2(\xmem_data[32][1] ), .B1(n28045), .B2(
        \xmem_data[33][1] ), .ZN(n17602) );
  AOI22_X1 U21660 ( .A1(n16974), .A2(\xmem_data[34][1] ), .B1(n29307), .B2(
        \xmem_data[35][1] ), .ZN(n17601) );
  AOI22_X1 U21661 ( .A1(n29308), .A2(\xmem_data[36][1] ), .B1(n13168), .B2(
        \xmem_data[37][1] ), .ZN(n17600) );
  AOI22_X1 U21662 ( .A1(n29310), .A2(\xmem_data[38][1] ), .B1(n29309), .B2(
        \xmem_data[39][1] ), .ZN(n17599) );
  NAND4_X1 U21663 ( .A1(n17602), .A2(n17601), .A3(n17600), .A4(n17599), .ZN(
        n17618) );
  AOI22_X1 U21664 ( .A1(n28053), .A2(\xmem_data[40][1] ), .B1(n27516), .B2(
        \xmem_data[41][1] ), .ZN(n17606) );
  AOI22_X1 U21665 ( .A1(n29317), .A2(\xmem_data[42][1] ), .B1(n29316), .B2(
        \xmem_data[43][1] ), .ZN(n17605) );
  AOI22_X1 U21666 ( .A1(n29319), .A2(\xmem_data[44][1] ), .B1(n29318), .B2(
        \xmem_data[45][1] ), .ZN(n17604) );
  AOI22_X1 U21667 ( .A1(n25717), .A2(\xmem_data[46][1] ), .B1(n17001), .B2(
        \xmem_data[47][1] ), .ZN(n17603) );
  NAND4_X1 U21668 ( .A1(n17606), .A2(n17605), .A3(n17604), .A4(n17603), .ZN(
        n17617) );
  AOI22_X1 U21669 ( .A1(n29324), .A2(\xmem_data[48][1] ), .B1(n14975), .B2(
        \xmem_data[49][1] ), .ZN(n17610) );
  AOI22_X1 U21670 ( .A1(n29325), .A2(\xmem_data[50][1] ), .B1(n27463), .B2(
        \xmem_data[51][1] ), .ZN(n17609) );
  AOI22_X1 U21671 ( .A1(n29327), .A2(\xmem_data[52][1] ), .B1(n29326), .B2(
        \xmem_data[53][1] ), .ZN(n17608) );
  AOI22_X1 U21672 ( .A1(n28076), .A2(\xmem_data[54][1] ), .B1(n29328), .B2(
        \xmem_data[55][1] ), .ZN(n17607) );
  NAND4_X1 U21673 ( .A1(n17610), .A2(n17609), .A3(n17608), .A4(n17607), .ZN(
        n17616) );
  AOI22_X1 U21674 ( .A1(n3383), .A2(\xmem_data[56][1] ), .B1(n25442), .B2(
        \xmem_data[57][1] ), .ZN(n17614) );
  AOI22_X1 U21675 ( .A1(n28082), .A2(\xmem_data[58][1] ), .B1(n3218), .B2(
        \xmem_data[59][1] ), .ZN(n17613) );
  AOI22_X1 U21676 ( .A1(n24139), .A2(\xmem_data[60][1] ), .B1(n23739), .B2(
        \xmem_data[61][1] ), .ZN(n17612) );
  AOI22_X1 U21677 ( .A1(n25416), .A2(\xmem_data[62][1] ), .B1(n28342), .B2(
        \xmem_data[63][1] ), .ZN(n17611) );
  NAND4_X1 U21678 ( .A1(n17614), .A2(n17613), .A3(n17612), .A4(n17611), .ZN(
        n17615) );
  OR4_X1 U21679 ( .A1(n17618), .A2(n17617), .A3(n17616), .A4(n17615), .ZN(
        n17619) );
  NAND2_X1 U21680 ( .A1(n17619), .A2(n29343), .ZN(n17648) );
  AOI22_X1 U21681 ( .A1(n25441), .A2(\xmem_data[22][1] ), .B1(n31309), .B2(
        \xmem_data[23][1] ), .ZN(n17620) );
  INV_X1 U21682 ( .A(n17620), .ZN(n17623) );
  AOI22_X1 U21683 ( .A1(n24443), .A2(\xmem_data[26][1] ), .B1(n3218), .B2(
        \xmem_data[27][1] ), .ZN(n17621) );
  INV_X1 U21684 ( .A(n17621), .ZN(n17622) );
  NOR2_X1 U21685 ( .A1(n17623), .A2(n17622), .ZN(n17645) );
  AOI22_X1 U21686 ( .A1(n29807), .A2(\xmem_data[8][1] ), .B1(n29279), .B2(
        \xmem_data[9][1] ), .ZN(n17627) );
  AOI22_X1 U21687 ( .A1(n25434), .A2(\xmem_data[10][1] ), .B1(n25398), .B2(
        \xmem_data[11][1] ), .ZN(n17626) );
  AOI22_X1 U21688 ( .A1(n29319), .A2(\xmem_data[12][1] ), .B1(n29280), .B2(
        \xmem_data[13][1] ), .ZN(n17625) );
  AOI22_X1 U21689 ( .A1(n28460), .A2(\xmem_data[14][1] ), .B1(n27856), .B2(
        \xmem_data[15][1] ), .ZN(n17624) );
  AOI22_X1 U21690 ( .A1(n29298), .A2(\xmem_data[20][1] ), .B1(n27957), .B2(
        \xmem_data[21][1] ), .ZN(n17644) );
  AOI22_X1 U21691 ( .A1(n28743), .A2(\xmem_data[4][1] ), .B1(n29232), .B2(
        \xmem_data[5][1] ), .ZN(n17630) );
  AOI22_X1 U21692 ( .A1(n29272), .A2(\xmem_data[6][1] ), .B1(n29271), .B2(
        \xmem_data[7][1] ), .ZN(n17629) );
  AOI22_X1 U21693 ( .A1(n24638), .A2(\xmem_data[2][1] ), .B1(n29307), .B2(
        \xmem_data[3][1] ), .ZN(n17628) );
  NAND3_X1 U21694 ( .A1(n17630), .A2(n17629), .A3(n17628), .ZN(n17642) );
  NAND2_X1 U21695 ( .A1(n28007), .A2(\xmem_data[1][1] ), .ZN(n17632) );
  AOI22_X1 U21696 ( .A1(n29297), .A2(\xmem_data[16][1] ), .B1(n29126), .B2(
        \xmem_data[17][1] ), .ZN(n17631) );
  NAND2_X1 U21697 ( .A1(n17632), .A2(n17631), .ZN(n17636) );
  AND2_X1 U21698 ( .A1(n29350), .A2(\xmem_data[0][1] ), .ZN(n17635) );
  AOI22_X1 U21699 ( .A1(n3335), .A2(\xmem_data[24][1] ), .B1(n29286), .B2(
        \xmem_data[25][1] ), .ZN(n17633) );
  INV_X1 U21700 ( .A(n17633), .ZN(n17634) );
  NOR3_X1 U21701 ( .A1(n17636), .A2(n17635), .A3(n17634), .ZN(n17640) );
  AOI22_X1 U21702 ( .A1(n29289), .A2(\xmem_data[30][1] ), .B1(n30882), .B2(
        \xmem_data[31][1] ), .ZN(n17639) );
  AOI22_X1 U21703 ( .A1(n29288), .A2(\xmem_data[28][1] ), .B1(n25509), .B2(
        \xmem_data[29][1] ), .ZN(n17638) );
  AOI22_X1 U21704 ( .A1(n24606), .A2(\xmem_data[18][1] ), .B1(n28468), .B2(
        \xmem_data[19][1] ), .ZN(n17637) );
  NAND4_X1 U21705 ( .A1(n17640), .A2(n17639), .A3(n17638), .A4(n17637), .ZN(
        n17641) );
  NOR2_X1 U21706 ( .A1(n17642), .A2(n17641), .ZN(n17643) );
  NAND4_X1 U21707 ( .A1(n17645), .A2(n3819), .A3(n17644), .A4(n17643), .ZN(
        n17646) );
  NAND2_X1 U21708 ( .A1(n17646), .A2(n25790), .ZN(n17647) );
  AOI22_X1 U21709 ( .A1(n28036), .A2(\xmem_data[116][0] ), .B1(n29248), .B2(
        \xmem_data[117][0] ), .ZN(n17652) );
  AOI22_X1 U21710 ( .A1(n29257), .A2(\xmem_data[126][0] ), .B1(n27903), .B2(
        \xmem_data[127][0] ), .ZN(n17651) );
  AOI22_X1 U21711 ( .A1(n29256), .A2(\xmem_data[124][0] ), .B1(n29255), .B2(
        \xmem_data[125][0] ), .ZN(n17650) );
  NAND3_X1 U21712 ( .A1(n17652), .A2(n17651), .A3(n17650), .ZN(n17655) );
  AOI22_X1 U21713 ( .A1(n3380), .A2(\xmem_data[118][0] ), .B1(n22752), .B2(
        \xmem_data[119][0] ), .ZN(n17653) );
  INV_X1 U21714 ( .A(n17653), .ZN(n17654) );
  AOI22_X1 U21715 ( .A1(n23795), .A2(\xmem_data[104][0] ), .B1(n20543), .B2(
        \xmem_data[105][0] ), .ZN(n17659) );
  AOI22_X1 U21716 ( .A1(n21007), .A2(\xmem_data[106][0] ), .B1(n17043), .B2(
        \xmem_data[107][0] ), .ZN(n17658) );
  AOI22_X1 U21717 ( .A1(n29239), .A2(\xmem_data[108][0] ), .B1(n29238), .B2(
        \xmem_data[109][0] ), .ZN(n17657) );
  AOI22_X1 U21718 ( .A1(n29240), .A2(\xmem_data[110][0] ), .B1(n25581), .B2(
        \xmem_data[111][0] ), .ZN(n17656) );
  NAND4_X1 U21719 ( .A1(n17659), .A2(n17658), .A3(n17657), .A4(n17656), .ZN(
        n17664) );
  AOI22_X1 U21720 ( .A1(n27542), .A2(\xmem_data[114][0] ), .B1(n29247), .B2(
        \xmem_data[115][0] ), .ZN(n17662) );
  AOI22_X1 U21721 ( .A1(n29246), .A2(\xmem_data[112][0] ), .B1(n29245), .B2(
        \xmem_data[113][0] ), .ZN(n17661) );
  AOI22_X1 U21722 ( .A1(n30864), .A2(\xmem_data[120][0] ), .B1(n29253), .B2(
        \xmem_data[121][0] ), .ZN(n17660) );
  NOR2_X1 U21723 ( .A1(n17664), .A2(n17663), .ZN(n17670) );
  AOI22_X1 U21724 ( .A1(n29254), .A2(\xmem_data[122][0] ), .B1(n3215), .B2(
        \xmem_data[123][0] ), .ZN(n17669) );
  AOI22_X1 U21725 ( .A1(n29231), .A2(\xmem_data[96][0] ), .B1(n13474), .B2(
        \xmem_data[97][0] ), .ZN(n17668) );
  AOI22_X1 U21726 ( .A1(n27447), .A2(\xmem_data[98][0] ), .B1(n28481), .B2(
        \xmem_data[99][0] ), .ZN(n17667) );
  AOI22_X1 U21727 ( .A1(n28089), .A2(\xmem_data[100][0] ), .B1(n29232), .B2(
        \xmem_data[101][0] ), .ZN(n17666) );
  AOI22_X1 U21728 ( .A1(n28980), .A2(\xmem_data[102][0] ), .B1(n20544), .B2(
        \xmem_data[103][0] ), .ZN(n17665) );
  OAI21_X1 U21729 ( .B1(n3991), .B2(n17671), .A(n29269), .ZN(n17742) );
  AND2_X1 U21730 ( .A1(n29326), .A2(\xmem_data[53][0] ), .ZN(n17672) );
  AOI21_X1 U21731 ( .B1(n29327), .B2(\xmem_data[52][0] ), .A(n17672), .ZN(
        n17673) );
  INV_X1 U21732 ( .A(n17673), .ZN(n17682) );
  AOI22_X1 U21733 ( .A1(n20807), .A2(\xmem_data[62][0] ), .B1(n20993), .B2(
        \xmem_data[63][0] ), .ZN(n17675) );
  AOI22_X1 U21734 ( .A1(n24139), .A2(\xmem_data[60][0] ), .B1(n22667), .B2(
        \xmem_data[61][0] ), .ZN(n17674) );
  NAND2_X1 U21735 ( .A1(n17675), .A2(n17674), .ZN(n17680) );
  AOI22_X1 U21736 ( .A1(n29325), .A2(\xmem_data[50][0] ), .B1(n29247), .B2(
        \xmem_data[51][0] ), .ZN(n17678) );
  AOI22_X1 U21737 ( .A1(n29324), .A2(\xmem_data[48][0] ), .B1(n14975), .B2(
        \xmem_data[49][0] ), .ZN(n17677) );
  AOI22_X1 U21738 ( .A1(n3383), .A2(\xmem_data[56][0] ), .B1(n28501), .B2(
        \xmem_data[57][0] ), .ZN(n17676) );
  NAND3_X1 U21739 ( .A1(n17678), .A2(n17677), .A3(n17676), .ZN(n17679) );
  AOI22_X1 U21740 ( .A1(n3281), .A2(\xmem_data[32][0] ), .B1(n23771), .B2(
        \xmem_data[33][0] ), .ZN(n17686) );
  AOI22_X1 U21741 ( .A1(n25707), .A2(\xmem_data[34][0] ), .B1(n29307), .B2(
        \xmem_data[35][0] ), .ZN(n17685) );
  AOI22_X1 U21742 ( .A1(n29308), .A2(\xmem_data[36][0] ), .B1(n13168), .B2(
        \xmem_data[37][0] ), .ZN(n17684) );
  AOI22_X1 U21743 ( .A1(n29310), .A2(\xmem_data[38][0] ), .B1(n29309), .B2(
        \xmem_data[39][0] ), .ZN(n17683) );
  AOI22_X1 U21744 ( .A1(n30909), .A2(\xmem_data[54][0] ), .B1(n29328), .B2(
        \xmem_data[55][0] ), .ZN(n17692) );
  AOI22_X1 U21745 ( .A1(n24694), .A2(\xmem_data[58][0] ), .B1(n3222), .B2(
        \xmem_data[59][0] ), .ZN(n17691) );
  AOI22_X1 U21746 ( .A1(n20776), .A2(\xmem_data[40][0] ), .B1(n27989), .B2(
        \xmem_data[41][0] ), .ZN(n17690) );
  AOI22_X1 U21747 ( .A1(n29317), .A2(\xmem_data[42][0] ), .B1(n29316), .B2(
        \xmem_data[43][0] ), .ZN(n17689) );
  AOI22_X1 U21748 ( .A1(n25717), .A2(\xmem_data[46][0] ), .B1(
        \xmem_data[47][0] ), .B2(n31361), .ZN(n17688) );
  AOI22_X1 U21749 ( .A1(n29319), .A2(\xmem_data[44][0] ), .B1(n29318), .B2(
        \xmem_data[45][0] ), .ZN(n17687) );
  NAND4_X1 U21750 ( .A1(n3912), .A2(n17692), .A3(n17691), .A4(n3511), .ZN(
        n17693) );
  AOI22_X1 U21751 ( .A1(n20770), .A2(\xmem_data[84][0] ), .B1(n29248), .B2(
        \xmem_data[85][0] ), .ZN(n17697) );
  AOI22_X1 U21752 ( .A1(n29257), .A2(\xmem_data[94][0] ), .B1(n31275), .B2(
        \xmem_data[95][0] ), .ZN(n17696) );
  AOI22_X1 U21753 ( .A1(n29256), .A2(\xmem_data[92][0] ), .B1(n29255), .B2(
        \xmem_data[93][0] ), .ZN(n17695) );
  NAND3_X1 U21754 ( .A1(n17697), .A2(n17696), .A3(n17695), .ZN(n17700) );
  AOI22_X1 U21755 ( .A1(n29124), .A2(\xmem_data[86][0] ), .B1(n27499), .B2(
        \xmem_data[87][0] ), .ZN(n17698) );
  INV_X1 U21756 ( .A(n17698), .ZN(n17699) );
  AOI22_X1 U21757 ( .A1(n29231), .A2(\xmem_data[64][0] ), .B1(n25514), .B2(
        \xmem_data[65][0] ), .ZN(n17704) );
  AOI22_X1 U21758 ( .A1(n27447), .A2(\xmem_data[66][0] ), .B1(n28373), .B2(
        \xmem_data[67][0] ), .ZN(n17703) );
  AOI22_X1 U21759 ( .A1(n20799), .A2(\xmem_data[68][0] ), .B1(n29232), .B2(
        \xmem_data[69][0] ), .ZN(n17702) );
  AOI22_X1 U21760 ( .A1(n3175), .A2(\xmem_data[70][0] ), .B1(n28517), .B2(
        \xmem_data[71][0] ), .ZN(n17701) );
  AOI22_X1 U21761 ( .A1(n27517), .A2(\xmem_data[72][0] ), .B1(n28299), .B2(
        \xmem_data[73][0] ), .ZN(n17708) );
  AOI22_X1 U21762 ( .A1(n24509), .A2(\xmem_data[74][0] ), .B1(n28058), .B2(
        \xmem_data[75][0] ), .ZN(n17707) );
  AOI22_X1 U21763 ( .A1(n29239), .A2(\xmem_data[76][0] ), .B1(n29238), .B2(
        \xmem_data[77][0] ), .ZN(n17706) );
  AOI22_X1 U21764 ( .A1(n29240), .A2(\xmem_data[78][0] ), .B1(n17001), .B2(
        \xmem_data[79][0] ), .ZN(n17705) );
  NAND4_X1 U21765 ( .A1(n17708), .A2(n17707), .A3(n17706), .A4(n17705), .ZN(
        n17713) );
  AOI22_X1 U21766 ( .A1(n28293), .A2(\xmem_data[82][0] ), .B1(n29247), .B2(
        \xmem_data[83][0] ), .ZN(n17711) );
  AOI22_X1 U21767 ( .A1(n29246), .A2(\xmem_data[80][0] ), .B1(n29245), .B2(
        \xmem_data[81][0] ), .ZN(n17710) );
  AOI22_X1 U21768 ( .A1(n22728), .A2(\xmem_data[88][0] ), .B1(n29253), .B2(
        \xmem_data[89][0] ), .ZN(n17709) );
  NOR2_X1 U21769 ( .A1(n17713), .A2(n17712), .ZN(n17715) );
  AOI22_X1 U21770 ( .A1(n29254), .A2(\xmem_data[90][0] ), .B1(n3218), .B2(
        \xmem_data[91][0] ), .ZN(n17714) );
  NAND3_X1 U21771 ( .A1(n3807), .A2(n17715), .A3(n17714), .ZN(n17716) );
  OAI21_X1 U21772 ( .B1(n17717), .B2(n17716), .A(n29267), .ZN(n17740) );
  AOI22_X1 U21773 ( .A1(n30295), .A2(\xmem_data[0][0] ), .B1(n15011), .B2(
        \xmem_data[1][0] ), .ZN(n17721) );
  AOI22_X1 U21774 ( .A1(n25422), .A2(\xmem_data[2][0] ), .B1(n28415), .B2(
        \xmem_data[3][0] ), .ZN(n17720) );
  AOI22_X1 U21775 ( .A1(n30886), .A2(\xmem_data[4][0] ), .B1(n28375), .B2(
        \xmem_data[5][0] ), .ZN(n17719) );
  AOI22_X1 U21776 ( .A1(n29272), .A2(\xmem_data[6][0] ), .B1(n29271), .B2(
        \xmem_data[7][0] ), .ZN(n17718) );
  NAND4_X1 U21777 ( .A1(n17721), .A2(n17720), .A3(n17719), .A4(n17718), .ZN(
        n17737) );
  AOI22_X1 U21778 ( .A1(n30746), .A2(\xmem_data[8][0] ), .B1(n29279), .B2(
        \xmem_data[9][0] ), .ZN(n17725) );
  AOI22_X1 U21779 ( .A1(n17020), .A2(\xmem_data[10][0] ), .B1(n29316), .B2(
        \xmem_data[11][0] ), .ZN(n17724) );
  AOI22_X1 U21780 ( .A1(n17021), .A2(\xmem_data[12][0] ), .B1(n29280), .B2(
        \xmem_data[13][0] ), .ZN(n17723) );
  AOI22_X1 U21781 ( .A1(n25575), .A2(\xmem_data[14][0] ), .B1(n27856), .B2(
        \xmem_data[15][0] ), .ZN(n17722) );
  NAND4_X1 U21782 ( .A1(n17725), .A2(n17724), .A3(n17723), .A4(n17722), .ZN(
        n17736) );
  AOI22_X1 U21783 ( .A1(n29297), .A2(\xmem_data[16][0] ), .B1(n14975), .B2(
        \xmem_data[17][0] ), .ZN(n17729) );
  AOI22_X1 U21784 ( .A1(n31316), .A2(\xmem_data[18][0] ), .B1(n27526), .B2(
        \xmem_data[19][0] ), .ZN(n17728) );
  AOI22_X1 U21785 ( .A1(n29298), .A2(\xmem_data[20][0] ), .B1(n30900), .B2(
        \xmem_data[21][0] ), .ZN(n17727) );
  AOI22_X1 U21786 ( .A1(n25686), .A2(\xmem_data[22][0] ), .B1(n22752), .B2(
        \xmem_data[23][0] ), .ZN(n17726) );
  NAND4_X1 U21787 ( .A1(n17729), .A2(n17728), .A3(n17727), .A4(n17726), .ZN(
        n17735) );
  AOI22_X1 U21788 ( .A1(n3335), .A2(\xmem_data[24][0] ), .B1(n29286), .B2(
        \xmem_data[25][0] ), .ZN(n17733) );
  AOI22_X1 U21789 ( .A1(n24532), .A2(\xmem_data[26][0] ), .B1(n3219), .B2(
        \xmem_data[27][0] ), .ZN(n17732) );
  AOI22_X1 U21790 ( .A1(n29288), .A2(\xmem_data[28][0] ), .B1(n30534), .B2(
        \xmem_data[29][0] ), .ZN(n17731) );
  AOI22_X1 U21791 ( .A1(n29289), .A2(\xmem_data[30][0] ), .B1(n27550), .B2(
        \xmem_data[31][0] ), .ZN(n17730) );
  NAND4_X1 U21792 ( .A1(n17733), .A2(n17732), .A3(n17731), .A4(n17730), .ZN(
        n17734) );
  OR4_X1 U21793 ( .A1(n17737), .A2(n17736), .A3(n17735), .A4(n17734), .ZN(
        n17738) );
  NAND2_X1 U21794 ( .A1(n17738), .A2(n25790), .ZN(n17739) );
  XNOR2_X1 U21795 ( .A(n34626), .B(\fmem_data[8][7] ), .ZN(n17744) );
  XOR2_X1 U21796 ( .A(\fmem_data[8][6] ), .B(\fmem_data[8][7] ), .Z(n17743) );
  XNOR2_X1 U21797 ( .A(n35258), .B(\fmem_data[23][1] ), .ZN(n32191) );
  INV_X1 U21798 ( .A(n17745), .ZN(n26802) );
  INV_X1 U21799 ( .A(n26797), .ZN(n17747) );
  NAND2_X1 U21800 ( .A1(n26794), .A2(n26795), .ZN(n17746) );
  OAI21_X1 U21801 ( .B1(n17748), .B2(n17747), .A(n17746), .ZN(n26266) );
  XNOR2_X1 U21802 ( .A(n17750), .B(n17749), .ZN(n17752) );
  XNOR2_X1 U21803 ( .A(n17752), .B(n17751), .ZN(n22155) );
  AOI22_X1 U21804 ( .A1(n28147), .A2(\xmem_data[20][1] ), .B1(n24460), .B2(
        \xmem_data[21][1] ), .ZN(n17760) );
  AOI22_X1 U21805 ( .A1(n30663), .A2(\xmem_data[12][1] ), .B1(n24448), .B2(
        \xmem_data[13][1] ), .ZN(n17759) );
  NAND2_X1 U21806 ( .A1(n27988), .A2(\xmem_data[11][1] ), .ZN(n17756) );
  NAND2_X1 U21807 ( .A1(n24458), .A2(\xmem_data[16][1] ), .ZN(n17755) );
  NAND2_X1 U21808 ( .A1(n17756), .A2(n17755), .ZN(n17757) );
  AOI21_X1 U21809 ( .B1(\xmem_data[15][1] ), .B2(n25606), .A(n17757), .ZN(
        n17758) );
  NAND3_X1 U21810 ( .A1(n17760), .A2(n17759), .A3(n17758), .ZN(n17771) );
  AOI22_X1 U21811 ( .A1(n3144), .A2(\xmem_data[0][1] ), .B1(n24439), .B2(
        \xmem_data[1][1] ), .ZN(n17764) );
  AOI22_X1 U21812 ( .A1(n24443), .A2(\xmem_data[2][1] ), .B1(n3221), .B2(
        \xmem_data[3][1] ), .ZN(n17763) );
  AOI22_X1 U21813 ( .A1(n30278), .A2(\xmem_data[4][1] ), .B1(n28508), .B2(
        \xmem_data[5][1] ), .ZN(n17762) );
  AOI22_X1 U21814 ( .A1(n24438), .A2(\xmem_data[6][1] ), .B1(n17061), .B2(
        \xmem_data[7][1] ), .ZN(n17761) );
  NAND4_X1 U21815 ( .A1(n17764), .A2(n17763), .A3(n17762), .A4(n17761), .ZN(
        n17770) );
  AOI22_X1 U21816 ( .A1(n3338), .A2(\xmem_data[24][1] ), .B1(n24521), .B2(
        \xmem_data[25][1] ), .ZN(n17768) );
  AOI22_X1 U21817 ( .A1(n24467), .A2(\xmem_data[26][1] ), .B1(n27981), .B2(
        \xmem_data[27][1] ), .ZN(n17767) );
  AOI22_X1 U21818 ( .A1(n20952), .A2(\xmem_data[28][1] ), .B1(n24468), .B2(
        \xmem_data[29][1] ), .ZN(n17766) );
  AOI22_X1 U21819 ( .A1(n30862), .A2(\xmem_data[30][1] ), .B1(n24470), .B2(
        \xmem_data[31][1] ), .ZN(n17765) );
  NAND4_X1 U21820 ( .A1(n17768), .A2(n17767), .A3(n17766), .A4(n17765), .ZN(
        n17769) );
  OR3_X1 U21821 ( .A1(n17771), .A2(n17770), .A3(n17769), .ZN(n17783) );
  AOI22_X1 U21822 ( .A1(n3178), .A2(\xmem_data[22][1] ), .B1(n25679), .B2(
        \xmem_data[23][1] ), .ZN(n17772) );
  INV_X1 U21823 ( .A(n17772), .ZN(n17779) );
  AOI22_X1 U21824 ( .A1(n24133), .A2(\xmem_data[18][1] ), .B1(n24459), .B2(
        \xmem_data[19][1] ), .ZN(n17773) );
  INV_X1 U21825 ( .A(n17773), .ZN(n17778) );
  NAND2_X1 U21826 ( .A1(n24450), .A2(\xmem_data[10][1] ), .ZN(n17776) );
  NAND2_X1 U21827 ( .A1(n25459), .A2(\xmem_data[14][1] ), .ZN(n17775) );
  NAND2_X1 U21828 ( .A1(n30698), .A2(\xmem_data[8][1] ), .ZN(n17774) );
  NAND3_X1 U21829 ( .A1(n17776), .A2(n17775), .A3(n17774), .ZN(n17777) );
  NOR3_X1 U21830 ( .A1(n17779), .A2(n17778), .A3(n17777), .ZN(n17781) );
  AOI21_X1 U21831 ( .B1(n25450), .B2(\xmem_data[9][1] ), .A(n17784), .ZN(
        n17850) );
  AOI22_X1 U21832 ( .A1(n20828), .A2(\xmem_data[96][1] ), .B1(n28501), .B2(
        \xmem_data[97][1] ), .ZN(n17788) );
  AOI22_X1 U21833 ( .A1(n24532), .A2(\xmem_data[98][1] ), .B1(n3222), .B2(
        \xmem_data[99][1] ), .ZN(n17787) );
  AOI22_X1 U21834 ( .A1(n24533), .A2(\xmem_data[100][1] ), .B1(n20787), .B2(
        \xmem_data[101][1] ), .ZN(n17786) );
  AOI22_X1 U21835 ( .A1(n24534), .A2(\xmem_data[102][1] ), .B1(n17061), .B2(
        \xmem_data[103][1] ), .ZN(n17785) );
  NAND4_X1 U21836 ( .A1(n17788), .A2(n17787), .A3(n17786), .A4(n17785), .ZN(
        n17804) );
  AOI22_X1 U21837 ( .A1(n29762), .A2(\xmem_data[104][1] ), .B1(n24657), .B2(
        \xmem_data[105][1] ), .ZN(n17792) );
  AOI22_X1 U21838 ( .A1(n27447), .A2(\xmem_data[106][1] ), .B1(n24130), .B2(
        \xmem_data[107][1] ), .ZN(n17791) );
  AOI22_X1 U21839 ( .A1(n20587), .A2(\xmem_data[108][1] ), .B1(n24516), .B2(
        \xmem_data[109][1] ), .ZN(n17790) );
  AOI22_X1 U21840 ( .A1(n28298), .A2(\xmem_data[110][1] ), .B1(n30541), .B2(
        \xmem_data[111][1] ), .ZN(n17789) );
  NAND4_X1 U21841 ( .A1(n17792), .A2(n17791), .A3(n17790), .A4(n17789), .ZN(
        n17803) );
  AOI22_X1 U21842 ( .A1(n23795), .A2(\xmem_data[112][1] ), .B1(n22742), .B2(
        \xmem_data[113][1] ), .ZN(n17796) );
  AOI22_X1 U21843 ( .A1(n24509), .A2(\xmem_data[114][1] ), .B1(n31355), .B2(
        \xmem_data[115][1] ), .ZN(n17795) );
  AOI22_X1 U21844 ( .A1(n21008), .A2(\xmem_data[116][1] ), .B1(n24510), .B2(
        \xmem_data[117][1] ), .ZN(n17794) );
  AOI22_X1 U21845 ( .A1(n24511), .A2(\xmem_data[118][1] ), .B1(n28429), .B2(
        \xmem_data[119][1] ), .ZN(n17793) );
  NAND4_X1 U21846 ( .A1(n17796), .A2(n17795), .A3(n17794), .A4(n17793), .ZN(
        n17802) );
  AOI22_X1 U21847 ( .A1(n24522), .A2(\xmem_data[120][1] ), .B1(n24521), .B2(
        \xmem_data[121][1] ), .ZN(n17800) );
  AOI22_X1 U21848 ( .A1(n3209), .A2(\xmem_data[122][1] ), .B1(n17003), .B2(
        \xmem_data[123][1] ), .ZN(n17799) );
  AOI22_X1 U21849 ( .A1(n20708), .A2(\xmem_data[124][1] ), .B1(n24524), .B2(
        \xmem_data[125][1] ), .ZN(n17798) );
  AOI22_X1 U21850 ( .A1(n24526), .A2(\xmem_data[126][1] ), .B1(n24525), .B2(
        \xmem_data[127][1] ), .ZN(n17797) );
  NAND4_X1 U21851 ( .A1(n17800), .A2(n17799), .A3(n17798), .A4(n17797), .ZN(
        n17801) );
  OR4_X1 U21852 ( .A1(n17804), .A2(n17803), .A3(n17802), .A4(n17801), .ZN(
        n17826) );
  AOI22_X1 U21853 ( .A1(n16980), .A2(\xmem_data[64][1] ), .B1(n3247), .B2(
        \xmem_data[65][1] ), .ZN(n17808) );
  AOI22_X1 U21854 ( .A1(n24532), .A2(\xmem_data[66][1] ), .B1(n3222), .B2(
        \xmem_data[67][1] ), .ZN(n17807) );
  AOI22_X1 U21855 ( .A1(n24533), .A2(\xmem_data[68][1] ), .B1(n27507), .B2(
        \xmem_data[69][1] ), .ZN(n17806) );
  AOI22_X1 U21856 ( .A1(n24534), .A2(\xmem_data[70][1] ), .B1(n21068), .B2(
        \xmem_data[71][1] ), .ZN(n17805) );
  NAND4_X1 U21857 ( .A1(n17808), .A2(n17807), .A3(n17806), .A4(n17805), .ZN(
        n17824) );
  AOI22_X1 U21858 ( .A1(n3345), .A2(\xmem_data[72][1] ), .B1(n30877), .B2(
        \xmem_data[73][1] ), .ZN(n17812) );
  AOI22_X1 U21859 ( .A1(n27447), .A2(\xmem_data[74][1] ), .B1(n20588), .B2(
        \xmem_data[75][1] ), .ZN(n17811) );
  AOI22_X1 U21860 ( .A1(n25457), .A2(\xmem_data[76][1] ), .B1(n24516), .B2(
        \xmem_data[77][1] ), .ZN(n17810) );
  AOI22_X1 U21861 ( .A1(n28334), .A2(\xmem_data[78][1] ), .B1(n30541), .B2(
        \xmem_data[79][1] ), .ZN(n17809) );
  NAND4_X1 U21862 ( .A1(n17812), .A2(n17811), .A3(n17810), .A4(n17809), .ZN(
        n17823) );
  AOI22_X1 U21863 ( .A1(n3466), .A2(\xmem_data[80][1] ), .B1(n15000), .B2(
        \xmem_data[81][1] ), .ZN(n17816) );
  AOI22_X1 U21864 ( .A1(n24509), .A2(\xmem_data[82][1] ), .B1(n20505), .B2(
        \xmem_data[83][1] ), .ZN(n17815) );
  AOI22_X1 U21865 ( .A1(n27855), .A2(\xmem_data[84][1] ), .B1(n24510), .B2(
        \xmem_data[85][1] ), .ZN(n17814) );
  AOI22_X1 U21866 ( .A1(n24511), .A2(\xmem_data[86][1] ), .B1(n30495), .B2(
        \xmem_data[87][1] ), .ZN(n17813) );
  NAND4_X1 U21867 ( .A1(n17816), .A2(n17815), .A3(n17814), .A4(n17813), .ZN(
        n17822) );
  AOI22_X1 U21868 ( .A1(n24522), .A2(\xmem_data[88][1] ), .B1(n24521), .B2(
        \xmem_data[89][1] ), .ZN(n17820) );
  AOI22_X1 U21869 ( .A1(n3209), .A2(\xmem_data[90][1] ), .B1(n25406), .B2(
        \xmem_data[91][1] ), .ZN(n17819) );
  AOI22_X1 U21870 ( .A1(n25407), .A2(\xmem_data[92][1] ), .B1(n24524), .B2(
        \xmem_data[93][1] ), .ZN(n17818) );
  AOI22_X1 U21871 ( .A1(n24526), .A2(\xmem_data[94][1] ), .B1(n24525), .B2(
        \xmem_data[95][1] ), .ZN(n17817) );
  NAND4_X1 U21872 ( .A1(n17820), .A2(n17819), .A3(n17818), .A4(n17817), .ZN(
        n17821) );
  OR4_X1 U21873 ( .A1(n17824), .A2(n17823), .A3(n17822), .A4(n17821), .ZN(
        n17825) );
  AOI22_X1 U21874 ( .A1(n24542), .A2(n17826), .B1(n24581), .B2(n17825), .ZN(
        n17849) );
  AOI22_X1 U21875 ( .A1(n3433), .A2(\xmem_data[32][1] ), .B1(n30589), .B2(
        \xmem_data[33][1] ), .ZN(n17830) );
  AOI22_X1 U21876 ( .A1(n24562), .A2(\xmem_data[34][1] ), .B1(n3219), .B2(
        \xmem_data[35][1] ), .ZN(n17829) );
  AOI22_X1 U21877 ( .A1(n24563), .A2(\xmem_data[36][1] ), .B1(n20787), .B2(
        \xmem_data[37][1] ), .ZN(n17828) );
  AOI22_X1 U21878 ( .A1(n24565), .A2(\xmem_data[38][1] ), .B1(n24564), .B2(
        \xmem_data[39][1] ), .ZN(n17827) );
  NAND4_X1 U21879 ( .A1(n17830), .A2(n17829), .A3(n17828), .A4(n17827), .ZN(
        n17846) );
  AOI22_X1 U21880 ( .A1(n25377), .A2(\xmem_data[40][1] ), .B1(n24553), .B2(
        \xmem_data[41][1] ), .ZN(n17834) );
  AOI22_X1 U21881 ( .A1(n24554), .A2(\xmem_data[42][1] ), .B1(n27863), .B2(
        \xmem_data[43][1] ), .ZN(n17833) );
  AOI22_X1 U21882 ( .A1(n24556), .A2(\xmem_data[44][1] ), .B1(n24555), .B2(
        \xmem_data[45][1] ), .ZN(n17832) );
  AOI22_X1 U21883 ( .A1(n28298), .A2(\xmem_data[46][1] ), .B1(n24597), .B2(
        \xmem_data[47][1] ), .ZN(n17831) );
  NAND4_X1 U21884 ( .A1(n17834), .A2(n17833), .A3(n17832), .A4(n17831), .ZN(
        n17845) );
  AOI22_X1 U21885 ( .A1(n24545), .A2(\xmem_data[48][1] ), .B1(n27454), .B2(
        \xmem_data[49][1] ), .ZN(n17838) );
  AOI22_X1 U21886 ( .A1(n24547), .A2(\xmem_data[50][1] ), .B1(n24546), .B2(
        \xmem_data[51][1] ), .ZN(n17837) );
  AOI22_X1 U21887 ( .A1(n21050), .A2(\xmem_data[52][1] ), .B1(n29238), .B2(
        \xmem_data[53][1] ), .ZN(n17836) );
  AOI22_X1 U21888 ( .A1(n30899), .A2(\xmem_data[54][1] ), .B1(n25581), .B2(
        \xmem_data[55][1] ), .ZN(n17835) );
  NAND4_X1 U21889 ( .A1(n17838), .A2(n17837), .A3(n17836), .A4(n17835), .ZN(
        n17844) );
  AOI22_X1 U21890 ( .A1(n24571), .A2(\xmem_data[56][1] ), .B1(n24570), .B2(
        \xmem_data[57][1] ), .ZN(n17842) );
  AOI22_X1 U21891 ( .A1(n24572), .A2(\xmem_data[58][1] ), .B1(n28500), .B2(
        \xmem_data[59][1] ), .ZN(n17841) );
  AOI22_X1 U21892 ( .A1(n31308), .A2(\xmem_data[60][1] ), .B1(n29248), .B2(
        \xmem_data[61][1] ), .ZN(n17840) );
  AOI22_X1 U21893 ( .A1(n30862), .A2(\xmem_data[62][1] ), .B1(n24573), .B2(
        \xmem_data[63][1] ), .ZN(n17839) );
  NAND4_X1 U21894 ( .A1(n17842), .A2(n17841), .A3(n17840), .A4(n17839), .ZN(
        n17843) );
  OR4_X1 U21895 ( .A1(n17846), .A2(n17845), .A3(n17844), .A4(n17843), .ZN(
        n17847) );
  NAND2_X1 U21896 ( .A1(n17847), .A2(n24508), .ZN(n17848) );
  AOI22_X1 U21897 ( .A1(n28468), .A2(\xmem_data[96][6] ), .B1(n20567), .B2(
        \xmem_data[97][6] ), .ZN(n17855) );
  AOI22_X1 U21898 ( .A1(n30524), .A2(\xmem_data[98][6] ), .B1(n27564), .B2(
        \xmem_data[99][6] ), .ZN(n17854) );
  AOI22_X1 U21899 ( .A1(n20578), .A2(\xmem_data[100][6] ), .B1(n24630), .B2(
        \xmem_data[101][6] ), .ZN(n17853) );
  AOI22_X1 U21900 ( .A1(n20568), .A2(\xmem_data[102][6] ), .B1(n28082), .B2(
        \xmem_data[103][6] ), .ZN(n17852) );
  NAND4_X1 U21901 ( .A1(n17855), .A2(n17854), .A3(n17853), .A4(n17852), .ZN(
        n17871) );
  AOI22_X1 U21902 ( .A1(n3218), .A2(\xmem_data[104][6] ), .B1(n29256), .B2(
        \xmem_data[105][6] ), .ZN(n17859) );
  AOI22_X1 U21903 ( .A1(n20558), .A2(\xmem_data[106][6] ), .B1(n24565), .B2(
        \xmem_data[107][6] ), .ZN(n17858) );
  AOI22_X1 U21904 ( .A1(n20559), .A2(\xmem_data[108][6] ), .B1(n3128), .B2(
        \xmem_data[109][6] ), .ZN(n17857) );
  AOI22_X1 U21905 ( .A1(n28343), .A2(\xmem_data[110][6] ), .B1(n25707), .B2(
        \xmem_data[111][6] ), .ZN(n17856) );
  NAND4_X1 U21906 ( .A1(n17859), .A2(n17858), .A3(n17857), .A4(n17856), .ZN(
        n17870) );
  AOI22_X1 U21907 ( .A1(n20546), .A2(\xmem_data[112][6] ), .B1(n20545), .B2(
        \xmem_data[113][6] ), .ZN(n17863) );
  AOI22_X1 U21908 ( .A1(n28345), .A2(\xmem_data[114][6] ), .B1(n30891), .B2(
        \xmem_data[115][6] ), .ZN(n17862) );
  AOI22_X1 U21909 ( .A1(n20544), .A2(\xmem_data[116][6] ), .B1(n21005), .B2(
        \xmem_data[117][6] ), .ZN(n17861) );
  AOI22_X1 U21910 ( .A1(n20543), .A2(\xmem_data[118][6] ), .B1(n20542), .B2(
        \xmem_data[119][6] ), .ZN(n17860) );
  NAND4_X1 U21911 ( .A1(n17863), .A2(n17862), .A3(n17861), .A4(n17860), .ZN(
        n17869) );
  AOI22_X1 U21912 ( .A1(n14970), .A2(\xmem_data[120][6] ), .B1(n20942), .B2(
        \xmem_data[121][6] ), .ZN(n17867) );
  AOI22_X1 U21913 ( .A1(n29318), .A2(\xmem_data[122][6] ), .B1(n28428), .B2(
        \xmem_data[123][6] ), .ZN(n17866) );
  AOI22_X1 U21914 ( .A1(n20551), .A2(\xmem_data[124][6] ), .B1(n29246), .B2(
        \xmem_data[125][6] ), .ZN(n17865) );
  AOI22_X1 U21915 ( .A1(n20553), .A2(\xmem_data[126][6] ), .B1(n20552), .B2(
        \xmem_data[127][6] ), .ZN(n17864) );
  NAND4_X1 U21916 ( .A1(n17867), .A2(n17866), .A3(n17865), .A4(n17864), .ZN(
        n17868) );
  OR4_X1 U21917 ( .A1(n17871), .A2(n17870), .A3(n17869), .A4(n17868), .ZN(
        n17895) );
  AND2_X1 U21918 ( .A1(n17003), .A2(\xmem_data[64][6] ), .ZN(n17872) );
  AOI21_X1 U21919 ( .B1(n20577), .B2(\xmem_data[65][6] ), .A(n17872), .ZN(
        n17877) );
  AOI22_X1 U21920 ( .A1(n20579), .A2(\xmem_data[66][6] ), .B1(n27925), .B2(
        \xmem_data[67][6] ), .ZN(n17876) );
  AOI22_X1 U21921 ( .A1(n20578), .A2(\xmem_data[68][6] ), .B1(n30864), .B2(
        \xmem_data[69][6] ), .ZN(n17875) );
  AND2_X1 U21922 ( .A1(n28501), .A2(\xmem_data[70][6] ), .ZN(n17873) );
  AOI21_X1 U21923 ( .B1(n20518), .B2(\xmem_data[71][6] ), .A(n17873), .ZN(
        n17874) );
  NAND4_X1 U21924 ( .A1(n17877), .A2(n17876), .A3(n17875), .A4(n17874), .ZN(
        n17893) );
  AOI22_X1 U21925 ( .A1(n20588), .A2(\xmem_data[80][6] ), .B1(n20587), .B2(
        \xmem_data[81][6] ), .ZN(n17881) );
  AOI22_X1 U21926 ( .A1(n31326), .A2(\xmem_data[82][6] ), .B1(n29272), .B2(
        \xmem_data[83][6] ), .ZN(n17880) );
  AOI22_X1 U21927 ( .A1(n20584), .A2(\xmem_data[84][6] ), .B1(n27818), .B2(
        \xmem_data[85][6] ), .ZN(n17879) );
  AOI22_X1 U21928 ( .A1(n20586), .A2(\xmem_data[86][6] ), .B1(n20585), .B2(
        \xmem_data[87][6] ), .ZN(n17878) );
  NAND4_X1 U21929 ( .A1(n17881), .A2(n17880), .A3(n17879), .A4(n17878), .ZN(
        n17892) );
  AOI22_X1 U21930 ( .A1(n21006), .A2(\xmem_data[88][6] ), .B1(n30617), .B2(
        \xmem_data[89][6] ), .ZN(n17885) );
  AOI22_X1 U21931 ( .A1(n21049), .A2(\xmem_data[90][6] ), .B1(n24220), .B2(
        \xmem_data[91][6] ), .ZN(n17884) );
  AOI22_X1 U21932 ( .A1(n27856), .A2(\xmem_data[92][6] ), .B1(n28955), .B2(
        \xmem_data[93][6] ), .ZN(n17883) );
  AOI22_X1 U21933 ( .A1(n14975), .A2(\xmem_data[94][6] ), .B1(n24166), .B2(
        \xmem_data[95][6] ), .ZN(n17882) );
  NAND4_X1 U21934 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        n17891) );
  AOI22_X1 U21935 ( .A1(n3222), .A2(\xmem_data[72][6] ), .B1(n29026), .B2(
        \xmem_data[73][6] ), .ZN(n17889) );
  AOI22_X1 U21936 ( .A1(n20598), .A2(\xmem_data[74][6] ), .B1(n29289), .B2(
        \xmem_data[75][6] ), .ZN(n17888) );
  AOI22_X1 U21937 ( .A1(n24140), .A2(\xmem_data[76][6] ), .B1(n17063), .B2(
        \xmem_data[77][6] ), .ZN(n17887) );
  AOI22_X1 U21938 ( .A1(n29103), .A2(\xmem_data[78][6] ), .B1(n24450), .B2(
        \xmem_data[79][6] ), .ZN(n17886) );
  NAND4_X1 U21939 ( .A1(n17889), .A2(n17888), .A3(n17887), .A4(n17886), .ZN(
        n17890) );
  AOI22_X1 U21940 ( .A1(n20538), .A2(n17895), .B1(n20573), .B2(n17894), .ZN(
        n17944) );
  AOI22_X1 U21941 ( .A1(n20488), .A2(\xmem_data[0][6] ), .B1(n21060), .B2(
        \xmem_data[1][6] ), .ZN(n17900) );
  AOI22_X1 U21942 ( .A1(n25440), .A2(\xmem_data[2][6] ), .B1(n25441), .B2(
        \xmem_data[3][6] ), .ZN(n17899) );
  AOI22_X1 U21943 ( .A1(n20489), .A2(\xmem_data[4][6] ), .B1(n3144), .B2(
        \xmem_data[5][6] ), .ZN(n17898) );
  AND2_X1 U21944 ( .A1(n23731), .A2(\xmem_data[6][6] ), .ZN(n17896) );
  AOI21_X1 U21945 ( .B1(n24443), .B2(\xmem_data[7][6] ), .A(n17896), .ZN(
        n17897) );
  NAND4_X1 U21946 ( .A1(n17900), .A2(n17899), .A3(n17898), .A4(n17897), .ZN(
        n17920) );
  AOI22_X1 U21947 ( .A1(n27863), .A2(\xmem_data[16][6] ), .B1(n20716), .B2(
        \xmem_data[17][6] ), .ZN(n17904) );
  AOI22_X1 U21948 ( .A1(n24639), .A2(\xmem_data[18][6] ), .B1(n24131), .B2(
        \xmem_data[19][6] ), .ZN(n17903) );
  AOI22_X1 U21949 ( .A1(n25606), .A2(\xmem_data[20][6] ), .B1(n29237), .B2(
        \xmem_data[21][6] ), .ZN(n17902) );
  AOI22_X1 U21950 ( .A1(n30542), .A2(\xmem_data[22][6] ), .B1(n24593), .B2(
        \xmem_data[23][6] ), .ZN(n17901) );
  NAND4_X1 U21951 ( .A1(n17904), .A2(n17903), .A3(n17902), .A4(n17901), .ZN(
        n17910) );
  AOI22_X1 U21952 ( .A1(n20505), .A2(\xmem_data[24][6] ), .B1(n28994), .B2(
        \xmem_data[25][6] ), .ZN(n17908) );
  AOI22_X1 U21953 ( .A1(n13481), .A2(\xmem_data[26][6] ), .B1(n28428), .B2(
        \xmem_data[27][6] ), .ZN(n17907) );
  AOI22_X1 U21954 ( .A1(n28429), .A2(\xmem_data[28][6] ), .B1(n25636), .B2(
        \xmem_data[29][6] ), .ZN(n17906) );
  AOI22_X1 U21955 ( .A1(n20507), .A2(\xmem_data[30][6] ), .B1(n29151), .B2(
        \xmem_data[31][6] ), .ZN(n17905) );
  NAND4_X1 U21956 ( .A1(n17908), .A2(n17907), .A3(n17906), .A4(n17905), .ZN(
        n17909) );
  OR3_X1 U21957 ( .A1(n17910), .A2(n17909), .A3(n3974), .ZN(n17919) );
  AOI22_X1 U21958 ( .A1(n13444), .A2(\xmem_data[12][6] ), .B1(n22668), .B2(
        \xmem_data[13][6] ), .ZN(n17917) );
  AOI22_X1 U21959 ( .A1(n3222), .A2(\xmem_data[8][6] ), .B1(n24563), .B2(
        \xmem_data[9][6] ), .ZN(n17911) );
  INV_X1 U21960 ( .A(n17911), .ZN(n17915) );
  AOI22_X1 U21961 ( .A1(n20500), .A2(\xmem_data[10][6] ), .B1(n24697), .B2(
        \xmem_data[11][6] ), .ZN(n17912) );
  INV_X1 U21962 ( .A(n17912), .ZN(n17914) );
  AND2_X1 U21963 ( .A1(n24450), .A2(\xmem_data[15][6] ), .ZN(n17913) );
  NOR3_X1 U21964 ( .A1(n17915), .A2(n17914), .A3(n17913), .ZN(n17916) );
  NAND2_X1 U21965 ( .A1(n17917), .A2(n17916), .ZN(n17918) );
  OAI21_X1 U21966 ( .B1(n17920), .B2(n4003), .A(n20515), .ZN(n17943) );
  AOI22_X1 U21967 ( .A1(n17003), .A2(\xmem_data[32][6] ), .B1(n20577), .B2(
        \xmem_data[33][6] ), .ZN(n17924) );
  AOI22_X1 U21968 ( .A1(n20579), .A2(\xmem_data[34][6] ), .B1(n27500), .B2(
        \xmem_data[35][6] ), .ZN(n17923) );
  AOI22_X1 U21969 ( .A1(n20578), .A2(\xmem_data[36][6] ), .B1(n3433), .B2(
        \xmem_data[37][6] ), .ZN(n17922) );
  AOI22_X1 U21970 ( .A1(n27437), .A2(\xmem_data[38][6] ), .B1(n20518), .B2(
        \xmem_data[39][6] ), .ZN(n17921) );
  NAND4_X1 U21971 ( .A1(n17924), .A2(n17923), .A3(n17922), .A4(n17921), .ZN(
        n17940) );
  AOI22_X1 U21972 ( .A1(n3222), .A2(\xmem_data[40][6] ), .B1(n28137), .B2(
        \xmem_data[41][6] ), .ZN(n17928) );
  AOI22_X1 U21973 ( .A1(n20598), .A2(\xmem_data[42][6] ), .B1(n3341), .B2(
        \xmem_data[43][6] ), .ZN(n17927) );
  AOI22_X1 U21974 ( .A1(n20806), .A2(\xmem_data[44][6] ), .B1(n3134), .B2(
        \xmem_data[45][6] ), .ZN(n17926) );
  AOI22_X1 U21975 ( .A1(n31252), .A2(\xmem_data[46][6] ), .B1(n16974), .B2(
        \xmem_data[47][6] ), .ZN(n17925) );
  NAND4_X1 U21976 ( .A1(n17928), .A2(n17927), .A3(n17926), .A4(n17925), .ZN(
        n17939) );
  AOI22_X1 U21977 ( .A1(n20588), .A2(\xmem_data[48][6] ), .B1(n20587), .B2(
        \xmem_data[49][6] ), .ZN(n17932) );
  AOI22_X1 U21978 ( .A1(n24448), .A2(\xmem_data[50][6] ), .B1(n31268), .B2(
        \xmem_data[51][6] ), .ZN(n17931) );
  AOI22_X1 U21979 ( .A1(n20584), .A2(\xmem_data[52][6] ), .B1(n29237), .B2(
        \xmem_data[53][6] ), .ZN(n17930) );
  AOI22_X1 U21980 ( .A1(n20586), .A2(\xmem_data[54][6] ), .B1(n20585), .B2(
        \xmem_data[55][6] ), .ZN(n17929) );
  NAND4_X1 U21981 ( .A1(n17932), .A2(n17931), .A3(n17930), .A4(n17929), .ZN(
        n17938) );
  AOI22_X1 U21982 ( .A1(n25520), .A2(\xmem_data[56][6] ), .B1(n25678), .B2(
        \xmem_data[57][6] ), .ZN(n17936) );
  AOI22_X1 U21983 ( .A1(n20941), .A2(\xmem_data[58][6] ), .B1(n28460), .B2(
        \xmem_data[59][6] ), .ZN(n17935) );
  AOI22_X1 U21984 ( .A1(n27461), .A2(\xmem_data[60][6] ), .B1(n20984), .B2(
        \xmem_data[61][6] ), .ZN(n17934) );
  AOI22_X1 U21985 ( .A1(n24570), .A2(\xmem_data[62][6] ), .B1(n3209), .B2(
        \xmem_data[63][6] ), .ZN(n17933) );
  NAND4_X1 U21986 ( .A1(n17936), .A2(n17935), .A3(n17934), .A4(n17933), .ZN(
        n17937) );
  OR4_X1 U21987 ( .A1(n17940), .A2(n17939), .A3(n17938), .A4(n17937), .ZN(
        n17941) );
  NAND2_X1 U21988 ( .A1(n17941), .A2(n20606), .ZN(n17942) );
  XNOR2_X1 U21989 ( .A(n31660), .B(\fmem_data[21][1] ), .ZN(n31883) );
  OAI22_X1 U21990 ( .A1(n31883), .A2(n34613), .B1(n3570), .B2(n31943), .ZN(
        n22782) );
  AOI22_X1 U21991 ( .A1(n3217), .A2(\xmem_data[32][3] ), .B1(n31368), .B2(
        \xmem_data[33][3] ), .ZN(n17948) );
  AOI22_X1 U21992 ( .A1(n24207), .A2(\xmem_data[34][3] ), .B1(n27904), .B2(
        \xmem_data[35][3] ), .ZN(n17947) );
  AOI22_X1 U21993 ( .A1(n31275), .A2(\xmem_data[36][3] ), .B1(n20808), .B2(
        \xmem_data[37][3] ), .ZN(n17946) );
  AOI22_X1 U21994 ( .A1(n28045), .A2(\xmem_data[38][3] ), .B1(n25604), .B2(
        \xmem_data[39][3] ), .ZN(n17945) );
  NAND4_X1 U21995 ( .A1(n17948), .A2(n17947), .A3(n17946), .A4(n17945), .ZN(
        n17965) );
  AOI22_X1 U21996 ( .A1(n20546), .A2(\xmem_data[40][3] ), .B1(n29451), .B2(
        \xmem_data[41][3] ), .ZN(n17952) );
  AOI22_X1 U21997 ( .A1(n24212), .A2(\xmem_data[42][3] ), .B1(n24131), .B2(
        \xmem_data[43][3] ), .ZN(n17951) );
  AOI22_X1 U21998 ( .A1(n28517), .A2(\xmem_data[44][3] ), .B1(n29396), .B2(
        \xmem_data[45][3] ), .ZN(n17950) );
  AOI22_X1 U21999 ( .A1(n29188), .A2(\xmem_data[46][3] ), .B1(n24214), .B2(
        \xmem_data[47][3] ), .ZN(n17949) );
  NAND4_X1 U22000 ( .A1(n17952), .A2(n17951), .A3(n17950), .A4(n17949), .ZN(
        n17964) );
  AOI22_X1 U22001 ( .A1(n24219), .A2(\xmem_data[48][3] ), .B1(n14971), .B2(
        \xmem_data[49][3] ), .ZN(n17956) );
  AOI22_X1 U22002 ( .A1(n24221), .A2(\xmem_data[50][3] ), .B1(n28460), .B2(
        \xmem_data[51][3] ), .ZN(n17955) );
  AOI22_X1 U22003 ( .A1(n24222), .A2(\xmem_data[52][3] ), .B1(n28202), .B2(
        \xmem_data[53][3] ), .ZN(n17954) );
  AOI22_X1 U22004 ( .A1(n24223), .A2(\xmem_data[54][3] ), .B1(n29325), .B2(
        \xmem_data[55][3] ), .ZN(n17953) );
  NAND4_X1 U22005 ( .A1(n17956), .A2(n17955), .A3(n17954), .A4(n17953), .ZN(
        n17963) );
  AOI22_X1 U22006 ( .A1(n17003), .A2(\xmem_data[56][3] ), .B1(n27568), .B2(
        \xmem_data[57][3] ), .ZN(n17961) );
  AOI22_X1 U22007 ( .A1(n20769), .A2(\xmem_data[58][3] ), .B1(n24607), .B2(
        \xmem_data[59][3] ), .ZN(n17960) );
  AOI22_X1 U22008 ( .A1(n3203), .A2(\xmem_data[60][3] ), .B1(n3333), .B2(
        \xmem_data[61][3] ), .ZN(n17959) );
  AND2_X1 U22009 ( .A1(n24439), .A2(\xmem_data[62][3] ), .ZN(n17957) );
  AOI21_X1 U22010 ( .B1(n28470), .B2(\xmem_data[63][3] ), .A(n17957), .ZN(
        n17958) );
  NAND4_X1 U22011 ( .A1(n17961), .A2(n17960), .A3(n17959), .A4(n17958), .ZN(
        n17962) );
  OR4_X1 U22012 ( .A1(n17965), .A2(n17964), .A3(n17963), .A4(n17962), .ZN(
        n17967) );
  NOR2_X1 U22013 ( .A1(n24151), .A2(n39012), .ZN(n17966) );
  AOI21_X1 U22014 ( .B1(n17967), .B2(n24236), .A(n3888), .ZN(n18042) );
  AOI22_X1 U22015 ( .A1(n3221), .A2(\xmem_data[96][3] ), .B1(n20805), .B2(
        \xmem_data[97][3] ), .ZN(n17971) );
  AOI22_X1 U22016 ( .A1(n30534), .A2(\xmem_data[98][3] ), .B1(n30883), .B2(
        \xmem_data[99][3] ), .ZN(n17970) );
  AOI22_X1 U22017 ( .A1(n29104), .A2(\xmem_data[100][3] ), .B1(n3375), .B2(
        \xmem_data[101][3] ), .ZN(n17969) );
  AOI22_X1 U22018 ( .A1(n25450), .A2(\xmem_data[102][3] ), .B1(n28374), .B2(
        \xmem_data[103][3] ), .ZN(n17968) );
  NAND4_X1 U22019 ( .A1(n17971), .A2(n17970), .A3(n17969), .A4(n17968), .ZN(
        n17988) );
  AOI22_X1 U22020 ( .A1(n24158), .A2(\xmem_data[104][3] ), .B1(n24157), .B2(
        \xmem_data[105][3] ), .ZN(n17975) );
  AOI22_X1 U22021 ( .A1(n24159), .A2(\xmem_data[106][3] ), .B1(n30514), .B2(
        \xmem_data[107][3] ), .ZN(n17974) );
  AOI22_X1 U22022 ( .A1(n24160), .A2(\xmem_data[108][3] ), .B1(n3158), .B2(
        \xmem_data[109][3] ), .ZN(n17973) );
  AOI22_X1 U22023 ( .A1(n27516), .A2(\xmem_data[110][3] ), .B1(n24214), .B2(
        \xmem_data[111][3] ), .ZN(n17972) );
  NAND4_X1 U22024 ( .A1(n17975), .A2(n17974), .A3(n17973), .A4(n17972), .ZN(
        n17987) );
  AOI22_X1 U22025 ( .A1(n24459), .A2(\xmem_data[112][3] ), .B1(n17021), .B2(
        \xmem_data[113][3] ), .ZN(n17979) );
  AOI22_X1 U22026 ( .A1(n24165), .A2(\xmem_data[114][3] ), .B1(n30557), .B2(
        \xmem_data[115][3] ), .ZN(n17978) );
  AOI22_X1 U22027 ( .A1(n29281), .A2(\xmem_data[116][3] ), .B1(n3307), .B2(
        \xmem_data[117][3] ), .ZN(n17977) );
  AOI22_X1 U22028 ( .A1(n24167), .A2(\xmem_data[118][3] ), .B1(n24166), .B2(
        \xmem_data[119][3] ), .ZN(n17976) );
  NAND4_X1 U22029 ( .A1(n17979), .A2(n17978), .A3(n17977), .A4(n17976), .ZN(
        n17986) );
  AOI22_X1 U22030 ( .A1(n27981), .A2(\xmem_data[120][3] ), .B1(n29298), .B2(
        \xmem_data[121][3] ), .ZN(n17984) );
  AOI22_X1 U22031 ( .A1(n31344), .A2(\xmem_data[122][3] ), .B1(n27925), .B2(
        \xmem_data[123][3] ), .ZN(n17983) );
  AOI22_X1 U22032 ( .A1(n21309), .A2(\xmem_data[124][3] ), .B1(n25725), .B2(
        \xmem_data[125][3] ), .ZN(n17982) );
  AND2_X1 U22033 ( .A1(n24172), .A2(\xmem_data[126][3] ), .ZN(n17980) );
  AOI21_X1 U22034 ( .B1(n24562), .B2(\xmem_data[127][3] ), .A(n17980), .ZN(
        n17981) );
  NAND4_X1 U22035 ( .A1(n17984), .A2(n17983), .A3(n17982), .A4(n17981), .ZN(
        n17985) );
  OR4_X1 U22036 ( .A1(n17988), .A2(n17987), .A3(n17986), .A4(n17985), .ZN(
        n18011) );
  AOI22_X1 U22037 ( .A1(n3221), .A2(\xmem_data[64][3] ), .B1(n29431), .B2(
        \xmem_data[65][3] ), .ZN(n17992) );
  AOI22_X1 U22038 ( .A1(n24695), .A2(\xmem_data[66][3] ), .B1(n20994), .B2(
        \xmem_data[67][3] ), .ZN(n17991) );
  AOI22_X1 U22039 ( .A1(n22669), .A2(\xmem_data[68][3] ), .B1(n25451), .B2(
        \xmem_data[69][3] ), .ZN(n17990) );
  AOI22_X1 U22040 ( .A1(n29045), .A2(\xmem_data[70][3] ), .B1(n28374), .B2(
        \xmem_data[71][3] ), .ZN(n17989) );
  NAND4_X1 U22041 ( .A1(n17992), .A2(n17991), .A3(n17990), .A4(n17989), .ZN(
        n18009) );
  AOI22_X1 U22042 ( .A1(n24158), .A2(\xmem_data[72][3] ), .B1(n24157), .B2(
        \xmem_data[73][3] ), .ZN(n17996) );
  AOI22_X1 U22043 ( .A1(n24159), .A2(\xmem_data[74][3] ), .B1(n30514), .B2(
        \xmem_data[75][3] ), .ZN(n17995) );
  AOI22_X1 U22044 ( .A1(n24160), .A2(\xmem_data[76][3] ), .B1(n17018), .B2(
        \xmem_data[77][3] ), .ZN(n17994) );
  AOI22_X1 U22045 ( .A1(n15000), .A2(\xmem_data[78][3] ), .B1(n21007), .B2(
        \xmem_data[79][3] ), .ZN(n17993) );
  NAND4_X1 U22046 ( .A1(n17996), .A2(n17995), .A3(n17994), .A4(n17993), .ZN(
        n18008) );
  AOI22_X1 U22047 ( .A1(n31270), .A2(\xmem_data[80][3] ), .B1(n22717), .B2(
        \xmem_data[81][3] ), .ZN(n18000) );
  AOI22_X1 U22048 ( .A1(n24165), .A2(\xmem_data[82][3] ), .B1(n25717), .B2(
        \xmem_data[83][3] ), .ZN(n17999) );
  AOI22_X1 U22049 ( .A1(n28327), .A2(\xmem_data[84][3] ), .B1(n30600), .B2(
        \xmem_data[85][3] ), .ZN(n17998) );
  AOI22_X1 U22050 ( .A1(n24167), .A2(\xmem_data[86][3] ), .B1(n24166), .B2(
        \xmem_data[87][3] ), .ZN(n17997) );
  NAND4_X1 U22051 ( .A1(n18000), .A2(n17999), .A3(n17998), .A4(n17997), .ZN(
        n18007) );
  AOI22_X1 U22052 ( .A1(n17049), .A2(\xmem_data[88][3] ), .B1(n25628), .B2(
        \xmem_data[89][3] ), .ZN(n18005) );
  AOI22_X1 U22053 ( .A1(n30524), .A2(\xmem_data[90][3] ), .B1(n25686), .B2(
        \xmem_data[91][3] ), .ZN(n18004) );
  AOI22_X1 U22054 ( .A1(n29118), .A2(\xmem_data[92][3] ), .B1(n3384), .B2(
        \xmem_data[93][3] ), .ZN(n18003) );
  AND2_X1 U22055 ( .A1(n24172), .A2(\xmem_data[94][3] ), .ZN(n18001) );
  AOI21_X1 U22056 ( .B1(n25730), .B2(\xmem_data[95][3] ), .A(n18001), .ZN(
        n18002) );
  NAND4_X1 U22057 ( .A1(n18005), .A2(n18004), .A3(n18003), .A4(n18002), .ZN(
        n18006) );
  OR4_X1 U22058 ( .A1(n18009), .A2(n18008), .A3(n18007), .A4(n18006), .ZN(
        n18010) );
  AOI22_X1 U22059 ( .A1(n24205), .A2(n18011), .B1(n24204), .B2(n18010), .ZN(
        n18041) );
  AOI22_X1 U22060 ( .A1(n3219), .A2(\xmem_data[0][3] ), .B1(n24139), .B2(
        \xmem_data[1][3] ), .ZN(n18018) );
  AOI22_X1 U22061 ( .A1(n24140), .A2(\xmem_data[4][3] ), .B1(n3282), .B2(
        \xmem_data[5][3] ), .ZN(n18012) );
  INV_X1 U22062 ( .A(n18012), .ZN(n18016) );
  AOI22_X1 U22063 ( .A1(n27869), .A2(\xmem_data[2][3] ), .B1(n24141), .B2(
        \xmem_data[3][3] ), .ZN(n18014) );
  NAND2_X1 U22064 ( .A1(n23813), .A2(\xmem_data[7][3] ), .ZN(n18013) );
  NAND2_X1 U22065 ( .A1(n18014), .A2(n18013), .ZN(n18015) );
  NOR2_X1 U22066 ( .A1(n18016), .A2(n18015), .ZN(n18017) );
  NAND2_X1 U22067 ( .A1(n18018), .A2(n18017), .ZN(n18024) );
  AOI22_X1 U22068 ( .A1(n24130), .A2(\xmem_data[8][3] ), .B1(n30943), .B2(
        \xmem_data[9][3] ), .ZN(n18022) );
  AOI22_X1 U22069 ( .A1(n24132), .A2(\xmem_data[10][3] ), .B1(n20495), .B2(
        \xmem_data[11][3] ), .ZN(n18021) );
  AOI22_X1 U22070 ( .A1(n25606), .A2(\xmem_data[12][3] ), .B1(n3157), .B2(
        \xmem_data[13][3] ), .ZN(n18020) );
  AOI22_X1 U22071 ( .A1(n24134), .A2(\xmem_data[14][3] ), .B1(n24133), .B2(
        \xmem_data[15][3] ), .ZN(n18019) );
  NAND4_X1 U22072 ( .A1(n18022), .A2(n18021), .A3(n18020), .A4(n18019), .ZN(
        n18023) );
  OR2_X1 U22073 ( .A1(n18024), .A2(n18023), .ZN(n18038) );
  NAND2_X1 U22074 ( .A1(n28192), .A2(\xmem_data[25][3] ), .ZN(n18026) );
  NAND2_X1 U22075 ( .A1(n11008), .A2(\xmem_data[24][3] ), .ZN(n18025) );
  NAND2_X1 U22076 ( .A1(n18026), .A2(n18025), .ZN(n18029) );
  AOI22_X1 U22077 ( .A1(n24122), .A2(\xmem_data[26][3] ), .B1(n20710), .B2(
        \xmem_data[27][3] ), .ZN(n18027) );
  INV_X1 U22078 ( .A(n18027), .ZN(n18028) );
  AOI22_X1 U22079 ( .A1(n30544), .A2(\xmem_data[16][3] ), .B1(n24115), .B2(
        \xmem_data[17][3] ), .ZN(n18033) );
  AOI22_X1 U22080 ( .A1(n24116), .A2(\xmem_data[18][3] ), .B1(n3325), .B2(
        \xmem_data[19][3] ), .ZN(n18032) );
  AOI22_X1 U22081 ( .A1(n24117), .A2(\xmem_data[20][3] ), .B1(n30600), .B2(
        \xmem_data[21][3] ), .ZN(n18031) );
  AOI22_X1 U22082 ( .A1(n20507), .A2(\xmem_data[22][3] ), .B1(n29151), .B2(
        \xmem_data[23][3] ), .ZN(n18030) );
  AOI22_X1 U22083 ( .A1(n29118), .A2(\xmem_data[28][3] ), .B1(n27813), .B2(
        \xmem_data[29][3] ), .ZN(n18035) );
  AOI22_X1 U22084 ( .A1(n30589), .A2(\xmem_data[30][3] ), .B1(n25354), .B2(
        \xmem_data[31][3] ), .ZN(n18034) );
  NOR3_X1 U22085 ( .A1(n18038), .A2(n3993), .A3(n18037), .ZN(n18039) );
  XNOR2_X1 U22086 ( .A(n30846), .B(\fmem_data[13][5] ), .ZN(n33164) );
  AOI22_X1 U22087 ( .A1(n3221), .A2(\xmem_data[0][2] ), .B1(n24139), .B2(
        \xmem_data[1][2] ), .ZN(n18049) );
  AOI22_X1 U22088 ( .A1(n24140), .A2(\xmem_data[4][2] ), .B1(n25377), .B2(
        \xmem_data[5][2] ), .ZN(n18043) );
  INV_X1 U22089 ( .A(n18043), .ZN(n18047) );
  AOI22_X1 U22090 ( .A1(n27507), .A2(\xmem_data[2][2] ), .B1(n24141), .B2(
        \xmem_data[3][2] ), .ZN(n18045) );
  NAND2_X1 U22091 ( .A1(n23813), .A2(\xmem_data[7][2] ), .ZN(n18044) );
  NAND2_X1 U22092 ( .A1(n18045), .A2(n18044), .ZN(n18046) );
  NOR2_X1 U22093 ( .A1(n18047), .A2(n18046), .ZN(n18048) );
  NAND2_X1 U22094 ( .A1(n18049), .A2(n18048), .ZN(n18055) );
  AOI22_X1 U22095 ( .A1(n24130), .A2(\xmem_data[8][2] ), .B1(n29403), .B2(
        \xmem_data[9][2] ), .ZN(n18053) );
  AOI22_X1 U22096 ( .A1(n24132), .A2(\xmem_data[10][2] ), .B1(n30891), .B2(
        \xmem_data[11][2] ), .ZN(n18052) );
  AOI22_X1 U22097 ( .A1(n23715), .A2(\xmem_data[12][2] ), .B1(n29315), .B2(
        \xmem_data[13][2] ), .ZN(n18051) );
  AOI22_X1 U22098 ( .A1(n24134), .A2(\xmem_data[14][2] ), .B1(n24133), .B2(
        \xmem_data[15][2] ), .ZN(n18050) );
  NAND4_X1 U22099 ( .A1(n18053), .A2(n18052), .A3(n18051), .A4(n18050), .ZN(
        n18054) );
  OR2_X1 U22100 ( .A1(n18055), .A2(n18054), .ZN(n18068) );
  AOI22_X1 U22101 ( .A1(n24117), .A2(\xmem_data[20][2] ), .B1(n24571), .B2(
        \xmem_data[21][2] ), .ZN(n18059) );
  AOI22_X1 U22102 ( .A1(n28062), .A2(\xmem_data[22][2] ), .B1(n24467), .B2(
        \xmem_data[23][2] ), .ZN(n18058) );
  AOI22_X1 U22103 ( .A1(n24459), .A2(\xmem_data[16][2] ), .B1(n24115), .B2(
        \xmem_data[17][2] ), .ZN(n18057) );
  AOI22_X1 U22104 ( .A1(n20593), .A2(\xmem_data[19][2] ), .B1(
        \xmem_data[18][2] ), .B2(n24116), .ZN(n18056) );
  AOI22_X1 U22105 ( .A1(n24122), .A2(\xmem_data[26][2] ), .B1(n27436), .B2(
        \xmem_data[27][2] ), .ZN(n18063) );
  NAND2_X1 U22106 ( .A1(n30589), .A2(\xmem_data[30][2] ), .ZN(n18062) );
  AND2_X1 U22107 ( .A1(n31256), .A2(\xmem_data[24][2] ), .ZN(n18060) );
  AOI21_X1 U22108 ( .B1(n29725), .B2(\xmem_data[25][2] ), .A(n18060), .ZN(
        n18061) );
  AOI22_X1 U22109 ( .A1(n20489), .A2(\xmem_data[28][2] ), .B1(n29661), .B2(
        \xmem_data[29][2] ), .ZN(n18065) );
  NAND2_X1 U22110 ( .A1(n28503), .A2(\xmem_data[31][2] ), .ZN(n18064) );
  NAND4_X1 U22111 ( .A1(n3841), .A2(n18066), .A3(n18065), .A4(n18064), .ZN(
        n18067) );
  NOR2_X1 U22112 ( .A1(n18068), .A2(n18067), .ZN(n18069) );
  AOI22_X1 U22113 ( .A1(n3220), .A2(\xmem_data[32][2] ), .B1(n30593), .B2(
        \xmem_data[33][2] ), .ZN(n18073) );
  AOI22_X1 U22114 ( .A1(n24207), .A2(\xmem_data[34][2] ), .B1(n22666), .B2(
        \xmem_data[35][2] ), .ZN(n18072) );
  AOI22_X1 U22115 ( .A1(n24633), .A2(\xmem_data[36][2] ), .B1(n3129), .B2(
        \xmem_data[37][2] ), .ZN(n18071) );
  AOI22_X1 U22116 ( .A1(n23771), .A2(\xmem_data[38][2] ), .B1(n25604), .B2(
        \xmem_data[39][2] ), .ZN(n18070) );
  NAND4_X1 U22117 ( .A1(n18073), .A2(n18072), .A3(n18071), .A4(n18070), .ZN(
        n18089) );
  AOI22_X1 U22118 ( .A1(n29180), .A2(\xmem_data[40][2] ), .B1(n27514), .B2(
        \xmem_data[41][2] ), .ZN(n18077) );
  AOI22_X1 U22119 ( .A1(n24212), .A2(\xmem_data[42][2] ), .B1(n31268), .B2(
        \xmem_data[43][2] ), .ZN(n18076) );
  AOI22_X1 U22120 ( .A1(n22674), .A2(\xmem_data[44][2] ), .B1(n27945), .B2(
        \xmem_data[45][2] ), .ZN(n18075) );
  AOI22_X1 U22121 ( .A1(n25574), .A2(\xmem_data[46][2] ), .B1(n24214), .B2(
        \xmem_data[47][2] ), .ZN(n18074) );
  NAND4_X1 U22122 ( .A1(n18077), .A2(n18076), .A3(n18075), .A4(n18074), .ZN(
        n18088) );
  AOI22_X1 U22123 ( .A1(n24219), .A2(\xmem_data[48][2] ), .B1(n30893), .B2(
        \xmem_data[49][2] ), .ZN(n18081) );
  AOI22_X1 U22124 ( .A1(n24221), .A2(\xmem_data[50][2] ), .B1(n3205), .B2(
        \xmem_data[51][2] ), .ZN(n18080) );
  AOI22_X1 U22125 ( .A1(n24222), .A2(\xmem_data[52][2] ), .B1(n28461), .B2(
        \xmem_data[53][2] ), .ZN(n18079) );
  AOI22_X1 U22126 ( .A1(n24223), .A2(\xmem_data[54][2] ), .B1(n20782), .B2(
        \xmem_data[55][2] ), .ZN(n18078) );
  NAND4_X1 U22127 ( .A1(n18081), .A2(n18080), .A3(n18079), .A4(n18078), .ZN(
        n18087) );
  AOI22_X1 U22128 ( .A1(n11008), .A2(\xmem_data[56][2] ), .B1(n27568), .B2(
        \xmem_data[57][2] ), .ZN(n18085) );
  AOI22_X1 U22129 ( .A1(n20579), .A2(\xmem_data[58][2] ), .B1(n25630), .B2(
        \xmem_data[59][2] ), .ZN(n18084) );
  AOI22_X1 U22130 ( .A1(n20489), .A2(\xmem_data[60][2] ), .B1(n3387), .B2(
        \xmem_data[61][2] ), .ZN(n18083) );
  AOI22_X1 U22131 ( .A1(n29173), .A2(\xmem_data[62][2] ), .B1(n25730), .B2(
        \xmem_data[63][2] ), .ZN(n18082) );
  NAND4_X1 U22132 ( .A1(n18085), .A2(n18084), .A3(n18083), .A4(n18082), .ZN(
        n18086) );
  OR4_X1 U22133 ( .A1(n18089), .A2(n18088), .A3(n18087), .A4(n18086), .ZN(
        n18091) );
  NOR2_X1 U22134 ( .A1(n24151), .A2(n39019), .ZN(n18090) );
  AOI21_X1 U22135 ( .B1(n18091), .B2(n24236), .A(n3889), .ZN(n18140) );
  AOI22_X1 U22136 ( .A1(n24158), .A2(\xmem_data[104][2] ), .B1(n24157), .B2(
        \xmem_data[105][2] ), .ZN(n18095) );
  AOI22_X1 U22137 ( .A1(n24159), .A2(\xmem_data[106][2] ), .B1(n3176), .B2(
        \xmem_data[107][2] ), .ZN(n18094) );
  AOI22_X1 U22138 ( .A1(n24160), .A2(\xmem_data[108][2] ), .B1(n3466), .B2(
        \xmem_data[109][2] ), .ZN(n18093) );
  AOI22_X1 U22139 ( .A1(n3207), .A2(\xmem_data[110][2] ), .B1(n25635), .B2(
        \xmem_data[111][2] ), .ZN(n18092) );
  NAND4_X1 U22140 ( .A1(n18095), .A2(n18094), .A3(n18093), .A4(n18092), .ZN(
        n18104) );
  AOI22_X1 U22141 ( .A1(n16989), .A2(\xmem_data[112][2] ), .B1(n23777), .B2(
        \xmem_data[113][2] ), .ZN(n18099) );
  AOI22_X1 U22142 ( .A1(n24165), .A2(\xmem_data[114][2] ), .B1(n20593), .B2(
        \xmem_data[115][2] ), .ZN(n18098) );
  AOI22_X1 U22143 ( .A1(n31361), .A2(\xmem_data[116][2] ), .B1(n23780), .B2(
        \xmem_data[117][2] ), .ZN(n18097) );
  AOI22_X1 U22144 ( .A1(n24167), .A2(\xmem_data[118][2] ), .B1(n24166), .B2(
        \xmem_data[119][2] ), .ZN(n18096) );
  NAND4_X1 U22145 ( .A1(n18099), .A2(n18098), .A3(n18097), .A4(n18096), .ZN(
        n18102) );
  AOI22_X1 U22146 ( .A1(n29326), .A2(\xmem_data[122][2] ), .B1(n27564), .B2(
        \xmem_data[123][2] ), .ZN(n18100) );
  INV_X1 U22147 ( .A(n18100), .ZN(n18101) );
  OR2_X1 U22148 ( .A1(n18102), .A2(n18101), .ZN(n18103) );
  NOR2_X1 U22149 ( .A1(n18104), .A2(n18103), .ZN(n18115) );
  AOI22_X1 U22150 ( .A1(n14981), .A2(\xmem_data[120][2] ), .B1(n29327), .B2(
        \xmem_data[121][2] ), .ZN(n18114) );
  AOI22_X1 U22151 ( .A1(n24172), .A2(\xmem_data[126][2] ), .B1(n27902), .B2(
        \xmem_data[127][2] ), .ZN(n18113) );
  AOI22_X1 U22152 ( .A1(n3220), .A2(\xmem_data[96][2] ), .B1(n20805), .B2(
        \xmem_data[97][2] ), .ZN(n18108) );
  AOI22_X1 U22153 ( .A1(n25509), .A2(\xmem_data[98][2] ), .B1(n25490), .B2(
        \xmem_data[99][2] ), .ZN(n18107) );
  AOI22_X1 U22154 ( .A1(n22759), .A2(\xmem_data[100][2] ), .B1(n3374), .B2(
        \xmem_data[101][2] ), .ZN(n18106) );
  AOI22_X1 U22155 ( .A1(n25492), .A2(\xmem_data[102][2] ), .B1(n28374), .B2(
        \xmem_data[103][2] ), .ZN(n18105) );
  NAND4_X1 U22156 ( .A1(n18108), .A2(n18107), .A3(n18106), .A4(n18105), .ZN(
        n18111) );
  AOI22_X1 U22157 ( .A1(n20578), .A2(\xmem_data[124][2] ), .B1(n3229), .B2(
        \xmem_data[125][2] ), .ZN(n18109) );
  INV_X1 U22158 ( .A(n18109), .ZN(n18110) );
  NOR2_X1 U22159 ( .A1(n18111), .A2(n18110), .ZN(n18112) );
  NAND4_X1 U22160 ( .A1(n18115), .A2(n18114), .A3(n18113), .A4(n18112), .ZN(
        n18138) );
  AOI22_X1 U22161 ( .A1(n20733), .A2(\xmem_data[88][2] ), .B1(n31345), .B2(
        \xmem_data[89][2] ), .ZN(n18120) );
  AOI22_X1 U22162 ( .A1(n24122), .A2(\xmem_data[90][2] ), .B1(n25358), .B2(
        \xmem_data[91][2] ), .ZN(n18119) );
  AOI22_X1 U22163 ( .A1(n25357), .A2(\xmem_data[92][2] ), .B1(n3229), .B2(
        \xmem_data[93][2] ), .ZN(n18118) );
  AND2_X1 U22164 ( .A1(n24172), .A2(\xmem_data[94][2] ), .ZN(n18116) );
  AOI21_X1 U22165 ( .B1(n20991), .B2(\xmem_data[95][2] ), .A(n18116), .ZN(
        n18117) );
  NAND4_X1 U22166 ( .A1(n18120), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18136) );
  AOI22_X1 U22167 ( .A1(n24158), .A2(\xmem_data[72][2] ), .B1(n24157), .B2(
        \xmem_data[73][2] ), .ZN(n18124) );
  AOI22_X1 U22168 ( .A1(n24159), .A2(\xmem_data[74][2] ), .B1(n30514), .B2(
        \xmem_data[75][2] ), .ZN(n18123) );
  AOI22_X1 U22169 ( .A1(n24160), .A2(\xmem_data[76][2] ), .B1(n27818), .B2(
        \xmem_data[77][2] ), .ZN(n18122) );
  AOI22_X1 U22170 ( .A1(n28299), .A2(\xmem_data[78][2] ), .B1(n25635), .B2(
        \xmem_data[79][2] ), .ZN(n18121) );
  NAND4_X1 U22171 ( .A1(n18124), .A2(n18123), .A3(n18122), .A4(n18121), .ZN(
        n18135) );
  AOI22_X1 U22172 ( .A1(n28058), .A2(\xmem_data[80][2] ), .B1(n31255), .B2(
        \xmem_data[81][2] ), .ZN(n18128) );
  AOI22_X1 U22173 ( .A1(n24165), .A2(\xmem_data[82][2] ), .B1(n29100), .B2(
        \xmem_data[83][2] ), .ZN(n18127) );
  AOI22_X1 U22174 ( .A1(n30955), .A2(\xmem_data[84][2] ), .B1(n28955), .B2(
        \xmem_data[85][2] ), .ZN(n18126) );
  AOI22_X1 U22175 ( .A1(n24167), .A2(\xmem_data[86][2] ), .B1(n24166), .B2(
        \xmem_data[87][2] ), .ZN(n18125) );
  NAND4_X1 U22176 ( .A1(n18128), .A2(n18127), .A3(n18126), .A4(n18125), .ZN(
        n18134) );
  AOI22_X1 U22177 ( .A1(n3218), .A2(\xmem_data[64][2] ), .B1(n24533), .B2(
        \xmem_data[65][2] ), .ZN(n18132) );
  AOI22_X1 U22178 ( .A1(n23739), .A2(\xmem_data[66][2] ), .B1(n23812), .B2(
        \xmem_data[67][2] ), .ZN(n18131) );
  AOI22_X1 U22179 ( .A1(n13444), .A2(\xmem_data[68][2] ), .B1(n28344), .B2(
        \xmem_data[69][2] ), .ZN(n18130) );
  AOI22_X1 U22180 ( .A1(n29045), .A2(\xmem_data[70][2] ), .B1(n28374), .B2(
        \xmem_data[71][2] ), .ZN(n18129) );
  NAND4_X1 U22181 ( .A1(n18132), .A2(n18131), .A3(n18130), .A4(n18129), .ZN(
        n18133) );
  AOI22_X1 U22182 ( .A1(n18138), .A2(n24205), .B1(n24204), .B2(n18137), .ZN(
        n18139) );
  XNOR2_X1 U22183 ( .A(n3295), .B(\fmem_data[13][5] ), .ZN(n30815) );
  XNOR2_X1 U22184 ( .A(n31658), .B(\fmem_data[30][3] ), .ZN(n31998) );
  XNOR2_X1 U22185 ( .A(n31655), .B(\fmem_data[30][3] ), .ZN(n32613) );
  XOR2_X1 U22186 ( .A(\fmem_data[30][3] ), .B(\fmem_data[30][2] ), .Z(n18142)
         );
  OAI22_X1 U22187 ( .A1(n31998), .A2(n34435), .B1(n32613), .B2(n34437), .ZN(
        n22780) );
  AOI22_X1 U22188 ( .A1(n29699), .A2(\xmem_data[34][2] ), .B1(n30292), .B2(
        \xmem_data[35][2] ), .ZN(n18146) );
  AOI22_X1 U22189 ( .A1(n27710), .A2(\xmem_data[32][2] ), .B1(n30775), .B2(
        \xmem_data[33][2] ), .ZN(n18145) );
  AOI22_X1 U22190 ( .A1(n30294), .A2(\xmem_data[36][2] ), .B1(n30217), .B2(
        \xmem_data[37][2] ), .ZN(n18144) );
  AOI22_X1 U22191 ( .A1(n30219), .A2(\xmem_data[38][2] ), .B1(n30295), .B2(
        \xmem_data[39][2] ), .ZN(n18143) );
  NAND4_X1 U22192 ( .A1(n18146), .A2(n18145), .A3(n18144), .A4(n18143), .ZN(
        n18152) );
  AOI22_X1 U22193 ( .A1(n3211), .A2(\xmem_data[56][2] ), .B1(n3193), .B2(
        \xmem_data[57][2] ), .ZN(n18150) );
  AOI22_X1 U22194 ( .A1(n30258), .A2(\xmem_data[58][2] ), .B1(n29820), .B2(
        \xmem_data[59][2] ), .ZN(n18149) );
  AOI22_X1 U22195 ( .A1(n30318), .A2(\xmem_data[60][2] ), .B1(n30317), .B2(
        \xmem_data[61][2] ), .ZN(n18148) );
  AOI22_X1 U22196 ( .A1(n30200), .A2(\xmem_data[62][2] ), .B1(n3153), .B2(
        \xmem_data[63][2] ), .ZN(n18147) );
  NAND4_X1 U22197 ( .A1(n18150), .A2(n18149), .A3(n18148), .A4(n18147), .ZN(
        n18151) );
  OR2_X1 U22198 ( .A1(n18152), .A2(n18151), .ZN(n18166) );
  AOI22_X1 U22199 ( .A1(n29590), .A2(\xmem_data[40][2] ), .B1(n30190), .B2(
        \xmem_data[41][2] ), .ZN(n18156) );
  AOI22_X1 U22200 ( .A1(n30300), .A2(\xmem_data[42][2] ), .B1(n17064), .B2(
        \xmem_data[43][2] ), .ZN(n18155) );
  AOI22_X1 U22201 ( .A1(n28779), .A2(\xmem_data[44][2] ), .B1(n28110), .B2(
        \xmem_data[45][2] ), .ZN(n18154) );
  AOI22_X1 U22202 ( .A1(n30304), .A2(\xmem_data[46][2] ), .B1(n20776), .B2(
        \xmem_data[47][2] ), .ZN(n18153) );
  AND4_X1 U22203 ( .A1(n18156), .A2(n18155), .A3(n18154), .A4(n18153), .ZN(
        n18164) );
  AOI22_X1 U22204 ( .A1(n28173), .A2(\xmem_data[52][2] ), .B1(n30765), .B2(
        \xmem_data[53][2] ), .ZN(n18157) );
  AOI22_X1 U22205 ( .A1(n28689), .A2(\xmem_data[50][2] ), .B1(n30309), .B2(
        \xmem_data[51][2] ), .ZN(n18160) );
  AOI22_X1 U22206 ( .A1(n3167), .A2(\xmem_data[48][2] ), .B1(n3183), .B2(
        \xmem_data[49][2] ), .ZN(n18159) );
  AOI22_X1 U22207 ( .A1(n30270), .A2(\xmem_data[54][2] ), .B1(n30311), .B2(
        \xmem_data[55][2] ), .ZN(n18158) );
  NAND3_X1 U22208 ( .A1(n18160), .A2(n18159), .A3(n18158), .ZN(n18161) );
  NOR2_X1 U22209 ( .A1(n18162), .A2(n18161), .ZN(n18163) );
  NAND2_X1 U22210 ( .A1(n18164), .A2(n18163), .ZN(n18165) );
  OAI21_X1 U22211 ( .B1(n18166), .B2(n18165), .A(n30329), .ZN(n18239) );
  AOI22_X1 U22212 ( .A1(n29602), .A2(\xmem_data[72][2] ), .B1(n27761), .B2(
        \xmem_data[73][2] ), .ZN(n18170) );
  AOI22_X1 U22213 ( .A1(n30300), .A2(\xmem_data[74][2] ), .B1(n23792), .B2(
        \xmem_data[75][2] ), .ZN(n18169) );
  AOI22_X1 U22214 ( .A1(n29604), .A2(\xmem_data[76][2] ), .B1(n27728), .B2(
        \xmem_data[77][2] ), .ZN(n18168) );
  AOI22_X1 U22215 ( .A1(n30251), .A2(\xmem_data[78][2] ), .B1(n28752), .B2(
        \xmem_data[79][2] ), .ZN(n18167) );
  AND4_X1 U22216 ( .A1(n18170), .A2(n18169), .A3(n18168), .A4(n18167), .ZN(
        n18184) );
  AOI22_X1 U22217 ( .A1(n3211), .A2(\xmem_data[88][2] ), .B1(n30256), .B2(
        \xmem_data[89][2] ), .ZN(n18174) );
  AOI22_X1 U22218 ( .A1(n30048), .A2(\xmem_data[90][2] ), .B1(n30257), .B2(
        \xmem_data[91][2] ), .ZN(n18173) );
  AOI22_X1 U22219 ( .A1(n30260), .A2(\xmem_data[92][2] ), .B1(n3421), .B2(
        \xmem_data[93][2] ), .ZN(n18172) );
  AOI22_X1 U22220 ( .A1(n30261), .A2(\xmem_data[94][2] ), .B1(n3351), .B2(
        \xmem_data[95][2] ), .ZN(n18171) );
  NAND2_X1 U22221 ( .A1(n30310), .A2(\xmem_data[82][2] ), .ZN(n18179) );
  AOI22_X1 U22222 ( .A1(n30270), .A2(\xmem_data[86][2] ), .B1(n30269), .B2(
        \xmem_data[87][2] ), .ZN(n18176) );
  NAND2_X1 U22223 ( .A1(n16990), .A2(\xmem_data[83][2] ), .ZN(n18175) );
  AOI22_X1 U22224 ( .A1(\xmem_data[80][2] ), .A2(n3162), .B1(n3186), .B2(
        \xmem_data[81][2] ), .ZN(n18177) );
  NAND4_X1 U22225 ( .A1(n3830), .A2(n18179), .A3(n18178), .A4(n18177), .ZN(
        n18182) );
  AOI22_X1 U22226 ( .A1(n29547), .A2(\xmem_data[84][2] ), .B1(n30716), .B2(
        \xmem_data[85][2] ), .ZN(n18180) );
  INV_X1 U22227 ( .A(n18180), .ZN(n18181) );
  NOR2_X1 U22228 ( .A1(n18182), .A2(n18181), .ZN(n18183) );
  NAND2_X1 U22229 ( .A1(n18184), .A2(n18183), .ZN(n18190) );
  AOI22_X1 U22230 ( .A1(n28734), .A2(\xmem_data[64][2] ), .B1(n27013), .B2(
        \xmem_data[65][2] ), .ZN(n18188) );
  AOI22_X1 U22231 ( .A1(n29628), .A2(\xmem_data[66][2] ), .B1(n30292), .B2(
        \xmem_data[67][2] ), .ZN(n18187) );
  AOI22_X1 U22232 ( .A1(n30280), .A2(\xmem_data[68][2] ), .B1(n3198), .B2(
        \xmem_data[69][2] ), .ZN(n18186) );
  AOI22_X1 U22233 ( .A1(n30282), .A2(\xmem_data[70][2] ), .B1(n3138), .B2(
        \xmem_data[71][2] ), .ZN(n18185) );
  NAND4_X1 U22234 ( .A1(n18188), .A2(n18187), .A3(n18186), .A4(n18185), .ZN(
        n18189) );
  OAI21_X1 U22235 ( .B1(n18190), .B2(n18189), .A(n30188), .ZN(n18238) );
  AOI22_X1 U22236 ( .A1(n30743), .A2(\xmem_data[104][2] ), .B1(n29589), .B2(
        \xmem_data[105][2] ), .ZN(n18194) );
  AOI22_X1 U22237 ( .A1(n30192), .A2(\xmem_data[106][2] ), .B1(n24640), .B2(
        \xmem_data[107][2] ), .ZN(n18193) );
  AOI22_X1 U22238 ( .A1(n30745), .A2(\xmem_data[108][2] ), .B1(n30249), .B2(
        \xmem_data[109][2] ), .ZN(n18192) );
  AOI22_X1 U22239 ( .A1(n30251), .A2(\xmem_data[110][2] ), .B1(n31354), .B2(
        \xmem_data[111][2] ), .ZN(n18191) );
  AND4_X1 U22240 ( .A1(n18194), .A2(n18193), .A3(n18192), .A4(n18191), .ZN(
        n18207) );
  AOI22_X1 U22241 ( .A1(n3210), .A2(\xmem_data[120][2] ), .B1(n30256), .B2(
        \xmem_data[121][2] ), .ZN(n18198) );
  AOI22_X1 U22242 ( .A1(n30048), .A2(\xmem_data[122][2] ), .B1(n30257), .B2(
        \xmem_data[123][2] ), .ZN(n18197) );
  AOI22_X1 U22243 ( .A1(n30260), .A2(\xmem_data[124][2] ), .B1(n3420), .B2(
        \xmem_data[125][2] ), .ZN(n18196) );
  NAND2_X1 U22244 ( .A1(n27031), .A2(\xmem_data[114][2] ), .ZN(n18202) );
  AOI22_X1 U22245 ( .A1(n30270), .A2(\xmem_data[118][2] ), .B1(n30269), .B2(
        \xmem_data[119][2] ), .ZN(n18200) );
  NAND2_X1 U22246 ( .A1(n27855), .A2(\xmem_data[115][2] ), .ZN(n18199) );
  AOI22_X1 U22247 ( .A1(\xmem_data[112][2] ), .A2(n3164), .B1(n3185), .B2(
        \xmem_data[113][2] ), .ZN(n18201) );
  NAND4_X1 U22248 ( .A1(n3544), .A2(n18202), .A3(n4008), .A4(n18201), .ZN(
        n18205) );
  AOI22_X1 U22249 ( .A1(n28680), .A2(\xmem_data[116][2] ), .B1(n29487), .B2(
        \xmem_data[117][2] ), .ZN(n18203) );
  INV_X1 U22250 ( .A(n18203), .ZN(n18204) );
  NOR2_X1 U22251 ( .A1(n18205), .A2(n18204), .ZN(n18206) );
  NAND2_X1 U22252 ( .A1(n18207), .A2(n18206), .ZN(n18213) );
  AOI22_X1 U22253 ( .A1(n30291), .A2(\xmem_data[96][2] ), .B1(n30182), .B2(
        \xmem_data[97][2] ), .ZN(n18211) );
  AOI22_X1 U22254 ( .A1(n29790), .A2(\xmem_data[98][2] ), .B1(n30278), .B2(
        \xmem_data[99][2] ), .ZN(n18210) );
  AOI22_X1 U22255 ( .A1(n30280), .A2(\xmem_data[100][2] ), .B1(n3198), .B2(
        \xmem_data[101][2] ), .ZN(n18209) );
  AOI22_X1 U22256 ( .A1(n30282), .A2(\xmem_data[102][2] ), .B1(n3137), .B2(
        \xmem_data[103][2] ), .ZN(n18208) );
  NAND4_X1 U22257 ( .A1(n18211), .A2(n18210), .A3(n18209), .A4(n18208), .ZN(
        n18212) );
  OAI21_X1 U22258 ( .B1(n18213), .B2(n18212), .A(n30287), .ZN(n18237) );
  AOI22_X1 U22259 ( .A1(n28739), .A2(\xmem_data[8][2] ), .B1(n29704), .B2(
        \xmem_data[9][2] ), .ZN(n18217) );
  AOI22_X1 U22260 ( .A1(n30300), .A2(\xmem_data[10][2] ), .B1(n29591), .B2(
        \xmem_data[11][2] ), .ZN(n18216) );
  AOI22_X1 U22261 ( .A1(n27754), .A2(\xmem_data[12][2] ), .B1(n28684), .B2(
        \xmem_data[13][2] ), .ZN(n18215) );
  AOI22_X1 U22262 ( .A1(n30304), .A2(\xmem_data[14][2] ), .B1(n3466), .B2(
        \xmem_data[15][2] ), .ZN(n18214) );
  AOI22_X1 U22263 ( .A1(n29716), .A2(\xmem_data[18][2] ), .B1(n28232), .B2(
        \xmem_data[19][2] ), .ZN(n18227) );
  AOI22_X1 U22264 ( .A1(n3163), .A2(\xmem_data[16][2] ), .B1(n3180), .B2(
        \xmem_data[17][2] ), .ZN(n18226) );
  AOI22_X1 U22265 ( .A1(n3211), .A2(\xmem_data[24][2] ), .B1(n6247), .B2(
        \xmem_data[25][2] ), .ZN(n18221) );
  AOI22_X1 U22266 ( .A1(n30048), .A2(\xmem_data[26][2] ), .B1(n29820), .B2(
        \xmem_data[27][2] ), .ZN(n18220) );
  AOI22_X1 U22267 ( .A1(n30199), .A2(\xmem_data[28][2] ), .B1(n30259), .B2(
        \xmem_data[29][2] ), .ZN(n18219) );
  AOI22_X1 U22268 ( .A1(n30261), .A2(\xmem_data[30][2] ), .B1(n29661), .B2(
        \xmem_data[31][2] ), .ZN(n18218) );
  NAND4_X1 U22269 ( .A1(n18221), .A2(n18220), .A3(n18219), .A4(n18218), .ZN(
        n18224) );
  AOI22_X1 U22270 ( .A1(n30205), .A2(\xmem_data[22][2] ), .B1(n29816), .B2(
        \xmem_data[23][2] ), .ZN(n18222) );
  INV_X1 U22271 ( .A(n18222), .ZN(n18223) );
  NOR2_X1 U22272 ( .A1(n18224), .A2(n18223), .ZN(n18225) );
  AOI22_X1 U22273 ( .A1(n30717), .A2(\xmem_data[20][2] ), .B1(n30266), .B2(
        \xmem_data[21][2] ), .ZN(n18228) );
  NAND3_X1 U22274 ( .A1(n18229), .A2(n3550), .A3(n18228), .ZN(n18235) );
  AOI22_X1 U22275 ( .A1(n28136), .A2(\xmem_data[0][2] ), .B1(n29432), .B2(
        \xmem_data[1][2] ), .ZN(n18233) );
  AOI22_X1 U22276 ( .A1(n28700), .A2(\xmem_data[2][2] ), .B1(n30278), .B2(
        \xmem_data[3][2] ), .ZN(n18232) );
  AOI22_X1 U22277 ( .A1(n30777), .A2(\xmem_data[4][2] ), .B1(n29629), .B2(
        \xmem_data[5][2] ), .ZN(n18231) );
  AOI22_X1 U22278 ( .A1(n30219), .A2(\xmem_data[6][2] ), .B1(n3131), .B2(
        \xmem_data[7][2] ), .ZN(n18230) );
  NAND4_X1 U22279 ( .A1(n18233), .A2(n18232), .A3(n18231), .A4(n18230), .ZN(
        n18234) );
  OAI21_X1 U22280 ( .B1(n18235), .B2(n18234), .A(n30228), .ZN(n18236) );
  XNOR2_X1 U22281 ( .A(n33939), .B(\fmem_data[15][7] ), .ZN(n30334) );
  AOI22_X1 U22282 ( .A1(n29810), .A2(\xmem_data[82][3] ), .B1(n14971), .B2(
        \xmem_data[83][3] ), .ZN(n18242) );
  AOI22_X1 U22283 ( .A1(n3164), .A2(\xmem_data[80][3] ), .B1(n3186), .B2(
        \xmem_data[81][3] ), .ZN(n18241) );
  AOI22_X1 U22284 ( .A1(n30270), .A2(\xmem_data[86][3] ), .B1(n30269), .B2(
        \xmem_data[87][3] ), .ZN(n18240) );
  NAND3_X1 U22285 ( .A1(n18242), .A2(n18241), .A3(n18240), .ZN(n18250) );
  AOI22_X1 U22286 ( .A1(n29488), .A2(\xmem_data[84][3] ), .B1(n30266), .B2(
        \xmem_data[85][3] ), .ZN(n18243) );
  INV_X1 U22287 ( .A(n18243), .ZN(n18249) );
  AOI22_X1 U22288 ( .A1(n3210), .A2(\xmem_data[88][3] ), .B1(n30256), .B2(
        \xmem_data[89][3] ), .ZN(n18247) );
  AOI22_X1 U22289 ( .A1(n30258), .A2(\xmem_data[90][3] ), .B1(n30257), .B2(
        \xmem_data[91][3] ), .ZN(n18246) );
  AOI22_X1 U22290 ( .A1(n30260), .A2(\xmem_data[92][3] ), .B1(n3421), .B2(
        \xmem_data[93][3] ), .ZN(n18245) );
  AOI22_X1 U22291 ( .A1(n30200), .A2(\xmem_data[94][3] ), .B1(n3332), .B2(
        \xmem_data[95][3] ), .ZN(n18244) );
  NAND4_X1 U22292 ( .A1(n18247), .A2(n18246), .A3(n18245), .A4(n18244), .ZN(
        n18248) );
  AOI22_X1 U22293 ( .A1(n30633), .A2(\xmem_data[72][3] ), .B1(n28665), .B2(
        \xmem_data[73][3] ), .ZN(n18254) );
  AOI22_X1 U22294 ( .A1(n30171), .A2(\xmem_data[74][3] ), .B1(n28671), .B2(
        \xmem_data[75][3] ), .ZN(n18253) );
  AOI22_X1 U22295 ( .A1(n30250), .A2(\xmem_data[76][3] ), .B1(n30634), .B2(
        \xmem_data[77][3] ), .ZN(n18252) );
  AOI22_X1 U22296 ( .A1(n30251), .A2(\xmem_data[78][3] ), .B1(n27755), .B2(
        \xmem_data[79][3] ), .ZN(n18251) );
  AND4_X1 U22297 ( .A1(n18254), .A2(n18253), .A3(n18252), .A4(n18251), .ZN(
        n18255) );
  NAND2_X1 U22298 ( .A1(n18256), .A2(n18255), .ZN(n18262) );
  AOI22_X1 U22299 ( .A1(n29433), .A2(\xmem_data[64][3] ), .B1(n30290), .B2(
        \xmem_data[65][3] ), .ZN(n18260) );
  AOI22_X1 U22300 ( .A1(n30279), .A2(\xmem_data[66][3] ), .B1(n30292), .B2(
        \xmem_data[67][3] ), .ZN(n18259) );
  AOI22_X1 U22301 ( .A1(n30280), .A2(\xmem_data[68][3] ), .B1(n3170), .B2(
        \xmem_data[69][3] ), .ZN(n18258) );
  AOI22_X1 U22302 ( .A1(n30282), .A2(\xmem_data[70][3] ), .B1(n3137), .B2(
        \xmem_data[71][3] ), .ZN(n18257) );
  NAND4_X1 U22303 ( .A1(n18260), .A2(n18259), .A3(n18258), .A4(n18257), .ZN(
        n18261) );
  OAI21_X1 U22304 ( .B1(n18262), .B2(n18261), .A(n30188), .ZN(n18345) );
  AOI22_X1 U22305 ( .A1(n29699), .A2(\xmem_data[98][3] ), .B1(n30278), .B2(
        \xmem_data[99][3] ), .ZN(n18263) );
  INV_X1 U22306 ( .A(n18263), .ZN(n18272) );
  AOI22_X1 U22307 ( .A1(n30270), .A2(\xmem_data[118][3] ), .B1(n30269), .B2(
        \xmem_data[119][3] ), .ZN(n18264) );
  INV_X1 U22308 ( .A(n18264), .ZN(n18265) );
  AOI21_X1 U22309 ( .B1(\xmem_data[105][3] ), .B2(n28738), .A(n18265), .ZN(
        n18270) );
  AOI22_X1 U22310 ( .A1(n3211), .A2(\xmem_data[120][3] ), .B1(n30256), .B2(
        \xmem_data[121][3] ), .ZN(n18269) );
  AOI22_X1 U22311 ( .A1(n30048), .A2(\xmem_data[122][3] ), .B1(n30257), .B2(
        \xmem_data[123][3] ), .ZN(n18268) );
  AOI22_X1 U22312 ( .A1(n30260), .A2(\xmem_data[124][3] ), .B1(n3421), .B2(
        \xmem_data[125][3] ), .ZN(n18267) );
  AOI22_X1 U22313 ( .A1(n30200), .A2(\xmem_data[126][3] ), .B1(n3412), .B2(
        \xmem_data[127][3] ), .ZN(n18266) );
  NAND2_X1 U22314 ( .A1(n18270), .A2(n3756), .ZN(n18271) );
  NOR2_X1 U22315 ( .A1(n18272), .A2(n18271), .ZN(n18290) );
  AOI22_X1 U22316 ( .A1(n29626), .A2(\xmem_data[96][3] ), .B1(n30100), .B2(
        \xmem_data[97][3] ), .ZN(n18273) );
  INV_X1 U22317 ( .A(n18273), .ZN(n18276) );
  AOI22_X1 U22318 ( .A1(n30280), .A2(\xmem_data[100][3] ), .B1(n3198), .B2(
        \xmem_data[101][3] ), .ZN(n18274) );
  INV_X1 U22319 ( .A(n18274), .ZN(n18275) );
  NOR2_X1 U22320 ( .A1(n18276), .A2(n18275), .ZN(n18289) );
  AOI22_X1 U22321 ( .A1(n3162), .A2(\xmem_data[112][3] ), .B1(n3187), .B2(
        \xmem_data[113][3] ), .ZN(n18278) );
  AOI22_X1 U22322 ( .A1(n30250), .A2(\xmem_data[108][3] ), .B1(n30084), .B2(
        \xmem_data[109][3] ), .ZN(n18277) );
  NAND2_X1 U22323 ( .A1(n18278), .A2(n18277), .ZN(n18284) );
  AOI22_X1 U22324 ( .A1(n30171), .A2(\xmem_data[106][3] ), .B1(n28233), .B2(
        \xmem_data[107][3] ), .ZN(n18279) );
  INV_X1 U22325 ( .A(n18279), .ZN(n18280) );
  AOI21_X1 U22326 ( .B1(n29647), .B2(\xmem_data[104][3] ), .A(n18280), .ZN(
        n18282) );
  AOI22_X1 U22327 ( .A1(n30062), .A2(\xmem_data[114][3] ), .B1(n23722), .B2(
        \xmem_data[115][3] ), .ZN(n18281) );
  NAND2_X1 U22328 ( .A1(n18282), .A2(n18281), .ZN(n18283) );
  NOR2_X1 U22329 ( .A1(n18284), .A2(n18283), .ZN(n18288) );
  AOI22_X1 U22330 ( .A1(n27713), .A2(\xmem_data[116][3] ), .B1(n30716), .B2(
        \xmem_data[117][3] ), .ZN(n18287) );
  AOI22_X1 U22331 ( .A1(n30251), .A2(\xmem_data[110][3] ), .B1(n20718), .B2(
        \xmem_data[111][3] ), .ZN(n18286) );
  AOI22_X1 U22332 ( .A1(n30282), .A2(\xmem_data[102][3] ), .B1(n3137), .B2(
        \xmem_data[103][3] ), .ZN(n18285) );
  NAND4_X1 U22333 ( .A1(n18290), .A2(n18289), .A3(n18288), .A4(n3900), .ZN(
        n18291) );
  NAND2_X1 U22334 ( .A1(n18291), .A2(n30287), .ZN(n18344) );
  AOI22_X1 U22335 ( .A1(n30745), .A2(\xmem_data[44][3] ), .B1(n30237), .B2(
        \xmem_data[45][3] ), .ZN(n18292) );
  INV_X1 U22336 ( .A(n18292), .ZN(n18296) );
  AOI22_X1 U22337 ( .A1(n30270), .A2(\xmem_data[54][3] ), .B1(n30311), .B2(
        \xmem_data[55][3] ), .ZN(n18294) );
  AOI22_X1 U22338 ( .A1(n30304), .A2(\xmem_data[46][3] ), .B1(n27517), .B2(
        \xmem_data[47][3] ), .ZN(n18293) );
  NAND2_X1 U22339 ( .A1(n18294), .A2(n18293), .ZN(n18295) );
  NOR2_X1 U22340 ( .A1(n18296), .A2(n18295), .ZN(n18306) );
  AOI22_X1 U22341 ( .A1(\xmem_data[40][3] ), .A2(n29446), .B1(n28689), .B2(
        \xmem_data[50][3] ), .ZN(n18298) );
  NAND2_X1 U22342 ( .A1(n29347), .A2(\xmem_data[41][3] ), .ZN(n18297) );
  AOI22_X1 U22343 ( .A1(n30766), .A2(\xmem_data[52][3] ), .B1(n29640), .B2(
        \xmem_data[53][3] ), .ZN(n18299) );
  AOI22_X1 U22344 ( .A1(n3163), .A2(\xmem_data[48][3] ), .B1(n3191), .B2(
        \xmem_data[49][3] ), .ZN(n18300) );
  INV_X1 U22345 ( .A(n18300), .ZN(n18303) );
  AOI22_X1 U22346 ( .A1(n30171), .A2(\xmem_data[42][3] ), .B1(n29591), .B2(
        \xmem_data[43][3] ), .ZN(n18301) );
  INV_X1 U22347 ( .A(n18301), .ZN(n18302) );
  NOR2_X1 U22348 ( .A1(n18303), .A2(n3995), .ZN(n18304) );
  NAND4_X1 U22349 ( .A1(n18306), .A2(n18305), .A3(n18299), .A4(n18304), .ZN(
        n18318) );
  AOI22_X1 U22350 ( .A1(n28136), .A2(\xmem_data[32][3] ), .B1(n29831), .B2(
        \xmem_data[33][3] ), .ZN(n18310) );
  AOI22_X1 U22351 ( .A1(n30279), .A2(\xmem_data[34][3] ), .B1(n30292), .B2(
        \xmem_data[35][3] ), .ZN(n18309) );
  AOI22_X1 U22352 ( .A1(n30294), .A2(\xmem_data[36][3] ), .B1(n30293), .B2(
        \xmem_data[37][3] ), .ZN(n18308) );
  AOI22_X1 U22353 ( .A1(n30219), .A2(\xmem_data[38][3] ), .B1(n30295), .B2(
        \xmem_data[39][3] ), .ZN(n18307) );
  NAND4_X1 U22354 ( .A1(n18310), .A2(n18309), .A3(n18308), .A4(n18307), .ZN(
        n18316) );
  AOI22_X1 U22355 ( .A1(n3210), .A2(\xmem_data[56][3] ), .B1(n3193), .B2(
        \xmem_data[57][3] ), .ZN(n18314) );
  AOI22_X1 U22356 ( .A1(n30258), .A2(\xmem_data[58][3] ), .B1(n27568), .B2(
        \xmem_data[59][3] ), .ZN(n18313) );
  AOI22_X1 U22357 ( .A1(n30318), .A2(\xmem_data[60][3] ), .B1(n30317), .B2(
        \xmem_data[61][3] ), .ZN(n18312) );
  AOI22_X1 U22358 ( .A1(n30200), .A2(\xmem_data[62][3] ), .B1(n3153), .B2(
        \xmem_data[63][3] ), .ZN(n18311) );
  NAND4_X1 U22359 ( .A1(n18314), .A2(n18313), .A3(n18312), .A4(n18311), .ZN(
        n18315) );
  OR2_X1 U22360 ( .A1(n18316), .A2(n18315), .ZN(n18317) );
  OAI21_X1 U22361 ( .B1(n18318), .B2(n18317), .A(n30329), .ZN(n18343) );
  AOI22_X1 U22362 ( .A1(n30764), .A2(\xmem_data[18][3] ), .B1(n28754), .B2(
        \xmem_data[19][3] ), .ZN(n18322) );
  AOI22_X1 U22363 ( .A1(n3168), .A2(\xmem_data[16][3] ), .B1(n3184), .B2(
        \xmem_data[17][3] ), .ZN(n18321) );
  AOI22_X1 U22364 ( .A1(n29547), .A2(\xmem_data[20][3] ), .B1(n30644), .B2(
        \xmem_data[21][3] ), .ZN(n18320) );
  AOI22_X1 U22365 ( .A1(n30205), .A2(\xmem_data[22][3] ), .B1(n30311), .B2(
        \xmem_data[23][3] ), .ZN(n18319) );
  NAND4_X1 U22366 ( .A1(n18322), .A2(n18321), .A3(n18320), .A4(n18319), .ZN(
        n18329) );
  AOI22_X1 U22367 ( .A1(n30199), .A2(\xmem_data[28][3] ), .B1(n3420), .B2(
        \xmem_data[29][3] ), .ZN(n18327) );
  AOI22_X1 U22368 ( .A1(n30320), .A2(\xmem_data[30][3] ), .B1(n3352), .B2(
        \xmem_data[31][3] ), .ZN(n18326) );
  AOI22_X1 U22369 ( .A1(n3210), .A2(\xmem_data[24][3] ), .B1(n3192), .B2(
        \xmem_data[25][3] ), .ZN(n18324) );
  AOI22_X1 U22370 ( .A1(n30048), .A2(\xmem_data[26][3] ), .B1(n14982), .B2(
        \xmem_data[27][3] ), .ZN(n18323) );
  AND2_X1 U22371 ( .A1(n18324), .A2(n18323), .ZN(n18325) );
  NAND3_X1 U22372 ( .A1(n18327), .A2(n18326), .A3(n18325), .ZN(n18328) );
  NOR2_X1 U22373 ( .A1(n18329), .A2(n18328), .ZN(n18340) );
  AOI22_X1 U22374 ( .A1(n30191), .A2(\xmem_data[8][3] ), .B1(n28738), .B2(
        \xmem_data[9][3] ), .ZN(n18333) );
  AOI22_X1 U22375 ( .A1(n30171), .A2(\xmem_data[10][3] ), .B1(n30083), .B2(
        \xmem_data[11][3] ), .ZN(n18332) );
  AOI22_X1 U22376 ( .A1(n29436), .A2(\xmem_data[12][3] ), .B1(n28684), .B2(
        \xmem_data[13][3] ), .ZN(n18331) );
  AOI22_X1 U22377 ( .A1(n30304), .A2(\xmem_data[14][3] ), .B1(n30666), .B2(
        \xmem_data[15][3] ), .ZN(n18330) );
  AND4_X1 U22378 ( .A1(n18333), .A2(n18332), .A3(n18331), .A4(n18330), .ZN(
        n18339) );
  AOI22_X1 U22379 ( .A1(n29433), .A2(\xmem_data[0][3] ), .B1(n30100), .B2(
        \xmem_data[1][3] ), .ZN(n18337) );
  AOI22_X1 U22380 ( .A1(n27740), .A2(\xmem_data[2][3] ), .B1(n29565), .B2(
        \xmem_data[3][3] ), .ZN(n18336) );
  AOI22_X1 U22381 ( .A1(n27771), .A2(\xmem_data[4][3] ), .B1(n28667), .B2(
        \xmem_data[5][3] ), .ZN(n18335) );
  AOI22_X1 U22382 ( .A1(n30219), .A2(\xmem_data[6][3] ), .B1(n3132), .B2(
        \xmem_data[7][3] ), .ZN(n18334) );
  AND4_X1 U22383 ( .A1(n18337), .A2(n18336), .A3(n18335), .A4(n18334), .ZN(
        n18338) );
  NAND3_X1 U22384 ( .A1(n18340), .A2(n18339), .A3(n18338), .ZN(n18341) );
  NAND2_X1 U22385 ( .A1(n18341), .A2(n30228), .ZN(n18342) );
  XNOR2_X1 U22386 ( .A(n3425), .B(\fmem_data[15][7] ), .ZN(n33234) );
  OAI22_X1 U22387 ( .A1(n30334), .A2(n35696), .B1(n33234), .B2(n35697), .ZN(
        n23602) );
  AOI22_X1 U22388 ( .A1(n29786), .A2(\xmem_data[32][4] ), .B1(n29785), .B2(
        \xmem_data[33][4] ), .ZN(n18349) );
  AOI22_X1 U22389 ( .A1(n29787), .A2(\xmem_data[34][4] ), .B1(n28039), .B2(
        \xmem_data[35][4] ), .ZN(n18348) );
  AOI22_X1 U22390 ( .A1(n27741), .A2(\xmem_data[36][4] ), .B1(n30290), .B2(
        \xmem_data[37][4] ), .ZN(n18347) );
  AOI22_X1 U22391 ( .A1(n29699), .A2(\xmem_data[38][4] ), .B1(n29789), .B2(
        \xmem_data[39][4] ), .ZN(n18346) );
  NAND4_X1 U22392 ( .A1(n18349), .A2(n18348), .A3(n18347), .A4(n18346), .ZN(
        n18365) );
  AOI22_X1 U22393 ( .A1(n28209), .A2(\xmem_data[40][4] ), .B1(n29798), .B2(
        \xmem_data[41][4] ), .ZN(n18353) );
  AOI22_X1 U22394 ( .A1(n29707), .A2(\xmem_data[42][4] ), .B1(n3375), .B2(
        \xmem_data[43][4] ), .ZN(n18352) );
  AOI22_X1 U22395 ( .A1(n29446), .A2(\xmem_data[44][4] ), .B1(n30190), .B2(
        \xmem_data[45][4] ), .ZN(n18351) );
  AOI22_X1 U22396 ( .A1(n29763), .A2(\xmem_data[46][4] ), .B1(n29308), .B2(
        \xmem_data[47][4] ), .ZN(n18350) );
  NAND4_X1 U22397 ( .A1(n18353), .A2(n18352), .A3(n18351), .A4(n18350), .ZN(
        n18364) );
  AOI22_X1 U22398 ( .A1(n30745), .A2(\xmem_data[48][4] ), .B1(n26884), .B2(
        \xmem_data[49][4] ), .ZN(n18357) );
  AOI22_X1 U22399 ( .A1(n29740), .A2(\xmem_data[50][4] ), .B1(n29605), .B2(
        \xmem_data[51][4] ), .ZN(n18356) );
  AOI22_X1 U22400 ( .A1(n3165), .A2(\xmem_data[52][4] ), .B1(n3191), .B2(
        \xmem_data[53][4] ), .ZN(n18355) );
  AOI22_X1 U22401 ( .A1(n26812), .A2(\xmem_data[54][4] ), .B1(n22717), .B2(
        \xmem_data[55][4] ), .ZN(n18354) );
  NAND4_X1 U22402 ( .A1(n18357), .A2(n18356), .A3(n18355), .A4(n18354), .ZN(
        n18363) );
  AOI22_X1 U22403 ( .A1(n27713), .A2(\xmem_data[56][4] ), .B1(n30644), .B2(
        \xmem_data[57][4] ), .ZN(n18361) );
  AOI22_X1 U22404 ( .A1(n3226), .A2(\xmem_data[58][4] ), .B1(n29816), .B2(
        \xmem_data[59][4] ), .ZN(n18360) );
  AOI22_X1 U22405 ( .A1(n29819), .A2(\xmem_data[60][4] ), .B1(n29818), .B2(
        \xmem_data[61][4] ), .ZN(n18359) );
  AOI22_X1 U22406 ( .A1(n29821), .A2(\xmem_data[62][4] ), .B1(n29820), .B2(
        \xmem_data[63][4] ), .ZN(n18358) );
  NAND4_X1 U22407 ( .A1(n18361), .A2(n18360), .A3(n18359), .A4(n18358), .ZN(
        n18362) );
  AOI22_X1 U22408 ( .A1(n29829), .A2(\xmem_data[0][4] ), .B1(n29695), .B2(
        \xmem_data[1][4] ), .ZN(n18369) );
  AOI22_X1 U22409 ( .A1(n29696), .A2(\xmem_data[2][4] ), .B1(n3153), .B2(
        \xmem_data[3][4] ), .ZN(n18368) );
  AOI22_X1 U22410 ( .A1(n30223), .A2(\xmem_data[4][4] ), .B1(n27832), .B2(
        \xmem_data[5][4] ), .ZN(n18367) );
  AOI22_X1 U22411 ( .A1(n30215), .A2(\xmem_data[6][4] ), .B1(n29698), .B2(
        \xmem_data[7][4] ), .ZN(n18366) );
  AOI22_X1 U22412 ( .A1(n27703), .A2(\xmem_data[12][4] ), .B1(n29704), .B2(
        \xmem_data[13][4] ), .ZN(n18373) );
  AOI22_X1 U22413 ( .A1(n29707), .A2(\xmem_data[10][4] ), .B1(n29706), .B2(
        \xmem_data[11][4] ), .ZN(n18372) );
  AOI22_X1 U22414 ( .A1(n29566), .A2(\xmem_data[8][4] ), .B1(n30293), .B2(
        \xmem_data[9][4] ), .ZN(n18371) );
  AOI22_X1 U22415 ( .A1(n29709), .A2(\xmem_data[14][4] ), .B1(n28152), .B2(
        \xmem_data[15][4] ), .ZN(n18370) );
  AOI22_X1 U22416 ( .A1(n28685), .A2(\xmem_data[16][4] ), .B1(n30634), .B2(
        \xmem_data[17][4] ), .ZN(n18377) );
  AOI22_X1 U22417 ( .A1(n29740), .A2(\xmem_data[18][4] ), .B1(n27818), .B2(
        \xmem_data[19][4] ), .ZN(n18376) );
  AOI22_X1 U22418 ( .A1(n3165), .A2(\xmem_data[20][4] ), .B1(n3191), .B2(
        \xmem_data[21][4] ), .ZN(n18375) );
  AOI22_X1 U22419 ( .A1(n29476), .A2(\xmem_data[22][4] ), .B1(n28147), .B2(
        \xmem_data[23][4] ), .ZN(n18374) );
  AOI22_X1 U22420 ( .A1(n28680), .A2(\xmem_data[24][4] ), .B1(n30765), .B2(
        \xmem_data[25][4] ), .ZN(n18381) );
  AOI22_X1 U22421 ( .A1(n3226), .A2(\xmem_data[26][4] ), .B1(n28461), .B2(
        \xmem_data[27][4] ), .ZN(n18380) );
  AOI22_X1 U22422 ( .A1(n29724), .A2(\xmem_data[28][4] ), .B1(n29723), .B2(
        \xmem_data[29][4] ), .ZN(n18379) );
  AOI22_X1 U22423 ( .A1(n29726), .A2(\xmem_data[30][4] ), .B1(n29725), .B2(
        \xmem_data[31][4] ), .ZN(n18378) );
  AOI22_X1 U22424 ( .A1(n29795), .A2(n18383), .B1(n29733), .B2(n18382), .ZN(
        n18428) );
  AOI22_X1 U22425 ( .A1(n29829), .A2(\xmem_data[96][4] ), .B1(n29785), .B2(
        \xmem_data[97][4] ), .ZN(n18387) );
  AOI22_X1 U22426 ( .A1(n29830), .A2(\xmem_data[98][4] ), .B1(n3144), .B2(
        \xmem_data[99][4] ), .ZN(n18386) );
  AOI22_X1 U22427 ( .A1(n29421), .A2(\xmem_data[100][4] ), .B1(n27013), .B2(
        \xmem_data[101][4] ), .ZN(n18385) );
  AOI22_X1 U22428 ( .A1(n30279), .A2(\xmem_data[102][4] ), .B1(n29832), .B2(
        \xmem_data[103][4] ), .ZN(n18384) );
  NAND4_X1 U22429 ( .A1(n18387), .A2(n18386), .A3(n18385), .A4(n18384), .ZN(
        n18403) );
  AOI22_X1 U22430 ( .A1(n29799), .A2(\xmem_data[104][4] ), .B1(n30776), .B2(
        \xmem_data[105][4] ), .ZN(n18391) );
  AOI22_X1 U22431 ( .A1(n29800), .A2(\xmem_data[106][4] ), .B1(n29706), .B2(
        \xmem_data[107][4] ), .ZN(n18390) );
  AOI22_X1 U22432 ( .A1(n28146), .A2(\xmem_data[108][4] ), .B1(n27761), .B2(
        \xmem_data[109][4] ), .ZN(n18389) );
  AOI22_X1 U22433 ( .A1(n29802), .A2(\xmem_data[110][4] ), .B1(n30744), .B2(
        \xmem_data[111][4] ), .ZN(n18388) );
  NAND4_X1 U22434 ( .A1(n18391), .A2(n18390), .A3(n18389), .A4(n18388), .ZN(
        n18402) );
  AOI22_X1 U22435 ( .A1(n27811), .A2(\xmem_data[112][4] ), .B1(n27753), .B2(
        \xmem_data[113][4] ), .ZN(n18395) );
  AOI22_X1 U22436 ( .A1(n29771), .A2(\xmem_data[114][4] ), .B1(n29807), .B2(
        \xmem_data[115][4] ), .ZN(n18394) );
  AOI22_X1 U22437 ( .A1(n3168), .A2(\xmem_data[116][4] ), .B1(n3182), .B2(
        \xmem_data[117][4] ), .ZN(n18393) );
  AOI22_X1 U22438 ( .A1(n30062), .A2(\xmem_data[118][4] ), .B1(n28994), .B2(
        \xmem_data[119][4] ), .ZN(n18392) );
  NAND4_X1 U22439 ( .A1(n18392), .A2(n18394), .A3(n18393), .A4(n18395), .ZN(
        n18401) );
  AOI22_X1 U22440 ( .A1(n29815), .A2(\xmem_data[120][4] ), .B1(n30170), .B2(
        \xmem_data[121][4] ), .ZN(n18399) );
  AOI22_X1 U22441 ( .A1(n29817), .A2(\xmem_data[122][4] ), .B1(n29324), .B2(
        \xmem_data[123][4] ), .ZN(n18398) );
  AOI22_X1 U22442 ( .A1(n29777), .A2(\xmem_data[124][4] ), .B1(n29723), .B2(
        \xmem_data[125][4] ), .ZN(n18397) );
  AOI22_X1 U22443 ( .A1(n29384), .A2(\xmem_data[126][4] ), .B1(n29725), .B2(
        \xmem_data[127][4] ), .ZN(n18396) );
  NAND4_X1 U22444 ( .A1(n18399), .A2(n18398), .A3(n18397), .A4(n18396), .ZN(
        n18400) );
  AOI22_X1 U22445 ( .A1(n28139), .A2(\xmem_data[72][4] ), .B1(n3197), .B2(
        \xmem_data[73][4] ), .ZN(n18407) );
  AOI22_X1 U22446 ( .A1(n29707), .A2(\xmem_data[74][4] ), .B1(n29762), .B2(
        \xmem_data[75][4] ), .ZN(n18406) );
  AOI22_X1 U22447 ( .A1(n28180), .A2(\xmem_data[76][4] ), .B1(n30190), .B2(
        \xmem_data[77][4] ), .ZN(n18405) );
  AOI22_X1 U22448 ( .A1(n29763), .A2(\xmem_data[78][4] ), .B1(n20799), .B2(
        \xmem_data[79][4] ), .ZN(n18404) );
  NAND4_X1 U22449 ( .A1(n18407), .A2(n18406), .A3(n18405), .A4(n18404), .ZN(
        n18424) );
  AOI22_X1 U22450 ( .A1(n28765), .A2(\xmem_data[64][4] ), .B1(n29785), .B2(
        \xmem_data[65][4] ), .ZN(n18411) );
  AOI22_X1 U22451 ( .A1(n29787), .A2(\xmem_data[66][4] ), .B1(n3413), .B2(
        \xmem_data[67][4] ), .ZN(n18410) );
  AOI22_X1 U22452 ( .A1(n27741), .A2(\xmem_data[68][4] ), .B1(n28206), .B2(
        \xmem_data[69][4] ), .ZN(n18409) );
  AOI22_X1 U22453 ( .A1(n3392), .A2(\xmem_data[70][4] ), .B1(n29789), .B2(
        \xmem_data[71][4] ), .ZN(n18408) );
  NAND4_X1 U22454 ( .A1(n18411), .A2(n18410), .A3(n18409), .A4(n18408), .ZN(
        n18423) );
  AOI22_X1 U22455 ( .A1(n30745), .A2(\xmem_data[80][4] ), .B1(n30090), .B2(
        \xmem_data[81][4] ), .ZN(n18416) );
  AOI22_X1 U22456 ( .A1(n29808), .A2(\xmem_data[82][4] ), .B1(n28053), .B2(
        \xmem_data[83][4] ), .ZN(n18415) );
  AOI22_X1 U22457 ( .A1(n3168), .A2(\xmem_data[84][4] ), .B1(n3181), .B2(
        \xmem_data[85][4] ), .ZN(n18414) );
  AND2_X1 U22458 ( .A1(n29410), .A2(\xmem_data[87][4] ), .ZN(n18412) );
  AOI21_X1 U22459 ( .B1(n27031), .B2(\xmem_data[86][4] ), .A(n18412), .ZN(
        n18413) );
  NAND4_X1 U22460 ( .A1(n18416), .A2(n18415), .A3(n18414), .A4(n18413), .ZN(
        n18422) );
  AOI22_X1 U22461 ( .A1(n30076), .A2(\xmem_data[88][4] ), .B1(n30644), .B2(
        \xmem_data[89][4] ), .ZN(n18420) );
  AOI22_X1 U22462 ( .A1(n3226), .A2(\xmem_data[90][4] ), .B1(n30311), .B2(
        \xmem_data[91][4] ), .ZN(n18419) );
  AOI22_X1 U22463 ( .A1(n29777), .A2(\xmem_data[92][4] ), .B1(n29776), .B2(
        \xmem_data[93][4] ), .ZN(n18418) );
  AOI22_X1 U22464 ( .A1(n27718), .A2(\xmem_data[94][4] ), .B1(n30674), .B2(
        \xmem_data[95][4] ), .ZN(n18417) );
  NAND4_X1 U22465 ( .A1(n18420), .A2(n18419), .A3(n18418), .A4(n18417), .ZN(
        n18421) );
  AOI22_X1 U22466 ( .A1(n18426), .A2(n29837), .B1(n18425), .B2(n29758), .ZN(
        n18427) );
  NAND2_X1 U22467 ( .A1(n18428), .A2(n18427), .ZN(n32727) );
  XNOR2_X1 U22468 ( .A(n32727), .B(\fmem_data[19][5] ), .ZN(n22454) );
  XOR2_X1 U22469 ( .A(\fmem_data[19][4] ), .B(\fmem_data[19][5] ), .Z(n18429)
         );
  AOI22_X1 U22470 ( .A1(n28765), .A2(\xmem_data[96][5] ), .B1(n29785), .B2(
        \xmem_data[97][5] ), .ZN(n18433) );
  AOI22_X1 U22471 ( .A1(n29830), .A2(\xmem_data[98][5] ), .B1(n3153), .B2(
        \xmem_data[99][5] ), .ZN(n18432) );
  AOI22_X1 U22472 ( .A1(n28734), .A2(\xmem_data[100][5] ), .B1(n30182), .B2(
        \xmem_data[101][5] ), .ZN(n18431) );
  AOI22_X1 U22473 ( .A1(n29790), .A2(\xmem_data[102][5] ), .B1(n29832), .B2(
        \xmem_data[103][5] ), .ZN(n18430) );
  NAND4_X1 U22474 ( .A1(n18433), .A2(n18432), .A3(n18431), .A4(n18430), .ZN(
        n18450) );
  AOI22_X1 U22475 ( .A1(n29799), .A2(\xmem_data[104][5] ), .B1(n29708), .B2(
        \xmem_data[105][5] ), .ZN(n18437) );
  AOI22_X1 U22476 ( .A1(n29800), .A2(\xmem_data[106][5] ), .B1(n3375), .B2(
        \xmem_data[107][5] ), .ZN(n18436) );
  AOI22_X1 U22477 ( .A1(n29602), .A2(\xmem_data[108][5] ), .B1(n27761), .B2(
        \xmem_data[109][5] ), .ZN(n18435) );
  AOI22_X1 U22478 ( .A1(n29802), .A2(\xmem_data[110][5] ), .B1(n28089), .B2(
        \xmem_data[111][5] ), .ZN(n18434) );
  NAND4_X1 U22479 ( .A1(n18437), .A2(n18436), .A3(n18435), .A4(n18434), .ZN(
        n18449) );
  AOI22_X1 U22480 ( .A1(n3164), .A2(\xmem_data[116][5] ), .B1(n3183), .B2(
        \xmem_data[117][5] ), .ZN(n18442) );
  AOI22_X1 U22481 ( .A1(n29808), .A2(\xmem_data[114][5] ), .B1(n29807), .B2(
        \xmem_data[115][5] ), .ZN(n18441) );
  AOI22_X1 U22482 ( .A1(n27811), .A2(\xmem_data[112][5] ), .B1(n28110), .B2(
        \xmem_data[113][5] ), .ZN(n18440) );
  AND2_X1 U22483 ( .A1(n28232), .A2(\xmem_data[119][5] ), .ZN(n18438) );
  AOI21_X1 U22484 ( .B1(n28755), .B2(\xmem_data[118][5] ), .A(n18438), .ZN(
        n18439) );
  NAND4_X1 U22485 ( .A1(n18442), .A2(n18441), .A3(n18440), .A4(n18439), .ZN(
        n18448) );
  AOI22_X1 U22486 ( .A1(n30063), .A2(\xmem_data[120][5] ), .B1(n30765), .B2(
        \xmem_data[121][5] ), .ZN(n18446) );
  AOI22_X1 U22487 ( .A1(n29817), .A2(\xmem_data[122][5] ), .B1(n29816), .B2(
        \xmem_data[123][5] ), .ZN(n18445) );
  AOI22_X1 U22488 ( .A1(n29819), .A2(\xmem_data[124][5] ), .B1(n29818), .B2(
        \xmem_data[125][5] ), .ZN(n18444) );
  AOI22_X1 U22489 ( .A1(n29821), .A2(\xmem_data[126][5] ), .B1(n29820), .B2(
        \xmem_data[127][5] ), .ZN(n18443) );
  NAND4_X1 U22490 ( .A1(n18446), .A2(n18445), .A3(n18444), .A4(n18443), .ZN(
        n18447) );
  NAND2_X1 U22491 ( .A1(n18451), .A2(n29837), .ZN(n18531) );
  AOI22_X1 U22492 ( .A1(n29786), .A2(\xmem_data[32][5] ), .B1(n29785), .B2(
        \xmem_data[33][5] ), .ZN(n18455) );
  AOI22_X1 U22493 ( .A1(n29787), .A2(\xmem_data[34][5] ), .B1(n22728), .B2(
        \xmem_data[35][5] ), .ZN(n18454) );
  AOI22_X1 U22494 ( .A1(n29626), .A2(\xmem_data[36][5] ), .B1(n30100), .B2(
        \xmem_data[37][5] ), .ZN(n18453) );
  AOI22_X1 U22495 ( .A1(n30279), .A2(\xmem_data[38][5] ), .B1(n29789), .B2(
        \xmem_data[39][5] ), .ZN(n18452) );
  AOI22_X1 U22496 ( .A1(n29384), .A2(\xmem_data[62][5] ), .B1(n28467), .B2(
        \xmem_data[63][5] ), .ZN(n18460) );
  AOI22_X1 U22497 ( .A1(n3226), .A2(\xmem_data[58][5] ), .B1(n29379), .B2(
        \xmem_data[59][5] ), .ZN(n18457) );
  AOI22_X1 U22498 ( .A1(n29777), .A2(\xmem_data[60][5] ), .B1(n29776), .B2(
        \xmem_data[61][5] ), .ZN(n18456) );
  NAND2_X1 U22499 ( .A1(n18457), .A2(n18456), .ZN(n18458) );
  AOI21_X1 U22500 ( .B1(n3249), .B2(\xmem_data[44][5] ), .A(n18458), .ZN(
        n18459) );
  AND2_X1 U22501 ( .A1(n18460), .A2(n18459), .ZN(n18463) );
  AOI22_X1 U22502 ( .A1(n3167), .A2(\xmem_data[52][5] ), .B1(n3186), .B2(
        \xmem_data[53][5] ), .ZN(n18462) );
  AOI22_X1 U22503 ( .A1(n30302), .A2(\xmem_data[48][5] ), .B1(n30301), .B2(
        \xmem_data[49][5] ), .ZN(n18461) );
  NAND4_X1 U22504 ( .A1(n3859), .A2(n18463), .A3(n18462), .A4(n18461), .ZN(
        n18479) );
  AOI22_X1 U22505 ( .A1(n29771), .A2(\xmem_data[50][5] ), .B1(n25607), .B2(
        \xmem_data[51][5] ), .ZN(n18466) );
  AOI21_X1 U22506 ( .B1(n30198), .B2(\xmem_data[56][5] ), .A(n18464), .ZN(
        n18465) );
  AND2_X1 U22507 ( .A1(n18466), .A2(n18465), .ZN(n18472) );
  AOI22_X1 U22508 ( .A1(n29763), .A2(\xmem_data[46][5] ), .B1(n25424), .B2(
        \xmem_data[47][5] ), .ZN(n18467) );
  INV_X1 U22509 ( .A(n18467), .ZN(n18468) );
  AOI21_X1 U22510 ( .B1(\xmem_data[57][5] ), .B2(n30765), .A(n18468), .ZN(
        n18471) );
  NAND2_X1 U22511 ( .A1(n30310), .A2(\xmem_data[54][5] ), .ZN(n18470) );
  NAND2_X1 U22512 ( .A1(n30217), .A2(\xmem_data[41][5] ), .ZN(n18469) );
  NAND4_X1 U22513 ( .A1(n18472), .A2(n18471), .A3(n18470), .A4(n18469), .ZN(
        n18477) );
  AOI22_X1 U22514 ( .A1(n29707), .A2(\xmem_data[42][5] ), .B1(n29762), .B2(
        \xmem_data[43][5] ), .ZN(n18474) );
  NAND3_X1 U22515 ( .A1(n18475), .A2(n18474), .A3(n18473), .ZN(n18476) );
  OR2_X1 U22516 ( .A1(n18477), .A2(n18476), .ZN(n18478) );
  OAI21_X1 U22517 ( .B1(n18479), .B2(n18478), .A(n29795), .ZN(n18530) );
  AOI22_X1 U22518 ( .A1(n29829), .A2(\xmem_data[64][5] ), .B1(n29785), .B2(
        \xmem_data[65][5] ), .ZN(n18483) );
  AOI22_X1 U22519 ( .A1(n29787), .A2(\xmem_data[66][5] ), .B1(n3412), .B2(
        \xmem_data[67][5] ), .ZN(n18482) );
  AOI22_X1 U22520 ( .A1(n29788), .A2(\xmem_data[68][5] ), .B1(n26616), .B2(
        \xmem_data[69][5] ), .ZN(n18481) );
  AOI22_X1 U22521 ( .A1(n30279), .A2(\xmem_data[70][5] ), .B1(n29789), .B2(
        \xmem_data[71][5] ), .ZN(n18480) );
  AOI22_X1 U22522 ( .A1(n28751), .A2(\xmem_data[80][5] ), .B1(n28778), .B2(
        \xmem_data[81][5] ), .ZN(n18488) );
  AOI22_X1 U22523 ( .A1(n29771), .A2(\xmem_data[82][5] ), .B1(n17018), .B2(
        \xmem_data[83][5] ), .ZN(n18487) );
  AOI22_X1 U22524 ( .A1(n3166), .A2(\xmem_data[84][5] ), .B1(n3185), .B2(
        \xmem_data[85][5] ), .ZN(n18486) );
  AND2_X1 U22525 ( .A1(n28781), .A2(\xmem_data[87][5] ), .ZN(n18484) );
  AOI21_X1 U22526 ( .B1(n29476), .B2(\xmem_data[86][5] ), .A(n18484), .ZN(
        n18485) );
  NAND4_X1 U22527 ( .A1(n18488), .A2(n18487), .A3(n18486), .A4(n18485), .ZN(
        n18494) );
  AOI22_X1 U22528 ( .A1(n28173), .A2(\xmem_data[88][5] ), .B1(n29640), .B2(
        \xmem_data[89][5] ), .ZN(n18492) );
  AOI22_X1 U22529 ( .A1(n3226), .A2(\xmem_data[90][5] ), .B1(n29379), .B2(
        \xmem_data[91][5] ), .ZN(n18491) );
  AOI22_X1 U22530 ( .A1(n29724), .A2(\xmem_data[92][5] ), .B1(n29723), .B2(
        \xmem_data[93][5] ), .ZN(n18490) );
  AOI22_X1 U22531 ( .A1(n29726), .A2(\xmem_data[94][5] ), .B1(n29725), .B2(
        \xmem_data[95][5] ), .ZN(n18489) );
  NAND4_X1 U22532 ( .A1(n18492), .A2(n18491), .A3(n18490), .A4(n18489), .ZN(
        n18493) );
  NOR2_X1 U22533 ( .A1(n18494), .A2(n18493), .ZN(n18503) );
  AOI22_X1 U22534 ( .A1(n30280), .A2(\xmem_data[72][5] ), .B1(n30217), .B2(
        \xmem_data[73][5] ), .ZN(n18502) );
  NAND2_X1 U22535 ( .A1(n28238), .A2(\xmem_data[77][5] ), .ZN(n18496) );
  NAND2_X1 U22536 ( .A1(n30191), .A2(\xmem_data[76][5] ), .ZN(n18495) );
  NAND2_X1 U22537 ( .A1(n18496), .A2(n18495), .ZN(n18500) );
  AOI22_X1 U22538 ( .A1(n29707), .A2(\xmem_data[74][5] ), .B1(n29706), .B2(
        \xmem_data[75][5] ), .ZN(n18498) );
  AOI22_X1 U22539 ( .A1(n29763), .A2(\xmem_data[78][5] ), .B1(n25457), .B2(
        \xmem_data[79][5] ), .ZN(n18497) );
  NAND2_X1 U22540 ( .A1(n18498), .A2(n18497), .ZN(n18499) );
  NOR2_X1 U22541 ( .A1(n18500), .A2(n18499), .ZN(n18501) );
  NAND4_X1 U22542 ( .A1(n3838), .A2(n18503), .A3(n18502), .A4(n18501), .ZN(
        n18504) );
  NAND2_X1 U22543 ( .A1(n18504), .A2(n29758), .ZN(n18529) );
  AOI22_X1 U22544 ( .A1(n28717), .A2(\xmem_data[0][5] ), .B1(n29695), .B2(
        \xmem_data[1][5] ), .ZN(n18508) );
  AOI22_X1 U22545 ( .A1(n29696), .A2(\xmem_data[2][5] ), .B1(n29661), .B2(
        \xmem_data[3][5] ), .ZN(n18507) );
  AOI22_X1 U22546 ( .A1(n30291), .A2(\xmem_data[4][5] ), .B1(n30775), .B2(
        \xmem_data[5][5] ), .ZN(n18506) );
  AOI22_X1 U22547 ( .A1(n3392), .A2(\xmem_data[6][5] ), .B1(n29698), .B2(
        \xmem_data[7][5] ), .ZN(n18505) );
  AND4_X1 U22548 ( .A1(n18508), .A2(n18507), .A3(n18506), .A4(n18505), .ZN(
        n18526) );
  AOI22_X1 U22549 ( .A1(n29390), .A2(\xmem_data[12][5] ), .B1(n30662), .B2(
        \xmem_data[13][5] ), .ZN(n18512) );
  AOI22_X1 U22550 ( .A1(n29707), .A2(\xmem_data[10][5] ), .B1(n3375), .B2(
        \xmem_data[11][5] ), .ZN(n18511) );
  AOI22_X1 U22551 ( .A1(n28787), .A2(\xmem_data[8][5] ), .B1(n29495), .B2(
        \xmem_data[9][5] ), .ZN(n18510) );
  AOI22_X1 U22552 ( .A1(n29709), .A2(\xmem_data[14][5] ), .B1(n20716), .B2(
        \xmem_data[15][5] ), .ZN(n18509) );
  AND4_X1 U22553 ( .A1(n18512), .A2(n18511), .A3(n18510), .A4(n18509), .ZN(
        n18525) );
  AOI22_X1 U22554 ( .A1(n3162), .A2(\xmem_data[20][5] ), .B1(n11426), .B2(
        \xmem_data[21][5] ), .ZN(n18517) );
  AOI22_X1 U22555 ( .A1(n29808), .A2(\xmem_data[18][5] ), .B1(n17018), .B2(
        \xmem_data[19][5] ), .ZN(n18516) );
  AOI22_X1 U22556 ( .A1(n29436), .A2(\xmem_data[16][5] ), .B1(n28778), .B2(
        \xmem_data[17][5] ), .ZN(n18515) );
  AND2_X1 U22557 ( .A1(n28781), .A2(\xmem_data[23][5] ), .ZN(n18513) );
  AOI21_X1 U22558 ( .B1(n26812), .B2(\xmem_data[22][5] ), .A(n18513), .ZN(
        n18514) );
  AND4_X1 U22559 ( .A1(n18517), .A2(n18516), .A3(n18515), .A4(n18514), .ZN(
        n18524) );
  AOI22_X1 U22560 ( .A1(n30766), .A2(\xmem_data[24][5] ), .B1(n18518), .B2(
        \xmem_data[25][5] ), .ZN(n18522) );
  AOI22_X1 U22561 ( .A1(n3226), .A2(\xmem_data[26][5] ), .B1(n29816), .B2(
        \xmem_data[27][5] ), .ZN(n18521) );
  AOI22_X1 U22562 ( .A1(n29819), .A2(\xmem_data[28][5] ), .B1(n29818), .B2(
        \xmem_data[29][5] ), .ZN(n18520) );
  AOI22_X1 U22563 ( .A1(n29821), .A2(\xmem_data[30][5] ), .B1(n29820), .B2(
        \xmem_data[31][5] ), .ZN(n18519) );
  AND4_X1 U22564 ( .A1(n18522), .A2(n18521), .A3(n18520), .A4(n18519), .ZN(
        n18523) );
  NAND4_X1 U22565 ( .A1(n18526), .A2(n18525), .A3(n18524), .A4(n18523), .ZN(
        n18527) );
  NAND2_X1 U22566 ( .A1(n18527), .A2(n29733), .ZN(n18528) );
  XNOR2_X1 U22567 ( .A(n3454), .B(\fmem_data[19][5] ), .ZN(n33218) );
  OAI22_X1 U22568 ( .A1(n22454), .A2(n34922), .B1(n33218), .B2(n34923), .ZN(
        n23601) );
  AOI22_X1 U22569 ( .A1(n30645), .A2(\xmem_data[96][5] ), .B1(n20507), .B2(
        \xmem_data[97][5] ), .ZN(n18535) );
  AOI22_X1 U22570 ( .A1(n24685), .A2(\xmem_data[98][5] ), .B1(n29136), .B2(
        \xmem_data[99][5] ), .ZN(n18534) );
  AOI22_X1 U22571 ( .A1(n24687), .A2(\xmem_data[100][5] ), .B1(n24686), .B2(
        \xmem_data[101][5] ), .ZN(n18533) );
  AOI22_X1 U22572 ( .A1(n24688), .A2(\xmem_data[102][5] ), .B1(n24470), .B2(
        \xmem_data[103][5] ), .ZN(n18532) );
  NAND4_X1 U22573 ( .A1(n18535), .A2(n18534), .A3(n18533), .A4(n18532), .ZN(
        n18551) );
  AOI22_X1 U22574 ( .A1(n24693), .A2(\xmem_data[104][5] ), .B1(n25360), .B2(
        \xmem_data[105][5] ), .ZN(n18539) );
  AOI22_X1 U22575 ( .A1(n24694), .A2(\xmem_data[106][5] ), .B1(n3219), .B2(
        \xmem_data[107][5] ), .ZN(n18538) );
  AOI22_X1 U22576 ( .A1(n24696), .A2(\xmem_data[108][5] ), .B1(n24695), .B2(
        \xmem_data[109][5] ), .ZN(n18537) );
  AOI22_X1 U22577 ( .A1(n24697), .A2(\xmem_data[110][5] ), .B1(n23811), .B2(
        \xmem_data[111][5] ), .ZN(n18536) );
  NAND4_X1 U22578 ( .A1(n18539), .A2(n18538), .A3(n18537), .A4(n18536), .ZN(
        n18550) );
  AOI22_X1 U22579 ( .A1(n24702), .A2(\xmem_data[112][5] ), .B1(n28307), .B2(
        \xmem_data[113][5] ), .ZN(n18543) );
  AOI22_X1 U22580 ( .A1(n23813), .A2(\xmem_data[114][5] ), .B1(n3358), .B2(
        \xmem_data[115][5] ), .ZN(n18542) );
  AOI22_X1 U22581 ( .A1(n28051), .A2(\xmem_data[116][5] ), .B1(n28345), .B2(
        \xmem_data[117][5] ), .ZN(n18541) );
  AOI22_X1 U22582 ( .A1(n20959), .A2(\xmem_data[118][5] ), .B1(n27536), .B2(
        \xmem_data[119][5] ), .ZN(n18540) );
  NAND4_X1 U22583 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        n18549) );
  AOI22_X1 U22584 ( .A1(n29315), .A2(\xmem_data[120][5] ), .B1(n30615), .B2(
        \xmem_data[121][5] ), .ZN(n18547) );
  AOI22_X1 U22585 ( .A1(n24708), .A2(\xmem_data[122][5] ), .B1(n24707), .B2(
        \xmem_data[123][5] ), .ZN(n18546) );
  AOI22_X1 U22586 ( .A1(n24710), .A2(\xmem_data[124][5] ), .B1(n24709), .B2(
        \xmem_data[125][5] ), .ZN(n18545) );
  AOI22_X1 U22587 ( .A1(n30956), .A2(\xmem_data[126][5] ), .B1(n25581), .B2(
        \xmem_data[127][5] ), .ZN(n18544) );
  NAND4_X1 U22588 ( .A1(n18547), .A2(n18546), .A3(n18545), .A4(n18544), .ZN(
        n18548) );
  OR4_X1 U22589 ( .A1(n18551), .A2(n18550), .A3(n18549), .A4(n18548), .ZN(
        n18573) );
  AOI22_X1 U22590 ( .A1(n24623), .A2(\xmem_data[64][5] ), .B1(n24622), .B2(
        \xmem_data[65][5] ), .ZN(n18555) );
  AOI22_X1 U22591 ( .A1(n25526), .A2(\xmem_data[66][5] ), .B1(n29247), .B2(
        \xmem_data[67][5] ), .ZN(n18554) );
  AOI22_X1 U22592 ( .A1(n17051), .A2(\xmem_data[68][5] ), .B1(n24624), .B2(
        \xmem_data[69][5] ), .ZN(n18553) );
  AOI22_X1 U22593 ( .A1(n17030), .A2(\xmem_data[70][5] ), .B1(n3203), .B2(
        \xmem_data[71][5] ), .ZN(n18552) );
  NAND4_X1 U22594 ( .A1(n18555), .A2(n18554), .A3(n18553), .A4(n18552), .ZN(
        n18571) );
  AOI22_X1 U22595 ( .A1(n24630), .A2(\xmem_data[72][5] ), .B1(n3247), .B2(
        \xmem_data[73][5] ), .ZN(n18559) );
  AOI22_X1 U22596 ( .A1(n24631), .A2(\xmem_data[74][5] ), .B1(n3222), .B2(
        \xmem_data[75][5] ), .ZN(n18558) );
  AOI22_X1 U22597 ( .A1(n24632), .A2(\xmem_data[76][5] ), .B1(n30963), .B2(
        \xmem_data[77][5] ), .ZN(n18557) );
  AOI22_X1 U22598 ( .A1(n3341), .A2(\xmem_data[78][5] ), .B1(n24633), .B2(
        \xmem_data[79][5] ), .ZN(n18556) );
  NAND4_X1 U22599 ( .A1(n18559), .A2(n18558), .A3(n18557), .A4(n18556), .ZN(
        n18570) );
  AOI22_X1 U22600 ( .A1(n3282), .A2(\xmem_data[80][5] ), .B1(n3231), .B2(
        \xmem_data[81][5] ), .ZN(n18563) );
  AOI22_X1 U22601 ( .A1(n24638), .A2(\xmem_data[82][5] ), .B1(n3358), .B2(
        \xmem_data[83][5] ), .ZN(n18562) );
  AOI22_X1 U22602 ( .A1(n24640), .A2(\xmem_data[84][5] ), .B1(n24639), .B2(
        \xmem_data[85][5] ), .ZN(n18561) );
  AOI22_X1 U22603 ( .A1(n25459), .A2(\xmem_data[86][5] ), .B1(n28517), .B2(
        \xmem_data[87][5] ), .ZN(n18560) );
  NAND4_X1 U22604 ( .A1(n18563), .A2(n18562), .A3(n18561), .A4(n18560), .ZN(
        n18569) );
  AOI22_X1 U22605 ( .A1(n25461), .A2(\xmem_data[88][5] ), .B1(n25383), .B2(
        \xmem_data[89][5] ), .ZN(n18567) );
  AOI22_X1 U22606 ( .A1(n20542), .A2(\xmem_data[90][5] ), .B1(n24645), .B2(
        \xmem_data[91][5] ), .ZN(n18566) );
  AOI22_X1 U22607 ( .A1(n14971), .A2(\xmem_data[92][5] ), .B1(n24646), .B2(
        \xmem_data[93][5] ), .ZN(n18565) );
  AOI22_X1 U22608 ( .A1(n24647), .A2(\xmem_data[94][5] ), .B1(n28462), .B2(
        \xmem_data[95][5] ), .ZN(n18564) );
  NAND4_X1 U22609 ( .A1(n18567), .A2(n18566), .A3(n18565), .A4(n18564), .ZN(
        n18568) );
  OR4_X1 U22610 ( .A1(n18571), .A2(n18570), .A3(n18569), .A4(n18568), .ZN(
        n18572) );
  AOI22_X1 U22611 ( .A1(n24722), .A2(n18573), .B1(n24720), .B2(n18572), .ZN(
        n18631) );
  AOI22_X1 U22612 ( .A1(n28233), .A2(\xmem_data[20][5] ), .B1(n13168), .B2(
        \xmem_data[21][5] ), .ZN(n18575) );
  AOI22_X1 U22613 ( .A1(n24597), .A2(\xmem_data[23][5] ), .B1(
        \xmem_data[19][5] ), .B2(n24590), .ZN(n18574) );
  NAND2_X1 U22614 ( .A1(n18575), .A2(n18574), .ZN(n18587) );
  AOI22_X1 U22615 ( .A1(n28164), .A2(\xmem_data[8][5] ), .B1(n3247), .B2(
        \xmem_data[9][5] ), .ZN(n18580) );
  AND2_X1 U22616 ( .A1(n3222), .A2(\xmem_data[11][5] ), .ZN(n18576) );
  AOI21_X1 U22617 ( .B1(n24443), .B2(\xmem_data[10][5] ), .A(n18576), .ZN(
        n18579) );
  AOI22_X1 U22618 ( .A1(n27708), .A2(\xmem_data[12][5] ), .B1(n24695), .B2(
        \xmem_data[13][5] ), .ZN(n18578) );
  AOI22_X1 U22619 ( .A1(n27904), .A2(\xmem_data[14][5] ), .B1(n30882), .B2(
        \xmem_data[15][5] ), .ZN(n18577) );
  NAND4_X1 U22620 ( .A1(n18580), .A2(n18579), .A3(n18578), .A4(n18577), .ZN(
        n18586) );
  AOI22_X1 U22621 ( .A1(n3300), .A2(\xmem_data[0][5] ), .B1(n28495), .B2(
        \xmem_data[1][5] ), .ZN(n18584) );
  AOI22_X1 U22622 ( .A1(n24606), .A2(\xmem_data[2][5] ), .B1(n28468), .B2(
        \xmem_data[3][5] ), .ZN(n18583) );
  AOI22_X1 U22623 ( .A1(n21060), .A2(\xmem_data[4][5] ), .B1(n25440), .B2(
        \xmem_data[5][5] ), .ZN(n18582) );
  AOI22_X1 U22624 ( .A1(n24607), .A2(\xmem_data[6][5] ), .B1(n20489), .B2(
        \xmem_data[7][5] ), .ZN(n18581) );
  NAND4_X1 U22625 ( .A1(n18584), .A2(n18583), .A3(n18582), .A4(n18581), .ZN(
        n18585) );
  OR3_X1 U22626 ( .A1(n18587), .A2(n18586), .A3(n18585), .ZN(n18599) );
  AOI22_X1 U22627 ( .A1(n16988), .A2(\xmem_data[24][5] ), .B1(n23716), .B2(
        \xmem_data[25][5] ), .ZN(n18591) );
  AOI22_X1 U22628 ( .A1(n24593), .A2(\xmem_data[26][5] ), .B1(n24459), .B2(
        \xmem_data[27][5] ), .ZN(n18590) );
  AOI22_X1 U22629 ( .A1(n29639), .A2(\xmem_data[28][5] ), .B1(n24592), .B2(
        \xmem_data[29][5] ), .ZN(n18589) );
  AOI22_X1 U22630 ( .A1(n3325), .A2(\xmem_data[30][5] ), .B1(n28494), .B2(
        \xmem_data[31][5] ), .ZN(n18588) );
  NAND4_X1 U22631 ( .A1(n18591), .A2(n18590), .A3(n18589), .A4(n18588), .ZN(
        n18597) );
  NAND2_X1 U22632 ( .A1(n24638), .A2(\xmem_data[18][5] ), .ZN(n18593) );
  NAND2_X1 U22633 ( .A1(n3345), .A2(\xmem_data[16][5] ), .ZN(n18592) );
  NAND2_X1 U22634 ( .A1(n18593), .A2(n18592), .ZN(n18595) );
  NOR2_X1 U22635 ( .A1(n18600), .A2(n24662), .ZN(n18629) );
  AOI22_X1 U22636 ( .A1(n30892), .A2(\xmem_data[56][5] ), .B1(n3207), .B2(
        \xmem_data[57][5] ), .ZN(n18604) );
  AOI22_X1 U22637 ( .A1(n22676), .A2(\xmem_data[58][5] ), .B1(n24645), .B2(
        \xmem_data[59][5] ), .ZN(n18603) );
  AOI22_X1 U22638 ( .A1(n29012), .A2(\xmem_data[60][5] ), .B1(n24646), .B2(
        \xmem_data[61][5] ), .ZN(n18602) );
  AOI22_X1 U22639 ( .A1(n24647), .A2(\xmem_data[62][5] ), .B1(n25581), .B2(
        \xmem_data[63][5] ), .ZN(n18601) );
  NAND4_X1 U22640 ( .A1(n18604), .A2(n18603), .A3(n18602), .A4(n18601), .ZN(
        n18611) );
  AOI22_X1 U22641 ( .A1(n24630), .A2(\xmem_data[40][5] ), .B1(n3247), .B2(
        \xmem_data[41][5] ), .ZN(n18609) );
  AND2_X1 U22642 ( .A1(n3221), .A2(\xmem_data[43][5] ), .ZN(n18605) );
  AOI21_X1 U22643 ( .B1(n24631), .B2(\xmem_data[42][5] ), .A(n18605), .ZN(
        n18608) );
  AOI22_X1 U22644 ( .A1(n24632), .A2(\xmem_data[44][5] ), .B1(n25562), .B2(
        \xmem_data[45][5] ), .ZN(n18607) );
  AOI22_X1 U22645 ( .A1(n3340), .A2(\xmem_data[46][5] ), .B1(n24633), .B2(
        \xmem_data[47][5] ), .ZN(n18606) );
  NAND4_X1 U22646 ( .A1(n18609), .A2(n18608), .A3(n18607), .A4(n18606), .ZN(
        n18610) );
  OR2_X1 U22647 ( .A1(n18611), .A2(n18610), .ZN(n18622) );
  AOI22_X1 U22648 ( .A1(n24623), .A2(\xmem_data[32][5] ), .B1(n24622), .B2(
        \xmem_data[33][5] ), .ZN(n18615) );
  AOI22_X1 U22649 ( .A1(n29325), .A2(\xmem_data[34][5] ), .B1(n25723), .B2(
        \xmem_data[35][5] ), .ZN(n18614) );
  AOI22_X1 U22650 ( .A1(n27852), .A2(\xmem_data[36][5] ), .B1(n24624), .B2(
        \xmem_data[37][5] ), .ZN(n18613) );
  AOI22_X1 U22651 ( .A1(n20827), .A2(\xmem_data[38][5] ), .B1(n3203), .B2(
        \xmem_data[39][5] ), .ZN(n18612) );
  NAND4_X1 U22652 ( .A1(n18615), .A2(n18614), .A3(n18613), .A4(n18612), .ZN(
        n18620) );
  AOI22_X1 U22653 ( .A1(n24640), .A2(\xmem_data[52][5] ), .B1(n24639), .B2(
        \xmem_data[53][5] ), .ZN(n18618) );
  AOI22_X1 U22654 ( .A1(n31268), .A2(\xmem_data[54][5] ), .B1(n20544), .B2(
        \xmem_data[55][5] ), .ZN(n18617) );
  AOI22_X1 U22655 ( .A1(n24638), .A2(\xmem_data[50][5] ), .B1(n27943), .B2(
        \xmem_data[51][5] ), .ZN(n18616) );
  NAND3_X1 U22656 ( .A1(n18618), .A2(n18617), .A3(n18616), .ZN(n18619) );
  OR2_X1 U22657 ( .A1(n18620), .A2(n18619), .ZN(n18621) );
  NOR2_X1 U22658 ( .A1(n18622), .A2(n18621), .ZN(n18625) );
  AOI22_X1 U22659 ( .A1(n3281), .A2(\xmem_data[48][5] ), .B1(n28007), .B2(
        \xmem_data[49][5] ), .ZN(n18624) );
  INV_X1 U22660 ( .A(n24659), .ZN(n18623) );
  AOI21_X1 U22661 ( .B1(n18625), .B2(n18624), .A(n18623), .ZN(n18628) );
  NOR2_X1 U22662 ( .A1(n24662), .A2(n39005), .ZN(n18626) );
  AND2_X1 U22663 ( .A1(n24657), .A2(n18626), .ZN(n18627) );
  NOR3_X1 U22664 ( .A1(n18629), .A2(n18628), .A3(n18627), .ZN(n18630) );
  AOI22_X1 U22665 ( .A1(n3270), .A2(\xmem_data[96][4] ), .B1(n29245), .B2(
        \xmem_data[97][4] ), .ZN(n18635) );
  AOI22_X1 U22666 ( .A1(n24685), .A2(\xmem_data[98][4] ), .B1(n29136), .B2(
        \xmem_data[99][4] ), .ZN(n18634) );
  AOI22_X1 U22667 ( .A1(n24687), .A2(\xmem_data[100][4] ), .B1(n24686), .B2(
        \xmem_data[101][4] ), .ZN(n18633) );
  AOI22_X1 U22668 ( .A1(n24688), .A2(\xmem_data[102][4] ), .B1(n29118), .B2(
        \xmem_data[103][4] ), .ZN(n18632) );
  NAND4_X1 U22669 ( .A1(n18635), .A2(n18634), .A3(n18633), .A4(n18632), .ZN(
        n18651) );
  AOI22_X1 U22670 ( .A1(n24693), .A2(\xmem_data[104][4] ), .B1(n25360), .B2(
        \xmem_data[105][4] ), .ZN(n18639) );
  AOI22_X1 U22671 ( .A1(n24694), .A2(\xmem_data[106][4] ), .B1(n3219), .B2(
        \xmem_data[107][4] ), .ZN(n18638) );
  AOI22_X1 U22672 ( .A1(n24696), .A2(\xmem_data[108][4] ), .B1(n24695), .B2(
        \xmem_data[109][4] ), .ZN(n18637) );
  AOI22_X1 U22673 ( .A1(n24697), .A2(\xmem_data[110][4] ), .B1(n20806), .B2(
        \xmem_data[111][4] ), .ZN(n18636) );
  NAND4_X1 U22674 ( .A1(n18639), .A2(n18638), .A3(n18637), .A4(n18636), .ZN(
        n18650) );
  AOI22_X1 U22675 ( .A1(n24702), .A2(\xmem_data[112][4] ), .B1(n29045), .B2(
        \xmem_data[113][4] ), .ZN(n18643) );
  AOI22_X1 U22676 ( .A1(n23813), .A2(\xmem_data[114][4] ), .B1(n27943), .B2(
        \xmem_data[115][4] ), .ZN(n18642) );
  AOI22_X1 U22677 ( .A1(n30886), .A2(\xmem_data[116][4] ), .B1(n29232), .B2(
        \xmem_data[117][4] ), .ZN(n18641) );
  AOI22_X1 U22678 ( .A1(n30891), .A2(\xmem_data[118][4] ), .B1(n22703), .B2(
        \xmem_data[119][4] ), .ZN(n18640) );
  NAND4_X1 U22679 ( .A1(n18643), .A2(n18642), .A3(n18641), .A4(n18640), .ZN(
        n18649) );
  AOI22_X1 U22680 ( .A1(n29237), .A2(\xmem_data[120][4] ), .B1(n27864), .B2(
        \xmem_data[121][4] ), .ZN(n18647) );
  AOI22_X1 U22681 ( .A1(n24708), .A2(\xmem_data[122][4] ), .B1(n24707), .B2(
        \xmem_data[123][4] ), .ZN(n18646) );
  AOI22_X1 U22682 ( .A1(n24710), .A2(\xmem_data[124][4] ), .B1(n24709), .B2(
        \xmem_data[125][4] ), .ZN(n18645) );
  AOI22_X1 U22683 ( .A1(n24647), .A2(\xmem_data[126][4] ), .B1(n29281), .B2(
        \xmem_data[127][4] ), .ZN(n18644) );
  NAND4_X1 U22684 ( .A1(n18647), .A2(n18646), .A3(n18645), .A4(n18644), .ZN(
        n18648) );
  OR4_X1 U22685 ( .A1(n18651), .A2(n18650), .A3(n18649), .A4(n18648), .ZN(
        n18673) );
  AOI22_X1 U22686 ( .A1(n24623), .A2(\xmem_data[64][4] ), .B1(n24622), .B2(
        \xmem_data[65][4] ), .ZN(n18655) );
  AOI22_X1 U22687 ( .A1(n20782), .A2(\xmem_data[66][4] ), .B1(n28979), .B2(
        \xmem_data[67][4] ), .ZN(n18654) );
  AOI22_X1 U22688 ( .A1(n23753), .A2(\xmem_data[68][4] ), .B1(n24624), .B2(
        \xmem_data[69][4] ), .ZN(n18653) );
  AOI22_X1 U22689 ( .A1(n20710), .A2(\xmem_data[70][4] ), .B1(n3203), .B2(
        \xmem_data[71][4] ), .ZN(n18652) );
  NAND4_X1 U22690 ( .A1(n18655), .A2(n18654), .A3(n18653), .A4(n18652), .ZN(
        n18671) );
  AOI22_X1 U22691 ( .A1(n24630), .A2(\xmem_data[72][4] ), .B1(n3247), .B2(
        \xmem_data[73][4] ), .ZN(n18659) );
  AOI22_X1 U22692 ( .A1(n24631), .A2(\xmem_data[74][4] ), .B1(n3220), .B2(
        \xmem_data[75][4] ), .ZN(n18658) );
  AOI22_X1 U22693 ( .A1(n24632), .A2(\xmem_data[76][4] ), .B1(n28319), .B2(
        \xmem_data[77][4] ), .ZN(n18657) );
  AOI22_X1 U22694 ( .A1(n3322), .A2(\xmem_data[78][4] ), .B1(n24633), .B2(
        \xmem_data[79][4] ), .ZN(n18656) );
  NAND4_X1 U22695 ( .A1(n18659), .A2(n18658), .A3(n18657), .A4(n18656), .ZN(
        n18670) );
  AOI22_X1 U22696 ( .A1(n3281), .A2(\xmem_data[80][4] ), .B1(n25514), .B2(
        \xmem_data[81][4] ), .ZN(n18663) );
  AOI22_X1 U22697 ( .A1(n24638), .A2(\xmem_data[82][4] ), .B1(n28373), .B2(
        \xmem_data[83][4] ), .ZN(n18662) );
  AOI22_X1 U22698 ( .A1(n24640), .A2(\xmem_data[84][4] ), .B1(n24639), .B2(
        \xmem_data[85][4] ), .ZN(n18661) );
  AOI22_X1 U22699 ( .A1(n20495), .A2(\xmem_data[86][4] ), .B1(n28090), .B2(
        \xmem_data[87][4] ), .ZN(n18660) );
  NAND4_X1 U22700 ( .A1(n18663), .A2(n18662), .A3(n18661), .A4(n18660), .ZN(
        n18669) );
  AOI22_X1 U22701 ( .A1(n27945), .A2(\xmem_data[88][4] ), .B1(n27989), .B2(
        \xmem_data[89][4] ), .ZN(n18667) );
  AOI22_X1 U22702 ( .A1(n24708), .A2(\xmem_data[90][4] ), .B1(n24645), .B2(
        \xmem_data[91][4] ), .ZN(n18666) );
  AOI22_X1 U22703 ( .A1(n22717), .A2(\xmem_data[92][4] ), .B1(n24646), .B2(
        \xmem_data[93][4] ), .ZN(n18665) );
  AOI22_X1 U22704 ( .A1(n24647), .A2(\xmem_data[94][4] ), .B1(n27461), .B2(
        \xmem_data[95][4] ), .ZN(n18664) );
  NAND4_X1 U22705 ( .A1(n18667), .A2(n18666), .A3(n18665), .A4(n18664), .ZN(
        n18668) );
  OR4_X1 U22706 ( .A1(n18671), .A2(n18670), .A3(n18669), .A4(n18668), .ZN(
        n18672) );
  AOI22_X1 U22707 ( .A1(n24722), .A2(n18673), .B1(n24720), .B2(n18672), .ZN(
        n18721) );
  AOI22_X1 U22708 ( .A1(n24623), .A2(\xmem_data[32][4] ), .B1(n24622), .B2(
        \xmem_data[33][4] ), .ZN(n18677) );
  AOI22_X1 U22709 ( .A1(n22684), .A2(\xmem_data[34][4] ), .B1(n11008), .B2(
        \xmem_data[35][4] ), .ZN(n18676) );
  AOI22_X1 U22710 ( .A1(n29327), .A2(\xmem_data[36][4] ), .B1(n24624), .B2(
        \xmem_data[37][4] ), .ZN(n18675) );
  AOI22_X1 U22711 ( .A1(n27436), .A2(\xmem_data[38][4] ), .B1(n3203), .B2(
        \xmem_data[39][4] ), .ZN(n18674) );
  NAND4_X1 U22712 ( .A1(n18677), .A2(n18676), .A3(n18675), .A4(n18674), .ZN(
        n18693) );
  AOI22_X1 U22713 ( .A1(n24630), .A2(\xmem_data[40][4] ), .B1(n3247), .B2(
        \xmem_data[41][4] ), .ZN(n18681) );
  AOI22_X1 U22714 ( .A1(n24631), .A2(\xmem_data[42][4] ), .B1(n3219), .B2(
        \xmem_data[43][4] ), .ZN(n18680) );
  AOI22_X1 U22715 ( .A1(n24632), .A2(\xmem_data[44][4] ), .B1(n25509), .B2(
        \xmem_data[45][4] ), .ZN(n18679) );
  AOI22_X1 U22716 ( .A1(n3342), .A2(\xmem_data[46][4] ), .B1(n24633), .B2(
        \xmem_data[47][4] ), .ZN(n18678) );
  NAND4_X1 U22717 ( .A1(n18681), .A2(n18680), .A3(n18679), .A4(n18678), .ZN(
        n18692) );
  AOI22_X1 U22718 ( .A1(n3281), .A2(\xmem_data[48][4] ), .B1(n30877), .B2(
        \xmem_data[49][4] ), .ZN(n18685) );
  AOI22_X1 U22719 ( .A1(n24638), .A2(\xmem_data[50][4] ), .B1(n28415), .B2(
        \xmem_data[51][4] ), .ZN(n18684) );
  AOI22_X1 U22720 ( .A1(n24640), .A2(\xmem_data[52][4] ), .B1(n24639), .B2(
        \xmem_data[53][4] ), .ZN(n18683) );
  AOI22_X1 U22721 ( .A1(n28298), .A2(\xmem_data[54][4] ), .B1(n20544), .B2(
        \xmem_data[55][4] ), .ZN(n18682) );
  NAND4_X1 U22722 ( .A1(n18685), .A2(n18684), .A3(n18683), .A4(n18682), .ZN(
        n18691) );
  AOI22_X1 U22723 ( .A1(n3465), .A2(\xmem_data[56][4] ), .B1(n28299), .B2(
        \xmem_data[57][4] ), .ZN(n18689) );
  AOI22_X1 U22724 ( .A1(n21007), .A2(\xmem_data[58][4] ), .B1(n24645), .B2(
        \xmem_data[59][4] ), .ZN(n18688) );
  AOI22_X1 U22725 ( .A1(n21008), .A2(\xmem_data[60][4] ), .B1(n24646), .B2(
        \xmem_data[61][4] ), .ZN(n18687) );
  AOI22_X1 U22726 ( .A1(n24647), .A2(\xmem_data[62][4] ), .B1(n29089), .B2(
        \xmem_data[63][4] ), .ZN(n18686) );
  NAND4_X1 U22727 ( .A1(n18689), .A2(n18688), .A3(n18687), .A4(n18686), .ZN(
        n18690) );
  OR4_X1 U22728 ( .A1(n18693), .A2(n18692), .A3(n18691), .A4(n18690), .ZN(
        n18694) );
  NAND2_X1 U22729 ( .A1(n18694), .A2(n24659), .ZN(n18720) );
  AOI22_X1 U22730 ( .A1(n28245), .A2(\xmem_data[8][4] ), .B1(n3247), .B2(
        \xmem_data[9][4] ), .ZN(n18699) );
  AND2_X1 U22731 ( .A1(n3219), .A2(\xmem_data[11][4] ), .ZN(n18695) );
  AOI21_X1 U22732 ( .B1(n27902), .B2(\xmem_data[10][4] ), .A(n18695), .ZN(
        n18698) );
  AOI22_X1 U22733 ( .A1(n28218), .A2(\xmem_data[12][4] ), .B1(n25491), .B2(
        \xmem_data[13][4] ), .ZN(n18697) );
  AOI22_X1 U22734 ( .A1(n29257), .A2(\xmem_data[14][4] ), .B1(n20993), .B2(
        \xmem_data[15][4] ), .ZN(n18696) );
  NAND4_X1 U22735 ( .A1(n18699), .A2(n18698), .A3(n18697), .A4(n18696), .ZN(
        n18716) );
  AOI22_X1 U22736 ( .A1(n29379), .A2(\xmem_data[0][4] ), .B1(n28495), .B2(
        \xmem_data[1][4] ), .ZN(n18703) );
  AOI22_X1 U22737 ( .A1(n24606), .A2(\xmem_data[2][4] ), .B1(n20488), .B2(
        \xmem_data[3][4] ), .ZN(n18702) );
  AOI22_X1 U22738 ( .A1(n29327), .A2(\xmem_data[4][4] ), .B1(n25440), .B2(
        \xmem_data[5][4] ), .ZN(n18701) );
  AOI22_X1 U22739 ( .A1(n24607), .A2(\xmem_data[6][4] ), .B1(n28075), .B2(
        \xmem_data[7][4] ), .ZN(n18700) );
  NAND4_X1 U22740 ( .A1(n18703), .A2(n18702), .A3(n18701), .A4(n18700), .ZN(
        n18715) );
  AOI22_X1 U22741 ( .A1(n28053), .A2(\xmem_data[24][4] ), .B1(n29279), .B2(
        \xmem_data[25][4] ), .ZN(n18707) );
  AOI22_X1 U22742 ( .A1(n24593), .A2(\xmem_data[26][4] ), .B1(n24645), .B2(
        \xmem_data[27][4] ), .ZN(n18706) );
  AOI22_X1 U22743 ( .A1(n30893), .A2(\xmem_data[28][4] ), .B1(n24592), .B2(
        \xmem_data[29][4] ), .ZN(n18705) );
  AOI22_X1 U22744 ( .A1(n24220), .A2(\xmem_data[30][4] ), .B1(n28462), .B2(
        \xmem_data[31][4] ), .ZN(n18704) );
  NAND4_X1 U22745 ( .A1(n18707), .A2(n18706), .A3(n18705), .A4(n18704), .ZN(
        n18714) );
  AOI22_X1 U22746 ( .A1(n20587), .A2(\xmem_data[20][4] ), .B1(n13168), .B2(
        \xmem_data[21][4] ), .ZN(n18710) );
  AOI22_X1 U22747 ( .A1(n16986), .A2(\xmem_data[22][4] ), .B1(n24597), .B2(
        \xmem_data[23][4] ), .ZN(n18709) );
  AOI22_X1 U22748 ( .A1(n27447), .A2(\xmem_data[18][4] ), .B1(n24590), .B2(
        \xmem_data[19][4] ), .ZN(n18708) );
  NAND3_X1 U22749 ( .A1(n18710), .A2(n18709), .A3(n18708), .ZN(n18712) );
  AND2_X1 U22750 ( .A1(n3147), .A2(\xmem_data[16][4] ), .ZN(n18711) );
  AOI21_X1 U22751 ( .B1(n25450), .B2(\xmem_data[17][4] ), .A(n18717), .ZN(
        n18718) );
  INV_X1 U22752 ( .A(n21278), .ZN(n24662) );
  OR2_X1 U22753 ( .A1(n18718), .A2(n24662), .ZN(n18719) );
  XNOR2_X1 U22754 ( .A(n32615), .B(\fmem_data[24][5] ), .ZN(n34040) );
  XOR2_X1 U22755 ( .A(\fmem_data[24][5] ), .B(\fmem_data[24][4] ), .Z(n18722)
         );
  OAI22_X1 U22756 ( .A1(n33215), .A2(n34039), .B1(n34040), .B2(n34041), .ZN(
        n23600) );
  OAI21_X1 U22757 ( .B1(n26266), .B2(n26263), .A(n26264), .ZN(n18724) );
  NAND2_X1 U22758 ( .A1(n26263), .A2(n26266), .ZN(n18723) );
  NAND2_X1 U22759 ( .A1(n18724), .A2(n18723), .ZN(n31852) );
  XNOR2_X1 U22760 ( .A(n18726), .B(n18725), .ZN(n18728) );
  XNOR2_X1 U22761 ( .A(n18727), .B(n18728), .ZN(n26262) );
  XNOR2_X1 U22762 ( .A(n35405), .B(\fmem_data[5][1] ), .ZN(n31968) );
  XNOR2_X1 U22763 ( .A(n35023), .B(\fmem_data[5][1] ), .ZN(n31886) );
  XNOR2_X1 U22764 ( .A(n31451), .B(\fmem_data[10][5] ), .ZN(n32000) );
  AOI22_X1 U22765 ( .A1(n30862), .A2(\xmem_data[24][2] ), .B1(n30861), .B2(
        \xmem_data[25][2] ), .ZN(n18732) );
  AOI22_X1 U22766 ( .A1(n30864), .A2(\xmem_data[26][2] ), .B1(n30863), .B2(
        \xmem_data[27][2] ), .ZN(n18731) );
  AOI22_X1 U22767 ( .A1(n20991), .A2(\xmem_data[28][2] ), .B1(n3220), .B2(
        \xmem_data[29][2] ), .ZN(n18730) );
  AOI22_X1 U22768 ( .A1(n25731), .A2(\xmem_data[30][2] ), .B1(n20723), .B2(
        \xmem_data[31][2] ), .ZN(n18729) );
  NAND4_X1 U22769 ( .A1(n18732), .A2(n18731), .A3(n18730), .A4(n18729), .ZN(
        n18751) );
  AOI22_X1 U22770 ( .A1(n30849), .A2(\xmem_data[16][2] ), .B1(n24117), .B2(
        \xmem_data[17][2] ), .ZN(n18736) );
  AOI22_X1 U22771 ( .A1(n24571), .A2(\xmem_data[18][2] ), .B1(n14975), .B2(
        \xmem_data[19][2] ), .ZN(n18735) );
  AOI22_X1 U22772 ( .A1(n29151), .A2(\xmem_data[20][2] ), .B1(n31256), .B2(
        \xmem_data[21][2] ), .ZN(n18734) );
  AOI22_X1 U22773 ( .A1(n28467), .A2(\xmem_data[22][2] ), .B1(n31261), .B2(
        \xmem_data[23][2] ), .ZN(n18733) );
  NAND4_X1 U22774 ( .A1(n18736), .A2(n18735), .A3(n18734), .A4(n18733), .ZN(
        n18749) );
  AOI22_X1 U22775 ( .A1(n25694), .A2(\xmem_data[0][2] ), .B1(n13444), .B2(
        \xmem_data[1][2] ), .ZN(n18738) );
  AOI22_X1 U22776 ( .A1(n28346), .A2(\xmem_data[6][2] ), .B1(n14998), .B2(
        \xmem_data[7][2] ), .ZN(n18737) );
  NAND2_X1 U22777 ( .A1(n18738), .A2(n18737), .ZN(n18742) );
  AOI22_X1 U22778 ( .A1(n23813), .A2(\xmem_data[4][2] ), .B1(n30854), .B2(
        \xmem_data[5][2] ), .ZN(n18740) );
  NAND2_X1 U22779 ( .A1(n29231), .A2(\xmem_data[2][2] ), .ZN(n18739) );
  NAND2_X1 U22780 ( .A1(n18740), .A2(n18739), .ZN(n18741) );
  OR2_X1 U22781 ( .A1(n18742), .A2(n18741), .ZN(n18748) );
  AOI22_X1 U22782 ( .A1(n16986), .A2(\xmem_data[8][2] ), .B1(n27536), .B2(
        \xmem_data[9][2] ), .ZN(n18746) );
  AOI22_X1 U22783 ( .A1(n25461), .A2(\xmem_data[10][2] ), .B1(n20586), .B2(
        \xmem_data[11][2] ), .ZN(n18745) );
  AOI22_X1 U22784 ( .A1(n23717), .A2(\xmem_data[12][2] ), .B1(n20505), .B2(
        \xmem_data[13][2] ), .ZN(n18744) );
  AOI22_X1 U22785 ( .A1(n30872), .A2(\xmem_data[14][2] ), .B1(n30871), .B2(
        \xmem_data[15][2] ), .ZN(n18743) );
  NAND4_X1 U22786 ( .A1(n18746), .A2(n18745), .A3(n18744), .A4(n18743), .ZN(
        n18747) );
  NOR2_X1 U22787 ( .A1(n18751), .A2(n18750), .ZN(n18753) );
  NAND2_X1 U22788 ( .A1(n25450), .A2(\xmem_data[3][2] ), .ZN(n18752) );
  AOI21_X1 U22789 ( .B1(n18753), .B2(n18752), .A(n30879), .ZN(n18776) );
  AOI22_X1 U22790 ( .A1(n3325), .A2(\xmem_data[48][2] ), .B1(n30898), .B2(
        \xmem_data[49][2] ), .ZN(n18757) );
  AOI22_X1 U22791 ( .A1(n3302), .A2(\xmem_data[50][2] ), .B1(n28062), .B2(
        \xmem_data[51][2] ), .ZN(n18756) );
  AOI22_X1 U22792 ( .A1(n20782), .A2(\xmem_data[52][2] ), .B1(n28328), .B2(
        \xmem_data[53][2] ), .ZN(n18755) );
  AOI22_X1 U22793 ( .A1(n30901), .A2(\xmem_data[54][2] ), .B1(n30900), .B2(
        \xmem_data[55][2] ), .ZN(n18754) );
  NAND4_X1 U22794 ( .A1(n18757), .A2(n18756), .A3(n18755), .A4(n18754), .ZN(
        n18773) );
  AOI22_X1 U22795 ( .A1(n30906), .A2(\xmem_data[60][2] ), .B1(n3222), .B2(
        \xmem_data[61][2] ), .ZN(n18761) );
  AOI22_X1 U22796 ( .A1(n3351), .A2(\xmem_data[58][2] ), .B1(n3247), .B2(
        \xmem_data[59][2] ), .ZN(n18760) );
  AOI22_X1 U22797 ( .A1(n30909), .A2(\xmem_data[56][2] ), .B1(n30908), .B2(
        \xmem_data[57][2] ), .ZN(n18759) );
  AOI22_X1 U22798 ( .A1(n30593), .A2(\xmem_data[62][2] ), .B1(n24695), .B2(
        \xmem_data[63][2] ), .ZN(n18758) );
  NAND4_X1 U22799 ( .A1(n18761), .A2(n18760), .A3(n18759), .A4(n18758), .ZN(
        n18772) );
  AOI22_X1 U22800 ( .A1(n30883), .A2(\xmem_data[32][2] ), .B1(n30882), .B2(
        \xmem_data[33][2] ), .ZN(n18765) );
  AOI22_X1 U22801 ( .A1(n25377), .A2(\xmem_data[34][2] ), .B1(n28007), .B2(
        \xmem_data[35][2] ), .ZN(n18764) );
  AOI22_X1 U22802 ( .A1(n30885), .A2(\xmem_data[36][2] ), .B1(n30884), .B2(
        \xmem_data[37][2] ), .ZN(n18763) );
  AOI22_X1 U22803 ( .A1(n30886), .A2(\xmem_data[38][2] ), .B1(n27452), .B2(
        \xmem_data[39][2] ), .ZN(n18762) );
  NAND4_X1 U22804 ( .A1(n18765), .A2(n18764), .A3(n18763), .A4(n18762), .ZN(
        n18771) );
  AOI22_X1 U22805 ( .A1(n20495), .A2(\xmem_data[40][2] ), .B1(n22703), .B2(
        \xmem_data[41][2] ), .ZN(n18769) );
  AOI22_X1 U22806 ( .A1(n25607), .A2(\xmem_data[42][2] ), .B1(n27516), .B2(
        \xmem_data[43][2] ), .ZN(n18768) );
  AOI22_X1 U22807 ( .A1(n23717), .A2(\xmem_data[44][2] ), .B1(n20940), .B2(
        \xmem_data[45][2] ), .ZN(n18767) );
  AOI22_X1 U22808 ( .A1(n30893), .A2(\xmem_data[46][2] ), .B1(n20941), .B2(
        \xmem_data[47][2] ), .ZN(n18766) );
  NAND4_X1 U22809 ( .A1(n18769), .A2(n18768), .A3(n18767), .A4(n18766), .ZN(
        n18770) );
  OR4_X1 U22810 ( .A1(n18773), .A2(n18772), .A3(n18771), .A4(n18770), .ZN(
        n18774) );
  AND2_X1 U22811 ( .A1(n18774), .A2(n30918), .ZN(n18775) );
  NOR2_X1 U22812 ( .A1(n18776), .A2(n18775), .ZN(n18820) );
  AOI22_X1 U22813 ( .A1(n17010), .A2(\xmem_data[96][2] ), .B1(n22759), .B2(
        \xmem_data[97][2] ), .ZN(n18780) );
  AOI22_X1 U22814 ( .A1(n3129), .A2(\xmem_data[98][2] ), .B1(n28307), .B2(
        \xmem_data[99][2] ), .ZN(n18779) );
  AOI22_X1 U22815 ( .A1(n27551), .A2(\xmem_data[100][2] ), .B1(n30884), .B2(
        \xmem_data[101][2] ), .ZN(n18778) );
  AOI22_X1 U22816 ( .A1(n30943), .A2(\xmem_data[102][2] ), .B1(n13168), .B2(
        \xmem_data[103][2] ), .ZN(n18777) );
  NAND4_X1 U22817 ( .A1(n18780), .A2(n18779), .A3(n18778), .A4(n18777), .ZN(
        n18796) );
  AOI22_X1 U22818 ( .A1(n27537), .A2(\xmem_data[104][2] ), .B1(n25709), .B2(
        \xmem_data[105][2] ), .ZN(n18784) );
  AOI22_X1 U22819 ( .A1(n30666), .A2(\xmem_data[106][2] ), .B1(n23716), .B2(
        \xmem_data[107][2] ), .ZN(n18783) );
  AOI22_X1 U22820 ( .A1(n30949), .A2(\xmem_data[108][2] ), .B1(n22718), .B2(
        \xmem_data[109][2] ), .ZN(n18782) );
  AOI22_X1 U22821 ( .A1(n30950), .A2(\xmem_data[110][2] ), .B1(n23776), .B2(
        \xmem_data[111][2] ), .ZN(n18781) );
  NAND4_X1 U22822 ( .A1(n18784), .A2(n18783), .A3(n18782), .A4(n18781), .ZN(
        n18795) );
  AOI22_X1 U22823 ( .A1(n30956), .A2(\xmem_data[112][2] ), .B1(n30955), .B2(
        \xmem_data[113][2] ), .ZN(n18788) );
  AOI22_X1 U22824 ( .A1(n24522), .A2(\xmem_data[114][2] ), .B1(n28983), .B2(
        \xmem_data[115][2] ), .ZN(n18787) );
  AOI22_X1 U22825 ( .A1(n25526), .A2(\xmem_data[116][2] ), .B1(n28500), .B2(
        \xmem_data[117][2] ), .ZN(n18786) );
  AOI22_X1 U22826 ( .A1(n31308), .A2(\xmem_data[118][2] ), .B1(n24122), .B2(
        \xmem_data[119][2] ), .ZN(n18785) );
  NAND4_X1 U22827 ( .A1(n18788), .A2(n18787), .A3(n18786), .A4(n18785), .ZN(
        n18794) );
  AOI22_X1 U22828 ( .A1(n25630), .A2(\xmem_data[120][2] ), .B1(n27563), .B2(
        \xmem_data[121][2] ), .ZN(n18792) );
  AOI22_X1 U22829 ( .A1(n3333), .A2(\xmem_data[122][2] ), .B1(n29173), .B2(
        \xmem_data[123][2] ), .ZN(n18791) );
  AOI22_X1 U22830 ( .A1(n30962), .A2(\xmem_data[124][2] ), .B1(n3219), .B2(
        \xmem_data[125][2] ), .ZN(n18790) );
  AOI22_X1 U22831 ( .A1(n30964), .A2(\xmem_data[126][2] ), .B1(n30963), .B2(
        \xmem_data[127][2] ), .ZN(n18789) );
  NAND4_X1 U22832 ( .A1(n18792), .A2(n18791), .A3(n18790), .A4(n18789), .ZN(
        n18793) );
  OR4_X1 U22833 ( .A1(n18796), .A2(n18795), .A3(n18794), .A4(n18793), .ZN(
        n18818) );
  AOI22_X1 U22834 ( .A1(n3322), .A2(\xmem_data[64][2] ), .B1(n21068), .B2(
        \xmem_data[65][2] ), .ZN(n18800) );
  AOI22_X1 U22835 ( .A1(n3128), .A2(\xmem_data[66][2] ), .B1(n28045), .B2(
        \xmem_data[67][2] ), .ZN(n18799) );
  AOI22_X1 U22836 ( .A1(n27551), .A2(\xmem_data[68][2] ), .B1(n27988), .B2(
        \xmem_data[69][2] ), .ZN(n18798) );
  AOI22_X1 U22837 ( .A1(n30943), .A2(\xmem_data[70][2] ), .B1(n13168), .B2(
        \xmem_data[71][2] ), .ZN(n18797) );
  NAND4_X1 U22838 ( .A1(n18800), .A2(n18799), .A3(n18798), .A4(n18797), .ZN(
        n18816) );
  AOI22_X1 U22839 ( .A1(n28298), .A2(\xmem_data[72][2] ), .B1(n29009), .B2(
        \xmem_data[73][2] ), .ZN(n18804) );
  AOI22_X1 U22840 ( .A1(n3158), .A2(\xmem_data[74][2] ), .B1(n13188), .B2(
        \xmem_data[75][2] ), .ZN(n18803) );
  AOI22_X1 U22841 ( .A1(n30949), .A2(\xmem_data[76][2] ), .B1(n17043), .B2(
        \xmem_data[77][2] ), .ZN(n18802) );
  AOI22_X1 U22842 ( .A1(n30950), .A2(\xmem_data[78][2] ), .B1(n30871), .B2(
        \xmem_data[79][2] ), .ZN(n18801) );
  NAND4_X1 U22843 ( .A1(n18804), .A2(n18803), .A3(n18802), .A4(n18801), .ZN(
        n18815) );
  AOI22_X1 U22844 ( .A1(n30956), .A2(\xmem_data[80][2] ), .B1(n30955), .B2(
        \xmem_data[81][2] ), .ZN(n18808) );
  AOI22_X1 U22845 ( .A1(n29054), .A2(\xmem_data[82][2] ), .B1(n24223), .B2(
        \xmem_data[83][2] ), .ZN(n18807) );
  AOI22_X1 U22846 ( .A1(n25582), .A2(\xmem_data[84][2] ), .B1(n28468), .B2(
        \xmem_data[85][2] ), .ZN(n18806) );
  AOI22_X1 U22847 ( .A1(n20985), .A2(\xmem_data[86][2] ), .B1(n24524), .B2(
        \xmem_data[87][2] ), .ZN(n18805) );
  NAND4_X1 U22848 ( .A1(n18808), .A2(n18807), .A3(n18806), .A4(n18805), .ZN(
        n18814) );
  AOI22_X1 U22849 ( .A1(n29124), .A2(\xmem_data[88][2] ), .B1(n27499), .B2(
        \xmem_data[89][2] ), .ZN(n18812) );
  AOI22_X1 U22850 ( .A1(n3332), .A2(\xmem_data[90][2] ), .B1(n25442), .B2(
        \xmem_data[91][2] ), .ZN(n18811) );
  AOI22_X1 U22851 ( .A1(n30962), .A2(\xmem_data[92][2] ), .B1(n3218), .B2(
        \xmem_data[93][2] ), .ZN(n18810) );
  AOI22_X1 U22852 ( .A1(n30964), .A2(\xmem_data[94][2] ), .B1(n30963), .B2(
        \xmem_data[95][2] ), .ZN(n18809) );
  NAND4_X1 U22853 ( .A1(n18812), .A2(n18811), .A3(n18810), .A4(n18809), .ZN(
        n18813) );
  OR4_X1 U22854 ( .A1(n18816), .A2(n18815), .A3(n18814), .A4(n18813), .ZN(
        n18817) );
  AOI22_X1 U22855 ( .A1(n30976), .A2(n18818), .B1(n30974), .B2(n18817), .ZN(
        n18819) );
  XNOR2_X1 U22856 ( .A(n31452), .B(\fmem_data[10][5] ), .ZN(n30800) );
  OAI22_X1 U22857 ( .A1(n32000), .A2(n35089), .B1(n30800), .B2(n35088), .ZN(
        n23590) );
  AOI22_X1 U22858 ( .A1(n25628), .A2(\xmem_data[18][1] ), .B1(n20769), .B2(
        \xmem_data[19][1] ), .ZN(n18834) );
  AOI22_X1 U22859 ( .A1(n3172), .A2(\xmem_data[16][1] ), .B1(n25359), .B2(
        \xmem_data[17][1] ), .ZN(n18821) );
  INV_X1 U22860 ( .A(n18821), .ZN(n18824) );
  AOI22_X1 U22861 ( .A1(n25624), .A2(\xmem_data[22][1] ), .B1(n30589), .B2(
        \xmem_data[23][1] ), .ZN(n18822) );
  INV_X1 U22862 ( .A(n18822), .ZN(n18823) );
  NOR2_X1 U22863 ( .A1(n18824), .A2(n18823), .ZN(n18833) );
  AOI22_X1 U22864 ( .A1(n25630), .A2(\xmem_data[20][1] ), .B1(n25629), .B2(
        \xmem_data[21][1] ), .ZN(n18832) );
  AOI22_X1 U22865 ( .A1(n25632), .A2(\xmem_data[12][1] ), .B1(n25581), .B2(
        \xmem_data[13][1] ), .ZN(n18825) );
  INV_X1 U22866 ( .A(n18825), .ZN(n18830) );
  AOI22_X1 U22867 ( .A1(n30893), .A2(\xmem_data[10][1] ), .B1(n20814), .B2(
        \xmem_data[11][1] ), .ZN(n18828) );
  AOI22_X1 U22868 ( .A1(n25635), .A2(\xmem_data[8][1] ), .B1(n20940), .B2(
        \xmem_data[9][1] ), .ZN(n18827) );
  AOI22_X1 U22869 ( .A1(n25636), .A2(\xmem_data[14][1] ), .B1(n27975), .B2(
        \xmem_data[15][1] ), .ZN(n18826) );
  NOR2_X1 U22870 ( .A1(n18830), .A2(n18829), .ZN(n18831) );
  NAND4_X1 U22871 ( .A1(n18834), .A2(n18833), .A3(n18832), .A4(n18831), .ZN(
        n18835) );
  NOR2_X1 U22872 ( .A1(n18835), .A2(n3886), .ZN(n18850) );
  AOI22_X1 U22873 ( .A1(n25612), .A2(\xmem_data[26][1] ), .B1(n29028), .B2(
        \xmem_data[27][1] ), .ZN(n18836) );
  INV_X1 U22874 ( .A(n18836), .ZN(n18842) );
  AOI22_X1 U22875 ( .A1(n25354), .A2(\xmem_data[24][1] ), .B1(n3221), .B2(
        \xmem_data[25][1] ), .ZN(n18837) );
  INV_X1 U22876 ( .A(n18837), .ZN(n18841) );
  AOI22_X1 U22877 ( .A1(n25617), .A2(\xmem_data[28][1] ), .B1(n25616), .B2(
        \xmem_data[29][1] ), .ZN(n18839) );
  NAND2_X1 U22878 ( .A1(n3375), .A2(\xmem_data[30][1] ), .ZN(n18838) );
  NAND2_X1 U22879 ( .A1(n18839), .A2(n18838), .ZN(n18840) );
  NOR3_X1 U22880 ( .A1(n18842), .A2(n18841), .A3(n18840), .ZN(n18848) );
  AOI22_X1 U22881 ( .A1(n25604), .A2(\xmem_data[0][1] ), .B1(n22739), .B2(
        \xmem_data[1][1] ), .ZN(n18846) );
  AOI22_X1 U22882 ( .A1(n28309), .A2(\xmem_data[2][1] ), .B1(n25605), .B2(
        \xmem_data[3][1] ), .ZN(n18845) );
  AOI22_X1 U22883 ( .A1(n13436), .A2(\xmem_data[4][1] ), .B1(n25606), .B2(
        \xmem_data[5][1] ), .ZN(n18844) );
  AOI22_X1 U22884 ( .A1(n30543), .A2(\xmem_data[6][1] ), .B1(n3213), .B2(
        \xmem_data[7][1] ), .ZN(n18843) );
  AND4_X1 U22885 ( .A1(n18846), .A2(n18845), .A3(n18844), .A4(n18843), .ZN(
        n18847) );
  AOI21_X1 U22886 ( .B1(n18850), .B2(n18849), .A(n25647), .ZN(n18851) );
  INV_X1 U22887 ( .A(n18851), .ZN(n18917) );
  AOI22_X1 U22888 ( .A1(n25670), .A2(\xmem_data[96][1] ), .B1(n22701), .B2(
        \xmem_data[97][1] ), .ZN(n18855) );
  AOI22_X1 U22889 ( .A1(n27453), .A2(\xmem_data[98][1] ), .B1(n20775), .B2(
        \xmem_data[99][1] ), .ZN(n18854) );
  AOI22_X1 U22890 ( .A1(n25459), .A2(\xmem_data[100][1] ), .B1(n25671), .B2(
        \xmem_data[101][1] ), .ZN(n18853) );
  AOI22_X1 U22891 ( .A1(n25672), .A2(\xmem_data[102][1] ), .B1(n3207), .B2(
        \xmem_data[103][1] ), .ZN(n18852) );
  NAND4_X1 U22892 ( .A1(n18855), .A2(n18854), .A3(n18853), .A4(n18852), .ZN(
        n18871) );
  AOI22_X1 U22893 ( .A1(n23717), .A2(\xmem_data[104][1] ), .B1(n25677), .B2(
        \xmem_data[105][1] ), .ZN(n18859) );
  AOI22_X1 U22894 ( .A1(n25678), .A2(\xmem_data[106][1] ), .B1(n25399), .B2(
        \xmem_data[107][1] ), .ZN(n18858) );
  AOI22_X1 U22895 ( .A1(n24548), .A2(\xmem_data[108][1] ), .B1(n21009), .B2(
        \xmem_data[109][1] ), .ZN(n18857) );
  AOI22_X1 U22896 ( .A1(n3269), .A2(\xmem_data[110][1] ), .B1(n28062), .B2(
        \xmem_data[111][1] ), .ZN(n18856) );
  NAND4_X1 U22897 ( .A1(n18859), .A2(n18858), .A3(n18857), .A4(n18856), .ZN(
        n18870) );
  AOI22_X1 U22898 ( .A1(n20552), .A2(\xmem_data[112][1] ), .B1(n27463), .B2(
        \xmem_data[113][1] ), .ZN(n18863) );
  AOI22_X1 U22899 ( .A1(n25684), .A2(\xmem_data[114][1] ), .B1(n30498), .B2(
        \xmem_data[115][1] ), .ZN(n18862) );
  AOI22_X1 U22900 ( .A1(n25686), .A2(\xmem_data[116][1] ), .B1(n25685), .B2(
        \xmem_data[117][1] ), .ZN(n18861) );
  AOI22_X1 U22901 ( .A1(n30864), .A2(\xmem_data[118][1] ), .B1(n25687), .B2(
        \xmem_data[119][1] ), .ZN(n18860) );
  NAND4_X1 U22902 ( .A1(n18863), .A2(n18862), .A3(n18861), .A4(n18860), .ZN(
        n18869) );
  AOI22_X1 U22903 ( .A1(n25692), .A2(\xmem_data[120][1] ), .B1(n3221), .B2(
        \xmem_data[121][1] ), .ZN(n18867) );
  AOI22_X1 U22904 ( .A1(n25693), .A2(\xmem_data[122][1] ), .B1(n28508), .B2(
        \xmem_data[123][1] ), .ZN(n18866) );
  AOI22_X1 U22905 ( .A1(n25694), .A2(\xmem_data[124][1] ), .B1(n13444), .B2(
        \xmem_data[125][1] ), .ZN(n18865) );
  AOI22_X1 U22906 ( .A1(n30710), .A2(\xmem_data[126][1] ), .B1(n30877), .B2(
        \xmem_data[127][1] ), .ZN(n18864) );
  NAND4_X1 U22907 ( .A1(n18867), .A2(n18866), .A3(n18865), .A4(n18864), .ZN(
        n18868) );
  OR4_X1 U22908 ( .A1(n18871), .A2(n18870), .A3(n18869), .A4(n18868), .ZN(
        n18893) );
  AOI22_X1 U22909 ( .A1(n25670), .A2(\xmem_data[64][1] ), .B1(n20588), .B2(
        \xmem_data[65][1] ), .ZN(n18875) );
  AOI22_X1 U22910 ( .A1(n27944), .A2(\xmem_data[66][1] ), .B1(n21015), .B2(
        \xmem_data[67][1] ), .ZN(n18874) );
  AOI22_X1 U22911 ( .A1(n29272), .A2(\xmem_data[68][1] ), .B1(n25671), .B2(
        \xmem_data[69][1] ), .ZN(n18873) );
  AOI22_X1 U22912 ( .A1(n25672), .A2(\xmem_data[70][1] ), .B1(n29188), .B2(
        \xmem_data[71][1] ), .ZN(n18872) );
  NAND4_X1 U22913 ( .A1(n18875), .A2(n18874), .A3(n18873), .A4(n18872), .ZN(
        n18891) );
  AOI22_X1 U22914 ( .A1(n24708), .A2(\xmem_data[72][1] ), .B1(n25677), .B2(
        \xmem_data[73][1] ), .ZN(n18879) );
  AOI22_X1 U22915 ( .A1(n25678), .A2(\xmem_data[74][1] ), .B1(n27460), .B2(
        \xmem_data[75][1] ), .ZN(n18878) );
  AOI22_X1 U22916 ( .A1(n29240), .A2(\xmem_data[76][1] ), .B1(n25679), .B2(
        \xmem_data[77][1] ), .ZN(n18877) );
  AOI22_X1 U22917 ( .A1(n3269), .A2(\xmem_data[78][1] ), .B1(n24622), .B2(
        \xmem_data[79][1] ), .ZN(n18876) );
  NAND4_X1 U22918 ( .A1(n18879), .A2(n18878), .A3(n18877), .A4(n18876), .ZN(
        n18890) );
  AOI22_X1 U22919 ( .A1(n3209), .A2(\xmem_data[80][1] ), .B1(n28468), .B2(
        \xmem_data[81][1] ), .ZN(n18883) );
  AOI22_X1 U22920 ( .A1(n25684), .A2(\xmem_data[82][1] ), .B1(n16999), .B2(
        \xmem_data[83][1] ), .ZN(n18882) );
  AOI22_X1 U22921 ( .A1(n25686), .A2(\xmem_data[84][1] ), .B1(n25685), .B2(
        \xmem_data[85][1] ), .ZN(n18881) );
  AOI22_X1 U22922 ( .A1(n16980), .A2(\xmem_data[86][1] ), .B1(n25687), .B2(
        \xmem_data[87][1] ), .ZN(n18880) );
  NAND4_X1 U22923 ( .A1(n18883), .A2(n18882), .A3(n18881), .A4(n18880), .ZN(
        n18889) );
  AOI22_X1 U22924 ( .A1(n25692), .A2(\xmem_data[88][1] ), .B1(n3222), .B2(
        \xmem_data[89][1] ), .ZN(n18887) );
  AOI22_X1 U22925 ( .A1(n25693), .A2(\xmem_data[90][1] ), .B1(n24695), .B2(
        \xmem_data[91][1] ), .ZN(n18886) );
  AOI22_X1 U22926 ( .A1(n25694), .A2(\xmem_data[92][1] ), .B1(n13444), .B2(
        \xmem_data[93][1] ), .ZN(n18885) );
  AOI22_X1 U22927 ( .A1(n25377), .A2(\xmem_data[94][1] ), .B1(n13474), .B2(
        \xmem_data[95][1] ), .ZN(n18884) );
  NAND4_X1 U22928 ( .A1(n18887), .A2(n18886), .A3(n18885), .A4(n18884), .ZN(
        n18888) );
  OR4_X1 U22929 ( .A1(n18891), .A2(n18890), .A3(n18889), .A4(n18888), .ZN(
        n18892) );
  AOI22_X1 U22930 ( .A1(n25706), .A2(n18893), .B1(n25704), .B2(n18892), .ZN(
        n18916) );
  AOI22_X1 U22931 ( .A1(n25707), .A2(\xmem_data[32][1] ), .B1(n27943), .B2(
        \xmem_data[33][1] ), .ZN(n18897) );
  AOI22_X1 U22932 ( .A1(n25708), .A2(\xmem_data[34][1] ), .B1(n25423), .B2(
        \xmem_data[35][1] ), .ZN(n18896) );
  AOI22_X1 U22933 ( .A1(n28980), .A2(\xmem_data[36][1] ), .B1(n25709), .B2(
        \xmem_data[37][1] ), .ZN(n18895) );
  AOI22_X1 U22934 ( .A1(n29237), .A2(\xmem_data[38][1] ), .B1(n23716), .B2(
        \xmem_data[39][1] ), .ZN(n18894) );
  NAND4_X1 U22935 ( .A1(n18897), .A2(n18896), .A3(n18895), .A4(n18894), .ZN(
        n18913) );
  AOI22_X1 U22936 ( .A1(n25573), .A2(\xmem_data[40][1] ), .B1(n25715), .B2(
        \xmem_data[41][1] ), .ZN(n18901) );
  AOI22_X1 U22937 ( .A1(n20942), .A2(\xmem_data[42][1] ), .B1(n29190), .B2(
        \xmem_data[43][1] ), .ZN(n18900) );
  AOI22_X1 U22938 ( .A1(n28460), .A2(\xmem_data[44][1] ), .B1(n30955), .B2(
        \xmem_data[45][1] ), .ZN(n18899) );
  AOI22_X1 U22939 ( .A1(n25718), .A2(\xmem_data[46][1] ), .B1(n25583), .B2(
        \xmem_data[47][1] ), .ZN(n18898) );
  NAND4_X1 U22940 ( .A1(n18901), .A2(n18900), .A3(n18899), .A4(n18898), .ZN(
        n18912) );
  AOI22_X1 U22941 ( .A1(n20734), .A2(\xmem_data[48][1] ), .B1(n25723), .B2(
        \xmem_data[49][1] ), .ZN(n18905) );
  AOI22_X1 U22942 ( .A1(n25628), .A2(\xmem_data[50][1] ), .B1(n25528), .B2(
        \xmem_data[51][1] ), .ZN(n18904) );
  AOI22_X1 U22943 ( .A1(n25724), .A2(\xmem_data[52][1] ), .B1(n28317), .B2(
        \xmem_data[53][1] ), .ZN(n18903) );
  AOI22_X1 U22944 ( .A1(n25725), .A2(\xmem_data[54][1] ), .B1(n25360), .B2(
        \xmem_data[55][1] ), .ZN(n18902) );
  NAND4_X1 U22945 ( .A1(n18905), .A2(n18904), .A3(n18903), .A4(n18902), .ZN(
        n18911) );
  AOI22_X1 U22946 ( .A1(n25730), .A2(\xmem_data[56][1] ), .B1(n3222), .B2(
        \xmem_data[57][1] ), .ZN(n18909) );
  AOI22_X1 U22947 ( .A1(n25731), .A2(\xmem_data[58][1] ), .B1(n27444), .B2(
        \xmem_data[59][1] ), .ZN(n18908) );
  AOI22_X1 U22948 ( .A1(n24438), .A2(\xmem_data[60][1] ), .B1(n31275), .B2(
        \xmem_data[61][1] ), .ZN(n18907) );
  AOI22_X1 U22949 ( .A1(n25732), .A2(\xmem_data[62][1] ), .B1(n24657), .B2(
        \xmem_data[63][1] ), .ZN(n18906) );
  NAND4_X1 U22950 ( .A1(n18909), .A2(n18908), .A3(n18907), .A4(n18906), .ZN(
        n18910) );
  OR4_X1 U22951 ( .A1(n18913), .A2(n18912), .A3(n18911), .A4(n18910), .ZN(
        n18914) );
  NAND2_X1 U22952 ( .A1(n18914), .A2(n25741), .ZN(n18915) );
  AOI22_X1 U22953 ( .A1(n3171), .A2(\xmem_data[80][0] ), .B1(n28500), .B2(
        \xmem_data[81][0] ), .ZN(n18923) );
  AND2_X1 U22954 ( .A1(n27957), .A2(\xmem_data[83][0] ), .ZN(n18918) );
  AOI21_X1 U22955 ( .B1(n25684), .B2(\xmem_data[82][0] ), .A(n18918), .ZN(
        n18922) );
  AND2_X1 U22956 ( .A1(n25686), .A2(\xmem_data[84][0] ), .ZN(n18919) );
  AOI21_X1 U22957 ( .B1(n25685), .B2(\xmem_data[85][0] ), .A(n18919), .ZN(
        n18921) );
  AOI22_X1 U22958 ( .A1(n28973), .A2(\xmem_data[86][0] ), .B1(n25687), .B2(
        \xmem_data[87][0] ), .ZN(n18920) );
  NAND4_X1 U22959 ( .A1(n18923), .A2(n18922), .A3(n18921), .A4(n18920), .ZN(
        n18943) );
  AND2_X1 U22960 ( .A1(n3222), .A2(\xmem_data[89][0] ), .ZN(n18924) );
  AOI21_X1 U22961 ( .B1(n25692), .B2(\xmem_data[88][0] ), .A(n18924), .ZN(
        n18931) );
  AOI22_X1 U22962 ( .A1(n25694), .A2(\xmem_data[92][0] ), .B1(n13444), .B2(
        \xmem_data[93][0] ), .ZN(n18925) );
  INV_X1 U22963 ( .A(n18925), .ZN(n18929) );
  AOI22_X1 U22964 ( .A1(n17063), .A2(\xmem_data[94][0] ), .B1(n13474), .B2(
        \xmem_data[95][0] ), .ZN(n18927) );
  AOI22_X1 U22965 ( .A1(n25693), .A2(\xmem_data[90][0] ), .B1(n30534), .B2(
        \xmem_data[91][0] ), .ZN(n18926) );
  NAND2_X1 U22966 ( .A1(n18927), .A2(n18926), .ZN(n18928) );
  NOR2_X1 U22967 ( .A1(n18929), .A2(n18928), .ZN(n18930) );
  NAND2_X1 U22968 ( .A1(n18931), .A2(n18930), .ZN(n18942) );
  AOI22_X1 U22969 ( .A1(n25670), .A2(\xmem_data[64][0] ), .B1(n30854), .B2(
        \xmem_data[65][0] ), .ZN(n18935) );
  AOI22_X1 U22970 ( .A1(n28346), .A2(\xmem_data[66][0] ), .B1(n24555), .B2(
        \xmem_data[67][0] ), .ZN(n18934) );
  AOI22_X1 U22971 ( .A1(n25425), .A2(\xmem_data[68][0] ), .B1(n25671), .B2(
        \xmem_data[69][0] ), .ZN(n18933) );
  AOI22_X1 U22972 ( .A1(n25672), .A2(\xmem_data[70][0] ), .B1(n30542), .B2(
        \xmem_data[71][0] ), .ZN(n18932) );
  NAND4_X1 U22973 ( .A1(n18935), .A2(n18934), .A3(n18933), .A4(n18932), .ZN(
        n18941) );
  AOI22_X1 U22974 ( .A1(n20800), .A2(\xmem_data[72][0] ), .B1(n25677), .B2(
        \xmem_data[73][0] ), .ZN(n18939) );
  AOI22_X1 U22975 ( .A1(n25678), .A2(\xmem_data[74][0] ), .B1(n28097), .B2(
        \xmem_data[75][0] ), .ZN(n18938) );
  AOI22_X1 U22976 ( .A1(n24647), .A2(\xmem_data[76][0] ), .B1(n25716), .B2(
        \xmem_data[77][0] ), .ZN(n18937) );
  AOI22_X1 U22977 ( .A1(n3269), .A2(\xmem_data[78][0] ), .B1(n20949), .B2(
        \xmem_data[79][0] ), .ZN(n18936) );
  NAND4_X1 U22978 ( .A1(n18939), .A2(n18938), .A3(n18937), .A4(n18936), .ZN(
        n18940) );
  OR4_X1 U22979 ( .A1(n18943), .A2(n18942), .A3(n18941), .A4(n18940), .ZN(
        n18944) );
  NAND2_X1 U22980 ( .A1(n18944), .A2(n25704), .ZN(n19023) );
  AOI22_X1 U22981 ( .A1(n22684), .A2(\xmem_data[112][0] ), .B1(n29247), .B2(
        \xmem_data[113][0] ), .ZN(n18950) );
  AND2_X1 U22982 ( .A1(n20579), .A2(\xmem_data[115][0] ), .ZN(n18945) );
  AOI21_X1 U22983 ( .B1(n25684), .B2(\xmem_data[114][0] ), .A(n18945), .ZN(
        n18949) );
  AND2_X1 U22984 ( .A1(n25686), .A2(\xmem_data[116][0] ), .ZN(n18946) );
  AOI21_X1 U22985 ( .B1(n25685), .B2(\xmem_data[117][0] ), .A(n18946), .ZN(
        n18948) );
  AOI22_X1 U22986 ( .A1(n27813), .A2(\xmem_data[118][0] ), .B1(n25687), .B2(
        \xmem_data[119][0] ), .ZN(n18947) );
  NAND4_X1 U22987 ( .A1(n18950), .A2(n18949), .A3(n18948), .A4(n18947), .ZN(
        n18970) );
  AND2_X1 U22988 ( .A1(n3220), .A2(\xmem_data[121][0] ), .ZN(n18951) );
  AOI21_X1 U22989 ( .B1(n25692), .B2(\xmem_data[120][0] ), .A(n18951), .ZN(
        n18958) );
  AOI22_X1 U22990 ( .A1(n25694), .A2(\xmem_data[124][0] ), .B1(n13444), .B2(
        \xmem_data[125][0] ), .ZN(n18952) );
  INV_X1 U22991 ( .A(n18952), .ZN(n18956) );
  AOI22_X1 U22992 ( .A1(n25693), .A2(\xmem_data[122][0] ), .B1(n14989), .B2(
        \xmem_data[123][0] ), .ZN(n18954) );
  AOI22_X1 U22993 ( .A1(n28952), .A2(\xmem_data[126][0] ), .B1(n24553), .B2(
        \xmem_data[127][0] ), .ZN(n18953) );
  NAND2_X1 U22994 ( .A1(n18954), .A2(n18953), .ZN(n18955) );
  NOR2_X1 U22995 ( .A1(n18956), .A2(n18955), .ZN(n18957) );
  NAND2_X1 U22996 ( .A1(n18958), .A2(n18957), .ZN(n18969) );
  AOI22_X1 U22997 ( .A1(n25670), .A2(\xmem_data[96][0] ), .B1(n22739), .B2(
        \xmem_data[97][0] ), .ZN(n18962) );
  AOI22_X1 U22998 ( .A1(n29403), .A2(\xmem_data[98][0] ), .B1(n21075), .B2(
        \xmem_data[99][0] ), .ZN(n18961) );
  AOI22_X1 U22999 ( .A1(n27537), .A2(\xmem_data[100][0] ), .B1(n25671), .B2(
        \xmem_data[101][0] ), .ZN(n18960) );
  AOI22_X1 U23000 ( .A1(n25672), .A2(\xmem_data[102][0] ), .B1(n27516), .B2(
        \xmem_data[103][0] ), .ZN(n18959) );
  NAND4_X1 U23001 ( .A1(n18962), .A2(n18961), .A3(n18960), .A4(n18959), .ZN(
        n18968) );
  AOI22_X1 U23002 ( .A1(n27919), .A2(\xmem_data[104][0] ), .B1(n25677), .B2(
        \xmem_data[105][0] ), .ZN(n18966) );
  AOI22_X1 U23003 ( .A1(n25678), .A2(\xmem_data[106][0] ), .B1(n21049), .B2(
        \xmem_data[107][0] ), .ZN(n18965) );
  AOI22_X1 U23004 ( .A1(n27462), .A2(\xmem_data[108][0] ), .B1(n25679), .B2(
        \xmem_data[109][0] ), .ZN(n18964) );
  AOI22_X1 U23005 ( .A1(n3269), .A2(\xmem_data[110][0] ), .B1(n20553), .B2(
        \xmem_data[111][0] ), .ZN(n18963) );
  NAND4_X1 U23006 ( .A1(n18966), .A2(n18965), .A3(n18964), .A4(n18963), .ZN(
        n18967) );
  OR4_X1 U23007 ( .A1(n18970), .A2(n18969), .A3(n18968), .A4(n18967), .ZN(
        n18971) );
  NAND2_X1 U23008 ( .A1(n18971), .A2(n25706), .ZN(n19022) );
  AOI22_X1 U23009 ( .A1(n3179), .A2(\xmem_data[48][0] ), .B1(n25723), .B2(
        \xmem_data[49][0] ), .ZN(n18976) );
  AND2_X1 U23010 ( .A1(n24624), .A2(\xmem_data[51][0] ), .ZN(n18972) );
  AOI21_X1 U23011 ( .B1(n30257), .B2(\xmem_data[50][0] ), .A(n18972), .ZN(
        n18975) );
  AOI22_X1 U23012 ( .A1(n25725), .A2(\xmem_data[54][0] ), .B1(n30589), .B2(
        \xmem_data[55][0] ), .ZN(n18973) );
  NAND4_X1 U23013 ( .A1(n18976), .A2(n18975), .A3(n18974), .A4(n18973), .ZN(
        n18996) );
  AND2_X1 U23014 ( .A1(n3219), .A2(\xmem_data[57][0] ), .ZN(n18977) );
  AOI21_X1 U23015 ( .B1(n25730), .B2(\xmem_data[56][0] ), .A(n18977), .ZN(
        n18984) );
  AOI22_X1 U23016 ( .A1(n27938), .A2(\xmem_data[60][0] ), .B1(n3255), .B2(
        \xmem_data[61][0] ), .ZN(n18978) );
  INV_X1 U23017 ( .A(n18978), .ZN(n18982) );
  AOI22_X1 U23018 ( .A1(n25731), .A2(\xmem_data[58][0] ), .B1(n13469), .B2(
        \xmem_data[59][0] ), .ZN(n18980) );
  AOI22_X1 U23019 ( .A1(n25732), .A2(\xmem_data[62][0] ), .B1(n13474), .B2(
        \xmem_data[63][0] ), .ZN(n18979) );
  NAND2_X1 U23020 ( .A1(n18980), .A2(n18979), .ZN(n18981) );
  NOR2_X1 U23021 ( .A1(n18982), .A2(n18981), .ZN(n18983) );
  NAND2_X1 U23022 ( .A1(n18984), .A2(n18983), .ZN(n18995) );
  AOI22_X1 U23023 ( .A1(n25707), .A2(\xmem_data[32][0] ), .B1(n25456), .B2(
        \xmem_data[33][0] ), .ZN(n18988) );
  AOI22_X1 U23024 ( .A1(n25708), .A2(\xmem_data[34][0] ), .B1(n21015), .B2(
        \xmem_data[35][0] ), .ZN(n18987) );
  AOI22_X1 U23025 ( .A1(n20541), .A2(\xmem_data[36][0] ), .B1(n25709), .B2(
        \xmem_data[37][0] ), .ZN(n18986) );
  AOI22_X1 U23026 ( .A1(n31328), .A2(\xmem_data[38][0] ), .B1(n25460), .B2(
        \xmem_data[39][0] ), .ZN(n18985) );
  NAND4_X1 U23027 ( .A1(n18988), .A2(n18987), .A3(n18986), .A4(n18985), .ZN(
        n18994) );
  AOI22_X1 U23028 ( .A1(n24133), .A2(\xmem_data[40][0] ), .B1(n25715), .B2(
        \xmem_data[41][0] ), .ZN(n18992) );
  AOI22_X1 U23029 ( .A1(n30617), .A2(\xmem_data[42][0] ), .B1(n29280), .B2(
        \xmem_data[43][0] ), .ZN(n18991) );
  AOI22_X1 U23030 ( .A1(n25717), .A2(\xmem_data[44][0] ), .B1(n28429), .B2(
        \xmem_data[45][0] ), .ZN(n18990) );
  AOI22_X1 U23031 ( .A1(n25718), .A2(\xmem_data[46][0] ), .B1(n22685), .B2(
        \xmem_data[47][0] ), .ZN(n18989) );
  NAND4_X1 U23032 ( .A1(n18992), .A2(n18991), .A3(n18990), .A4(n18989), .ZN(
        n18993) );
  OR4_X1 U23033 ( .A1(n18996), .A2(n18995), .A3(n18994), .A4(n18993), .ZN(
        n18997) );
  NAND2_X1 U23034 ( .A1(n18997), .A2(n25741), .ZN(n19021) );
  AOI22_X1 U23035 ( .A1(n20782), .A2(\xmem_data[16][0] ), .B1(n29136), .B2(
        \xmem_data[17][0] ), .ZN(n19001) );
  AOI22_X1 U23036 ( .A1(n25628), .A2(\xmem_data[18][0] ), .B1(n25528), .B2(
        \xmem_data[19][0] ), .ZN(n19000) );
  AOI22_X1 U23037 ( .A1(n25630), .A2(\xmem_data[20][0] ), .B1(n25629), .B2(
        \xmem_data[21][0] ), .ZN(n18999) );
  AOI22_X1 U23038 ( .A1(n25624), .A2(\xmem_data[22][0] ), .B1(n30589), .B2(
        \xmem_data[23][0] ), .ZN(n18998) );
  NAND4_X1 U23039 ( .A1(n19001), .A2(n19000), .A3(n18999), .A4(n18998), .ZN(
        n19017) );
  AOI22_X1 U23040 ( .A1(n30962), .A2(\xmem_data[24][0] ), .B1(n3222), .B2(
        \xmem_data[25][0] ), .ZN(n19005) );
  AOI22_X1 U23041 ( .A1(n25612), .A2(\xmem_data[26][0] ), .B1(n20723), .B2(
        \xmem_data[27][0] ), .ZN(n19004) );
  AOI22_X1 U23042 ( .A1(n25617), .A2(\xmem_data[28][0] ), .B1(n25616), .B2(
        \xmem_data[29][0] ), .ZN(n19003) );
  AOI22_X1 U23043 ( .A1(n3281), .A2(\xmem_data[30][0] ), .B1(n25514), .B2(
        \xmem_data[31][0] ), .ZN(n19002) );
  NAND4_X1 U23044 ( .A1(n19005), .A2(n19004), .A3(n19003), .A4(n19002), .ZN(
        n19016) );
  AOI22_X1 U23045 ( .A1(n25604), .A2(\xmem_data[0][0] ), .B1(n3357), .B2(
        \xmem_data[1][0] ), .ZN(n19009) );
  AOI22_X1 U23046 ( .A1(n28089), .A2(\xmem_data[2][0] ), .B1(n25605), .B2(
        \xmem_data[3][0] ), .ZN(n19008) );
  AOI22_X1 U23047 ( .A1(n29023), .A2(\xmem_data[4][0] ), .B1(n25606), .B2(
        \xmem_data[5][0] ), .ZN(n19007) );
  AOI22_X1 U23048 ( .A1(n3120), .A2(\xmem_data[6][0] ), .B1(n30615), .B2(
        \xmem_data[7][0] ), .ZN(n19006) );
  NAND4_X1 U23049 ( .A1(n19009), .A2(n19008), .A3(n19007), .A4(n19006), .ZN(
        n19015) );
  AOI22_X1 U23050 ( .A1(n25635), .A2(\xmem_data[8][0] ), .B1(n31355), .B2(
        \xmem_data[9][0] ), .ZN(n19013) );
  AOI22_X1 U23051 ( .A1(n31255), .A2(\xmem_data[10][0] ), .B1(n25367), .B2(
        \xmem_data[11][0] ), .ZN(n19012) );
  AOI22_X1 U23052 ( .A1(n25632), .A2(\xmem_data[12][0] ), .B1(n28429), .B2(
        \xmem_data[13][0] ), .ZN(n19011) );
  AOI22_X1 U23053 ( .A1(n25636), .A2(\xmem_data[14][0] ), .B1(n27975), .B2(
        \xmem_data[15][0] ), .ZN(n19010) );
  NAND4_X1 U23054 ( .A1(n19013), .A2(n19012), .A3(n19011), .A4(n19010), .ZN(
        n19014) );
  OR4_X1 U23055 ( .A1(n19017), .A2(n19016), .A3(n19015), .A4(n19014), .ZN(
        n19019) );
  NAND2_X1 U23056 ( .A1(n19019), .A2(n19018), .ZN(n19020) );
  INV_X1 U23057 ( .A(n23171), .ZN(n19509) );
  XNOR2_X1 U23058 ( .A(n32586), .B(\fmem_data[12][3] ), .ZN(n27583) );
  OAI22_X1 U23059 ( .A1(n33274), .A2(n34340), .B1(n27583), .B2(n33582), .ZN(
        n23577) );
  AOI22_X1 U23060 ( .A1(n25561), .A2(\xmem_data[32][0] ), .B1(n25725), .B2(
        \xmem_data[33][0] ), .ZN(n19028) );
  AOI22_X1 U23061 ( .A1(n25485), .A2(\xmem_data[34][0] ), .B1(n30592), .B2(
        \xmem_data[35][0] ), .ZN(n19027) );
  AOI22_X1 U23062 ( .A1(n3219), .A2(\xmem_data[36][0] ), .B1(n20805), .B2(
        \xmem_data[37][0] ), .ZN(n19026) );
  AOI22_X1 U23063 ( .A1(n25562), .A2(\xmem_data[38][0] ), .B1(n3341), .B2(
        \xmem_data[39][0] ), .ZN(n19025) );
  NAND4_X1 U23064 ( .A1(n19028), .A2(n19027), .A3(n19026), .A4(n19025), .ZN(
        n19046) );
  AOI22_X1 U23065 ( .A1(n3372), .A2(\xmem_data[56][0] ), .B1(n24522), .B2(
        \xmem_data[57][0] ), .ZN(n19033) );
  AOI22_X1 U23066 ( .A1(n25583), .A2(\xmem_data[58][0] ), .B1(n25582), .B2(
        \xmem_data[59][0] ), .ZN(n19032) );
  AND2_X1 U23067 ( .A1(n30496), .A2(\xmem_data[60][0] ), .ZN(n19029) );
  AOI21_X1 U23068 ( .B1(n25584), .B2(\xmem_data[61][0] ), .A(n19029), .ZN(
        n19031) );
  AOI22_X1 U23069 ( .A1(n20769), .A2(\xmem_data[62][0] ), .B1(n24607), .B2(
        \xmem_data[63][0] ), .ZN(n19030) );
  NAND4_X1 U23070 ( .A1(n19033), .A2(n19032), .A3(n19031), .A4(n19030), .ZN(
        n19044) );
  AOI22_X1 U23071 ( .A1(n25572), .A2(\xmem_data[48][0] ), .B1(n25519), .B2(
        \xmem_data[49][0] ), .ZN(n19037) );
  AOI22_X1 U23072 ( .A1(n25574), .A2(\xmem_data[50][0] ), .B1(n25573), .B2(
        \xmem_data[51][0] ), .ZN(n19036) );
  AOI22_X1 U23073 ( .A1(n20940), .A2(\xmem_data[52][0] ), .B1(n30617), .B2(
        \xmem_data[53][0] ), .ZN(n19035) );
  AOI22_X1 U23074 ( .A1(n25576), .A2(\xmem_data[54][0] ), .B1(n25575), .B2(
        \xmem_data[55][0] ), .ZN(n19034) );
  NAND4_X1 U23075 ( .A1(n19037), .A2(n19036), .A3(n19035), .A4(n19034), .ZN(
        n19043) );
  AOI22_X1 U23076 ( .A1(n25486), .A2(\xmem_data[40][0] ), .B1(n3146), .B2(
        \xmem_data[41][0] ), .ZN(n19041) );
  AOI22_X1 U23077 ( .A1(n25514), .A2(\xmem_data[42][0] ), .B1(n24638), .B2(
        \xmem_data[43][0] ), .ZN(n19040) );
  AOI22_X1 U23078 ( .A1(n13475), .A2(\xmem_data[44][0] ), .B1(n23762), .B2(
        \xmem_data[45][0] ), .ZN(n19039) );
  AOI22_X1 U23079 ( .A1(n24212), .A2(\xmem_data[46][0] ), .B1(n25567), .B2(
        \xmem_data[47][0] ), .ZN(n19038) );
  NAND4_X1 U23080 ( .A1(n19041), .A2(n19040), .A3(n19039), .A4(n19038), .ZN(
        n19042) );
  OR3_X1 U23081 ( .A1(n19044), .A2(n19043), .A3(n19042), .ZN(n19045) );
  OAI21_X1 U23082 ( .B1(n19046), .B2(n19045), .A(n25593), .ZN(n19115) );
  AOI22_X1 U23083 ( .A1(n29118), .A2(\xmem_data[64][0] ), .B1(n24630), .B2(
        \xmem_data[65][0] ), .ZN(n19050) );
  AOI22_X1 U23084 ( .A1(n25360), .A2(\xmem_data[66][0] ), .B1(n25508), .B2(
        \xmem_data[67][0] ), .ZN(n19049) );
  AOI22_X1 U23085 ( .A1(n3221), .A2(\xmem_data[68][0] ), .B1(n29026), .B2(
        \xmem_data[69][0] ), .ZN(n19048) );
  AOI22_X1 U23086 ( .A1(n25509), .A2(\xmem_data[70][0] ), .B1(n27904), .B2(
        \xmem_data[71][0] ), .ZN(n19047) );
  NAND4_X1 U23087 ( .A1(n19050), .A2(n19049), .A3(n19048), .A4(n19047), .ZN(
        n19068) );
  AOI22_X1 U23088 ( .A1(n28462), .A2(\xmem_data[88][0] ), .B1(n3270), .B2(
        \xmem_data[89][0] ), .ZN(n19055) );
  AOI22_X1 U23089 ( .A1(n24622), .A2(\xmem_data[90][0] ), .B1(n25526), .B2(
        \xmem_data[91][0] ), .ZN(n19054) );
  AND2_X1 U23090 ( .A1(n25527), .A2(\xmem_data[92][0] ), .ZN(n19051) );
  AOI21_X1 U23091 ( .B1(n14982), .B2(\xmem_data[93][0] ), .A(n19051), .ZN(
        n19053) );
  AOI22_X1 U23092 ( .A1(n25528), .A2(\xmem_data[94][0] ), .B1(n25441), .B2(
        \xmem_data[95][0] ), .ZN(n19052) );
  NAND4_X1 U23093 ( .A1(n19055), .A2(n19054), .A3(n19053), .A4(n19052), .ZN(
        n19066) );
  AOI22_X1 U23094 ( .A1(n25606), .A2(\xmem_data[80][0] ), .B1(n25519), .B2(
        \xmem_data[81][0] ), .ZN(n19059) );
  AOI22_X1 U23095 ( .A1(n29162), .A2(\xmem_data[82][0] ), .B1(n23717), .B2(
        \xmem_data[83][0] ), .ZN(n19058) );
  AOI22_X1 U23096 ( .A1(n25520), .A2(\xmem_data[84][0] ), .B1(n31255), .B2(
        \xmem_data[85][0] ), .ZN(n19057) );
  AOI22_X1 U23097 ( .A1(n25435), .A2(\xmem_data[86][0] ), .B1(n25521), .B2(
        \xmem_data[87][0] ), .ZN(n19056) );
  NAND4_X1 U23098 ( .A1(n19059), .A2(n19058), .A3(n19057), .A4(n19056), .ZN(
        n19065) );
  AOI22_X1 U23099 ( .A1(n29181), .A2(\xmem_data[72][0] ), .B1(n25377), .B2(
        \xmem_data[73][0] ), .ZN(n19063) );
  AOI22_X1 U23100 ( .A1(n25514), .A2(\xmem_data[74][0] ), .B1(n30551), .B2(
        \xmem_data[75][0] ), .ZN(n19062) );
  AOI22_X1 U23101 ( .A1(n3358), .A2(\xmem_data[76][0] ), .B1(n17064), .B2(
        \xmem_data[77][0] ), .ZN(n19061) );
  AOI22_X1 U23102 ( .A1(n27452), .A2(\xmem_data[78][0] ), .B1(n30891), .B2(
        \xmem_data[79][0] ), .ZN(n19060) );
  NAND4_X1 U23103 ( .A1(n19063), .A2(n19062), .A3(n19061), .A4(n19060), .ZN(
        n19064) );
  OR3_X1 U23104 ( .A1(n19066), .A2(n19065), .A3(n19064), .ZN(n19067) );
  OAI21_X1 U23105 ( .B1(n19068), .B2(n19067), .A(n25558), .ZN(n19114) );
  AOI22_X1 U23106 ( .A1(n30861), .A2(\xmem_data[96][0] ), .B1(n3333), .B2(
        \xmem_data[97][0] ), .ZN(n19072) );
  AOI22_X1 U23107 ( .A1(n25485), .A2(\xmem_data[98][0] ), .B1(n25508), .B2(
        \xmem_data[99][0] ), .ZN(n19071) );
  AOI22_X1 U23108 ( .A1(n3219), .A2(\xmem_data[100][0] ), .B1(n27445), .B2(
        \xmem_data[101][0] ), .ZN(n19070) );
  AOI22_X1 U23109 ( .A1(n25509), .A2(\xmem_data[102][0] ), .B1(n28083), .B2(
        \xmem_data[103][0] ), .ZN(n19069) );
  NAND4_X1 U23110 ( .A1(n19072), .A2(n19071), .A3(n19070), .A4(n19069), .ZN(
        n19089) );
  AOI22_X1 U23111 ( .A1(n25364), .A2(\xmem_data[120][0] ), .B1(n25718), .B2(
        \xmem_data[121][0] ), .ZN(n19076) );
  AOI22_X1 U23112 ( .A1(n24622), .A2(\xmem_data[122][0] ), .B1(n25526), .B2(
        \xmem_data[123][0] ), .ZN(n19075) );
  AOI22_X1 U23113 ( .A1(n25527), .A2(\xmem_data[124][0] ), .B1(n27852), .B2(
        \xmem_data[125][0] ), .ZN(n19074) );
  AOI22_X1 U23114 ( .A1(n25528), .A2(\xmem_data[126][0] ), .B1(n25408), .B2(
        \xmem_data[127][0] ), .ZN(n19073) );
  NAND4_X1 U23115 ( .A1(n19076), .A2(n19075), .A3(n19074), .A4(n19073), .ZN(
        n19087) );
  AOI22_X1 U23116 ( .A1(n20544), .A2(\xmem_data[112][0] ), .B1(n25519), .B2(
        \xmem_data[113][0] ), .ZN(n19080) );
  AOI22_X1 U23117 ( .A1(n27454), .A2(\xmem_data[114][0] ), .B1(n28337), .B2(
        \xmem_data[115][0] ), .ZN(n19079) );
  AOI22_X1 U23118 ( .A1(n25520), .A2(\xmem_data[116][0] ), .B1(n29047), .B2(
        \xmem_data[117][0] ), .ZN(n19078) );
  AOI22_X1 U23119 ( .A1(n29049), .A2(\xmem_data[118][0] ), .B1(n25521), .B2(
        \xmem_data[119][0] ), .ZN(n19077) );
  NAND4_X1 U23120 ( .A1(n19080), .A2(n19079), .A3(n19078), .A4(n19077), .ZN(
        n19086) );
  AOI22_X1 U23121 ( .A1(n20993), .A2(\xmem_data[104][0] ), .B1(n3131), .B2(
        \xmem_data[105][0] ), .ZN(n19084) );
  AOI22_X1 U23122 ( .A1(n25514), .A2(\xmem_data[106][0] ), .B1(n30551), .B2(
        \xmem_data[107][0] ), .ZN(n19083) );
  AOI22_X1 U23123 ( .A1(n27943), .A2(\xmem_data[108][0] ), .B1(n22738), .B2(
        \xmem_data[109][0] ), .ZN(n19082) );
  AOI22_X1 U23124 ( .A1(n13168), .A2(\xmem_data[110][0] ), .B1(n30891), .B2(
        \xmem_data[111][0] ), .ZN(n19081) );
  NAND4_X1 U23125 ( .A1(n19084), .A2(n19083), .A3(n19082), .A4(n19081), .ZN(
        n19085) );
  OR3_X1 U23126 ( .A1(n19087), .A2(n19086), .A3(n19085), .ZN(n19088) );
  OAI21_X1 U23127 ( .B1(n19089), .B2(n19088), .A(n25560), .ZN(n19113) );
  AOI22_X1 U23128 ( .A1(n25485), .A2(\xmem_data[2][0] ), .B1(n20576), .B2(
        \xmem_data[3][0] ), .ZN(n19093) );
  AOI22_X1 U23129 ( .A1(n12471), .A2(\xmem_data[0][0] ), .B1(n3229), .B2(
        \xmem_data[1][0] ), .ZN(n19092) );
  AOI22_X1 U23130 ( .A1(n3217), .A2(\xmem_data[4][0] ), .B1(n29494), .B2(
        \xmem_data[5][0] ), .ZN(n19091) );
  AOI22_X1 U23131 ( .A1(n25491), .A2(\xmem_data[6][0] ), .B1(n25490), .B2(
        \xmem_data[7][0] ), .ZN(n19090) );
  NAND4_X1 U23132 ( .A1(n19093), .A2(n19092), .A3(n19091), .A4(n19090), .ZN(
        n19109) );
  AOI22_X1 U23133 ( .A1(n25486), .A2(\xmem_data[8][0] ), .B1(n23742), .B2(
        \xmem_data[9][0] ), .ZN(n19097) );
  AOI22_X1 U23134 ( .A1(n25492), .A2(\xmem_data[10][0] ), .B1(n27447), .B2(
        \xmem_data[11][0] ), .ZN(n19096) );
  AOI22_X1 U23135 ( .A1(n25481), .A2(\xmem_data[12][0] ), .B1(n17013), .B2(
        \xmem_data[13][0] ), .ZN(n19095) );
  AOI22_X1 U23136 ( .A1(n17012), .A2(\xmem_data[14][0] ), .B1(n29272), .B2(
        \xmem_data[15][0] ), .ZN(n19094) );
  NAND4_X1 U23137 ( .A1(n19097), .A2(n19096), .A3(n19095), .A4(n19094), .ZN(
        n19108) );
  AOI22_X1 U23138 ( .A1(n25572), .A2(\xmem_data[16][0] ), .B1(n29315), .B2(
        \xmem_data[17][0] ), .ZN(n19101) );
  AOI22_X1 U23139 ( .A1(n20938), .A2(\xmem_data[18][0] ), .B1(n25635), .B2(
        \xmem_data[19][0] ), .ZN(n19100) );
  AOI22_X1 U23140 ( .A1(n16989), .A2(\xmem_data[20][0] ), .B1(n28994), .B2(
        \xmem_data[21][0] ), .ZN(n19099) );
  AOI22_X1 U23141 ( .A1(n28301), .A2(\xmem_data[22][0] ), .B1(n28385), .B2(
        \xmem_data[23][0] ), .ZN(n19098) );
  NAND4_X1 U23142 ( .A1(n19101), .A2(n19100), .A3(n19099), .A4(n19098), .ZN(
        n19107) );
  AOI22_X1 U23143 ( .A1(n25716), .A2(\xmem_data[24][0] ), .B1(n28955), .B2(
        \xmem_data[25][0] ), .ZN(n19105) );
  AOI22_X1 U23144 ( .A1(n20507), .A2(\xmem_data[26][0] ), .B1(n27847), .B2(
        \xmem_data[27][0] ), .ZN(n19104) );
  AOI22_X1 U23145 ( .A1(n20733), .A2(\xmem_data[28][0] ), .B1(n25584), .B2(
        \xmem_data[29][0] ), .ZN(n19103) );
  AOI22_X1 U23146 ( .A1(n27957), .A2(\xmem_data[30][0] ), .B1(n17056), .B2(
        \xmem_data[31][0] ), .ZN(n19102) );
  NAND4_X1 U23147 ( .A1(n19105), .A2(n19104), .A3(n19103), .A4(n19102), .ZN(
        n19106) );
  OR4_X1 U23148 ( .A1(n19109), .A2(n19108), .A3(n19107), .A4(n19106), .ZN(
        n19111) );
  XNOR2_X1 U23149 ( .A(n33751), .B(\fmem_data[17][7] ), .ZN(n19210) );
  AOI22_X1 U23150 ( .A1(n25561), .A2(\xmem_data[32][1] ), .B1(n28245), .B2(
        \xmem_data[33][1] ), .ZN(n19119) );
  AOI22_X1 U23151 ( .A1(n27437), .A2(\xmem_data[34][1] ), .B1(n30503), .B2(
        \xmem_data[35][1] ), .ZN(n19118) );
  AOI22_X1 U23152 ( .A1(n3219), .A2(\xmem_data[36][1] ), .B1(n28733), .B2(
        \xmem_data[37][1] ), .ZN(n19117) );
  AOI22_X1 U23153 ( .A1(n25562), .A2(\xmem_data[38][1] ), .B1(n3341), .B2(
        \xmem_data[39][1] ), .ZN(n19116) );
  NAND4_X1 U23154 ( .A1(n19119), .A2(n19118), .A3(n19117), .A4(n19116), .ZN(
        n19135) );
  AOI22_X1 U23155 ( .A1(n28342), .A2(\xmem_data[40][1] ), .B1(n3375), .B2(
        \xmem_data[41][1] ), .ZN(n19123) );
  AOI22_X1 U23156 ( .A1(n3231), .A2(\xmem_data[42][1] ), .B1(n25422), .B2(
        \xmem_data[43][1] ), .ZN(n19122) );
  AOI22_X1 U23157 ( .A1(n3358), .A2(\xmem_data[44][1] ), .B1(n30886), .B2(
        \xmem_data[45][1] ), .ZN(n19121) );
  AOI22_X1 U23158 ( .A1(n27452), .A2(\xmem_data[46][1] ), .B1(n25567), .B2(
        \xmem_data[47][1] ), .ZN(n19120) );
  NAND4_X1 U23159 ( .A1(n19123), .A2(n19122), .A3(n19121), .A4(n19120), .ZN(
        n19134) );
  AOI22_X1 U23160 ( .A1(n24160), .A2(\xmem_data[48][1] ), .B1(n20718), .B2(
        \xmem_data[49][1] ), .ZN(n19127) );
  AOI22_X1 U23161 ( .A1(n25574), .A2(\xmem_data[50][1] ), .B1(n25573), .B2(
        \xmem_data[51][1] ), .ZN(n19126) );
  AOI22_X1 U23162 ( .A1(n25398), .A2(\xmem_data[52][1] ), .B1(n24115), .B2(
        \xmem_data[53][1] ), .ZN(n19125) );
  AOI22_X1 U23163 ( .A1(n25576), .A2(\xmem_data[54][1] ), .B1(n25575), .B2(
        \xmem_data[55][1] ), .ZN(n19124) );
  NAND4_X1 U23164 ( .A1(n19127), .A2(n19126), .A3(n19125), .A4(n19124), .ZN(
        n19133) );
  AOI22_X1 U23165 ( .A1(n20816), .A2(\xmem_data[56][1] ), .B1(n28955), .B2(
        \xmem_data[57][1] ), .ZN(n19131) );
  AOI22_X1 U23166 ( .A1(n25583), .A2(\xmem_data[58][1] ), .B1(n25582), .B2(
        \xmem_data[59][1] ), .ZN(n19130) );
  AOI22_X1 U23167 ( .A1(n28500), .A2(\xmem_data[60][1] ), .B1(n25584), .B2(
        \xmem_data[61][1] ), .ZN(n19129) );
  AOI22_X1 U23168 ( .A1(n25528), .A2(\xmem_data[62][1] ), .B1(n17030), .B2(
        \xmem_data[63][1] ), .ZN(n19128) );
  NAND4_X1 U23169 ( .A1(n19131), .A2(n19130), .A3(n19129), .A4(n19128), .ZN(
        n19132) );
  OR4_X1 U23170 ( .A1(n19135), .A2(n19134), .A3(n19133), .A4(n19132), .ZN(
        n19163) );
  AOI22_X1 U23171 ( .A1(n22674), .A2(\xmem_data[16][1] ), .B1(n28336), .B2(
        \xmem_data[17][1] ), .ZN(n19139) );
  AOI22_X1 U23172 ( .A1(n3208), .A2(\xmem_data[18][1] ), .B1(n25434), .B2(
        \xmem_data[19][1] ), .ZN(n19138) );
  AOI22_X1 U23173 ( .A1(n29048), .A2(\xmem_data[20][1] ), .B1(n30950), .B2(
        \xmem_data[21][1] ), .ZN(n19137) );
  AOI22_X1 U23174 ( .A1(n29238), .A2(\xmem_data[22][1] ), .B1(n25575), .B2(
        \xmem_data[23][1] ), .ZN(n19136) );
  NAND4_X1 U23175 ( .A1(n19139), .A2(n19138), .A3(n19137), .A4(n19136), .ZN(
        n19146) );
  AOI22_X1 U23176 ( .A1(n25481), .A2(\xmem_data[12][1] ), .B1(n23792), .B2(
        \xmem_data[13][1] ), .ZN(n19140) );
  INV_X1 U23177 ( .A(n19140), .ZN(n19145) );
  AOI22_X1 U23178 ( .A1(n25486), .A2(\xmem_data[8][1] ), .B1(n3281), .B2(
        \xmem_data[9][1] ), .ZN(n19143) );
  AOI22_X1 U23179 ( .A1(n24639), .A2(\xmem_data[14][1] ), .B1(n29023), .B2(
        \xmem_data[15][1] ), .ZN(n19142) );
  NAND2_X1 U23180 ( .A1(n27551), .A2(\xmem_data[11][1] ), .ZN(n19141) );
  NAND3_X1 U23181 ( .A1(n19143), .A2(n19142), .A3(n19141), .ZN(n19144) );
  NOR2_X1 U23182 ( .A1(n19146), .A2(n3979), .ZN(n19161) );
  AOI22_X1 U23183 ( .A1(n3220), .A2(\xmem_data[4][1] ), .B1(n29698), .B2(
        \xmem_data[5][1] ), .ZN(n19149) );
  NAND2_X1 U23184 ( .A1(n25485), .A2(\xmem_data[2][1] ), .ZN(n19148) );
  AOI22_X1 U23185 ( .A1(n25491), .A2(\xmem_data[6][1] ), .B1(n25490), .B2(
        \xmem_data[7][1] ), .ZN(n19147) );
  NAND2_X1 U23186 ( .A1(n27502), .A2(\xmem_data[3][1] ), .ZN(n19151) );
  AOI22_X1 U23187 ( .A1(n29118), .A2(\xmem_data[0][1] ), .B1(n3228), .B2(
        \xmem_data[1][1] ), .ZN(n19150) );
  NAND2_X1 U23188 ( .A1(n19151), .A2(n19150), .ZN(n19159) );
  AND2_X1 U23189 ( .A1(n23781), .A2(\xmem_data[28][1] ), .ZN(n19152) );
  AOI21_X1 U23190 ( .B1(n29298), .B2(\xmem_data[29][1] ), .A(n19152), .ZN(
        n19153) );
  INV_X1 U23191 ( .A(n19153), .ZN(n19158) );
  AOI22_X1 U23192 ( .A1(n29281), .A2(\xmem_data[24][1] ), .B1(n25636), .B2(
        \xmem_data[25][1] ), .ZN(n19156) );
  AOI22_X1 U23193 ( .A1(n29125), .A2(\xmem_data[30][1] ), .B1(n17056), .B2(
        \xmem_data[31][1] ), .ZN(n19155) );
  AOI22_X1 U23194 ( .A1(n30599), .A2(\xmem_data[26][1] ), .B1(n20734), .B2(
        \xmem_data[27][1] ), .ZN(n19154) );
  NOR4_X1 U23195 ( .A1(n3988), .A2(n19159), .A3(n19158), .A4(n19157), .ZN(
        n19160) );
  AOI21_X1 U23196 ( .B1(n19161), .B2(n19160), .A(n25505), .ZN(n19162) );
  AOI21_X1 U23197 ( .B1(n19163), .B2(n25593), .A(n19162), .ZN(n19209) );
  AOI22_X1 U23198 ( .A1(n25485), .A2(\xmem_data[66][1] ), .B1(n25508), .B2(
        \xmem_data[67][1] ), .ZN(n19167) );
  AOI22_X1 U23199 ( .A1(n28075), .A2(\xmem_data[64][1] ), .B1(n20828), .B2(
        \xmem_data[65][1] ), .ZN(n19166) );
  AOI22_X1 U23200 ( .A1(n3222), .A2(\xmem_data[68][1] ), .B1(n24696), .B2(
        \xmem_data[69][1] ), .ZN(n19165) );
  AOI22_X1 U23201 ( .A1(n25509), .A2(\xmem_data[70][1] ), .B1(n24438), .B2(
        \xmem_data[71][1] ), .ZN(n19164) );
  NAND4_X1 U23202 ( .A1(n19167), .A2(n19166), .A3(n19165), .A4(n19164), .ZN(
        n19183) );
  AOI22_X1 U23203 ( .A1(n30882), .A2(\xmem_data[72][1] ), .B1(n30698), .B2(
        \xmem_data[73][1] ), .ZN(n19171) );
  AOI22_X1 U23204 ( .A1(n25514), .A2(\xmem_data[74][1] ), .B1(n27447), .B2(
        \xmem_data[75][1] ), .ZN(n19170) );
  AOI22_X1 U23205 ( .A1(n28373), .A2(\xmem_data[76][1] ), .B1(n23792), .B2(
        \xmem_data[77][1] ), .ZN(n19169) );
  AOI22_X1 U23206 ( .A1(n14998), .A2(\xmem_data[78][1] ), .B1(n30891), .B2(
        \xmem_data[79][1] ), .ZN(n19168) );
  NAND4_X1 U23207 ( .A1(n19171), .A2(n19170), .A3(n19169), .A4(n19168), .ZN(
        n19182) );
  AOI22_X1 U23208 ( .A1(n29046), .A2(\xmem_data[80][1] ), .B1(n25519), .B2(
        \xmem_data[81][1] ), .ZN(n19175) );
  AOI22_X1 U23209 ( .A1(n28335), .A2(\xmem_data[82][1] ), .B1(n23717), .B2(
        \xmem_data[83][1] ), .ZN(n19174) );
  AOI22_X1 U23210 ( .A1(n25520), .A2(\xmem_data[84][1] ), .B1(n29012), .B2(
        \xmem_data[85][1] ), .ZN(n19173) );
  AOI22_X1 U23211 ( .A1(n25435), .A2(\xmem_data[86][1] ), .B1(n25521), .B2(
        \xmem_data[87][1] ), .ZN(n19172) );
  NAND4_X1 U23212 ( .A1(n19175), .A2(n19174), .A3(n19173), .A4(n19172), .ZN(
        n19181) );
  AOI22_X1 U23213 ( .A1(n29055), .A2(\xmem_data[88][1] ), .B1(n29297), .B2(
        \xmem_data[89][1] ), .ZN(n19179) );
  AOI22_X1 U23214 ( .A1(n20507), .A2(\xmem_data[90][1] ), .B1(n25526), .B2(
        \xmem_data[91][1] ), .ZN(n19178) );
  AOI22_X1 U23215 ( .A1(n25527), .A2(\xmem_data[92][1] ), .B1(n21060), .B2(
        \xmem_data[93][1] ), .ZN(n19177) );
  AOI22_X1 U23216 ( .A1(n25528), .A2(\xmem_data[94][1] ), .B1(n21061), .B2(
        \xmem_data[95][1] ), .ZN(n19176) );
  NAND4_X1 U23217 ( .A1(n19179), .A2(n19178), .A3(n19177), .A4(n19176), .ZN(
        n19180) );
  OR4_X1 U23218 ( .A1(n19183), .A2(n19182), .A3(n19181), .A4(n19180), .ZN(
        n19185) );
  NOR2_X1 U23219 ( .A1(n25505), .A2(n39033), .ZN(n19184) );
  AOI21_X1 U23220 ( .B1(n19185), .B2(n25558), .A(n3901), .ZN(n19208) );
  AOI22_X1 U23221 ( .A1(n25561), .A2(\xmem_data[96][1] ), .B1(n28677), .B2(
        \xmem_data[97][1] ), .ZN(n19189) );
  AOI22_X1 U23222 ( .A1(n27437), .A2(\xmem_data[98][1] ), .B1(n25508), .B2(
        \xmem_data[99][1] ), .ZN(n19188) );
  AOI22_X1 U23223 ( .A1(n3220), .A2(\xmem_data[100][1] ), .B1(n25448), .B2(
        \xmem_data[101][1] ), .ZN(n19187) );
  AOI22_X1 U23224 ( .A1(n25509), .A2(\xmem_data[102][1] ), .B1(n24697), .B2(
        \xmem_data[103][1] ), .ZN(n19186) );
  NAND4_X1 U23225 ( .A1(n19189), .A2(n19188), .A3(n19187), .A4(n19186), .ZN(
        n19205) );
  AOI22_X1 U23226 ( .A1(n28372), .A2(\xmem_data[104][1] ), .B1(n3375), .B2(
        \xmem_data[105][1] ), .ZN(n19193) );
  AOI22_X1 U23227 ( .A1(n25514), .A2(\xmem_data[106][1] ), .B1(n27551), .B2(
        \xmem_data[107][1] ), .ZN(n19192) );
  AOI22_X1 U23228 ( .A1(n29307), .A2(\xmem_data[108][1] ), .B1(n29403), .B2(
        \xmem_data[109][1] ), .ZN(n19191) );
  AOI22_X1 U23229 ( .A1(n24448), .A2(\xmem_data[110][1] ), .B1(n16986), .B2(
        \xmem_data[111][1] ), .ZN(n19190) );
  NAND4_X1 U23230 ( .A1(n19193), .A2(n19192), .A3(n19191), .A4(n19190), .ZN(
        n19204) );
  AOI22_X1 U23231 ( .A1(n24597), .A2(\xmem_data[112][1] ), .B1(n25519), .B2(
        \xmem_data[113][1] ), .ZN(n19197) );
  AOI22_X1 U23232 ( .A1(n29279), .A2(\xmem_data[114][1] ), .B1(n24509), .B2(
        \xmem_data[115][1] ), .ZN(n19196) );
  AOI22_X1 U23233 ( .A1(n25520), .A2(\xmem_data[116][1] ), .B1(n21008), .B2(
        \xmem_data[117][1] ), .ZN(n19195) );
  AOI22_X1 U23234 ( .A1(n25399), .A2(\xmem_data[118][1] ), .B1(n25521), .B2(
        \xmem_data[119][1] ), .ZN(n19194) );
  NAND4_X1 U23235 ( .A1(n19197), .A2(n19196), .A3(n19195), .A4(n19194), .ZN(
        n19203) );
  AOI22_X1 U23236 ( .A1(n29055), .A2(\xmem_data[120][1] ), .B1(n30645), .B2(
        \xmem_data[121][1] ), .ZN(n19201) );
  AOI22_X1 U23237 ( .A1(n14883), .A2(\xmem_data[122][1] ), .B1(n25526), .B2(
        \xmem_data[123][1] ), .ZN(n19200) );
  AOI22_X1 U23238 ( .A1(n25527), .A2(\xmem_data[124][1] ), .B1(n24687), .B2(
        \xmem_data[125][1] ), .ZN(n19199) );
  AOI22_X1 U23239 ( .A1(n25528), .A2(\xmem_data[126][1] ), .B1(n27959), .B2(
        \xmem_data[127][1] ), .ZN(n19198) );
  NAND4_X1 U23240 ( .A1(n19201), .A2(n19200), .A3(n19199), .A4(n19198), .ZN(
        n19202) );
  OR4_X1 U23241 ( .A1(n19205), .A2(n19204), .A3(n19203), .A4(n19202), .ZN(
        n19206) );
  NAND2_X1 U23242 ( .A1(n19206), .A2(n25560), .ZN(n19207) );
  XNOR2_X1 U23243 ( .A(n33750), .B(\fmem_data[17][7] ), .ZN(n31988) );
  OAI22_X1 U23244 ( .A1(n19210), .A2(n35580), .B1(n35581), .B2(n31988), .ZN(
        n23574) );
  AOI22_X1 U23245 ( .A1(n28492), .A2(\xmem_data[96][2] ), .B1(n21050), .B2(
        \xmem_data[97][2] ), .ZN(n19214) );
  AOI22_X1 U23246 ( .A1(n29190), .A2(\xmem_data[98][2] ), .B1(n28493), .B2(
        \xmem_data[99][2] ), .ZN(n19213) );
  AOI22_X1 U23247 ( .A1(n28494), .A2(\xmem_data[100][2] ), .B1(n29379), .B2(
        \xmem_data[101][2] ), .ZN(n19212) );
  AOI22_X1 U23248 ( .A1(n28495), .A2(\xmem_data[102][2] ), .B1(n31316), .B2(
        \xmem_data[103][2] ), .ZN(n19211) );
  NAND4_X1 U23249 ( .A1(n19214), .A2(n19213), .A3(n19212), .A4(n19211), .ZN(
        n19230) );
  AOI22_X1 U23250 ( .A1(n28500), .A2(\xmem_data[104][2] ), .B1(n30257), .B2(
        \xmem_data[105][2] ), .ZN(n19218) );
  AOI22_X1 U23251 ( .A1(n25388), .A2(\xmem_data[106][2] ), .B1(n27925), .B2(
        \xmem_data[107][2] ), .ZN(n19217) );
  AOI22_X1 U23252 ( .A1(n31309), .A2(\xmem_data[108][2] ), .B1(n3334), .B2(
        \xmem_data[109][2] ), .ZN(n19216) );
  AOI22_X1 U23253 ( .A1(n28501), .A2(\xmem_data[110][2] ), .B1(n28503), .B2(
        \xmem_data[111][2] ), .ZN(n19215) );
  NAND4_X1 U23254 ( .A1(n19218), .A2(n19217), .A3(n19216), .A4(n19215), .ZN(
        n19229) );
  AOI22_X1 U23255 ( .A1(n3221), .A2(\xmem_data[112][2] ), .B1(n28733), .B2(
        \xmem_data[113][2] ), .ZN(n19222) );
  AOI22_X1 U23256 ( .A1(n28508), .A2(\xmem_data[114][2] ), .B1(n3342), .B2(
        \xmem_data[115][2] ), .ZN(n19221) );
  AOI22_X1 U23257 ( .A1(n28509), .A2(\xmem_data[116][2] ), .B1(n3344), .B2(
        \xmem_data[117][2] ), .ZN(n19220) );
  AOI22_X1 U23258 ( .A1(n28007), .A2(\xmem_data[118][2] ), .B1(n28374), .B2(
        \xmem_data[119][2] ), .ZN(n19219) );
  NAND4_X1 U23259 ( .A1(n19222), .A2(n19221), .A3(n19220), .A4(n19219), .ZN(
        n19228) );
  AOI22_X1 U23260 ( .A1(n3357), .A2(\xmem_data[120][2] ), .B1(n27763), .B2(
        \xmem_data[121][2] ), .ZN(n19226) );
  AOI22_X1 U23261 ( .A1(n28515), .A2(\xmem_data[122][2] ), .B1(n3175), .B2(
        \xmem_data[123][2] ), .ZN(n19225) );
  AOI22_X1 U23262 ( .A1(n28517), .A2(\xmem_data[124][2] ), .B1(n29396), .B2(
        \xmem_data[125][2] ), .ZN(n19224) );
  AOI22_X1 U23263 ( .A1(n3208), .A2(\xmem_data[126][2] ), .B1(n28096), .B2(
        \xmem_data[127][2] ), .ZN(n19223) );
  NAND4_X1 U23264 ( .A1(n19226), .A2(n19225), .A3(n19224), .A4(n19223), .ZN(
        n19227) );
  OR4_X1 U23265 ( .A1(n19230), .A2(n19229), .A3(n19228), .A4(n19227), .ZN(
        n19253) );
  AOI22_X1 U23266 ( .A1(n28492), .A2(\xmem_data[64][2] ), .B1(n30950), .B2(
        \xmem_data[65][2] ), .ZN(n19234) );
  AOI22_X1 U23267 ( .A1(n24592), .A2(\xmem_data[66][2] ), .B1(n28493), .B2(
        \xmem_data[67][2] ), .ZN(n19233) );
  AOI22_X1 U23268 ( .A1(n28494), .A2(\xmem_data[68][2] ), .B1(n3269), .B2(
        \xmem_data[69][2] ), .ZN(n19232) );
  AOI22_X1 U23269 ( .A1(n28495), .A2(\xmem_data[70][2] ), .B1(n13486), .B2(
        \xmem_data[71][2] ), .ZN(n19231) );
  NAND4_X1 U23270 ( .A1(n19234), .A2(n19233), .A3(n19232), .A4(n19231), .ZN(
        n19251) );
  AOI22_X1 U23271 ( .A1(n28500), .A2(\xmem_data[72][2] ), .B1(n27568), .B2(
        \xmem_data[73][2] ), .ZN(n19239) );
  AOI22_X1 U23272 ( .A1(n25388), .A2(\xmem_data[74][2] ), .B1(n24607), .B2(
        \xmem_data[75][2] ), .ZN(n19238) );
  AOI22_X1 U23273 ( .A1(n30861), .A2(\xmem_data[76][2] ), .B1(n20828), .B2(
        \xmem_data[77][2] ), .ZN(n19237) );
  AND2_X1 U23274 ( .A1(n28501), .A2(\xmem_data[78][2] ), .ZN(n19235) );
  AOI21_X1 U23275 ( .B1(n28503), .B2(\xmem_data[79][2] ), .A(n19235), .ZN(
        n19236) );
  NAND4_X1 U23276 ( .A1(n19239), .A2(n19238), .A3(n19237), .A4(n19236), .ZN(
        n19250) );
  AOI22_X1 U23277 ( .A1(n3220), .A2(\xmem_data[80][2] ), .B1(n29494), .B2(
        \xmem_data[81][2] ), .ZN(n19243) );
  AOI22_X1 U23278 ( .A1(n28508), .A2(\xmem_data[82][2] ), .B1(n3322), .B2(
        \xmem_data[83][2] ), .ZN(n19242) );
  AOI22_X1 U23279 ( .A1(n28509), .A2(\xmem_data[84][2] ), .B1(n29762), .B2(
        \xmem_data[85][2] ), .ZN(n19241) );
  AOI22_X1 U23280 ( .A1(n25450), .A2(\xmem_data[86][2] ), .B1(n28374), .B2(
        \xmem_data[87][2] ), .ZN(n19240) );
  NAND4_X1 U23281 ( .A1(n19243), .A2(n19242), .A3(n19241), .A4(n19240), .ZN(
        n19249) );
  AOI22_X1 U23282 ( .A1(n22701), .A2(\xmem_data[88][2] ), .B1(n20799), .B2(
        \xmem_data[89][2] ), .ZN(n19247) );
  AOI22_X1 U23283 ( .A1(n28515), .A2(\xmem_data[90][2] ), .B1(n29023), .B2(
        \xmem_data[91][2] ), .ZN(n19246) );
  AOI22_X1 U23284 ( .A1(n28517), .A2(\xmem_data[92][2] ), .B1(n3465), .B2(
        \xmem_data[93][2] ), .ZN(n19245) );
  AOI22_X1 U23285 ( .A1(n3208), .A2(\xmem_data[94][2] ), .B1(n29010), .B2(
        \xmem_data[95][2] ), .ZN(n19244) );
  NAND4_X1 U23286 ( .A1(n19247), .A2(n19246), .A3(n19245), .A4(n19244), .ZN(
        n19248) );
  OR4_X1 U23287 ( .A1(n19251), .A2(n19250), .A3(n19249), .A4(n19248), .ZN(
        n19252) );
  AOI22_X1 U23288 ( .A1(n28458), .A2(n19253), .B1(n28526), .B2(n19252), .ZN(
        n19303) );
  NOR2_X1 U23289 ( .A1(n15043), .A2(n39003), .ZN(n19254) );
  NAND2_X1 U23290 ( .A1(n29103), .A2(n19254), .ZN(n19302) );
  AOI22_X1 U23291 ( .A1(n24707), .A2(\xmem_data[32][2] ), .B1(n27855), .B2(
        \xmem_data[33][2] ), .ZN(n19258) );
  AOI22_X1 U23292 ( .A1(n24592), .A2(\xmem_data[34][2] ), .B1(n29100), .B2(
        \xmem_data[35][2] ), .ZN(n19257) );
  AOI22_X1 U23293 ( .A1(n28462), .A2(\xmem_data[36][2] ), .B1(n28461), .B2(
        \xmem_data[37][2] ), .ZN(n19256) );
  AOI22_X1 U23294 ( .A1(n20949), .A2(\xmem_data[38][2] ), .B1(n20782), .B2(
        \xmem_data[39][2] ), .ZN(n19255) );
  NAND4_X1 U23295 ( .A1(n19258), .A2(n19257), .A3(n19256), .A4(n19255), .ZN(
        n19274) );
  AOI22_X1 U23296 ( .A1(n28468), .A2(\xmem_data[40][2] ), .B1(n28467), .B2(
        \xmem_data[41][2] ), .ZN(n19262) );
  AOI22_X1 U23297 ( .A1(n22727), .A2(\xmem_data[42][2] ), .B1(n28354), .B2(
        \xmem_data[43][2] ), .ZN(n19261) );
  AOI22_X1 U23298 ( .A1(n22729), .A2(\xmem_data[44][2] ), .B1(n28164), .B2(
        \xmem_data[45][2] ), .ZN(n19260) );
  AOI22_X1 U23299 ( .A1(n20711), .A2(\xmem_data[46][2] ), .B1(n28470), .B2(
        \xmem_data[47][2] ), .ZN(n19259) );
  NAND4_X1 U23300 ( .A1(n19262), .A2(n19261), .A3(n19260), .A4(n19259), .ZN(
        n19273) );
  AOI22_X1 U23301 ( .A1(n3220), .A2(\xmem_data[48][2] ), .B1(n29789), .B2(
        \xmem_data[49][2] ), .ZN(n19266) );
  AOI22_X1 U23302 ( .A1(n28476), .A2(\xmem_data[50][2] ), .B1(n28475), .B2(
        \xmem_data[51][2] ), .ZN(n19265) );
  AOI22_X1 U23303 ( .A1(n27903), .A2(\xmem_data[52][2] ), .B1(n3135), .B2(
        \xmem_data[53][2] ), .ZN(n19264) );
  AOI22_X1 U23304 ( .A1(n27547), .A2(\xmem_data[54][2] ), .B1(n27508), .B2(
        \xmem_data[55][2] ), .ZN(n19263) );
  NAND4_X1 U23305 ( .A1(n19266), .A2(n19265), .A3(n19264), .A4(n19263), .ZN(
        n19272) );
  AOI22_X1 U23306 ( .A1(n28481), .A2(\xmem_data[56][2] ), .B1(n28309), .B2(
        \xmem_data[57][2] ), .ZN(n19270) );
  AOI22_X1 U23307 ( .A1(n30552), .A2(\xmem_data[58][2] ), .B1(n17041), .B2(
        \xmem_data[59][2] ), .ZN(n19269) );
  AOI22_X1 U23308 ( .A1(n27912), .A2(\xmem_data[60][2] ), .B1(n28231), .B2(
        \xmem_data[61][2] ), .ZN(n19268) );
  AOI22_X1 U23309 ( .A1(n22742), .A2(\xmem_data[62][2] ), .B1(n27919), .B2(
        \xmem_data[63][2] ), .ZN(n19267) );
  NAND4_X1 U23310 ( .A1(n19270), .A2(n19269), .A3(n19268), .A4(n19267), .ZN(
        n19271) );
  OR4_X1 U23311 ( .A1(n19274), .A2(n19273), .A3(n19272), .A4(n19271), .ZN(
        n19300) );
  AOI22_X1 U23312 ( .A1(n29017), .A2(\xmem_data[8][2] ), .B1(n21060), .B2(
        \xmem_data[9][2] ), .ZN(n19278) );
  AOI22_X1 U23313 ( .A1(n27567), .A2(\xmem_data[10][2] ), .B1(n30862), .B2(
        \xmem_data[11][2] ), .ZN(n19277) );
  AOI22_X1 U23314 ( .A1(n31262), .A2(\xmem_data[12][2] ), .B1(n24693), .B2(
        \xmem_data[13][2] ), .ZN(n19276) );
  AOI22_X1 U23315 ( .A1(n30589), .A2(\xmem_data[14][2] ), .B1(n25508), .B2(
        \xmem_data[15][2] ), .ZN(n19275) );
  NAND4_X1 U23316 ( .A1(n19278), .A2(n19277), .A3(n19276), .A4(n19275), .ZN(
        n19297) );
  AOI22_X1 U23317 ( .A1(n28373), .A2(\xmem_data[24][2] ), .B1(n28743), .B2(
        \xmem_data[25][2] ), .ZN(n19282) );
  AOI22_X1 U23318 ( .A1(n28416), .A2(\xmem_data[26][2] ), .B1(n20959), .B2(
        \xmem_data[27][2] ), .ZN(n19281) );
  AOI22_X1 U23319 ( .A1(n20798), .A2(\xmem_data[28][2] ), .B1(n3120), .B2(
        \xmem_data[29][2] ), .ZN(n19280) );
  AOI22_X1 U23320 ( .A1(n27989), .A2(\xmem_data[30][2] ), .B1(n24593), .B2(
        \xmem_data[31][2] ), .ZN(n19279) );
  NAND4_X1 U23321 ( .A1(n19282), .A2(n19281), .A3(n19280), .A4(n19279), .ZN(
        n19296) );
  AOI22_X1 U23322 ( .A1(n24140), .A2(\xmem_data[20][2] ), .B1(n29706), .B2(
        \xmem_data[21][2] ), .ZN(n19289) );
  AOI22_X1 U23323 ( .A1(n3222), .A2(\xmem_data[16][2] ), .B1(n25612), .B2(
        \xmem_data[17][2] ), .ZN(n19283) );
  INV_X1 U23324 ( .A(n19283), .ZN(n19287) );
  AOI22_X1 U23325 ( .A1(n20992), .A2(\xmem_data[18][2] ), .B1(n14990), .B2(
        \xmem_data[19][2] ), .ZN(n19284) );
  INV_X1 U23326 ( .A(n19284), .ZN(n19286) );
  AND2_X1 U23327 ( .A1(n25422), .A2(\xmem_data[23][2] ), .ZN(n19285) );
  NOR3_X1 U23328 ( .A1(n19287), .A2(n19286), .A3(n19285), .ZN(n19288) );
  NAND2_X1 U23329 ( .A1(n19289), .A2(n19288), .ZN(n19295) );
  AOI22_X1 U23330 ( .A1(n28427), .A2(\xmem_data[0][2] ), .B1(n30950), .B2(
        \xmem_data[1][2] ), .ZN(n19293) );
  AOI22_X1 U23331 ( .A1(n24592), .A2(\xmem_data[2][2] ), .B1(n28428), .B2(
        \xmem_data[3][2] ), .ZN(n19292) );
  AOI22_X1 U23332 ( .A1(n30598), .A2(\xmem_data[4][2] ), .B1(n3329), .B2(
        \xmem_data[5][2] ), .ZN(n19291) );
  AOI22_X1 U23333 ( .A1(n20983), .A2(\xmem_data[6][2] ), .B1(n22719), .B2(
        \xmem_data[7][2] ), .ZN(n19290) );
  NAND4_X1 U23334 ( .A1(n19293), .A2(n19292), .A3(n19291), .A4(n19290), .ZN(
        n19294) );
  NOR4_X1 U23335 ( .A1(n19297), .A2(n19296), .A3(n19295), .A4(n19294), .ZN(
        n19298) );
  NOR2_X1 U23336 ( .A1(n19298), .A2(n15043), .ZN(n19299) );
  AOI21_X1 U23337 ( .B1(n19300), .B2(n28490), .A(n19299), .ZN(n19301) );
  XNOR2_X1 U23338 ( .A(n32528), .B(\fmem_data[29][5] ), .ZN(n26370) );
  OAI21_X1 U23339 ( .B1(n23577), .B2(n23574), .A(n23575), .ZN(n19305) );
  NAND2_X1 U23340 ( .A1(n19305), .A2(n19304), .ZN(n23170) );
  AOI22_X1 U23341 ( .A1(n23717), .A2(\xmem_data[22][1] ), .B1(n28492), .B2(
        \xmem_data[23][1] ), .ZN(n19307) );
  AOI22_X1 U23342 ( .A1(n27542), .A2(\xmem_data[30][1] ), .B1(n11008), .B2(
        \xmem_data[31][1] ), .ZN(n19306) );
  NAND2_X1 U23343 ( .A1(n19307), .A2(n19306), .ZN(n19312) );
  AOI22_X1 U23344 ( .A1(n23795), .A2(\xmem_data[20][1] ), .B1(n27454), .B2(
        \xmem_data[21][1] ), .ZN(n19310) );
  AOI22_X1 U23345 ( .A1(n28701), .A2(\xmem_data[28][1] ), .B1(n27365), .B2(
        \xmem_data[29][1] ), .ZN(n19309) );
  AOI22_X1 U23346 ( .A1(n27536), .A2(\xmem_data[19][1] ), .B1(n28060), .B2(
        \xmem_data[27][1] ), .ZN(n19308) );
  NAND3_X1 U23347 ( .A1(n19310), .A2(n19309), .A3(n19308), .ZN(n19311) );
  NOR2_X1 U23348 ( .A1(n19312), .A2(n19311), .ZN(n19323) );
  NAND2_X1 U23349 ( .A1(n28980), .A2(\xmem_data[18][1] ), .ZN(n19314) );
  NAND2_X1 U23350 ( .A1(n22683), .A2(\xmem_data[26][1] ), .ZN(n19313) );
  NAND2_X1 U23351 ( .A1(n19314), .A2(n19313), .ZN(n19318) );
  AOI22_X1 U23352 ( .A1(n24640), .A2(\xmem_data[16][1] ), .B1(n27535), .B2(
        \xmem_data[17][1] ), .ZN(n19316) );
  AOI22_X1 U23353 ( .A1(n20730), .A2(\xmem_data[24][1] ), .B1(n13452), .B2(
        \xmem_data[25][1] ), .ZN(n19315) );
  AOI22_X1 U23354 ( .A1(n29494), .A2(\xmem_data[8][1] ), .B1(n25562), .B2(
        \xmem_data[9][1] ), .ZN(n19321) );
  AOI22_X1 U23355 ( .A1(n27551), .A2(\xmem_data[14][1] ), .B1(n28373), .B2(
        \xmem_data[15][1] ), .ZN(n19320) );
  AOI22_X1 U23356 ( .A1(n24697), .A2(\xmem_data[10][1] ), .B1(n27550), .B2(
        \xmem_data[11][1] ), .ZN(n19319) );
  NAND3_X1 U23357 ( .A1(n19323), .A2(n19322), .A3(n3952), .ZN(n19329) );
  AOI22_X1 U23358 ( .A1(n27568), .A2(\xmem_data[0][1] ), .B1(n27567), .B2(
        \xmem_data[1][1] ), .ZN(n19327) );
  AOI22_X1 U23359 ( .A1(n27564), .A2(\xmem_data[2][1] ), .B1(n27563), .B2(
        \xmem_data[3][1] ), .ZN(n19326) );
  AOI22_X1 U23360 ( .A1(n3153), .A2(\xmem_data[4][1] ), .B1(n30589), .B2(
        \xmem_data[5][1] ), .ZN(n19325) );
  AOI22_X1 U23361 ( .A1(n28318), .A2(\xmem_data[6][1] ), .B1(n3221), .B2(
        \xmem_data[7][1] ), .ZN(n19324) );
  NAND4_X1 U23362 ( .A1(n19327), .A2(n19326), .A3(n19325), .A4(n19324), .ZN(
        n19328) );
  AND2_X1 U23363 ( .A1(n30295), .A2(\xmem_data[12][1] ), .ZN(n19330) );
  OR2_X1 U23364 ( .A1(n19331), .A2(n19330), .ZN(n19354) );
  AOI22_X1 U23365 ( .A1(n24687), .A2(\xmem_data[64][1] ), .B1(n27435), .B2(
        \xmem_data[65][1] ), .ZN(n19335) );
  AOI22_X1 U23366 ( .A1(n27436), .A2(\xmem_data[66][1] ), .B1(n24470), .B2(
        \xmem_data[67][1] ), .ZN(n19334) );
  AOI22_X1 U23367 ( .A1(n24693), .A2(\xmem_data[68][1] ), .B1(n27437), .B2(
        \xmem_data[69][1] ), .ZN(n19333) );
  AOI22_X1 U23368 ( .A1(n27439), .A2(\xmem_data[70][1] ), .B1(n3217), .B2(
        \xmem_data[71][1] ), .ZN(n19332) );
  NAND4_X1 U23369 ( .A1(n19335), .A2(n19334), .A3(n19333), .A4(n19332), .ZN(
        n19351) );
  AOI22_X1 U23370 ( .A1(n27445), .A2(\xmem_data[72][1] ), .B1(n27444), .B2(
        \xmem_data[73][1] ), .ZN(n19339) );
  AOI22_X1 U23371 ( .A1(n20725), .A2(\xmem_data[74][1] ), .B1(n17061), .B2(
        \xmem_data[75][1] ), .ZN(n19338) );
  AOI22_X1 U23372 ( .A1(n28344), .A2(\xmem_data[76][1] ), .B1(n27446), .B2(
        \xmem_data[77][1] ), .ZN(n19337) );
  AOI22_X1 U23373 ( .A1(n27447), .A2(\xmem_data[78][1] ), .B1(n20982), .B2(
        \xmem_data[79][1] ), .ZN(n19336) );
  NAND4_X1 U23374 ( .A1(n19339), .A2(n19338), .A3(n19337), .A4(n19336), .ZN(
        n19350) );
  AOI22_X1 U23375 ( .A1(n27453), .A2(\xmem_data[80][1] ), .B1(n27452), .B2(
        \xmem_data[81][1] ), .ZN(n19343) );
  AOI22_X1 U23376 ( .A1(n25710), .A2(\xmem_data[82][1] ), .B1(n29271), .B2(
        \xmem_data[83][1] ), .ZN(n19342) );
  AOI22_X1 U23377 ( .A1(n28752), .A2(\xmem_data[84][1] ), .B1(n27454), .B2(
        \xmem_data[85][1] ), .ZN(n19341) );
  AOI22_X1 U23378 ( .A1(n13149), .A2(\xmem_data[86][1] ), .B1(n31329), .B2(
        \xmem_data[87][1] ), .ZN(n19340) );
  NAND4_X1 U23379 ( .A1(n19343), .A2(n19342), .A3(n19341), .A4(n19340), .ZN(
        n19349) );
  AOI22_X1 U23380 ( .A1(n21008), .A2(\xmem_data[88][1] ), .B1(n27460), .B2(
        \xmem_data[89][1] ), .ZN(n19347) );
  AOI22_X1 U23381 ( .A1(n27462), .A2(\xmem_data[90][1] ), .B1(n27461), .B2(
        \xmem_data[91][1] ), .ZN(n19346) );
  AOI22_X1 U23382 ( .A1(n24571), .A2(\xmem_data[92][1] ), .B1(n24622), .B2(
        \xmem_data[93][1] ), .ZN(n19345) );
  AOI22_X1 U23383 ( .A1(n22719), .A2(\xmem_data[94][1] ), .B1(n27463), .B2(
        \xmem_data[95][1] ), .ZN(n19344) );
  NAND4_X1 U23384 ( .A1(n19347), .A2(n19346), .A3(n19345), .A4(n19344), .ZN(
        n19348) );
  OR4_X1 U23385 ( .A1(n19351), .A2(n19350), .A3(n19349), .A4(n19348), .ZN(
        n19352) );
  AND2_X1 U23386 ( .A1(n19352), .A2(n27494), .ZN(n19353) );
  NAND2_X1 U23387 ( .A1(n27446), .A2(\xmem_data[109][1] ), .ZN(n19380) );
  AOI22_X1 U23388 ( .A1(n24115), .A2(\xmem_data[120][1] ), .B1(n27460), .B2(
        \xmem_data[121][1] ), .ZN(n19358) );
  AOI22_X1 U23389 ( .A1(n27462), .A2(\xmem_data[122][1] ), .B1(n27461), .B2(
        \xmem_data[123][1] ), .ZN(n19357) );
  AOI22_X1 U23390 ( .A1(n28461), .A2(\xmem_data[124][1] ), .B1(n27525), .B2(
        \xmem_data[125][1] ), .ZN(n19356) );
  AOI22_X1 U23391 ( .A1(n25582), .A2(\xmem_data[126][1] ), .B1(n27463), .B2(
        \xmem_data[127][1] ), .ZN(n19355) );
  NAND4_X1 U23392 ( .A1(n19358), .A2(n19357), .A3(n19356), .A4(n19355), .ZN(
        n19377) );
  AOI22_X1 U23393 ( .A1(n23753), .A2(\xmem_data[96][1] ), .B1(n27435), .B2(
        \xmem_data[97][1] ), .ZN(n19362) );
  AOI22_X1 U23394 ( .A1(n27436), .A2(\xmem_data[98][1] ), .B1(n22752), .B2(
        \xmem_data[99][1] ), .ZN(n19361) );
  AOI22_X1 U23395 ( .A1(n3434), .A2(\xmem_data[100][1] ), .B1(n27437), .B2(
        \xmem_data[101][1] ), .ZN(n19360) );
  AOI22_X1 U23396 ( .A1(n27439), .A2(\xmem_data[102][1] ), .B1(n3222), .B2(
        \xmem_data[103][1] ), .ZN(n19359) );
  NAND4_X1 U23397 ( .A1(n19362), .A2(n19361), .A3(n19360), .A4(n19359), .ZN(
        n19376) );
  AOI22_X1 U23398 ( .A1(n27453), .A2(\xmem_data[112][1] ), .B1(n27452), .B2(
        \xmem_data[113][1] ), .ZN(n19366) );
  AOI22_X1 U23399 ( .A1(n16986), .A2(\xmem_data[114][1] ), .B1(n30613), .B2(
        \xmem_data[115][1] ), .ZN(n19365) );
  AOI22_X1 U23400 ( .A1(n27455), .A2(\xmem_data[116][1] ), .B1(n27454), .B2(
        \xmem_data[117][1] ), .ZN(n19364) );
  AOI22_X1 U23401 ( .A1(n14937), .A2(\xmem_data[118][1] ), .B1(n25677), .B2(
        \xmem_data[119][1] ), .ZN(n19363) );
  NAND4_X1 U23402 ( .A1(n19366), .A2(n19365), .A3(n19364), .A4(n19363), .ZN(
        n19375) );
  AOI22_X1 U23403 ( .A1(n27447), .A2(\xmem_data[110][1] ), .B1(n3357), .B2(
        \xmem_data[111][1] ), .ZN(n19367) );
  INV_X1 U23404 ( .A(n19367), .ZN(n19371) );
  AOI22_X1 U23405 ( .A1(n27445), .A2(\xmem_data[104][1] ), .B1(n27444), .B2(
        \xmem_data[105][1] ), .ZN(n19368) );
  INV_X1 U23406 ( .A(n19368), .ZN(n19370) );
  AND2_X1 U23407 ( .A1(n29762), .A2(\xmem_data[108][1] ), .ZN(n19369) );
  NOR3_X1 U23408 ( .A1(n19371), .A2(n19370), .A3(n19369), .ZN(n19373) );
  AOI22_X1 U23409 ( .A1(n24565), .A2(\xmem_data[106][1] ), .B1(n27994), .B2(
        \xmem_data[107][1] ), .ZN(n19372) );
  NAND2_X1 U23410 ( .A1(n19373), .A2(n19372), .ZN(n19374) );
  NOR4_X1 U23411 ( .A1(n19377), .A2(n19376), .A3(n19375), .A4(n19374), .ZN(
        n19379) );
  INV_X1 U23412 ( .A(n27496), .ZN(n19378) );
  AOI21_X1 U23413 ( .B1(n19380), .B2(n19379), .A(n19378), .ZN(n19381) );
  INV_X1 U23414 ( .A(n19381), .ZN(n19414) );
  NAND2_X1 U23415 ( .A1(n29306), .A2(\xmem_data[45][1] ), .ZN(n19408) );
  AOI22_X1 U23416 ( .A1(n27498), .A2(\xmem_data[32][1] ), .B1(n22727), .B2(
        \xmem_data[33][1] ), .ZN(n19385) );
  AOI22_X1 U23417 ( .A1(n27500), .A2(\xmem_data[34][1] ), .B1(n27499), .B2(
        \xmem_data[35][1] ), .ZN(n19384) );
  AOI22_X1 U23418 ( .A1(n3387), .A2(\xmem_data[36][1] ), .B1(n27501), .B2(
        \xmem_data[37][1] ), .ZN(n19383) );
  AOI22_X1 U23419 ( .A1(n27502), .A2(\xmem_data[38][1] ), .B1(n3220), .B2(
        \xmem_data[39][1] ), .ZN(n19382) );
  NAND4_X1 U23420 ( .A1(n19385), .A2(n19384), .A3(n19383), .A4(n19382), .ZN(
        n19405) );
  AOI22_X1 U23421 ( .A1(n27508), .A2(\xmem_data[46][1] ), .B1(n28415), .B2(
        \xmem_data[47][1] ), .ZN(n19386) );
  INV_X1 U23422 ( .A(n19386), .ZN(n19390) );
  AOI22_X1 U23423 ( .A1(n27445), .A2(\xmem_data[40][1] ), .B1(n27507), .B2(
        \xmem_data[41][1] ), .ZN(n19387) );
  INV_X1 U23424 ( .A(n19387), .ZN(n19389) );
  AND2_X1 U23425 ( .A1(n20962), .A2(\xmem_data[44][1] ), .ZN(n19388) );
  NOR3_X1 U23426 ( .A1(n19390), .A2(n19389), .A3(n19388), .ZN(n19392) );
  AOI22_X1 U23427 ( .A1(n30606), .A2(\xmem_data[42][1] ), .B1(n13444), .B2(
        \xmem_data[43][1] ), .ZN(n19391) );
  NAND2_X1 U23428 ( .A1(n19392), .A2(n19391), .ZN(n19403) );
  AOI22_X1 U23429 ( .A1(n27514), .A2(\xmem_data[48][1] ), .B1(n27513), .B2(
        \xmem_data[49][1] ), .ZN(n19396) );
  AOI22_X1 U23430 ( .A1(n27515), .A2(\xmem_data[50][1] ), .B1(n24597), .B2(
        \xmem_data[51][1] ), .ZN(n19395) );
  AOI22_X1 U23431 ( .A1(n20718), .A2(\xmem_data[52][1] ), .B1(n27516), .B2(
        \xmem_data[53][1] ), .ZN(n19394) );
  AOI22_X1 U23432 ( .A1(n24133), .A2(\xmem_data[54][1] ), .B1(n27518), .B2(
        \xmem_data[55][1] ), .ZN(n19393) );
  NAND4_X1 U23433 ( .A1(n19396), .A2(n19395), .A3(n19394), .A4(n19393), .ZN(
        n19402) );
  AOI22_X1 U23434 ( .A1(n30893), .A2(\xmem_data[56][1] ), .B1(n27523), .B2(
        \xmem_data[57][1] ), .ZN(n19400) );
  AOI22_X1 U23435 ( .A1(n27524), .A2(\xmem_data[58][1] ), .B1(n29089), .B2(
        \xmem_data[59][1] ), .ZN(n19399) );
  AOI22_X1 U23436 ( .A1(n28955), .A2(\xmem_data[60][1] ), .B1(n27525), .B2(
        \xmem_data[61][1] ), .ZN(n19398) );
  AOI22_X1 U23437 ( .A1(n3209), .A2(\xmem_data[62][1] ), .B1(n27526), .B2(
        \xmem_data[63][1] ), .ZN(n19397) );
  NAND4_X1 U23438 ( .A1(n19400), .A2(n19399), .A3(n19398), .A4(n19397), .ZN(
        n19401) );
  OR3_X1 U23439 ( .A1(n19403), .A2(n19402), .A3(n19401), .ZN(n19404) );
  NOR2_X1 U23440 ( .A1(n19405), .A2(n19404), .ZN(n19407) );
  AOI21_X1 U23441 ( .B1(n19408), .B2(n19407), .A(n19406), .ZN(n19409) );
  INV_X1 U23442 ( .A(n19409), .ZN(n19413) );
  AND2_X1 U23443 ( .A1(n19410), .A2(\xmem_data[13][1] ), .ZN(n19411) );
  NAND2_X1 U23444 ( .A1(n24657), .A2(n19411), .ZN(n19412) );
  AOI22_X1 U23445 ( .A1(n20577), .A2(\xmem_data[96][2] ), .B1(n27435), .B2(
        \xmem_data[97][2] ), .ZN(n19419) );
  AOI22_X1 U23446 ( .A1(n27436), .A2(\xmem_data[98][2] ), .B1(n22752), .B2(
        \xmem_data[99][2] ), .ZN(n19418) );
  AOI22_X1 U23447 ( .A1(n3245), .A2(\xmem_data[100][2] ), .B1(n27437), .B2(
        \xmem_data[101][2] ), .ZN(n19417) );
  AOI22_X1 U23448 ( .A1(n27439), .A2(\xmem_data[102][2] ), .B1(n3221), .B2(
        \xmem_data[103][2] ), .ZN(n19416) );
  NAND4_X1 U23449 ( .A1(n19419), .A2(n19418), .A3(n19417), .A4(n19416), .ZN(
        n19436) );
  AOI22_X1 U23450 ( .A1(n27453), .A2(\xmem_data[112][2] ), .B1(n27452), .B2(
        \xmem_data[113][2] ), .ZN(n19423) );
  AOI22_X1 U23451 ( .A1(n29310), .A2(\xmem_data[114][2] ), .B1(n25572), .B2(
        \xmem_data[115][2] ), .ZN(n19422) );
  AOI22_X1 U23452 ( .A1(n27455), .A2(\xmem_data[116][2] ), .B1(n27454), .B2(
        \xmem_data[117][2] ), .ZN(n19421) );
  AOI22_X1 U23453 ( .A1(n24509), .A2(\xmem_data[118][2] ), .B1(n14912), .B2(
        \xmem_data[119][2] ), .ZN(n19420) );
  NAND4_X1 U23454 ( .A1(n19423), .A2(n19422), .A3(n19421), .A4(n19420), .ZN(
        n19434) );
  AOI22_X1 U23455 ( .A1(n27825), .A2(\xmem_data[120][2] ), .B1(n27460), .B2(
        \xmem_data[121][2] ), .ZN(n19427) );
  AOI22_X1 U23456 ( .A1(n27462), .A2(\xmem_data[122][2] ), .B1(n27461), .B2(
        \xmem_data[123][2] ), .ZN(n19426) );
  AOI22_X1 U23457 ( .A1(n3338), .A2(\xmem_data[124][2] ), .B1(n31314), .B2(
        \xmem_data[125][2] ), .ZN(n19425) );
  AOI22_X1 U23458 ( .A1(n28293), .A2(\xmem_data[126][2] ), .B1(n27463), .B2(
        \xmem_data[127][2] ), .ZN(n19424) );
  NAND4_X1 U23459 ( .A1(n19427), .A2(n19426), .A3(n19425), .A4(n19424), .ZN(
        n19433) );
  AOI22_X1 U23460 ( .A1(n27445), .A2(\xmem_data[104][2] ), .B1(n27444), .B2(
        \xmem_data[105][2] ), .ZN(n19431) );
  AOI22_X1 U23461 ( .A1(n30883), .A2(\xmem_data[106][2] ), .B1(n24633), .B2(
        \xmem_data[107][2] ), .ZN(n19430) );
  AOI22_X1 U23462 ( .A1(n23742), .A2(\xmem_data[108][2] ), .B1(n27446), .B2(
        \xmem_data[109][2] ), .ZN(n19429) );
  AOI22_X1 U23463 ( .A1(n27447), .A2(\xmem_data[110][2] ), .B1(n25481), .B2(
        \xmem_data[111][2] ), .ZN(n19428) );
  NAND4_X1 U23464 ( .A1(n19431), .A2(n19430), .A3(n19429), .A4(n19428), .ZN(
        n19432) );
  OR3_X1 U23465 ( .A1(n19434), .A2(n19433), .A3(n19432), .ZN(n19435) );
  OAI21_X1 U23466 ( .B1(n19436), .B2(n19435), .A(n27496), .ZN(n19506) );
  AOI22_X1 U23467 ( .A1(n27852), .A2(\xmem_data[64][2] ), .B1(n27435), .B2(
        \xmem_data[65][2] ), .ZN(n19441) );
  AOI22_X1 U23468 ( .A1(n27436), .A2(\xmem_data[66][2] ), .B1(n31346), .B2(
        \xmem_data[67][2] ), .ZN(n19440) );
  AOI22_X1 U23469 ( .A1(n3332), .A2(\xmem_data[68][2] ), .B1(n27437), .B2(
        \xmem_data[69][2] ), .ZN(n19439) );
  AND2_X1 U23470 ( .A1(n3220), .A2(\xmem_data[71][2] ), .ZN(n19437) );
  AOI21_X1 U23471 ( .B1(n27439), .B2(\xmem_data[70][2] ), .A(n19437), .ZN(
        n19438) );
  NAND4_X1 U23472 ( .A1(n19441), .A2(n19440), .A3(n19439), .A4(n19438), .ZN(
        n19458) );
  AOI22_X1 U23473 ( .A1(n27453), .A2(\xmem_data[80][2] ), .B1(n27452), .B2(
        \xmem_data[81][2] ), .ZN(n19445) );
  AOI22_X1 U23474 ( .A1(n24131), .A2(\xmem_data[82][2] ), .B1(n20798), .B2(
        \xmem_data[83][2] ), .ZN(n19444) );
  AOI22_X1 U23475 ( .A1(n25607), .A2(\xmem_data[84][2] ), .B1(n27454), .B2(
        \xmem_data[85][2] ), .ZN(n19443) );
  AOI22_X1 U23476 ( .A1(n24593), .A2(\xmem_data[86][2] ), .B1(n24707), .B2(
        \xmem_data[87][2] ), .ZN(n19442) );
  NAND4_X1 U23477 ( .A1(n19445), .A2(n19444), .A3(n19443), .A4(n19442), .ZN(
        n19456) );
  AOI22_X1 U23478 ( .A1(n29012), .A2(\xmem_data[88][2] ), .B1(n27460), .B2(
        \xmem_data[89][2] ), .ZN(n19449) );
  AOI22_X1 U23479 ( .A1(n27462), .A2(\xmem_data[90][2] ), .B1(n27461), .B2(
        \xmem_data[91][2] ), .ZN(n19448) );
  AOI22_X1 U23480 ( .A1(n25718), .A2(\xmem_data[92][2] ), .B1(n23779), .B2(
        \xmem_data[93][2] ), .ZN(n19447) );
  AOI22_X1 U23481 ( .A1(n20734), .A2(\xmem_data[94][2] ), .B1(n27463), .B2(
        \xmem_data[95][2] ), .ZN(n19446) );
  NAND4_X1 U23482 ( .A1(n19449), .A2(n19448), .A3(n19447), .A4(n19446), .ZN(
        n19455) );
  AOI22_X1 U23483 ( .A1(n27445), .A2(\xmem_data[72][2] ), .B1(n27444), .B2(
        \xmem_data[73][2] ), .ZN(n19453) );
  AOI22_X1 U23484 ( .A1(n29289), .A2(\xmem_data[74][2] ), .B1(n27903), .B2(
        \xmem_data[75][2] ), .ZN(n19452) );
  AOI22_X1 U23485 ( .A1(n3374), .A2(\xmem_data[76][2] ), .B1(n27446), .B2(
        \xmem_data[77][2] ), .ZN(n19451) );
  AOI22_X1 U23486 ( .A1(n27447), .A2(\xmem_data[78][2] ), .B1(n20546), .B2(
        \xmem_data[79][2] ), .ZN(n19450) );
  NAND4_X1 U23487 ( .A1(n19453), .A2(n19452), .A3(n19451), .A4(n19450), .ZN(
        n19454) );
  OR3_X1 U23488 ( .A1(n19456), .A2(n19455), .A3(n19454), .ZN(n19457) );
  OAI21_X1 U23489 ( .B1(n19458), .B2(n19457), .A(n27494), .ZN(n19505) );
  AOI22_X1 U23490 ( .A1(n27498), .A2(\xmem_data[32][2] ), .B1(n28035), .B2(
        \xmem_data[33][2] ), .ZN(n19462) );
  AOI22_X1 U23491 ( .A1(n27500), .A2(\xmem_data[34][2] ), .B1(n27499), .B2(
        \xmem_data[35][2] ), .ZN(n19461) );
  AOI22_X1 U23492 ( .A1(n3386), .A2(\xmem_data[36][2] ), .B1(n27501), .B2(
        \xmem_data[37][2] ), .ZN(n19460) );
  AOI22_X1 U23493 ( .A1(n27502), .A2(\xmem_data[38][2] ), .B1(n3218), .B2(
        \xmem_data[39][2] ), .ZN(n19459) );
  NAND4_X1 U23494 ( .A1(n19462), .A2(n19461), .A3(n19460), .A4(n19459), .ZN(
        n19479) );
  AOI22_X1 U23495 ( .A1(n20942), .A2(\xmem_data[56][2] ), .B1(n27523), .B2(
        \xmem_data[57][2] ), .ZN(n19466) );
  AOI22_X1 U23496 ( .A1(n27524), .A2(\xmem_data[58][2] ), .B1(n20551), .B2(
        \xmem_data[59][2] ), .ZN(n19465) );
  AOI22_X1 U23497 ( .A1(n24623), .A2(\xmem_data[60][2] ), .B1(n27525), .B2(
        \xmem_data[61][2] ), .ZN(n19464) );
  AOI22_X1 U23498 ( .A1(n25526), .A2(\xmem_data[62][2] ), .B1(n27526), .B2(
        \xmem_data[63][2] ), .ZN(n19463) );
  NAND4_X1 U23499 ( .A1(n19466), .A2(n19465), .A3(n19464), .A4(n19463), .ZN(
        n19477) );
  AOI22_X1 U23500 ( .A1(n27514), .A2(\xmem_data[48][2] ), .B1(n27513), .B2(
        \xmem_data[49][2] ), .ZN(n19470) );
  AOI22_X1 U23501 ( .A1(n27515), .A2(\xmem_data[50][2] ), .B1(n29046), .B2(
        \xmem_data[51][2] ), .ZN(n19469) );
  AOI22_X1 U23502 ( .A1(n23795), .A2(\xmem_data[52][2] ), .B1(n27516), .B2(
        \xmem_data[53][2] ), .ZN(n19468) );
  AOI22_X1 U23503 ( .A1(n31330), .A2(\xmem_data[54][2] ), .B1(n27518), .B2(
        \xmem_data[55][2] ), .ZN(n19467) );
  NAND4_X1 U23504 ( .A1(n19470), .A2(n19469), .A3(n19468), .A4(n19467), .ZN(
        n19476) );
  AOI22_X1 U23505 ( .A1(n20724), .A2(\xmem_data[40][2] ), .B1(n27507), .B2(
        \xmem_data[41][2] ), .ZN(n19474) );
  AOI22_X1 U23506 ( .A1(n25449), .A2(\xmem_data[42][2] ), .B1(n13444), .B2(
        \xmem_data[43][2] ), .ZN(n19473) );
  AOI22_X1 U23507 ( .A1(n3138), .A2(\xmem_data[44][2] ), .B1(n31252), .B2(
        \xmem_data[45][2] ), .ZN(n19472) );
  AOI22_X1 U23508 ( .A1(n27508), .A2(\xmem_data[46][2] ), .B1(n28415), .B2(
        \xmem_data[47][2] ), .ZN(n19471) );
  NAND4_X1 U23509 ( .A1(n19474), .A2(n19473), .A3(n19472), .A4(n19471), .ZN(
        n19475) );
  OR3_X1 U23510 ( .A1(n19477), .A2(n19476), .A3(n19475), .ZN(n19478) );
  OAI21_X1 U23511 ( .B1(n19479), .B2(n19478), .A(n27577), .ZN(n19504) );
  AOI22_X1 U23512 ( .A1(n27568), .A2(\xmem_data[0][2] ), .B1(n27567), .B2(
        \xmem_data[1][2] ), .ZN(n19484) );
  AOI22_X1 U23513 ( .A1(n27564), .A2(\xmem_data[2][2] ), .B1(n27563), .B2(
        \xmem_data[3][2] ), .ZN(n19483) );
  AOI22_X1 U23514 ( .A1(n28245), .A2(\xmem_data[4][2] ), .B1(n25360), .B2(
        \xmem_data[5][2] ), .ZN(n19482) );
  AND2_X1 U23515 ( .A1(n3222), .A2(\xmem_data[7][2] ), .ZN(n19480) );
  AOI21_X1 U23516 ( .B1(n30503), .B2(\xmem_data[6][2] ), .A(n19480), .ZN(
        n19481) );
  NAND4_X1 U23517 ( .A1(n19484), .A2(n19483), .A3(n19482), .A4(n19481), .ZN(
        n19502) );
  AOI22_X1 U23518 ( .A1(n30744), .A2(\xmem_data[16][2] ), .B1(n27535), .B2(
        \xmem_data[17][2] ), .ZN(n19488) );
  AOI22_X1 U23519 ( .A1(n25710), .A2(\xmem_data[18][2] ), .B1(n27536), .B2(
        \xmem_data[19][2] ), .ZN(n19487) );
  AOI22_X1 U23520 ( .A1(n25672), .A2(\xmem_data[20][2] ), .B1(n25460), .B2(
        \xmem_data[21][2] ), .ZN(n19486) );
  AOI22_X1 U23521 ( .A1(n28096), .A2(\xmem_data[22][2] ), .B1(n25520), .B2(
        \xmem_data[23][2] ), .ZN(n19485) );
  NAND4_X1 U23522 ( .A1(n19488), .A2(n19487), .A3(n19486), .A4(n19485), .ZN(
        n19500) );
  AOI22_X1 U23523 ( .A1(n3375), .A2(\xmem_data[12][2] ), .B1(n28510), .B2(
        \xmem_data[13][2] ), .ZN(n19489) );
  INV_X1 U23524 ( .A(n19489), .ZN(n19499) );
  AOI22_X1 U23525 ( .A1(n3342), .A2(\xmem_data[10][2] ), .B1(n27550), .B2(
        \xmem_data[11][2] ), .ZN(n19492) );
  AOI22_X1 U23526 ( .A1(n27551), .A2(\xmem_data[14][2] ), .B1(n20588), .B2(
        \xmem_data[15][2] ), .ZN(n19491) );
  AOI22_X1 U23527 ( .A1(n29494), .A2(\xmem_data[8][2] ), .B1(n25509), .B2(
        \xmem_data[9][2] ), .ZN(n19490) );
  NAND3_X1 U23528 ( .A1(n19492), .A2(n19491), .A3(n19490), .ZN(n19498) );
  AOI22_X1 U23529 ( .A1(n25678), .A2(\xmem_data[24][2] ), .B1(n13452), .B2(
        \xmem_data[25][2] ), .ZN(n19496) );
  AOI22_X1 U23530 ( .A1(n30849), .A2(\xmem_data[26][2] ), .B1(n30598), .B2(
        \xmem_data[27][2] ), .ZN(n19495) );
  AOI22_X1 U23531 ( .A1(n3328), .A2(\xmem_data[28][2] ), .B1(n24622), .B2(
        \xmem_data[29][2] ), .ZN(n19494) );
  AOI22_X1 U23532 ( .A1(n27542), .A2(\xmem_data[30][2] ), .B1(n11008), .B2(
        \xmem_data[31][2] ), .ZN(n19493) );
  NAND4_X1 U23533 ( .A1(n19496), .A2(n19495), .A3(n19494), .A4(n19493), .ZN(
        n19497) );
  XNOR2_X1 U23534 ( .A(n32127), .B(\fmem_data[20][7] ), .ZN(n30458) );
  OAI22_X1 U23535 ( .A1(n30795), .A2(n35740), .B1(n30458), .B2(n35739), .ZN(
        n23169) );
  NOR2_X1 U23536 ( .A1(n23170), .A2(n23169), .ZN(n19508) );
  NAND2_X1 U23537 ( .A1(n23170), .A2(n23169), .ZN(n19507) );
  OAI21_X1 U23538 ( .B1(n19509), .B2(n19508), .A(n19507), .ZN(n23186) );
  FA_X1 U23539 ( .A(n19512), .B(n19511), .CI(n19510), .CO(n16354), .S(n23185)
         );
  XNOR2_X1 U23540 ( .A(n35122), .B(\fmem_data[12][1] ), .ZN(n30828) );
  AOI22_X1 U23541 ( .A1(n20730), .A2(\xmem_data[96][1] ), .B1(n29049), .B2(
        \xmem_data[97][1] ), .ZN(n19516) );
  AOI22_X1 U23542 ( .A1(n20731), .A2(\xmem_data[98][1] ), .B1(n21009), .B2(
        \xmem_data[99][1] ), .ZN(n19515) );
  AOI22_X1 U23543 ( .A1(n20732), .A2(\xmem_data[100][1] ), .B1(n23723), .B2(
        \xmem_data[101][1] ), .ZN(n19514) );
  AOI22_X1 U23544 ( .A1(n20734), .A2(\xmem_data[102][1] ), .B1(n20733), .B2(
        \xmem_data[103][1] ), .ZN(n19513) );
  NAND4_X1 U23545 ( .A1(n19516), .A2(n19515), .A3(n19514), .A4(n19513), .ZN(
        n19532) );
  AOI22_X1 U23546 ( .A1(n20708), .A2(\xmem_data[104][1] ), .B1(n20707), .B2(
        \xmem_data[105][1] ), .ZN(n19520) );
  AOI22_X1 U23547 ( .A1(n20710), .A2(\xmem_data[106][1] ), .B1(n20709), .B2(
        \xmem_data[107][1] ), .ZN(n19519) );
  AOI22_X1 U23548 ( .A1(n3414), .A2(\xmem_data[108][1] ), .B1(n20711), .B2(
        \xmem_data[109][1] ), .ZN(n19518) );
  AOI22_X1 U23549 ( .A1(n28044), .A2(\xmem_data[110][1] ), .B1(n3222), .B2(
        \xmem_data[111][1] ), .ZN(n19517) );
  NAND4_X1 U23550 ( .A1(n19520), .A2(n19519), .A3(n19518), .A4(n19517), .ZN(
        n19531) );
  AOI22_X1 U23551 ( .A1(n20724), .A2(\xmem_data[112][1] ), .B1(n20723), .B2(
        \xmem_data[113][1] ), .ZN(n19524) );
  AOI22_X1 U23552 ( .A1(n20725), .A2(\xmem_data[114][1] ), .B1(n30882), .B2(
        \xmem_data[115][1] ), .ZN(n19523) );
  AOI22_X1 U23553 ( .A1(n30295), .A2(\xmem_data[116][1] ), .B1(n27547), .B2(
        \xmem_data[117][1] ), .ZN(n19522) );
  AOI22_X1 U23554 ( .A1(n30885), .A2(\xmem_data[118][1] ), .B1(n25481), .B2(
        \xmem_data[119][1] ), .ZN(n19521) );
  NAND4_X1 U23555 ( .A1(n19524), .A2(n19523), .A3(n19522), .A4(n19521), .ZN(
        n19530) );
  AOI22_X1 U23556 ( .A1(n20716), .A2(\xmem_data[120][1] ), .B1(n21015), .B2(
        \xmem_data[121][1] ), .ZN(n19528) );
  AOI22_X1 U23557 ( .A1(n25459), .A2(\xmem_data[122][1] ), .B1(n20717), .B2(
        \xmem_data[123][1] ), .ZN(n19527) );
  AOI22_X1 U23558 ( .A1(n29396), .A2(\xmem_data[124][1] ), .B1(n25574), .B2(
        \xmem_data[125][1] ), .ZN(n19526) );
  AOI22_X1 U23559 ( .A1(n24214), .A2(\xmem_data[126][1] ), .B1(n14912), .B2(
        \xmem_data[127][1] ), .ZN(n19525) );
  NAND4_X1 U23560 ( .A1(n19528), .A2(n19527), .A3(n19526), .A4(n19525), .ZN(
        n19529) );
  OR4_X1 U23561 ( .A1(n19532), .A2(n19531), .A3(n19530), .A4(n19529), .ZN(
        n19555) );
  AOI22_X1 U23562 ( .A1(n20730), .A2(\xmem_data[64][1] ), .B1(n28380), .B2(
        \xmem_data[65][1] ), .ZN(n19536) );
  AOI22_X1 U23563 ( .A1(n20731), .A2(\xmem_data[66][1] ), .B1(n27856), .B2(
        \xmem_data[67][1] ), .ZN(n19535) );
  AOI22_X1 U23564 ( .A1(n20732), .A2(\xmem_data[68][1] ), .B1(n24521), .B2(
        \xmem_data[69][1] ), .ZN(n19534) );
  AOI22_X1 U23565 ( .A1(n20734), .A2(\xmem_data[70][1] ), .B1(n20733), .B2(
        \xmem_data[71][1] ), .ZN(n19533) );
  NAND4_X1 U23566 ( .A1(n19536), .A2(n19535), .A3(n19534), .A4(n19533), .ZN(
        n19553) );
  AOI22_X1 U23567 ( .A1(n20708), .A2(\xmem_data[72][1] ), .B1(n20707), .B2(
        \xmem_data[73][1] ), .ZN(n19541) );
  AOI22_X1 U23568 ( .A1(n20710), .A2(\xmem_data[74][1] ), .B1(n20709), .B2(
        \xmem_data[75][1] ), .ZN(n19540) );
  AOI22_X1 U23569 ( .A1(n3306), .A2(\xmem_data[76][1] ), .B1(n20711), .B2(
        \xmem_data[77][1] ), .ZN(n19539) );
  AND2_X1 U23570 ( .A1(n3220), .A2(\xmem_data[79][1] ), .ZN(n19537) );
  AOI21_X1 U23571 ( .B1(n25508), .B2(\xmem_data[78][1] ), .A(n19537), .ZN(
        n19538) );
  NAND4_X1 U23572 ( .A1(n19541), .A2(n19540), .A3(n19539), .A4(n19538), .ZN(
        n19552) );
  AOI22_X1 U23573 ( .A1(n20724), .A2(\xmem_data[80][1] ), .B1(n20723), .B2(
        \xmem_data[81][1] ), .ZN(n19545) );
  AOI22_X1 U23574 ( .A1(n20725), .A2(\xmem_data[82][1] ), .B1(n25415), .B2(
        \xmem_data[83][1] ), .ZN(n19544) );
  AOI22_X1 U23575 ( .A1(n25732), .A2(\xmem_data[84][1] ), .B1(n28045), .B2(
        \xmem_data[85][1] ), .ZN(n19543) );
  AOI22_X1 U23576 ( .A1(n25422), .A2(\xmem_data[86][1] ), .B1(n13475), .B2(
        \xmem_data[87][1] ), .ZN(n19542) );
  NAND4_X1 U23577 ( .A1(n19545), .A2(n19544), .A3(n19543), .A4(n19542), .ZN(
        n19551) );
  AOI22_X1 U23578 ( .A1(n20716), .A2(\xmem_data[88][1] ), .B1(n24448), .B2(
        \xmem_data[89][1] ), .ZN(n19549) );
  AOI22_X1 U23579 ( .A1(n20541), .A2(\xmem_data[90][1] ), .B1(n20717), .B2(
        \xmem_data[91][1] ), .ZN(n19548) );
  AOI22_X1 U23580 ( .A1(n27755), .A2(\xmem_data[92][1] ), .B1(n27516), .B2(
        \xmem_data[93][1] ), .ZN(n19547) );
  AOI22_X1 U23581 ( .A1(n24509), .A2(\xmem_data[94][1] ), .B1(n22718), .B2(
        \xmem_data[95][1] ), .ZN(n19546) );
  NAND4_X1 U23582 ( .A1(n19549), .A2(n19548), .A3(n19547), .A4(n19546), .ZN(
        n19550) );
  OR4_X1 U23583 ( .A1(n19553), .A2(n19552), .A3(n19551), .A4(n19550), .ZN(
        n19554) );
  AOI22_X1 U23584 ( .A1(n20742), .A2(n19555), .B1(n20833), .B2(n19554), .ZN(
        n19608) );
  AOI22_X1 U23585 ( .A1(n27825), .A2(\xmem_data[0][1] ), .B1(n28380), .B2(
        \xmem_data[1][1] ), .ZN(n19559) );
  AOI22_X1 U23586 ( .A1(n25632), .A2(\xmem_data[2][1] ), .B1(n25716), .B2(
        \xmem_data[3][1] ), .ZN(n19558) );
  AOI22_X1 U23587 ( .A1(n23780), .A2(\xmem_data[4][1] ), .B1(n20781), .B2(
        \xmem_data[5][1] ), .ZN(n19557) );
  AOI22_X1 U23588 ( .A1(n20782), .A2(\xmem_data[6][1] ), .B1(n22751), .B2(
        \xmem_data[7][1] ), .ZN(n19556) );
  NAND4_X1 U23589 ( .A1(n19559), .A2(n19558), .A3(n19557), .A4(n19556), .ZN(
        n19562) );
  AOI22_X1 U23590 ( .A1(n3333), .A2(\xmem_data[12][1] ), .B1(n29253), .B2(
        \xmem_data[13][1] ), .ZN(n19560) );
  INV_X1 U23591 ( .A(n19560), .ZN(n19561) );
  NOR2_X1 U23592 ( .A1(n19562), .A2(n19561), .ZN(n19566) );
  AOI22_X1 U23593 ( .A1(n27439), .A2(\xmem_data[14][1] ), .B1(n3220), .B2(
        \xmem_data[15][1] ), .ZN(n19565) );
  AOI22_X1 U23594 ( .A1(n27500), .A2(\xmem_data[10][1] ), .B1(n28317), .B2(
        \xmem_data[11][1] ), .ZN(n19564) );
  AOI22_X1 U23595 ( .A1(n20770), .A2(\xmem_data[8][1] ), .B1(n20769), .B2(
        \xmem_data[9][1] ), .ZN(n19563) );
  NAND4_X1 U23596 ( .A1(n19566), .A2(n19565), .A3(n19564), .A4(n19563), .ZN(
        n19581) );
  AOI22_X1 U23597 ( .A1(n29494), .A2(\xmem_data[16][1] ), .B1(n20787), .B2(
        \xmem_data[17][1] ), .ZN(n19567) );
  AOI22_X1 U23598 ( .A1(n25422), .A2(\xmem_data[22][1] ), .B1(n28415), .B2(
        \xmem_data[23][1] ), .ZN(n19569) );
  NAND2_X1 U23599 ( .A1(n29762), .A2(\xmem_data[20][1] ), .ZN(n19568) );
  NAND2_X1 U23600 ( .A1(n19569), .A2(n19568), .ZN(n19572) );
  AOI22_X1 U23601 ( .A1(n25490), .A2(\xmem_data[18][1] ), .B1(n13444), .B2(
        \xmem_data[19][1] ), .ZN(n19570) );
  INV_X1 U23602 ( .A(n19570), .ZN(n19571) );
  OR3_X1 U23603 ( .A1(n19573), .A2(n19572), .A3(n19571), .ZN(n19579) );
  AOI22_X1 U23604 ( .A1(n30943), .A2(\xmem_data[24][1] ), .B1(n20775), .B2(
        \xmem_data[25][1] ), .ZN(n19577) );
  AOI22_X1 U23605 ( .A1(n29109), .A2(\xmem_data[26][1] ), .B1(n24597), .B2(
        \xmem_data[27][1] ), .ZN(n19576) );
  AOI22_X1 U23606 ( .A1(n28091), .A2(\xmem_data[28][1] ), .B1(n27864), .B2(
        \xmem_data[29][1] ), .ZN(n19575) );
  AOI22_X1 U23607 ( .A1(n28059), .A2(\xmem_data[30][1] ), .B1(n24219), .B2(
        \xmem_data[31][1] ), .ZN(n19574) );
  NAND4_X1 U23608 ( .A1(n19577), .A2(n19576), .A3(n19575), .A4(n19574), .ZN(
        n19578) );
  OR2_X1 U23609 ( .A1(n19579), .A2(n19578), .ZN(n19580) );
  NOR2_X1 U23610 ( .A1(n19581), .A2(n19580), .ZN(n19583) );
  NAND2_X1 U23611 ( .A1(n25514), .A2(\xmem_data[21][1] ), .ZN(n19582) );
  AOI21_X1 U23612 ( .B1(n19583), .B2(n19582), .A(n20188), .ZN(n19584) );
  INV_X1 U23613 ( .A(n19584), .ZN(n19607) );
  AOI22_X1 U23614 ( .A1(n20815), .A2(\xmem_data[32][1] ), .B1(n20814), .B2(
        \xmem_data[33][1] ), .ZN(n19588) );
  AOI22_X1 U23615 ( .A1(n30557), .A2(\xmem_data[34][1] ), .B1(n25364), .B2(
        \xmem_data[35][1] ), .ZN(n19587) );
  AOI22_X1 U23616 ( .A1(n20817), .A2(\xmem_data[36][1] ), .B1(n31314), .B2(
        \xmem_data[37][1] ), .ZN(n19586) );
  AOI22_X1 U23617 ( .A1(n20818), .A2(\xmem_data[38][1] ), .B1(n22751), .B2(
        \xmem_data[39][1] ), .ZN(n19585) );
  NAND4_X1 U23618 ( .A1(n19588), .A2(n19587), .A3(n19586), .A4(n19585), .ZN(
        n19604) );
  AOI22_X1 U23619 ( .A1(n20826), .A2(\xmem_data[40][1] ), .B1(n25388), .B2(
        \xmem_data[41][1] ), .ZN(n19592) );
  AOI22_X1 U23620 ( .A1(n20827), .A2(\xmem_data[42][1] ), .B1(n29328), .B2(
        \xmem_data[43][1] ), .ZN(n19591) );
  AOI22_X1 U23621 ( .A1(n20828), .A2(\xmem_data[44][1] ), .B1(n30863), .B2(
        \xmem_data[45][1] ), .ZN(n19590) );
  AOI22_X1 U23622 ( .A1(n27439), .A2(\xmem_data[46][1] ), .B1(n3222), .B2(
        \xmem_data[47][1] ), .ZN(n19589) );
  NAND4_X1 U23623 ( .A1(n19592), .A2(n19591), .A3(n19590), .A4(n19589), .ZN(
        n19603) );
  AOI22_X1 U23624 ( .A1(n20805), .A2(\xmem_data[48][1] ), .B1(n24207), .B2(
        \xmem_data[49][1] ), .ZN(n19596) );
  AOI22_X1 U23625 ( .A1(n20807), .A2(\xmem_data[50][1] ), .B1(n20806), .B2(
        \xmem_data[51][1] ), .ZN(n19595) );
  AOI22_X1 U23626 ( .A1(n20808), .A2(\xmem_data[52][1] ), .B1(n27446), .B2(
        \xmem_data[53][1] ), .ZN(n19594) );
  AOI22_X1 U23627 ( .A1(n20809), .A2(\xmem_data[54][1] ), .B1(n14933), .B2(
        \xmem_data[55][1] ), .ZN(n19593) );
  NAND4_X1 U23628 ( .A1(n19596), .A2(n19595), .A3(n19594), .A4(n19593), .ZN(
        n19602) );
  AOI22_X1 U23629 ( .A1(n20799), .A2(\xmem_data[56][1] ), .B1(n20958), .B2(
        \xmem_data[57][1] ), .ZN(n19600) );
  AOI22_X1 U23630 ( .A1(n29310), .A2(\xmem_data[58][1] ), .B1(n20798), .B2(
        \xmem_data[59][1] ), .ZN(n19599) );
  AOI22_X1 U23631 ( .A1(n29605), .A2(\xmem_data[60][1] ), .B1(n25383), .B2(
        \xmem_data[61][1] ), .ZN(n19598) );
  AOI22_X1 U23632 ( .A1(n20800), .A2(\xmem_data[62][1] ), .B1(n23796), .B2(
        \xmem_data[63][1] ), .ZN(n19597) );
  NAND4_X1 U23633 ( .A1(n19600), .A2(n19599), .A3(n19598), .A4(n19597), .ZN(
        n19601) );
  OR4_X1 U23634 ( .A1(n19604), .A2(n19603), .A3(n19602), .A4(n19601), .ZN(
        n19605) );
  NAND2_X1 U23635 ( .A1(n19605), .A2(n20765), .ZN(n19606) );
  XOR2_X1 U23636 ( .A(\fmem_data[28][6] ), .B(\fmem_data[28][7] ), .Z(n19609)
         );
  AOI22_X1 U23637 ( .A1(n20730), .A2(\xmem_data[96][0] ), .B1(n28097), .B2(
        \xmem_data[97][0] ), .ZN(n19613) );
  AOI22_X1 U23638 ( .A1(n20731), .A2(\xmem_data[98][0] ), .B1(n25716), .B2(
        \xmem_data[99][0] ), .ZN(n19612) );
  AOI22_X1 U23639 ( .A1(n20732), .A2(\xmem_data[100][0] ), .B1(n14883), .B2(
        \xmem_data[101][0] ), .ZN(n19611) );
  AOI22_X1 U23640 ( .A1(n20734), .A2(\xmem_data[102][0] ), .B1(n20733), .B2(
        \xmem_data[103][0] ), .ZN(n19610) );
  NAND4_X1 U23641 ( .A1(n19613), .A2(n19612), .A3(n19611), .A4(n19610), .ZN(
        n19630) );
  AOI22_X1 U23642 ( .A1(n20708), .A2(\xmem_data[104][0] ), .B1(n20707), .B2(
        \xmem_data[105][0] ), .ZN(n19618) );
  AOI22_X1 U23643 ( .A1(n20710), .A2(\xmem_data[106][0] ), .B1(n20709), .B2(
        \xmem_data[107][0] ), .ZN(n19617) );
  AOI22_X1 U23644 ( .A1(n3386), .A2(\xmem_data[108][0] ), .B1(n20711), .B2(
        \xmem_data[109][0] ), .ZN(n19616) );
  AND2_X1 U23645 ( .A1(n3217), .A2(\xmem_data[111][0] ), .ZN(n19614) );
  AOI21_X1 U23646 ( .B1(n27902), .B2(\xmem_data[110][0] ), .A(n19614), .ZN(
        n19615) );
  NAND4_X1 U23647 ( .A1(n19618), .A2(n19617), .A3(n19616), .A4(n19615), .ZN(
        n19629) );
  AOI22_X1 U23648 ( .A1(n20724), .A2(\xmem_data[112][0] ), .B1(n20723), .B2(
        \xmem_data[113][0] ), .ZN(n19622) );
  AOI22_X1 U23649 ( .A1(n20725), .A2(\xmem_data[114][0] ), .B1(n20993), .B2(
        \xmem_data[115][0] ), .ZN(n19621) );
  AOI22_X1 U23650 ( .A1(n25377), .A2(\xmem_data[116][0] ), .B1(n25450), .B2(
        \xmem_data[117][0] ), .ZN(n19620) );
  AOI22_X1 U23651 ( .A1(n30607), .A2(\xmem_data[118][0] ), .B1(n22739), .B2(
        \xmem_data[119][0] ), .ZN(n19619) );
  NAND4_X1 U23652 ( .A1(n19622), .A2(n19621), .A3(n19620), .A4(n19619), .ZN(
        n19628) );
  AOI22_X1 U23653 ( .A1(n28752), .A2(\xmem_data[124][0] ), .B1(n30542), .B2(
        \xmem_data[125][0] ), .ZN(n19626) );
  AOI22_X1 U23654 ( .A1(n23763), .A2(\xmem_data[122][0] ), .B1(n20717), .B2(
        \xmem_data[123][0] ), .ZN(n19625) );
  AOI22_X1 U23655 ( .A1(n20716), .A2(\xmem_data[120][0] ), .B1(n30552), .B2(
        \xmem_data[121][0] ), .ZN(n19624) );
  AOI22_X1 U23656 ( .A1(n23717), .A2(\xmem_data[126][0] ), .B1(n21006), .B2(
        \xmem_data[127][0] ), .ZN(n19623) );
  NAND4_X1 U23657 ( .A1(n19626), .A2(n19625), .A3(n19624), .A4(n19623), .ZN(
        n19627) );
  OR4_X1 U23658 ( .A1(n19630), .A2(n19629), .A3(n19628), .A4(n19627), .ZN(
        n19631) );
  NAND2_X1 U23659 ( .A1(n19631), .A2(n20742), .ZN(n19705) );
  AOI22_X1 U23660 ( .A1(n20815), .A2(\xmem_data[32][0] ), .B1(n20814), .B2(
        \xmem_data[33][0] ), .ZN(n19635) );
  AOI22_X1 U23661 ( .A1(n30557), .A2(\xmem_data[34][0] ), .B1(n28327), .B2(
        \xmem_data[35][0] ), .ZN(n19634) );
  AOI22_X1 U23662 ( .A1(n20817), .A2(\xmem_data[36][0] ), .B1(n23779), .B2(
        \xmem_data[37][0] ), .ZN(n19633) );
  AOI22_X1 U23663 ( .A1(n20818), .A2(\xmem_data[38][0] ), .B1(n17049), .B2(
        \xmem_data[39][0] ), .ZN(n19632) );
  NAND4_X1 U23664 ( .A1(n19635), .A2(n19634), .A3(n19633), .A4(n19632), .ZN(
        n19652) );
  AOI22_X1 U23665 ( .A1(n20826), .A2(\xmem_data[40][0] ), .B1(n30524), .B2(
        \xmem_data[41][0] ), .ZN(n19640) );
  AOI22_X1 U23666 ( .A1(n20827), .A2(\xmem_data[42][0] ), .B1(n29118), .B2(
        \xmem_data[43][0] ), .ZN(n19639) );
  AOI22_X1 U23667 ( .A1(n20828), .A2(\xmem_data[44][0] ), .B1(n30863), .B2(
        \xmem_data[45][0] ), .ZN(n19638) );
  AND2_X1 U23668 ( .A1(n3221), .A2(\xmem_data[47][0] ), .ZN(n19636) );
  AOI21_X1 U23669 ( .B1(n24562), .B2(\xmem_data[46][0] ), .A(n19636), .ZN(
        n19637) );
  NAND4_X1 U23670 ( .A1(n19640), .A2(n19639), .A3(n19638), .A4(n19637), .ZN(
        n19651) );
  AOI22_X1 U23671 ( .A1(n20805), .A2(\xmem_data[48][0] ), .B1(n24695), .B2(
        \xmem_data[49][0] ), .ZN(n19644) );
  AOI22_X1 U23672 ( .A1(n20807), .A2(\xmem_data[50][0] ), .B1(n20806), .B2(
        \xmem_data[51][0] ), .ZN(n19643) );
  AOI22_X1 U23673 ( .A1(n20808), .A2(\xmem_data[52][0] ), .B1(n15011), .B2(
        \xmem_data[53][0] ), .ZN(n19642) );
  AOI22_X1 U23674 ( .A1(n20809), .A2(\xmem_data[54][0] ), .B1(n27943), .B2(
        \xmem_data[55][0] ), .ZN(n19641) );
  NAND4_X1 U23675 ( .A1(n19644), .A2(n19643), .A3(n19642), .A4(n19641), .ZN(
        n19650) );
  AOI22_X1 U23676 ( .A1(n17018), .A2(\xmem_data[60][0] ), .B1(n27516), .B2(
        \xmem_data[61][0] ), .ZN(n19648) );
  AOI22_X1 U23677 ( .A1(n25567), .A2(\xmem_data[58][0] ), .B1(n20798), .B2(
        \xmem_data[59][0] ), .ZN(n19647) );
  AOI22_X1 U23678 ( .A1(n20799), .A2(\xmem_data[56][0] ), .B1(n21015), .B2(
        \xmem_data[57][0] ), .ZN(n19646) );
  AOI22_X1 U23679 ( .A1(n20800), .A2(\xmem_data[62][0] ), .B1(n29048), .B2(
        \xmem_data[63][0] ), .ZN(n19645) );
  NAND4_X1 U23680 ( .A1(n19648), .A2(n19647), .A3(n19646), .A4(n19645), .ZN(
        n19649) );
  OR4_X1 U23681 ( .A1(n19652), .A2(n19651), .A3(n19650), .A4(n19649), .ZN(
        n19653) );
  NAND2_X1 U23682 ( .A1(n19653), .A2(n20765), .ZN(n19704) );
  AOI22_X1 U23683 ( .A1(n20708), .A2(\xmem_data[72][0] ), .B1(n20707), .B2(
        \xmem_data[73][0] ), .ZN(n19658) );
  AOI22_X1 U23684 ( .A1(n20710), .A2(\xmem_data[74][0] ), .B1(n20709), .B2(
        \xmem_data[75][0] ), .ZN(n19657) );
  AOI22_X1 U23685 ( .A1(n3424), .A2(\xmem_data[76][0] ), .B1(n20711), .B2(
        \xmem_data[77][0] ), .ZN(n19656) );
  AND2_X1 U23686 ( .A1(n3218), .A2(\xmem_data[79][0] ), .ZN(n19654) );
  AOI21_X1 U23687 ( .B1(n28355), .B2(\xmem_data[78][0] ), .A(n19654), .ZN(
        n19655) );
  NAND4_X1 U23688 ( .A1(n19658), .A2(n19657), .A3(n19656), .A4(n19655), .ZN(
        n19674) );
  AOI22_X1 U23689 ( .A1(n20716), .A2(\xmem_data[88][0] ), .B1(n27535), .B2(
        \xmem_data[89][0] ), .ZN(n19662) );
  AOI22_X1 U23690 ( .A1(n28980), .A2(\xmem_data[90][0] ), .B1(n20717), .B2(
        \xmem_data[91][0] ), .ZN(n19661) );
  AOI22_X1 U23691 ( .A1(n3120), .A2(\xmem_data[92][0] ), .B1(n29162), .B2(
        \xmem_data[93][0] ), .ZN(n19660) );
  AOI22_X1 U23692 ( .A1(n21007), .A2(\xmem_data[94][0] ), .B1(n28492), .B2(
        \xmem_data[95][0] ), .ZN(n19659) );
  NAND4_X1 U23693 ( .A1(n19662), .A2(n19661), .A3(n19660), .A4(n19659), .ZN(
        n19673) );
  AOI22_X1 U23694 ( .A1(n20724), .A2(\xmem_data[80][0] ), .B1(n20723), .B2(
        \xmem_data[81][0] ), .ZN(n19666) );
  AOI22_X1 U23695 ( .A1(n20725), .A2(\xmem_data[82][0] ), .B1(n25616), .B2(
        \xmem_data[83][0] ), .ZN(n19665) );
  AOI22_X1 U23696 ( .A1(n27396), .A2(\xmem_data[84][0] ), .B1(n27547), .B2(
        \xmem_data[85][0] ), .ZN(n19664) );
  AOI22_X1 U23697 ( .A1(n27447), .A2(\xmem_data[86][0] ), .B1(n13475), .B2(
        \xmem_data[87][0] ), .ZN(n19663) );
  NAND4_X1 U23698 ( .A1(n19666), .A2(n19665), .A3(n19664), .A4(n19663), .ZN(
        n19672) );
  AOI22_X1 U23699 ( .A1(n20730), .A2(\xmem_data[64][0] ), .B1(n28301), .B2(
        \xmem_data[65][0] ), .ZN(n19670) );
  AOI22_X1 U23700 ( .A1(n20731), .A2(\xmem_data[66][0] ), .B1(n21009), .B2(
        \xmem_data[67][0] ), .ZN(n19669) );
  AOI22_X1 U23701 ( .A1(n20732), .A2(\xmem_data[68][0] ), .B1(n20949), .B2(
        \xmem_data[69][0] ), .ZN(n19668) );
  AOI22_X1 U23702 ( .A1(n20734), .A2(\xmem_data[70][0] ), .B1(n20733), .B2(
        \xmem_data[71][0] ), .ZN(n19667) );
  NAND4_X1 U23703 ( .A1(n19670), .A2(n19669), .A3(n19668), .A4(n19667), .ZN(
        n19671) );
  OR4_X1 U23704 ( .A1(n19674), .A2(n19673), .A3(n19672), .A4(n19671), .ZN(
        n19675) );
  NAND2_X1 U23705 ( .A1(n19675), .A2(n20833), .ZN(n19703) );
  AOI22_X1 U23706 ( .A1(n20770), .A2(\xmem_data[8][0] ), .B1(n20769), .B2(
        \xmem_data[9][0] ), .ZN(n19679) );
  AOI22_X1 U23707 ( .A1(n28038), .A2(\xmem_data[10][0] ), .B1(n22729), .B2(
        \xmem_data[11][0] ), .ZN(n19678) );
  AOI22_X1 U23708 ( .A1(n22728), .A2(\xmem_data[12][0] ), .B1(n30589), .B2(
        \xmem_data[13][0] ), .ZN(n19677) );
  AOI22_X1 U23709 ( .A1(n25508), .A2(\xmem_data[14][0] ), .B1(n3217), .B2(
        \xmem_data[15][0] ), .ZN(n19676) );
  AOI22_X1 U23710 ( .A1(n28754), .A2(\xmem_data[0][0] ), .B1(n25435), .B2(
        \xmem_data[1][0] ), .ZN(n19683) );
  AOI22_X1 U23711 ( .A1(n25632), .A2(\xmem_data[2][0] ), .B1(n21051), .B2(
        \xmem_data[3][0] ), .ZN(n19682) );
  AOI22_X1 U23712 ( .A1(n29816), .A2(\xmem_data[4][0] ), .B1(n20781), .B2(
        \xmem_data[5][0] ), .ZN(n19681) );
  AOI22_X1 U23713 ( .A1(n20782), .A2(\xmem_data[6][0] ), .B1(n28468), .B2(
        \xmem_data[7][0] ), .ZN(n19680) );
  NAND4_X1 U23714 ( .A1(n19683), .A2(n19682), .A3(n19681), .A4(n19680), .ZN(
        n19686) );
  AOI22_X1 U23715 ( .A1(n30883), .A2(\xmem_data[18][0] ), .B1(n25616), .B2(
        \xmem_data[19][0] ), .ZN(n19684) );
  INV_X1 U23716 ( .A(n19684), .ZN(n19685) );
  NOR2_X1 U23717 ( .A1(n19686), .A2(n19685), .ZN(n19700) );
  AOI22_X1 U23718 ( .A1(n25422), .A2(\xmem_data[22][0] ), .B1(n3358), .B2(
        \xmem_data[23][0] ), .ZN(n19687) );
  INV_X1 U23719 ( .A(n19687), .ZN(n19692) );
  AND2_X1 U23720 ( .A1(n3138), .A2(\xmem_data[20][0] ), .ZN(n19691) );
  NAND2_X1 U23721 ( .A1(n20787), .A2(\xmem_data[17][0] ), .ZN(n19689) );
  NAND2_X1 U23722 ( .A1(n29431), .A2(\xmem_data[16][0] ), .ZN(n19688) );
  NAND2_X1 U23723 ( .A1(n19689), .A2(n19688), .ZN(n19690) );
  NOR3_X1 U23724 ( .A1(n19692), .A2(n19691), .A3(n19690), .ZN(n19699) );
  AOI22_X1 U23725 ( .A1(n27944), .A2(\xmem_data[24][0] ), .B1(n20775), .B2(
        \xmem_data[25][0] ), .ZN(n19696) );
  AOI22_X1 U23726 ( .A1(n20495), .A2(\xmem_data[26][0] ), .B1(n20798), .B2(
        \xmem_data[27][0] ), .ZN(n19695) );
  AOI22_X1 U23727 ( .A1(n3158), .A2(\xmem_data[28][0] ), .B1(n3208), .B2(
        \xmem_data[29][0] ), .ZN(n19694) );
  AOI22_X1 U23728 ( .A1(n20800), .A2(\xmem_data[30][0] ), .B1(n17043), .B2(
        \xmem_data[31][0] ), .ZN(n19693) );
  NAND4_X1 U23729 ( .A1(n19696), .A2(n19695), .A3(n19694), .A4(n19693), .ZN(
        n19697) );
  NAND4_X1 U23730 ( .A1(n3825), .A2(n19700), .A3(n19699), .A4(n19698), .ZN(
        n19701) );
  NAND2_X1 U23731 ( .A1(n19701), .A2(n20795), .ZN(n19702) );
  XNOR2_X1 U23732 ( .A(n34624), .B(\fmem_data[28][7] ), .ZN(n19706) );
  OAI22_X1 U23733 ( .A1(n31951), .A2(n35761), .B1(n35760), .B2(n19706), .ZN(
        n23167) );
  XNOR2_X1 U23734 ( .A(n31673), .B(\fmem_data[10][3] ), .ZN(n31949) );
  XNOR2_X1 U23735 ( .A(n35399), .B(\fmem_data[28][1] ), .ZN(n31959) );
  XNOR2_X1 U23736 ( .A(n31657), .B(\fmem_data[28][1] ), .ZN(n30981) );
  OAI22_X1 U23737 ( .A1(n31959), .A2(n3562), .B1(n30981), .B2(n34745), .ZN(
        n23588) );
  AOI22_X1 U23738 ( .A1(n28500), .A2(\xmem_data[32][3] ), .B1(n20577), .B2(
        \xmem_data[33][3] ), .ZN(n19710) );
  AOI22_X1 U23739 ( .A1(n20579), .A2(\xmem_data[34][3] ), .B1(n25686), .B2(
        \xmem_data[35][3] ), .ZN(n19709) );
  AOI22_X1 U23740 ( .A1(n20578), .A2(\xmem_data[36][3] ), .B1(n3153), .B2(
        \xmem_data[37][3] ), .ZN(n19708) );
  AOI22_X1 U23741 ( .A1(n3247), .A2(\xmem_data[38][3] ), .B1(n20576), .B2(
        \xmem_data[39][3] ), .ZN(n19707) );
  NAND4_X1 U23742 ( .A1(n19710), .A2(n19709), .A3(n19708), .A4(n19707), .ZN(
        n19727) );
  AOI22_X1 U23743 ( .A1(n20588), .A2(\xmem_data[48][3] ), .B1(n20587), .B2(
        \xmem_data[49][3] ), .ZN(n19714) );
  AOI22_X1 U23744 ( .A1(n22740), .A2(\xmem_data[50][3] ), .B1(n31268), .B2(
        \xmem_data[51][3] ), .ZN(n19713) );
  AOI22_X1 U23745 ( .A1(n20584), .A2(\xmem_data[52][3] ), .B1(n29807), .B2(
        \xmem_data[53][3] ), .ZN(n19712) );
  AOI22_X1 U23746 ( .A1(n20586), .A2(\xmem_data[54][3] ), .B1(n20585), .B2(
        \xmem_data[55][3] ), .ZN(n19711) );
  NAND4_X1 U23747 ( .A1(n19714), .A2(n19713), .A3(n19712), .A4(n19711), .ZN(
        n19725) );
  AOI22_X1 U23748 ( .A1(n24707), .A2(\xmem_data[56][3] ), .B1(n30950), .B2(
        \xmem_data[57][3] ), .ZN(n19718) );
  AOI22_X1 U23749 ( .A1(n20814), .A2(\xmem_data[58][3] ), .B1(n3326), .B2(
        \xmem_data[59][3] ), .ZN(n19717) );
  AOI22_X1 U23750 ( .A1(n30898), .A2(\xmem_data[60][3] ), .B1(n3307), .B2(
        \xmem_data[61][3] ), .ZN(n19716) );
  AOI22_X1 U23751 ( .A1(n24570), .A2(\xmem_data[62][3] ), .B1(n28293), .B2(
        \xmem_data[63][3] ), .ZN(n19715) );
  NAND4_X1 U23752 ( .A1(n19718), .A2(n19717), .A3(n19716), .A4(n19715), .ZN(
        n19724) );
  AOI22_X1 U23753 ( .A1(n3221), .A2(\xmem_data[40][3] ), .B1(n25414), .B2(
        \xmem_data[41][3] ), .ZN(n19722) );
  AOI22_X1 U23754 ( .A1(n20598), .A2(\xmem_data[42][3] ), .B1(n20725), .B2(
        \xmem_data[43][3] ), .ZN(n19721) );
  AOI22_X1 U23755 ( .A1(n29181), .A2(\xmem_data[44][3] ), .B1(n20808), .B2(
        \xmem_data[45][3] ), .ZN(n19720) );
  AOI22_X1 U23756 ( .A1(n25514), .A2(\xmem_data[46][3] ), .B1(n25422), .B2(
        \xmem_data[47][3] ), .ZN(n19719) );
  NAND4_X1 U23757 ( .A1(n19722), .A2(n19721), .A3(n19720), .A4(n19719), .ZN(
        n19723) );
  OR3_X1 U23758 ( .A1(n19725), .A2(n19724), .A3(n19723), .ZN(n19726) );
  OAI21_X1 U23759 ( .B1(n19727), .B2(n19726), .A(n20606), .ZN(n19810) );
  AOI22_X1 U23760 ( .A1(n30861), .A2(\xmem_data[68][3] ), .B1(n3414), .B2(
        \xmem_data[69][3] ), .ZN(n19730) );
  AND2_X1 U23761 ( .A1(n20568), .A2(\xmem_data[70][3] ), .ZN(n19728) );
  AOI21_X1 U23762 ( .B1(n25508), .B2(\xmem_data[71][3] ), .A(n19728), .ZN(
        n19729) );
  AOI22_X1 U23763 ( .A1(n3219), .A2(\xmem_data[72][3] ), .B1(n24632), .B2(
        \xmem_data[73][3] ), .ZN(n19734) );
  AOI22_X1 U23764 ( .A1(n20558), .A2(\xmem_data[74][3] ), .B1(n20725), .B2(
        \xmem_data[75][3] ), .ZN(n19733) );
  AOI22_X1 U23765 ( .A1(n20559), .A2(\xmem_data[76][3] ), .B1(n29231), .B2(
        \xmem_data[77][3] ), .ZN(n19732) );
  AOI22_X1 U23766 ( .A1(n27446), .A2(\xmem_data[78][3] ), .B1(n25422), .B2(
        \xmem_data[79][3] ), .ZN(n19731) );
  NAND4_X1 U23767 ( .A1(n19734), .A2(n19733), .A3(n19732), .A4(n19731), .ZN(
        n19741) );
  AOI22_X1 U23768 ( .A1(n20553), .A2(\xmem_data[94][3] ), .B1(n20552), .B2(
        \xmem_data[95][3] ), .ZN(n19736) );
  AOI22_X1 U23769 ( .A1(n29048), .A2(\xmem_data[88][3] ), .B1(n30617), .B2(
        \xmem_data[89][3] ), .ZN(n19735) );
  AOI22_X1 U23770 ( .A1(n20551), .A2(\xmem_data[92][3] ), .B1(n24623), .B2(
        \xmem_data[93][3] ), .ZN(n19738) );
  AOI22_X1 U23771 ( .A1(n27920), .A2(\xmem_data[90][3] ), .B1(n30956), .B2(
        \xmem_data[91][3] ), .ZN(n19737) );
  NAND3_X1 U23772 ( .A1(n19739), .A2(n19738), .A3(n19737), .ZN(n19740) );
  NOR2_X1 U23773 ( .A1(n19741), .A2(n19740), .ZN(n19752) );
  AOI22_X1 U23774 ( .A1(n29136), .A2(\xmem_data[64][3] ), .B1(n20567), .B2(
        \xmem_data[65][3] ), .ZN(n19751) );
  AOI22_X1 U23775 ( .A1(n24448), .A2(\xmem_data[82][3] ), .B1(n24131), .B2(
        \xmem_data[83][3] ), .ZN(n19743) );
  AOI22_X1 U23776 ( .A1(n20544), .A2(\xmem_data[84][3] ), .B1(n27818), .B2(
        \xmem_data[85][3] ), .ZN(n19742) );
  NAND2_X1 U23777 ( .A1(n19743), .A2(n19742), .ZN(n19749) );
  AOI22_X1 U23778 ( .A1(n20543), .A2(\xmem_data[86][3] ), .B1(n20542), .B2(
        \xmem_data[87][3] ), .ZN(n19744) );
  INV_X1 U23779 ( .A(n19744), .ZN(n19748) );
  AOI22_X1 U23780 ( .A1(n20546), .A2(\xmem_data[80][3] ), .B1(n20545), .B2(
        \xmem_data[81][3] ), .ZN(n19746) );
  AOI22_X1 U23781 ( .A1(n21059), .A2(\xmem_data[66][3] ), .B1(n30909), .B2(
        \xmem_data[67][3] ), .ZN(n19745) );
  NAND2_X1 U23782 ( .A1(n19746), .A2(n19745), .ZN(n19747) );
  NOR3_X1 U23783 ( .A1(n19749), .A2(n19748), .A3(n19747), .ZN(n19750) );
  NAND4_X1 U23784 ( .A1(n19753), .A2(n19752), .A3(n19751), .A4(n19750), .ZN(
        n19755) );
  NOR2_X1 U23785 ( .A1(n3232), .A2(n39022), .ZN(n19754) );
  AOI21_X1 U23786 ( .B1(n19755), .B2(n20573), .A(n3891), .ZN(n19809) );
  AOI22_X1 U23787 ( .A1(n3218), .A2(\xmem_data[8][3] ), .B1(n29422), .B2(
        \xmem_data[9][3] ), .ZN(n19762) );
  AOI22_X1 U23788 ( .A1(n20993), .A2(\xmem_data[12][3] ), .B1(n27396), .B2(
        \xmem_data[13][3] ), .ZN(n19756) );
  INV_X1 U23789 ( .A(n19756), .ZN(n19760) );
  AOI22_X1 U23790 ( .A1(n20500), .A2(\xmem_data[10][3] ), .B1(n22758), .B2(
        \xmem_data[11][3] ), .ZN(n19758) );
  NAND2_X1 U23791 ( .A1(n24450), .A2(\xmem_data[15][3] ), .ZN(n19757) );
  NAND2_X1 U23792 ( .A1(n19758), .A2(n19757), .ZN(n19759) );
  NOR2_X1 U23793 ( .A1(n19760), .A2(n19759), .ZN(n19761) );
  NAND2_X1 U23794 ( .A1(n19762), .A2(n19761), .ZN(n19773) );
  AOI22_X1 U23795 ( .A1(n20505), .A2(\xmem_data[24][3] ), .B1(n28687), .B2(
        \xmem_data[25][3] ), .ZN(n19766) );
  AOI22_X1 U23796 ( .A1(n13481), .A2(\xmem_data[26][3] ), .B1(n3325), .B2(
        \xmem_data[27][3] ), .ZN(n19765) );
  AOI22_X1 U23797 ( .A1(n30598), .A2(\xmem_data[28][3] ), .B1(n30686), .B2(
        \xmem_data[29][3] ), .ZN(n19764) );
  AOI22_X1 U23798 ( .A1(n20507), .A2(\xmem_data[30][3] ), .B1(n30497), .B2(
        \xmem_data[31][3] ), .ZN(n19763) );
  NAND4_X1 U23799 ( .A1(n19766), .A2(n19765), .A3(n19764), .A4(n19763), .ZN(
        n19772) );
  AOI22_X1 U23800 ( .A1(n30854), .A2(\xmem_data[16][3] ), .B1(n28051), .B2(
        \xmem_data[17][3] ), .ZN(n19770) );
  AOI22_X1 U23801 ( .A1(n24132), .A2(\xmem_data[18][3] ), .B1(n20541), .B2(
        \xmem_data[19][3] ), .ZN(n19769) );
  AOI22_X1 U23802 ( .A1(n25606), .A2(\xmem_data[20][3] ), .B1(n20939), .B2(
        \xmem_data[21][3] ), .ZN(n19768) );
  AOI22_X1 U23803 ( .A1(n28993), .A2(\xmem_data[22][3] ), .B1(n27919), .B2(
        \xmem_data[23][3] ), .ZN(n19767) );
  NAND4_X1 U23804 ( .A1(n19770), .A2(n19769), .A3(n19768), .A4(n19767), .ZN(
        n19771) );
  OR3_X1 U23805 ( .A1(n19773), .A2(n19772), .A3(n19771), .ZN(n19781) );
  AOI22_X1 U23806 ( .A1(n20488), .A2(\xmem_data[0][3] ), .B1(n27717), .B2(
        \xmem_data[1][3] ), .ZN(n19779) );
  AOI22_X1 U23807 ( .A1(n20489), .A2(\xmem_data[4][3] ), .B1(n3144), .B2(
        \xmem_data[5][3] ), .ZN(n19778) );
  AND2_X1 U23808 ( .A1(n20711), .A2(\xmem_data[6][3] ), .ZN(n19776) );
  AOI22_X1 U23809 ( .A1(n29125), .A2(\xmem_data[2][3] ), .B1(n24526), .B2(
        \xmem_data[3][3] ), .ZN(n19774) );
  INV_X1 U23810 ( .A(n19774), .ZN(n19775) );
  AOI211_X1 U23811 ( .C1(n20518), .C2(\xmem_data[7][3] ), .A(n19776), .B(
        n19775), .ZN(n19777) );
  NAND3_X1 U23812 ( .A1(n19779), .A2(n19778), .A3(n19777), .ZN(n19780) );
  OAI21_X1 U23813 ( .B1(n19781), .B2(n19780), .A(n20515), .ZN(n19808) );
  AOI22_X1 U23814 ( .A1(n3219), .A2(\xmem_data[104][3] ), .B1(n29789), .B2(
        \xmem_data[105][3] ), .ZN(n19785) );
  AOI22_X1 U23815 ( .A1(n20558), .A2(\xmem_data[106][3] ), .B1(n20725), .B2(
        \xmem_data[107][3] ), .ZN(n19784) );
  AOI22_X1 U23816 ( .A1(n20559), .A2(\xmem_data[108][3] ), .B1(n3281), .B2(
        \xmem_data[109][3] ), .ZN(n19783) );
  AOI22_X1 U23817 ( .A1(n25450), .A2(\xmem_data[110][3] ), .B1(n30551), .B2(
        \xmem_data[111][3] ), .ZN(n19782) );
  AOI22_X1 U23818 ( .A1(n25357), .A2(\xmem_data[100][3] ), .B1(n24693), .B2(
        \xmem_data[101][3] ), .ZN(n19802) );
  AOI22_X1 U23819 ( .A1(n24592), .A2(\xmem_data[122][3] ), .B1(n27974), .B2(
        \xmem_data[123][3] ), .ZN(n19786) );
  INV_X1 U23820 ( .A(n19786), .ZN(n19791) );
  AOI22_X1 U23821 ( .A1(n20551), .A2(\xmem_data[124][3] ), .B1(n30600), .B2(
        \xmem_data[125][3] ), .ZN(n19789) );
  AOI22_X1 U23822 ( .A1(n20553), .A2(\xmem_data[126][3] ), .B1(n20552), .B2(
        \xmem_data[127][3] ), .ZN(n19788) );
  AOI22_X1 U23823 ( .A1(n20505), .A2(\xmem_data[120][3] ), .B1(n29047), .B2(
        \xmem_data[121][3] ), .ZN(n19787) );
  NOR2_X1 U23824 ( .A1(n19791), .A2(n19790), .ZN(n19801) );
  AOI22_X1 U23825 ( .A1(n27452), .A2(\xmem_data[114][3] ), .B1(n30891), .B2(
        \xmem_data[115][3] ), .ZN(n19793) );
  AOI22_X1 U23826 ( .A1(n20544), .A2(\xmem_data[116][3] ), .B1(n25607), .B2(
        \xmem_data[117][3] ), .ZN(n19792) );
  NAND2_X1 U23827 ( .A1(n19793), .A2(n19792), .ZN(n19799) );
  AOI22_X1 U23828 ( .A1(n20543), .A2(\xmem_data[118][3] ), .B1(n20542), .B2(
        \xmem_data[119][3] ), .ZN(n19794) );
  INV_X1 U23829 ( .A(n19794), .ZN(n19798) );
  AOI22_X1 U23830 ( .A1(n20546), .A2(\xmem_data[112][3] ), .B1(n20545), .B2(
        \xmem_data[113][3] ), .ZN(n19796) );
  AOI22_X1 U23831 ( .A1(n27435), .A2(\xmem_data[98][3] ), .B1(n24688), .B2(
        \xmem_data[99][3] ), .ZN(n19795) );
  NAND2_X1 U23832 ( .A1(n19796), .A2(n19795), .ZN(n19797) );
  NOR3_X1 U23833 ( .A1(n19799), .A2(n19798), .A3(n19797), .ZN(n19800) );
  NAND4_X1 U23834 ( .A1(n3853), .A2(n19802), .A3(n19801), .A4(n19800), .ZN(
        n19806) );
  AOI22_X1 U23835 ( .A1(n20568), .A2(\xmem_data[102][3] ), .B1(n20518), .B2(
        \xmem_data[103][3] ), .ZN(n19804) );
  AOI22_X1 U23836 ( .A1(n28979), .A2(\xmem_data[96][3] ), .B1(n20567), .B2(
        \xmem_data[97][3] ), .ZN(n19803) );
  NAND2_X1 U23837 ( .A1(n19804), .A2(n19803), .ZN(n19805) );
  OAI21_X1 U23838 ( .B1(n19806), .B2(n19805), .A(n20538), .ZN(n19807) );
  NAND4_X1 U23839 ( .A1(n19810), .A2(n19809), .A3(n19808), .A4(n19807), .ZN(
        n32115) );
  XNOR2_X1 U23840 ( .A(n32115), .B(\fmem_data[21][5] ), .ZN(n33270) );
  AOI22_X1 U23841 ( .A1(n30496), .A2(\xmem_data[32][2] ), .B1(n20577), .B2(
        \xmem_data[33][2] ), .ZN(n19814) );
  AOI22_X1 U23842 ( .A1(n20579), .A2(\xmem_data[34][2] ), .B1(n24607), .B2(
        \xmem_data[35][2] ), .ZN(n19813) );
  AOI22_X1 U23843 ( .A1(n20578), .A2(\xmem_data[36][2] ), .B1(n3142), .B2(
        \xmem_data[37][2] ), .ZN(n19812) );
  AOI22_X1 U23844 ( .A1(n30589), .A2(\xmem_data[38][2] ), .B1(n20576), .B2(
        \xmem_data[39][2] ), .ZN(n19811) );
  NAND4_X1 U23845 ( .A1(n19814), .A2(n19813), .A3(n19812), .A4(n19811), .ZN(
        n19830) );
  AOI22_X1 U23846 ( .A1(n3218), .A2(\xmem_data[40][2] ), .B1(n29422), .B2(
        \xmem_data[41][2] ), .ZN(n19818) );
  AOI22_X1 U23847 ( .A1(n20598), .A2(\xmem_data[42][2] ), .B1(n23741), .B2(
        \xmem_data[43][2] ), .ZN(n19817) );
  AOI22_X1 U23848 ( .A1(n28372), .A2(\xmem_data[44][2] ), .B1(n3147), .B2(
        \xmem_data[45][2] ), .ZN(n19816) );
  AOI22_X1 U23849 ( .A1(n28007), .A2(\xmem_data[46][2] ), .B1(n24554), .B2(
        \xmem_data[47][2] ), .ZN(n19815) );
  NAND4_X1 U23850 ( .A1(n19818), .A2(n19817), .A3(n19816), .A4(n19815), .ZN(
        n19829) );
  AOI22_X1 U23851 ( .A1(n20588), .A2(\xmem_data[48][2] ), .B1(n20587), .B2(
        \xmem_data[49][2] ), .ZN(n19822) );
  AOI22_X1 U23852 ( .A1(n24212), .A2(\xmem_data[50][2] ), .B1(n28980), .B2(
        \xmem_data[51][2] ), .ZN(n19821) );
  AOI22_X1 U23853 ( .A1(n20584), .A2(\xmem_data[52][2] ), .B1(n28091), .B2(
        \xmem_data[53][2] ), .ZN(n19820) );
  AOI22_X1 U23854 ( .A1(n20586), .A2(\xmem_data[54][2] ), .B1(n20585), .B2(
        \xmem_data[55][2] ), .ZN(n19819) );
  NAND4_X1 U23855 ( .A1(n19822), .A2(n19821), .A3(n19820), .A4(n19819), .ZN(
        n19828) );
  AOI22_X1 U23856 ( .A1(n24459), .A2(\xmem_data[56][2] ), .B1(n21008), .B2(
        \xmem_data[57][2] ), .ZN(n19826) );
  AOI22_X1 U23857 ( .A1(n29101), .A2(\xmem_data[58][2] ), .B1(n24220), .B2(
        \xmem_data[59][2] ), .ZN(n19825) );
  AOI22_X1 U23858 ( .A1(n27856), .A2(\xmem_data[60][2] ), .B1(n28461), .B2(
        \xmem_data[61][2] ), .ZN(n19824) );
  AOI22_X1 U23859 ( .A1(n31362), .A2(\xmem_data[62][2] ), .B1(n13486), .B2(
        \xmem_data[63][2] ), .ZN(n19823) );
  NAND4_X1 U23860 ( .A1(n19826), .A2(n19825), .A3(n19824), .A4(n19823), .ZN(
        n19827) );
  OR4_X1 U23861 ( .A1(n19830), .A2(n19829), .A3(n19828), .A4(n19827), .ZN(
        n19857) );
  AOI22_X1 U23862 ( .A1(n20488), .A2(\xmem_data[0][2] ), .B1(n28772), .B2(
        \xmem_data[1][2] ), .ZN(n19835) );
  AOI22_X1 U23863 ( .A1(n30900), .A2(\xmem_data[2][2] ), .B1(n24607), .B2(
        \xmem_data[3][2] ), .ZN(n19834) );
  AOI22_X1 U23864 ( .A1(n20489), .A2(\xmem_data[4][2] ), .B1(n3229), .B2(
        \xmem_data[5][2] ), .ZN(n19833) );
  AND2_X1 U23865 ( .A1(n24439), .A2(\xmem_data[6][2] ), .ZN(n19831) );
  AOI21_X1 U23866 ( .B1(n20518), .B2(\xmem_data[7][2] ), .A(n19831), .ZN(
        n19832) );
  AOI22_X1 U23867 ( .A1(n30882), .A2(\xmem_data[12][2] ), .B1(n30295), .B2(
        \xmem_data[13][2] ), .ZN(n19842) );
  AOI22_X1 U23868 ( .A1(n3221), .A2(\xmem_data[8][2] ), .B1(n23740), .B2(
        \xmem_data[9][2] ), .ZN(n19836) );
  INV_X1 U23869 ( .A(n19836), .ZN(n19840) );
  AOI22_X1 U23870 ( .A1(n20500), .A2(\xmem_data[10][2] ), .B1(n20994), .B2(
        \xmem_data[11][2] ), .ZN(n19837) );
  INV_X1 U23871 ( .A(n19837), .ZN(n19839) );
  AND2_X1 U23872 ( .A1(n20961), .A2(\xmem_data[15][2] ), .ZN(n19838) );
  NOR3_X1 U23873 ( .A1(n19840), .A2(n19839), .A3(n19838), .ZN(n19841) );
  NAND2_X1 U23874 ( .A1(n19842), .A2(n19841), .ZN(n19854) );
  AOI22_X1 U23875 ( .A1(n30854), .A2(\xmem_data[16][2] ), .B1(n25424), .B2(
        \xmem_data[17][2] ), .ZN(n19846) );
  AOI22_X1 U23876 ( .A1(n31326), .A2(\xmem_data[18][2] ), .B1(n29023), .B2(
        \xmem_data[19][2] ), .ZN(n19845) );
  AOI22_X1 U23877 ( .A1(n24597), .A2(\xmem_data[20][2] ), .B1(n25519), .B2(
        \xmem_data[21][2] ), .ZN(n19844) );
  AOI22_X1 U23878 ( .A1(n3213), .A2(\xmem_data[22][2] ), .B1(n29010), .B2(
        \xmem_data[23][2] ), .ZN(n19843) );
  NAND4_X1 U23879 ( .A1(n19846), .A2(n19845), .A3(n19844), .A4(n19843), .ZN(
        n19852) );
  AOI22_X1 U23880 ( .A1(n27856), .A2(\xmem_data[28][2] ), .B1(n25636), .B2(
        \xmem_data[29][2] ), .ZN(n19850) );
  AOI22_X1 U23881 ( .A1(n20505), .A2(\xmem_data[24][2] ), .B1(n28994), .B2(
        \xmem_data[25][2] ), .ZN(n19849) );
  AOI22_X1 U23882 ( .A1(n20507), .A2(\xmem_data[30][2] ), .B1(n22684), .B2(
        \xmem_data[31][2] ), .ZN(n19848) );
  AOI22_X1 U23883 ( .A1(n3324), .A2(\xmem_data[27][2] ), .B1(n13481), .B2(
        \xmem_data[26][2] ), .ZN(n19847) );
  NAND4_X1 U23884 ( .A1(n19850), .A2(n19849), .A3(n19848), .A4(n19847), .ZN(
        n19851) );
  OR3_X1 U23885 ( .A1(n19852), .A2(n3914), .A3(n19851), .ZN(n19853) );
  NOR2_X1 U23886 ( .A1(n19854), .A2(n19853), .ZN(n19855) );
  AOI21_X1 U23887 ( .B1(n3758), .B2(n19855), .A(n3232), .ZN(n19856) );
  AOI21_X1 U23888 ( .B1(n19857), .B2(n20606), .A(n19856), .ZN(n19904) );
  AOI22_X1 U23889 ( .A1(n11008), .A2(\xmem_data[96][2] ), .B1(n20567), .B2(
        \xmem_data[97][2] ), .ZN(n19862) );
  AOI22_X1 U23890 ( .A1(n13487), .A2(\xmem_data[98][2] ), .B1(n27959), .B2(
        \xmem_data[99][2] ), .ZN(n19861) );
  AOI22_X1 U23891 ( .A1(n29118), .A2(\xmem_data[100][2] ), .B1(n25725), .B2(
        \xmem_data[101][2] ), .ZN(n19860) );
  AOI21_X1 U23892 ( .B1(n20518), .B2(\xmem_data[103][2] ), .A(n19858), .ZN(
        n19859) );
  NAND4_X1 U23893 ( .A1(n19862), .A2(n19861), .A3(n19860), .A4(n19859), .ZN(
        n19878) );
  AOI22_X1 U23894 ( .A1(n3222), .A2(\xmem_data[104][2] ), .B1(n28733), .B2(
        \xmem_data[105][2] ), .ZN(n19866) );
  AOI22_X1 U23895 ( .A1(n20558), .A2(\xmem_data[106][2] ), .B1(n25694), .B2(
        \xmem_data[107][2] ), .ZN(n19865) );
  AOI22_X1 U23896 ( .A1(n20559), .A2(\xmem_data[108][2] ), .B1(n3140), .B2(
        \xmem_data[109][2] ), .ZN(n19864) );
  AOI22_X1 U23897 ( .A1(n25450), .A2(\xmem_data[110][2] ), .B1(n25670), .B2(
        \xmem_data[111][2] ), .ZN(n19863) );
  NAND4_X1 U23898 ( .A1(n19866), .A2(n19865), .A3(n19864), .A4(n19863), .ZN(
        n19877) );
  AOI22_X1 U23899 ( .A1(n20546), .A2(\xmem_data[112][2] ), .B1(n20545), .B2(
        \xmem_data[113][2] ), .ZN(n19870) );
  AOI22_X1 U23900 ( .A1(n24516), .A2(\xmem_data[114][2] ), .B1(n28980), .B2(
        \xmem_data[115][2] ), .ZN(n19869) );
  AOI22_X1 U23901 ( .A1(n20544), .A2(\xmem_data[116][2] ), .B1(n30892), .B2(
        \xmem_data[117][2] ), .ZN(n19868) );
  AOI22_X1 U23902 ( .A1(n20543), .A2(\xmem_data[118][2] ), .B1(n20542), .B2(
        \xmem_data[119][2] ), .ZN(n19867) );
  NAND4_X1 U23903 ( .A1(n19870), .A2(n19869), .A3(n19868), .A4(n19867), .ZN(
        n19876) );
  AOI22_X1 U23904 ( .A1(n30544), .A2(\xmem_data[120][2] ), .B1(n16990), .B2(
        \xmem_data[121][2] ), .ZN(n19874) );
  AOI22_X1 U23905 ( .A1(n28301), .A2(\xmem_data[122][2] ), .B1(n24511), .B2(
        \xmem_data[123][2] ), .ZN(n19873) );
  AOI22_X1 U23906 ( .A1(n20551), .A2(\xmem_data[124][2] ), .B1(n3329), .B2(
        \xmem_data[125][2] ), .ZN(n19872) );
  AOI22_X1 U23907 ( .A1(n20553), .A2(\xmem_data[126][2] ), .B1(n20552), .B2(
        \xmem_data[127][2] ), .ZN(n19871) );
  NAND4_X1 U23908 ( .A1(n19874), .A2(n19873), .A3(n19872), .A4(n19871), .ZN(
        n19875) );
  OR4_X1 U23909 ( .A1(n19878), .A2(n19877), .A3(n19876), .A4(n19875), .ZN(
        n19902) );
  AND2_X1 U23910 ( .A1(n17049), .A2(\xmem_data[64][2] ), .ZN(n19879) );
  AOI21_X1 U23911 ( .B1(n20567), .B2(\xmem_data[65][2] ), .A(n19879), .ZN(
        n19884) );
  AOI22_X1 U23912 ( .A1(n31344), .A2(\xmem_data[66][2] ), .B1(n28076), .B2(
        \xmem_data[67][2] ), .ZN(n19883) );
  AOI22_X1 U23913 ( .A1(n30861), .A2(\xmem_data[68][2] ), .B1(n28039), .B2(
        \xmem_data[69][2] ), .ZN(n19882) );
  AND2_X1 U23914 ( .A1(n20568), .A2(\xmem_data[70][2] ), .ZN(n19880) );
  AOI21_X1 U23915 ( .B1(n20518), .B2(\xmem_data[71][2] ), .A(n19880), .ZN(
        n19881) );
  NAND4_X1 U23916 ( .A1(n19884), .A2(n19883), .A3(n19882), .A4(n19881), .ZN(
        n19900) );
  AOI22_X1 U23917 ( .A1(n3222), .A2(\xmem_data[72][2] ), .B1(n30964), .B2(
        \xmem_data[73][2] ), .ZN(n19888) );
  AOI22_X1 U23918 ( .A1(n20558), .A2(\xmem_data[74][2] ), .B1(n3322), .B2(
        \xmem_data[75][2] ), .ZN(n19887) );
  AOI22_X1 U23919 ( .A1(n20559), .A2(\xmem_data[76][2] ), .B1(n29350), .B2(
        \xmem_data[77][2] ), .ZN(n19886) );
  AOI22_X1 U23920 ( .A1(n25450), .A2(\xmem_data[78][2] ), .B1(n20961), .B2(
        \xmem_data[79][2] ), .ZN(n19885) );
  NAND4_X1 U23921 ( .A1(n19888), .A2(n19887), .A3(n19886), .A4(n19885), .ZN(
        n19899) );
  AOI22_X1 U23922 ( .A1(n20546), .A2(\xmem_data[80][2] ), .B1(n20545), .B2(
        \xmem_data[81][2] ), .ZN(n19892) );
  AOI22_X1 U23923 ( .A1(n25423), .A2(\xmem_data[82][2] ), .B1(n30891), .B2(
        \xmem_data[83][2] ), .ZN(n19891) );
  AOI22_X1 U23924 ( .A1(n20544), .A2(\xmem_data[84][2] ), .B1(n29237), .B2(
        \xmem_data[85][2] ), .ZN(n19890) );
  AOI22_X1 U23925 ( .A1(n20543), .A2(\xmem_data[86][2] ), .B1(n20542), .B2(
        \xmem_data[87][2] ), .ZN(n19889) );
  NAND4_X1 U23926 ( .A1(n19892), .A2(n19891), .A3(n19890), .A4(n19889), .ZN(
        n19898) );
  AOI22_X1 U23927 ( .A1(n30544), .A2(\xmem_data[88][2] ), .B1(n21008), .B2(
        \xmem_data[89][2] ), .ZN(n19896) );
  AOI22_X1 U23928 ( .A1(n30545), .A2(\xmem_data[90][2] ), .B1(n30849), .B2(
        \xmem_data[91][2] ), .ZN(n19895) );
  AOI22_X1 U23929 ( .A1(n20551), .A2(\xmem_data[92][2] ), .B1(n29054), .B2(
        \xmem_data[93][2] ), .ZN(n19894) );
  AOI22_X1 U23930 ( .A1(n20553), .A2(\xmem_data[94][2] ), .B1(n20552), .B2(
        \xmem_data[95][2] ), .ZN(n19893) );
  NAND4_X1 U23931 ( .A1(n19896), .A2(n19895), .A3(n19894), .A4(n19893), .ZN(
        n19897) );
  OR4_X1 U23932 ( .A1(n19900), .A2(n19899), .A3(n19898), .A4(n19897), .ZN(
        n19901) );
  AOI22_X1 U23933 ( .A1(n20538), .A2(n19902), .B1(n20573), .B2(n19901), .ZN(
        n19903) );
  XNOR2_X1 U23934 ( .A(n32057), .B(\fmem_data[21][5] ), .ZN(n32221) );
  OAI22_X1 U23935 ( .A1(n33270), .A2(n34195), .B1(n32221), .B2(n34194), .ZN(
        n23587) );
  NAND2_X1 U23936 ( .A1(n25514), .A2(\xmem_data[25][6] ), .ZN(n19938) );
  AOI22_X1 U23937 ( .A1(n3176), .A2(\xmem_data[30][6] ), .B1(n30513), .B2(
        \xmem_data[31][6] ), .ZN(n19906) );
  INV_X1 U23938 ( .A(n19906), .ZN(n19910) );
  AOI22_X1 U23939 ( .A1(n25422), .A2(\xmem_data[26][6] ), .B1(n20982), .B2(
        \xmem_data[27][6] ), .ZN(n19908) );
  NAND2_X1 U23940 ( .A1(n29350), .A2(\xmem_data[24][6] ), .ZN(n19907) );
  NAND2_X1 U23941 ( .A1(n19908), .A2(n19907), .ZN(n19909) );
  NOR2_X1 U23942 ( .A1(n19910), .A2(n19909), .ZN(n19919) );
  NAND2_X1 U23943 ( .A1(n20985), .A2(\xmem_data[12][6] ), .ZN(n19918) );
  AOI22_X1 U23944 ( .A1(n27453), .A2(\xmem_data[28][6] ), .B1(n21015), .B2(
        \xmem_data[29][6] ), .ZN(n19911) );
  INV_X1 U23945 ( .A(n19911), .ZN(n19916) );
  NAND2_X1 U23946 ( .A1(n16999), .A2(\xmem_data[13][6] ), .ZN(n19914) );
  AND2_X1 U23947 ( .A1(n20986), .A2(\xmem_data[14][6] ), .ZN(n19912) );
  AOI21_X1 U23948 ( .B1(n3217), .B2(\xmem_data[19][6] ), .A(n19912), .ZN(
        n19913) );
  NAND2_X1 U23949 ( .A1(n19914), .A2(n19913), .ZN(n19915) );
  NOR2_X1 U23950 ( .A1(n19916), .A2(n19915), .ZN(n19917) );
  AOI22_X1 U23951 ( .A1(n21005), .A2(\xmem_data[0][6] ), .B1(n25574), .B2(
        \xmem_data[1][6] ), .ZN(n19923) );
  AOI22_X1 U23952 ( .A1(n21007), .A2(\xmem_data[2][6] ), .B1(n21006), .B2(
        \xmem_data[3][6] ), .ZN(n19922) );
  AOI22_X1 U23953 ( .A1(n21008), .A2(\xmem_data[4][6] ), .B1(n25576), .B2(
        \xmem_data[5][6] ), .ZN(n19921) );
  AOI22_X1 U23954 ( .A1(n21010), .A2(\xmem_data[6][6] ), .B1(n21051), .B2(
        \xmem_data[7][6] ), .ZN(n19920) );
  AOI22_X1 U23955 ( .A1(n24563), .A2(\xmem_data[20][6] ), .B1(n20992), .B2(
        \xmem_data[21][6] ), .ZN(n19926) );
  AOI22_X1 U23956 ( .A1(n24606), .A2(\xmem_data[10][6] ), .B1(n21057), .B2(
        \xmem_data[11][6] ), .ZN(n19925) );
  AOI22_X1 U23957 ( .A1(n3317), .A2(\xmem_data[16][6] ), .B1(n22753), .B2(
        \xmem_data[17][6] ), .ZN(n19924) );
  AOI22_X1 U23958 ( .A1(n20994), .A2(\xmem_data[22][6] ), .B1(n20993), .B2(
        \xmem_data[23][6] ), .ZN(n19927) );
  INV_X1 U23959 ( .A(n19927), .ZN(n19928) );
  NOR2_X1 U23960 ( .A1(n19929), .A2(n19928), .ZN(n19934) );
  NAND2_X1 U23961 ( .A1(n20991), .A2(\xmem_data[18][6] ), .ZN(n19933) );
  NAND2_X1 U23962 ( .A1(n24525), .A2(\xmem_data[15][6] ), .ZN(n19931) );
  AOI22_X1 U23963 ( .A1(n20984), .A2(\xmem_data[8][6] ), .B1(n20983), .B2(
        \xmem_data[9][6] ), .ZN(n19930) );
  NOR3_X1 U23964 ( .A1(n19936), .A2(n3989), .A3(n19935), .ZN(n19937) );
  AOI21_X1 U23965 ( .B1(n19938), .B2(n19937), .A(n20386), .ZN(n19939) );
  INV_X1 U23966 ( .A(n19939), .ZN(n20005) );
  AOI22_X1 U23967 ( .A1(n21048), .A2(\xmem_data[96][6] ), .B1(n24457), .B2(
        \xmem_data[97][6] ), .ZN(n19943) );
  AOI22_X1 U23968 ( .A1(n21007), .A2(\xmem_data[98][6] ), .B1(n28058), .B2(
        \xmem_data[99][6] ), .ZN(n19942) );
  AOI22_X1 U23969 ( .A1(n21050), .A2(\xmem_data[100][6] ), .B1(n21049), .B2(
        \xmem_data[101][6] ), .ZN(n19941) );
  AOI22_X1 U23970 ( .A1(n30557), .A2(\xmem_data[102][6] ), .B1(n25679), .B2(
        \xmem_data[103][6] ), .ZN(n19940) );
  NAND4_X1 U23971 ( .A1(n19943), .A2(n19942), .A3(n19941), .A4(n19940), .ZN(
        n19959) );
  AOI22_X1 U23972 ( .A1(n21056), .A2(\xmem_data[104][6] ), .B1(n28098), .B2(
        \xmem_data[105][6] ), .ZN(n19947) );
  AOI22_X1 U23973 ( .A1(n21058), .A2(\xmem_data[106][6] ), .B1(n21057), .B2(
        \xmem_data[107][6] ), .ZN(n19946) );
  AOI22_X1 U23974 ( .A1(n21060), .A2(\xmem_data[108][6] ), .B1(n21059), .B2(
        \xmem_data[109][6] ), .ZN(n19945) );
  AOI22_X1 U23975 ( .A1(n21061), .A2(\xmem_data[110][6] ), .B1(n28075), .B2(
        \xmem_data[111][6] ), .ZN(n19944) );
  NAND4_X1 U23976 ( .A1(n19947), .A2(n19946), .A3(n19945), .A4(n19944), .ZN(
        n19958) );
  AOI22_X1 U23977 ( .A1(n30864), .A2(\xmem_data[112][6] ), .B1(n30863), .B2(
        \xmem_data[113][6] ), .ZN(n19951) );
  AOI22_X1 U23978 ( .A1(n21066), .A2(\xmem_data[114][6] ), .B1(n3219), .B2(
        \xmem_data[115][6] ), .ZN(n19950) );
  AOI22_X1 U23979 ( .A1(n21067), .A2(\xmem_data[116][6] ), .B1(n24207), .B2(
        \xmem_data[117][6] ), .ZN(n19949) );
  AOI22_X1 U23980 ( .A1(n21069), .A2(\xmem_data[118][6] ), .B1(n21068), .B2(
        \xmem_data[119][6] ), .ZN(n19948) );
  NAND4_X1 U23981 ( .A1(n19951), .A2(n19950), .A3(n19949), .A4(n19948), .ZN(
        n19957) );
  AOI22_X1 U23982 ( .A1(n21074), .A2(\xmem_data[120][6] ), .B1(n25514), .B2(
        \xmem_data[121][6] ), .ZN(n19955) );
  AOI22_X1 U23983 ( .A1(n28972), .A2(\xmem_data[122][6] ), .B1(n25456), .B2(
        \xmem_data[123][6] ), .ZN(n19954) );
  AOI22_X1 U23984 ( .A1(n28671), .A2(\xmem_data[124][6] ), .B1(n21075), .B2(
        \xmem_data[125][6] ), .ZN(n19953) );
  AOI22_X1 U23985 ( .A1(n16986), .A2(\xmem_data[126][6] ), .B1(n21076), .B2(
        \xmem_data[127][6] ), .ZN(n19952) );
  NAND4_X1 U23986 ( .A1(n19955), .A2(n19954), .A3(n19953), .A4(n19952), .ZN(
        n19956) );
  OR4_X1 U23987 ( .A1(n19959), .A2(n19958), .A3(n19957), .A4(n19956), .ZN(
        n19981) );
  AOI22_X1 U23988 ( .A1(n20939), .A2(\xmem_data[64][6] ), .B1(n20938), .B2(
        \xmem_data[65][6] ), .ZN(n19963) );
  AOI22_X1 U23989 ( .A1(n28059), .A2(n20682), .B1(n20940), .B2(
        \xmem_data[67][6] ), .ZN(n19962) );
  AOI22_X1 U23990 ( .A1(n20942), .A2(\xmem_data[68][6] ), .B1(n20941), .B2(
        \xmem_data[69][6] ), .ZN(n19961) );
  AOI22_X1 U23991 ( .A1(n25632), .A2(\xmem_data[70][6] ), .B1(n20943), .B2(
        \xmem_data[71][6] ), .ZN(n19960) );
  NAND4_X1 U23992 ( .A1(n19963), .A2(n19962), .A3(n19961), .A4(n19960), .ZN(
        n19979) );
  AOI22_X1 U23993 ( .A1(n20950), .A2(\xmem_data[72][6] ), .B1(n20949), .B2(
        \xmem_data[73][6] ), .ZN(n19967) );
  AOI22_X1 U23994 ( .A1(n20782), .A2(\xmem_data[74][6] ), .B1(n28500), .B2(
        \xmem_data[75][6] ), .ZN(n19966) );
  AOI22_X1 U23995 ( .A1(n20952), .A2(\xmem_data[76][6] ), .B1(n20951), .B2(
        \xmem_data[77][6] ), .ZN(n19965) );
  AOI22_X1 U23996 ( .A1(n20953), .A2(\xmem_data[78][6] ), .B1(n31262), .B2(
        \xmem_data[79][6] ), .ZN(n19964) );
  NAND4_X1 U23997 ( .A1(n19967), .A2(n19966), .A3(n19965), .A4(n19964), .ZN(
        n19978) );
  AOI22_X1 U23998 ( .A1(n3388), .A2(\xmem_data[80][6] ), .B1(n20568), .B2(
        \xmem_data[81][6] ), .ZN(n19971) );
  AOI22_X1 U23999 ( .A1(n28503), .A2(\xmem_data[82][6] ), .B1(n3220), .B2(
        \xmem_data[83][6] ), .ZN(n19970) );
  AOI22_X1 U24000 ( .A1(n20724), .A2(\xmem_data[84][6] ), .B1(n23739), .B2(
        \xmem_data[85][6] ), .ZN(n19969) );
  AOI22_X1 U24001 ( .A1(n20969), .A2(\xmem_data[86][6] ), .B1(n25486), .B2(
        \xmem_data[87][6] ), .ZN(n19968) );
  NAND4_X1 U24002 ( .A1(n19971), .A2(n19970), .A3(n19969), .A4(n19968), .ZN(
        n19977) );
  AOI22_X1 U24003 ( .A1(n20962), .A2(\xmem_data[88][6] ), .B1(n28510), .B2(
        \xmem_data[89][6] ), .ZN(n19975) );
  AOI22_X1 U24004 ( .A1(n20961), .A2(\xmem_data[90][6] ), .B1(n24590), .B2(
        \xmem_data[91][6] ), .ZN(n19974) );
  AOI22_X1 U24005 ( .A1(n28671), .A2(\xmem_data[92][6] ), .B1(n20958), .B2(
        \xmem_data[93][6] ), .ZN(n19973) );
  AOI22_X1 U24006 ( .A1(n20959), .A2(\xmem_data[94][6] ), .B1(n28052), .B2(
        \xmem_data[95][6] ), .ZN(n19972) );
  NAND4_X1 U24007 ( .A1(n19975), .A2(n19974), .A3(n19973), .A4(n19972), .ZN(
        n19976) );
  OR4_X1 U24008 ( .A1(n19979), .A2(n19978), .A3(n19977), .A4(n19976), .ZN(
        n19980) );
  AOI22_X1 U24009 ( .A1(n21088), .A2(n19981), .B1(n21086), .B2(n19980), .ZN(
        n20004) );
  AOI22_X1 U24010 ( .A1(n20939), .A2(\xmem_data[32][6] ), .B1(n20938), .B2(
        \xmem_data[33][6] ), .ZN(n19985) );
  AOI22_X1 U24011 ( .A1(n24708), .A2(\xmem_data[34][6] ), .B1(n20940), .B2(
        \xmem_data[35][6] ), .ZN(n19984) );
  AOI22_X1 U24012 ( .A1(n20942), .A2(\xmem_data[36][6] ), .B1(n20941), .B2(
        \xmem_data[37][6] ), .ZN(n19983) );
  AOI22_X1 U24013 ( .A1(n25575), .A2(\xmem_data[38][6] ), .B1(n20943), .B2(
        \xmem_data[39][6] ), .ZN(n19982) );
  NAND4_X1 U24014 ( .A1(n19985), .A2(n19984), .A3(n19983), .A4(n19982), .ZN(
        n20001) );
  AOI22_X1 U24015 ( .A1(n20950), .A2(\xmem_data[40][6] ), .B1(n20949), .B2(
        \xmem_data[41][6] ), .ZN(n19989) );
  AOI22_X1 U24016 ( .A1(n20734), .A2(\xmem_data[42][6] ), .B1(n29247), .B2(
        \xmem_data[43][6] ), .ZN(n19988) );
  AOI22_X1 U24017 ( .A1(n20952), .A2(\xmem_data[44][6] ), .B1(n20951), .B2(
        \xmem_data[45][6] ), .ZN(n19987) );
  AOI22_X1 U24018 ( .A1(n20953), .A2(\xmem_data[46][6] ), .B1(n25629), .B2(
        \xmem_data[47][6] ), .ZN(n19986) );
  NAND4_X1 U24019 ( .A1(n19989), .A2(n19988), .A3(n19987), .A4(n19986), .ZN(
        n20000) );
  AOI22_X1 U24020 ( .A1(n3384), .A2(\xmem_data[48][6] ), .B1(n31347), .B2(
        \xmem_data[49][6] ), .ZN(n19993) );
  AOI22_X1 U24021 ( .A1(n25508), .A2(\xmem_data[50][6] ), .B1(n3217), .B2(
        \xmem_data[51][6] ), .ZN(n19992) );
  AOI22_X1 U24022 ( .A1(n29288), .A2(\xmem_data[52][6] ), .B1(n25562), .B2(
        \xmem_data[53][6] ), .ZN(n19991) );
  AOI22_X1 U24023 ( .A1(n20969), .A2(\xmem_data[54][6] ), .B1(n22759), .B2(
        \xmem_data[55][6] ), .ZN(n19990) );
  NAND4_X1 U24024 ( .A1(n19993), .A2(n19992), .A3(n19991), .A4(n19990), .ZN(
        n19999) );
  AOI22_X1 U24025 ( .A1(n20962), .A2(\xmem_data[56][6] ), .B1(n25514), .B2(
        \xmem_data[57][6] ), .ZN(n19997) );
  AOI22_X1 U24026 ( .A1(n20961), .A2(\xmem_data[58][6] ), .B1(n20546), .B2(
        \xmem_data[59][6] ), .ZN(n19996) );
  AOI22_X1 U24027 ( .A1(n27514), .A2(\xmem_data[60][6] ), .B1(n20958), .B2(
        \xmem_data[61][6] ), .ZN(n19995) );
  AOI22_X1 U24028 ( .A1(n20959), .A2(\xmem_data[62][6] ), .B1(n30613), .B2(
        \xmem_data[63][6] ), .ZN(n19994) );
  NAND4_X1 U24029 ( .A1(n19997), .A2(n19996), .A3(n19995), .A4(n19994), .ZN(
        n19998) );
  OR4_X1 U24030 ( .A1(n20001), .A2(n20000), .A3(n19999), .A4(n19998), .ZN(
        n20002) );
  NAND2_X1 U24031 ( .A1(n20002), .A2(n20311), .ZN(n20003) );
  XNOR2_X1 U24032 ( .A(n33039), .B(\fmem_data[0][1] ), .ZN(n23573) );
  OAI22_X1 U24033 ( .A1(n23573), .A2(n36295), .B1(n31966), .B2(n3564), .ZN(
        n23586) );
  XNOR2_X1 U24034 ( .A(n35395), .B(\fmem_data[24][1] ), .ZN(n32029) );
  AOI22_X1 U24035 ( .A1(n24630), .A2(\xmem_data[72][6] ), .B1(n3247), .B2(
        \xmem_data[73][6] ), .ZN(n20009) );
  AOI22_X1 U24036 ( .A1(n24631), .A2(\xmem_data[74][6] ), .B1(n3219), .B2(
        \xmem_data[75][6] ), .ZN(n20008) );
  AOI22_X1 U24037 ( .A1(n24632), .A2(\xmem_data[76][6] ), .B1(n25562), .B2(
        \xmem_data[77][6] ), .ZN(n20007) );
  AOI22_X1 U24038 ( .A1(n3340), .A2(\xmem_data[78][6] ), .B1(n24633), .B2(
        \xmem_data[79][6] ), .ZN(n20006) );
  NAND4_X1 U24039 ( .A1(n20009), .A2(n20008), .A3(n20007), .A4(n20006), .ZN(
        n20025) );
  AOI22_X1 U24040 ( .A1(n24623), .A2(\xmem_data[64][6] ), .B1(n24622), .B2(
        \xmem_data[65][6] ), .ZN(n20013) );
  AOI22_X1 U24041 ( .A1(n29325), .A2(n20682), .B1(n29247), .B2(
        \xmem_data[67][6] ), .ZN(n20012) );
  AOI22_X1 U24042 ( .A1(n29298), .A2(\xmem_data[68][6] ), .B1(n24624), .B2(
        \xmem_data[69][6] ), .ZN(n20011) );
  AOI22_X1 U24043 ( .A1(n24688), .A2(\xmem_data[70][6] ), .B1(n3203), .B2(
        \xmem_data[71][6] ), .ZN(n20010) );
  NAND4_X1 U24044 ( .A1(n20013), .A2(n20012), .A3(n20011), .A4(n20010), .ZN(
        n20024) );
  AOI22_X1 U24045 ( .A1(n3281), .A2(\xmem_data[80][6] ), .B1(n25450), .B2(
        \xmem_data[81][6] ), .ZN(n20017) );
  AOI22_X1 U24046 ( .A1(n24638), .A2(\xmem_data[82][6] ), .B1(n3358), .B2(
        \xmem_data[83][6] ), .ZN(n20016) );
  AOI22_X1 U24047 ( .A1(n24640), .A2(\xmem_data[84][6] ), .B1(n24639), .B2(
        \xmem_data[85][6] ), .ZN(n20015) );
  AOI22_X1 U24048 ( .A1(n29109), .A2(\xmem_data[86][6] ), .B1(n25458), .B2(
        \xmem_data[87][6] ), .ZN(n20014) );
  NAND4_X1 U24049 ( .A1(n20017), .A2(n20016), .A3(n20015), .A4(n20014), .ZN(
        n20023) );
  AOI22_X1 U24050 ( .A1(n20776), .A2(\xmem_data[88][6] ), .B1(n22742), .B2(
        \xmem_data[89][6] ), .ZN(n20021) );
  AOI22_X1 U24051 ( .A1(n21007), .A2(\xmem_data[90][6] ), .B1(n24645), .B2(
        \xmem_data[91][6] ), .ZN(n20020) );
  AOI22_X1 U24052 ( .A1(n20815), .A2(\xmem_data[92][6] ), .B1(n24646), .B2(
        \xmem_data[93][6] ), .ZN(n20019) );
  AOI22_X1 U24053 ( .A1(n24647), .A2(\xmem_data[94][6] ), .B1(n28060), .B2(
        \xmem_data[95][6] ), .ZN(n20018) );
  NAND4_X1 U24054 ( .A1(n20021), .A2(n20020), .A3(n20019), .A4(n20018), .ZN(
        n20022) );
  OR4_X1 U24055 ( .A1(n20025), .A2(n20024), .A3(n20023), .A4(n20022), .ZN(
        n20026) );
  NAND2_X1 U24056 ( .A1(n20026), .A2(n24720), .ZN(n20094) );
  AOI22_X1 U24057 ( .A1(n24630), .A2(\xmem_data[40][6] ), .B1(n3247), .B2(
        \xmem_data[41][6] ), .ZN(n20030) );
  AOI22_X1 U24058 ( .A1(n24631), .A2(\xmem_data[42][6] ), .B1(n3218), .B2(
        \xmem_data[43][6] ), .ZN(n20029) );
  AOI22_X1 U24059 ( .A1(n24632), .A2(\xmem_data[44][6] ), .B1(n25562), .B2(
        \xmem_data[45][6] ), .ZN(n20028) );
  AOI22_X1 U24060 ( .A1(n3340), .A2(\xmem_data[46][6] ), .B1(n24633), .B2(
        \xmem_data[47][6] ), .ZN(n20027) );
  NAND4_X1 U24061 ( .A1(n20030), .A2(n20029), .A3(n20028), .A4(n20027), .ZN(
        n20046) );
  AOI22_X1 U24062 ( .A1(n24623), .A2(\xmem_data[32][6] ), .B1(n24622), .B2(
        \xmem_data[33][6] ), .ZN(n20034) );
  AOI22_X1 U24063 ( .A1(n20782), .A2(\xmem_data[34][6] ), .B1(n29136), .B2(
        \xmem_data[35][6] ), .ZN(n20033) );
  AOI22_X1 U24064 ( .A1(n21060), .A2(\xmem_data[36][6] ), .B1(n24624), .B2(
        \xmem_data[37][6] ), .ZN(n20032) );
  AOI22_X1 U24065 ( .A1(n30588), .A2(\xmem_data[38][6] ), .B1(n3203), .B2(
        \xmem_data[39][6] ), .ZN(n20031) );
  NAND4_X1 U24066 ( .A1(n20034), .A2(n20033), .A3(n20032), .A4(n20031), .ZN(
        n20045) );
  AOI22_X1 U24067 ( .A1(n3281), .A2(\xmem_data[48][6] ), .B1(n24657), .B2(
        \xmem_data[49][6] ), .ZN(n20038) );
  AOI22_X1 U24068 ( .A1(n24638), .A2(\xmem_data[50][6] ), .B1(n27988), .B2(
        \xmem_data[51][6] ), .ZN(n20037) );
  AOI22_X1 U24069 ( .A1(n24640), .A2(\xmem_data[52][6] ), .B1(n24639), .B2(
        \xmem_data[53][6] ), .ZN(n20036) );
  AOI22_X1 U24070 ( .A1(n17041), .A2(\xmem_data[54][6] ), .B1(n25606), .B2(
        \xmem_data[55][6] ), .ZN(n20035) );
  NAND4_X1 U24071 ( .A1(n20038), .A2(n20037), .A3(n20036), .A4(n20035), .ZN(
        n20044) );
  AOI22_X1 U24072 ( .A1(n30666), .A2(\xmem_data[56][6] ), .B1(n25383), .B2(
        \xmem_data[57][6] ), .ZN(n20042) );
  AOI22_X1 U24073 ( .A1(n14937), .A2(\xmem_data[58][6] ), .B1(n24645), .B2(
        \xmem_data[59][6] ), .ZN(n20041) );
  AOI22_X1 U24074 ( .A1(n17044), .A2(\xmem_data[60][6] ), .B1(n24646), .B2(
        \xmem_data[61][6] ), .ZN(n20040) );
  AOI22_X1 U24075 ( .A1(n24647), .A2(\xmem_data[62][6] ), .B1(n28327), .B2(
        \xmem_data[63][6] ), .ZN(n20039) );
  NAND4_X1 U24076 ( .A1(n20042), .A2(n20041), .A3(n20040), .A4(n20039), .ZN(
        n20043) );
  OR4_X1 U24077 ( .A1(n20046), .A2(n20045), .A3(n20044), .A4(n20043), .ZN(
        n20047) );
  NAND2_X1 U24078 ( .A1(n20047), .A2(n24659), .ZN(n20093) );
  AOI22_X1 U24079 ( .A1(n24693), .A2(\xmem_data[104][6] ), .B1(n25360), .B2(
        \xmem_data[105][6] ), .ZN(n20052) );
  AND2_X1 U24080 ( .A1(n3219), .A2(\xmem_data[107][6] ), .ZN(n20048) );
  AOI21_X1 U24081 ( .B1(n24694), .B2(\xmem_data[106][6] ), .A(n20048), .ZN(
        n20051) );
  AOI22_X1 U24082 ( .A1(n24696), .A2(\xmem_data[108][6] ), .B1(n24695), .B2(
        \xmem_data[109][6] ), .ZN(n20050) );
  AOI22_X1 U24083 ( .A1(n24697), .A2(\xmem_data[110][6] ), .B1(n3256), .B2(
        \xmem_data[111][6] ), .ZN(n20049) );
  NAND4_X1 U24084 ( .A1(n20052), .A2(n20051), .A3(n20050), .A4(n20049), .ZN(
        n20068) );
  AOI22_X1 U24085 ( .A1(n20984), .A2(\xmem_data[96][6] ), .B1(n22685), .B2(
        \xmem_data[97][6] ), .ZN(n20056) );
  AOI22_X1 U24086 ( .A1(n24685), .A2(\xmem_data[98][6] ), .B1(n25359), .B2(
        \xmem_data[99][6] ), .ZN(n20055) );
  AOI22_X1 U24087 ( .A1(n24687), .A2(\xmem_data[100][6] ), .B1(n24686), .B2(
        \xmem_data[101][6] ), .ZN(n20054) );
  AOI22_X1 U24088 ( .A1(n24688), .A2(\xmem_data[102][6] ), .B1(n27499), .B2(
        \xmem_data[103][6] ), .ZN(n20053) );
  NAND4_X1 U24089 ( .A1(n20056), .A2(n20055), .A3(n20054), .A4(n20053), .ZN(
        n20067) );
  AOI22_X1 U24090 ( .A1(n24702), .A2(\xmem_data[112][6] ), .B1(n15011), .B2(
        \xmem_data[113][6] ), .ZN(n20060) );
  AOI22_X1 U24091 ( .A1(n23813), .A2(\xmem_data[114][6] ), .B1(n13475), .B2(
        \xmem_data[115][6] ), .ZN(n20059) );
  AOI22_X1 U24092 ( .A1(n24556), .A2(\xmem_data[116][6] ), .B1(n13168), .B2(
        \xmem_data[117][6] ), .ZN(n20058) );
  AOI22_X1 U24093 ( .A1(n30614), .A2(\xmem_data[118][6] ), .B1(n28052), .B2(
        \xmem_data[119][6] ), .ZN(n20057) );
  NAND4_X1 U24094 ( .A1(n20060), .A2(n20059), .A3(n20058), .A4(n20057), .ZN(
        n20066) );
  AOI22_X1 U24095 ( .A1(n30666), .A2(\xmem_data[120][6] ), .B1(n20586), .B2(
        \xmem_data[121][6] ), .ZN(n20064) );
  AOI22_X1 U24096 ( .A1(n24708), .A2(\xmem_data[122][6] ), .B1(n24707), .B2(
        \xmem_data[123][6] ), .ZN(n20063) );
  AOI22_X1 U24097 ( .A1(n24710), .A2(\xmem_data[124][6] ), .B1(n24709), .B2(
        \xmem_data[125][6] ), .ZN(n20062) );
  AOI22_X1 U24098 ( .A1(n30956), .A2(\xmem_data[126][6] ), .B1(n20506), .B2(
        \xmem_data[127][6] ), .ZN(n20061) );
  NAND4_X1 U24099 ( .A1(n20064), .A2(n20063), .A3(n20062), .A4(n20061), .ZN(
        n20065) );
  OR4_X1 U24100 ( .A1(n20068), .A2(n20067), .A3(n20066), .A4(n20065), .ZN(
        n20069) );
  NAND2_X1 U24101 ( .A1(n20069), .A2(n24722), .ZN(n20092) );
  AOI22_X1 U24102 ( .A1(n30311), .A2(\xmem_data[0][6] ), .B1(n24622), .B2(
        \xmem_data[1][6] ), .ZN(n20073) );
  AOI22_X1 U24103 ( .A1(n24606), .A2(\xmem_data[2][6] ), .B1(n27526), .B2(
        \xmem_data[3][6] ), .ZN(n20072) );
  AOI22_X1 U24104 ( .A1(n20708), .A2(\xmem_data[4][6] ), .B1(n30900), .B2(
        \xmem_data[5][6] ), .ZN(n20071) );
  AOI22_X1 U24105 ( .A1(n24607), .A2(\xmem_data[6][6] ), .B1(n28317), .B2(
        \xmem_data[7][6] ), .ZN(n20070) );
  NAND4_X1 U24106 ( .A1(n20073), .A2(n20072), .A3(n20071), .A4(n20070), .ZN(
        n20089) );
  AOI22_X1 U24107 ( .A1(n28677), .A2(\xmem_data[8][6] ), .B1(n3247), .B2(
        \xmem_data[9][6] ), .ZN(n20077) );
  AOI22_X1 U24108 ( .A1(n27902), .A2(\xmem_data[10][6] ), .B1(n3220), .B2(
        \xmem_data[11][6] ), .ZN(n20076) );
  AOI22_X1 U24109 ( .A1(n28137), .A2(\xmem_data[12][6] ), .B1(n25562), .B2(
        \xmem_data[13][6] ), .ZN(n20075) );
  AOI22_X1 U24110 ( .A1(n3341), .A2(\xmem_data[14][6] ), .B1(n24633), .B2(
        \xmem_data[15][6] ), .ZN(n20074) );
  NAND4_X1 U24111 ( .A1(n20077), .A2(n20076), .A3(n20075), .A4(n20074), .ZN(
        n20088) );
  AOI22_X1 U24112 ( .A1(n3128), .A2(\xmem_data[16][6] ), .B1(n28007), .B2(
        \xmem_data[17][6] ), .ZN(n20081) );
  AOI22_X1 U24113 ( .A1(n22712), .A2(\xmem_data[18][6] ), .B1(n24590), .B2(
        \xmem_data[19][6] ), .ZN(n20080) );
  AOI22_X1 U24114 ( .A1(n28671), .A2(\xmem_data[20][6] ), .B1(n13168), .B2(
        \xmem_data[21][6] ), .ZN(n20079) );
  AOI22_X1 U24115 ( .A1(n28334), .A2(\xmem_data[22][6] ), .B1(n24597), .B2(
        \xmem_data[23][6] ), .ZN(n20078) );
  NAND4_X1 U24116 ( .A1(n20081), .A2(n20080), .A3(n20079), .A4(n20078), .ZN(
        n20087) );
  AOI22_X1 U24117 ( .A1(n24458), .A2(\xmem_data[24][6] ), .B1(n3208), .B2(
        \xmem_data[25][6] ), .ZN(n20085) );
  AOI22_X1 U24118 ( .A1(n24593), .A2(\xmem_data[26][6] ), .B1(n25715), .B2(
        \xmem_data[27][6] ), .ZN(n20084) );
  AOI22_X1 U24119 ( .A1(n29012), .A2(\xmem_data[28][6] ), .B1(n24592), .B2(
        \xmem_data[29][6] ), .ZN(n20083) );
  AOI22_X1 U24120 ( .A1(n28460), .A2(\xmem_data[30][6] ), .B1(n25364), .B2(
        \xmem_data[31][6] ), .ZN(n20082) );
  NAND4_X1 U24121 ( .A1(n20085), .A2(n20084), .A3(n20083), .A4(n20082), .ZN(
        n20086) );
  OR4_X1 U24122 ( .A1(n20089), .A2(n20088), .A3(n20087), .A4(n20086), .ZN(
        n20090) );
  NAND2_X1 U24123 ( .A1(n20090), .A2(n21278), .ZN(n20091) );
  XNOR2_X1 U24124 ( .A(n33214), .B(\fmem_data[24][1] ), .ZN(n26806) );
  OAI22_X1 U24125 ( .A1(n32029), .A2(n3565), .B1(n26806), .B2(n36100), .ZN(
        n23189) );
  AOI22_X1 U24126 ( .A1(n28137), .A2(\xmem_data[16][3] ), .B1(n20787), .B2(
        \xmem_data[17][3] ), .ZN(n20095) );
  AOI22_X1 U24127 ( .A1(n20809), .A2(\xmem_data[22][3] ), .B1(n25456), .B2(
        \xmem_data[23][3] ), .ZN(n20097) );
  NAND2_X1 U24128 ( .A1(n3126), .A2(\xmem_data[20][3] ), .ZN(n20096) );
  NAND2_X1 U24129 ( .A1(n20097), .A2(n20096), .ZN(n20100) );
  AOI22_X1 U24130 ( .A1(n25490), .A2(\xmem_data[18][3] ), .B1(n29181), .B2(
        \xmem_data[19][3] ), .ZN(n20098) );
  INV_X1 U24131 ( .A(n20098), .ZN(n20099) );
  OR3_X1 U24132 ( .A1(n20101), .A2(n20100), .A3(n20099), .ZN(n20107) );
  AOI22_X1 U24133 ( .A1(n29639), .A2(\xmem_data[0][3] ), .B1(n29238), .B2(
        \xmem_data[1][3] ), .ZN(n20105) );
  AOI22_X1 U24134 ( .A1(n25575), .A2(\xmem_data[2][3] ), .B1(n31361), .B2(
        \xmem_data[3][3] ), .ZN(n20104) );
  AOI22_X1 U24135 ( .A1(n3269), .A2(\xmem_data[4][3] ), .B1(n20781), .B2(
        \xmem_data[5][3] ), .ZN(n20103) );
  AOI22_X1 U24136 ( .A1(n20782), .A2(\xmem_data[6][3] ), .B1(n27526), .B2(
        \xmem_data[7][3] ), .ZN(n20102) );
  NAND4_X1 U24137 ( .A1(n20105), .A2(n20104), .A3(n20103), .A4(n20102), .ZN(
        n20106) );
  NOR2_X1 U24138 ( .A1(n20107), .A2(n20106), .ZN(n20123) );
  AOI22_X1 U24139 ( .A1(n25724), .A2(\xmem_data[10][3] ), .B1(n28037), .B2(
        \xmem_data[11][3] ), .ZN(n20117) );
  AOI22_X1 U24140 ( .A1(n29437), .A2(\xmem_data[28][3] ), .B1(n3212), .B2(
        \xmem_data[29][3] ), .ZN(n20116) );
  AOI22_X1 U24141 ( .A1(n21308), .A2(\xmem_data[12][3] ), .B1(n25360), .B2(
        \xmem_data[13][3] ), .ZN(n20108) );
  INV_X1 U24142 ( .A(n20108), .ZN(n20114) );
  AOI22_X1 U24143 ( .A1(n29310), .A2(\xmem_data[26][3] ), .B1(n14999), .B2(
        \xmem_data[27][3] ), .ZN(n20109) );
  INV_X1 U24144 ( .A(n20109), .ZN(n20113) );
  AOI22_X1 U24145 ( .A1(n22738), .A2(\xmem_data[24][3] ), .B1(n20775), .B2(
        \xmem_data[25][3] ), .ZN(n20111) );
  AOI22_X1 U24146 ( .A1(n21007), .A2(\xmem_data[30][3] ), .B1(n20940), .B2(
        \xmem_data[31][3] ), .ZN(n20110) );
  NAND2_X1 U24147 ( .A1(n20111), .A2(n20110), .ZN(n20112) );
  NOR3_X1 U24148 ( .A1(n20114), .A2(n20113), .A3(n20112), .ZN(n20115) );
  AOI22_X1 U24149 ( .A1(n24443), .A2(\xmem_data[14][3] ), .B1(n3222), .B2(
        \xmem_data[15][3] ), .ZN(n20119) );
  AOI22_X1 U24150 ( .A1(n20770), .A2(\xmem_data[8][3] ), .B1(n20769), .B2(
        \xmem_data[9][3] ), .ZN(n20118) );
  NAND2_X1 U24151 ( .A1(n20119), .A2(n20118), .ZN(n20120) );
  NOR2_X1 U24152 ( .A1(n20121), .A2(n20120), .ZN(n20122) );
  AOI21_X1 U24153 ( .B1(n20123), .B2(n20122), .A(n20188), .ZN(n20124) );
  INV_X1 U24154 ( .A(n20124), .ZN(n20193) );
  AOI22_X1 U24155 ( .A1(n20730), .A2(\xmem_data[96][3] ), .B1(n23801), .B2(
        \xmem_data[97][3] ), .ZN(n20128) );
  AOI22_X1 U24156 ( .A1(n20731), .A2(\xmem_data[98][3] ), .B1(n29281), .B2(
        \xmem_data[99][3] ), .ZN(n20127) );
  AOI22_X1 U24157 ( .A1(n20732), .A2(\xmem_data[100][3] ), .B1(n24167), .B2(
        \xmem_data[101][3] ), .ZN(n20126) );
  AOI22_X1 U24158 ( .A1(n20734), .A2(\xmem_data[102][3] ), .B1(n20733), .B2(
        \xmem_data[103][3] ), .ZN(n20125) );
  NAND4_X1 U24159 ( .A1(n20128), .A2(n20127), .A3(n20126), .A4(n20125), .ZN(
        n20144) );
  AOI22_X1 U24160 ( .A1(n20708), .A2(\xmem_data[104][3] ), .B1(n20707), .B2(
        \xmem_data[105][3] ), .ZN(n20132) );
  AOI22_X1 U24161 ( .A1(n20710), .A2(\xmem_data[106][3] ), .B1(n20709), .B2(
        \xmem_data[107][3] ), .ZN(n20131) );
  AOI22_X1 U24162 ( .A1(n3384), .A2(\xmem_data[108][3] ), .B1(n20711), .B2(
        \xmem_data[109][3] ), .ZN(n20130) );
  AOI22_X1 U24163 ( .A1(n23756), .A2(\xmem_data[110][3] ), .B1(n3222), .B2(
        \xmem_data[111][3] ), .ZN(n20129) );
  NAND4_X1 U24164 ( .A1(n20132), .A2(n20131), .A3(n20130), .A4(n20129), .ZN(
        n20143) );
  AOI22_X1 U24165 ( .A1(n20724), .A2(\xmem_data[112][3] ), .B1(n20723), .B2(
        \xmem_data[113][3] ), .ZN(n20136) );
  AOI22_X1 U24166 ( .A1(n20725), .A2(\xmem_data[114][3] ), .B1(n29181), .B2(
        \xmem_data[115][3] ), .ZN(n20135) );
  AOI22_X1 U24167 ( .A1(n3281), .A2(\xmem_data[116][3] ), .B1(n25514), .B2(
        \xmem_data[117][3] ), .ZN(n20134) );
  AOI22_X1 U24168 ( .A1(n22712), .A2(\xmem_data[118][3] ), .B1(n20546), .B2(
        \xmem_data[119][3] ), .ZN(n20133) );
  NAND4_X1 U24169 ( .A1(n20136), .A2(n20135), .A3(n20134), .A4(n20133), .ZN(
        n20142) );
  AOI22_X1 U24170 ( .A1(n20716), .A2(\xmem_data[120][3] ), .B1(n22702), .B2(
        \xmem_data[121][3] ), .ZN(n20140) );
  AOI22_X1 U24171 ( .A1(n30614), .A2(\xmem_data[122][3] ), .B1(n20717), .B2(
        \xmem_data[123][3] ), .ZN(n20139) );
  AOI22_X1 U24172 ( .A1(n24213), .A2(\xmem_data[124][3] ), .B1(n22742), .B2(
        \xmem_data[125][3] ), .ZN(n20138) );
  AOI22_X1 U24173 ( .A1(n20542), .A2(\xmem_data[126][3] ), .B1(n25677), .B2(
        \xmem_data[127][3] ), .ZN(n20137) );
  NAND4_X1 U24174 ( .A1(n20140), .A2(n20139), .A3(n20138), .A4(n20137), .ZN(
        n20141) );
  OR4_X1 U24175 ( .A1(n20144), .A2(n20143), .A3(n20142), .A4(n20141), .ZN(
        n20167) );
  AOI22_X1 U24176 ( .A1(n20716), .A2(\xmem_data[88][3] ), .B1(n21015), .B2(
        \xmem_data[89][3] ), .ZN(n20148) );
  AOI22_X1 U24177 ( .A1(n23763), .A2(\xmem_data[90][3] ), .B1(n20717), .B2(
        \xmem_data[91][3] ), .ZN(n20147) );
  AOI22_X1 U24178 ( .A1(n29605), .A2(\xmem_data[92][3] ), .B1(n22677), .B2(
        \xmem_data[93][3] ), .ZN(n20146) );
  AOI22_X1 U24179 ( .A1(n20585), .A2(\xmem_data[94][3] ), .B1(n24219), .B2(
        \xmem_data[95][3] ), .ZN(n20145) );
  NAND4_X1 U24180 ( .A1(n20148), .A2(n20147), .A3(n20146), .A4(n20145), .ZN(
        n20159) );
  AOI22_X1 U24181 ( .A1(n20724), .A2(\xmem_data[80][3] ), .B1(n20723), .B2(
        \xmem_data[81][3] ), .ZN(n20152) );
  AOI22_X1 U24182 ( .A1(n20725), .A2(\xmem_data[82][3] ), .B1(n17061), .B2(
        \xmem_data[83][3] ), .ZN(n20151) );
  AOI22_X1 U24183 ( .A1(n3374), .A2(\xmem_data[84][3] ), .B1(n28007), .B2(
        \xmem_data[85][3] ), .ZN(n20150) );
  AOI22_X1 U24184 ( .A1(n27508), .A2(\xmem_data[86][3] ), .B1(n24130), .B2(
        \xmem_data[87][3] ), .ZN(n20149) );
  NAND4_X1 U24185 ( .A1(n20152), .A2(n20151), .A3(n20150), .A4(n20149), .ZN(
        n20158) );
  AOI22_X1 U24186 ( .A1(n20730), .A2(\xmem_data[64][3] ), .B1(n25435), .B2(
        \xmem_data[65][3] ), .ZN(n20156) );
  AOI22_X1 U24187 ( .A1(n20731), .A2(\xmem_data[66][3] ), .B1(n27856), .B2(
        \xmem_data[67][3] ), .ZN(n20155) );
  AOI22_X1 U24188 ( .A1(n20732), .A2(\xmem_data[68][3] ), .B1(n20553), .B2(
        \xmem_data[69][3] ), .ZN(n20154) );
  AOI22_X1 U24189 ( .A1(n20734), .A2(\xmem_data[70][3] ), .B1(n20733), .B2(
        \xmem_data[71][3] ), .ZN(n20153) );
  NAND4_X1 U24190 ( .A1(n20156), .A2(n20155), .A3(n20154), .A4(n20153), .ZN(
        n20157) );
  OR3_X1 U24191 ( .A1(n20157), .A2(n20158), .A3(n20159), .ZN(n20165) );
  AOI22_X1 U24192 ( .A1(n20708), .A2(\xmem_data[72][3] ), .B1(n20707), .B2(
        \xmem_data[73][3] ), .ZN(n20163) );
  AOI22_X1 U24193 ( .A1(n20710), .A2(\xmem_data[74][3] ), .B1(n20709), .B2(
        \xmem_data[75][3] ), .ZN(n20162) );
  AOI22_X1 U24194 ( .A1(n3434), .A2(\xmem_data[76][3] ), .B1(n20711), .B2(
        \xmem_data[77][3] ), .ZN(n20161) );
  AOI22_X1 U24195 ( .A1(n28364), .A2(\xmem_data[78][3] ), .B1(n3222), .B2(
        \xmem_data[79][3] ), .ZN(n20160) );
  NAND4_X1 U24196 ( .A1(n20163), .A2(n20162), .A3(n20161), .A4(n20160), .ZN(
        n20164) );
  OR2_X1 U24197 ( .A1(n20165), .A2(n20164), .ZN(n20166) );
  AOI22_X1 U24198 ( .A1(n20167), .A2(n20742), .B1(n20166), .B2(n20833), .ZN(
        n20192) );
  AOI22_X1 U24199 ( .A1(n20815), .A2(\xmem_data[32][3] ), .B1(n20814), .B2(
        \xmem_data[33][3] ), .ZN(n20171) );
  AOI22_X1 U24200 ( .A1(n3178), .A2(\xmem_data[34][3] ), .B1(n28327), .B2(
        \xmem_data[35][3] ), .ZN(n20170) );
  AOI22_X1 U24201 ( .A1(n20817), .A2(\xmem_data[36][3] ), .B1(n20781), .B2(
        \xmem_data[37][3] ), .ZN(n20169) );
  AOI22_X1 U24202 ( .A1(n20818), .A2(\xmem_data[38][3] ), .B1(n27526), .B2(
        \xmem_data[39][3] ), .ZN(n20168) );
  NAND4_X1 U24203 ( .A1(n20171), .A2(n20170), .A3(n20169), .A4(n20168), .ZN(
        n20187) );
  AOI22_X1 U24204 ( .A1(n20826), .A2(\xmem_data[40][3] ), .B1(n20707), .B2(
        \xmem_data[41][3] ), .ZN(n20175) );
  AOI22_X1 U24205 ( .A1(n20827), .A2(\xmem_data[42][3] ), .B1(n27958), .B2(
        \xmem_data[43][3] ), .ZN(n20174) );
  AOI22_X1 U24206 ( .A1(n20828), .A2(\xmem_data[44][3] ), .B1(n27437), .B2(
        \xmem_data[45][3] ), .ZN(n20173) );
  AOI22_X1 U24207 ( .A1(n30503), .A2(\xmem_data[46][3] ), .B1(n3222), .B2(
        \xmem_data[47][3] ), .ZN(n20172) );
  NAND4_X1 U24208 ( .A1(n20175), .A2(n20174), .A3(n20173), .A4(n20172), .ZN(
        n20186) );
  AOI22_X1 U24209 ( .A1(n20805), .A2(\xmem_data[48][3] ), .B1(n24695), .B2(
        \xmem_data[49][3] ), .ZN(n20179) );
  AOI22_X1 U24210 ( .A1(n20807), .A2(\xmem_data[50][3] ), .B1(n20806), .B2(
        \xmem_data[51][3] ), .ZN(n20178) );
  AOI22_X1 U24211 ( .A1(n20808), .A2(\xmem_data[52][3] ), .B1(n29103), .B2(
        \xmem_data[53][3] ), .ZN(n20177) );
  AOI22_X1 U24212 ( .A1(n20809), .A2(\xmem_data[54][3] ), .B1(n3358), .B2(
        \xmem_data[55][3] ), .ZN(n20176) );
  NAND4_X1 U24213 ( .A1(n20179), .A2(n20178), .A3(n20177), .A4(n20176), .ZN(
        n20185) );
  AOI22_X1 U24214 ( .A1(n20799), .A2(\xmem_data[56][3] ), .B1(n25423), .B2(
        \xmem_data[57][3] ), .ZN(n20183) );
  AOI22_X1 U24215 ( .A1(n28298), .A2(\xmem_data[58][3] ), .B1(n20798), .B2(
        \xmem_data[59][3] ), .ZN(n20182) );
  AOI22_X1 U24216 ( .A1(n29807), .A2(\xmem_data[60][3] ), .B1(n3213), .B2(
        \xmem_data[61][3] ), .ZN(n20181) );
  AOI22_X1 U24217 ( .A1(n20800), .A2(\xmem_data[62][3] ), .B1(n28427), .B2(
        \xmem_data[63][3] ), .ZN(n20180) );
  NAND4_X1 U24218 ( .A1(n20183), .A2(n20182), .A3(n20181), .A4(n20180), .ZN(
        n20184) );
  OR4_X1 U24219 ( .A1(n20187), .A2(n20186), .A3(n20185), .A4(n20184), .ZN(
        n20190) );
  NOR2_X1 U24220 ( .A1(n20188), .A2(n39008), .ZN(n20189) );
  AOI21_X1 U24221 ( .B1(n20190), .B2(n20765), .A(n3896), .ZN(n20191) );
  NAND3_X1 U24222 ( .A1(n20193), .A2(n20192), .A3(n20191), .ZN(n31897) );
  XNOR2_X1 U24223 ( .A(n31897), .B(\fmem_data[28][5] ), .ZN(n32755) );
  AOI22_X1 U24224 ( .A1(n28232), .A2(\xmem_data[0][2] ), .B1(n23776), .B2(
        \xmem_data[1][2] ), .ZN(n20197) );
  AOI22_X1 U24225 ( .A1(n25575), .A2(\xmem_data[2][2] ), .B1(n21051), .B2(
        \xmem_data[3][2] ), .ZN(n20196) );
  AOI22_X1 U24226 ( .A1(n20732), .A2(\xmem_data[4][2] ), .B1(n20781), .B2(
        \xmem_data[5][2] ), .ZN(n20195) );
  AOI22_X1 U24227 ( .A1(n20782), .A2(\xmem_data[6][2] ), .B1(n25406), .B2(
        \xmem_data[7][2] ), .ZN(n20194) );
  NAND4_X1 U24228 ( .A1(n20197), .A2(n20196), .A3(n20195), .A4(n20194), .ZN(
        n20203) );
  AOI22_X1 U24229 ( .A1(n20770), .A2(\xmem_data[8][2] ), .B1(n20769), .B2(
        \xmem_data[9][2] ), .ZN(n20201) );
  AOI22_X1 U24230 ( .A1(n28076), .A2(\xmem_data[10][2] ), .B1(n20489), .B2(
        \xmem_data[11][2] ), .ZN(n20200) );
  AOI22_X1 U24231 ( .A1(n28677), .A2(\xmem_data[12][2] ), .B1(n20568), .B2(
        \xmem_data[13][2] ), .ZN(n20199) );
  AOI22_X1 U24232 ( .A1(n30906), .A2(\xmem_data[14][2] ), .B1(n3219), .B2(
        \xmem_data[15][2] ), .ZN(n20198) );
  NAND4_X1 U24233 ( .A1(n20201), .A2(n20200), .A3(n20199), .A4(n20198), .ZN(
        n20202) );
  AOI22_X1 U24234 ( .A1(n27763), .A2(\xmem_data[24][2] ), .B1(n20775), .B2(
        \xmem_data[25][2] ), .ZN(n20207) );
  AOI22_X1 U24235 ( .A1(n30891), .A2(\xmem_data[26][2] ), .B1(n22674), .B2(
        \xmem_data[27][2] ), .ZN(n20206) );
  AOI22_X1 U24236 ( .A1(n29437), .A2(\xmem_data[28][2] ), .B1(n27516), .B2(
        \xmem_data[29][2] ), .ZN(n20205) );
  AOI22_X1 U24237 ( .A1(n21007), .A2(\xmem_data[30][2] ), .B1(n24459), .B2(
        \xmem_data[31][2] ), .ZN(n20204) );
  AND4_X1 U24238 ( .A1(n20207), .A2(n20206), .A3(n20205), .A4(n20204), .ZN(
        n20216) );
  AOI22_X1 U24239 ( .A1(n29627), .A2(\xmem_data[16][2] ), .B1(n20787), .B2(
        \xmem_data[17][2] ), .ZN(n20208) );
  INV_X1 U24240 ( .A(n20208), .ZN(n20213) );
  AOI22_X1 U24241 ( .A1(n29027), .A2(\xmem_data[18][2] ), .B1(n22669), .B2(
        \xmem_data[19][2] ), .ZN(n20211) );
  AOI22_X1 U24242 ( .A1(n25707), .A2(\xmem_data[22][2] ), .B1(n3357), .B2(
        \xmem_data[23][2] ), .ZN(n20210) );
  NAND2_X1 U24243 ( .A1(n3345), .A2(\xmem_data[20][2] ), .ZN(n20209) );
  NAND3_X1 U24244 ( .A1(n20211), .A2(n20210), .A3(n20209), .ZN(n20212) );
  NOR2_X1 U24245 ( .A1(n20213), .A2(n20212), .ZN(n20215) );
  NAND2_X1 U24246 ( .A1(n29306), .A2(\xmem_data[21][2] ), .ZN(n20214) );
  OAI21_X1 U24247 ( .B1(n3964), .B2(n20217), .A(n20795), .ZN(n20285) );
  AOI22_X1 U24248 ( .A1(n20708), .A2(\xmem_data[72][2] ), .B1(n20707), .B2(
        \xmem_data[73][2] ), .ZN(n20222) );
  AOI22_X1 U24249 ( .A1(n20710), .A2(\xmem_data[74][2] ), .B1(n20709), .B2(
        \xmem_data[75][2] ), .ZN(n20221) );
  AOI22_X1 U24250 ( .A1(n3333), .A2(\xmem_data[76][2] ), .B1(n20711), .B2(
        \xmem_data[77][2] ), .ZN(n20220) );
  AND2_X1 U24251 ( .A1(n3222), .A2(\xmem_data[79][2] ), .ZN(n20218) );
  AOI21_X1 U24252 ( .B1(n25730), .B2(\xmem_data[78][2] ), .A(n20218), .ZN(
        n20219) );
  NAND4_X1 U24253 ( .A1(n20222), .A2(n20221), .A3(n20220), .A4(n20219), .ZN(
        n20239) );
  AOI22_X1 U24254 ( .A1(n20716), .A2(\xmem_data[88][2] ), .B1(n30552), .B2(
        \xmem_data[89][2] ), .ZN(n20226) );
  AOI22_X1 U24255 ( .A1(n28980), .A2(\xmem_data[90][2] ), .B1(n20717), .B2(
        \xmem_data[91][2] ), .ZN(n20225) );
  AOI22_X1 U24256 ( .A1(n31354), .A2(\xmem_data[92][2] ), .B1(n20543), .B2(
        \xmem_data[93][2] ), .ZN(n20224) );
  AOI22_X1 U24257 ( .A1(n20585), .A2(\xmem_data[94][2] ), .B1(n24707), .B2(
        \xmem_data[95][2] ), .ZN(n20223) );
  NAND4_X1 U24258 ( .A1(n20226), .A2(n20225), .A3(n20224), .A4(n20223), .ZN(
        n20237) );
  AOI22_X1 U24259 ( .A1(n20724), .A2(\xmem_data[80][2] ), .B1(n20723), .B2(
        \xmem_data[81][2] ), .ZN(n20230) );
  AOI22_X1 U24260 ( .A1(n20725), .A2(\xmem_data[82][2] ), .B1(n24633), .B2(
        \xmem_data[83][2] ), .ZN(n20229) );
  AOI22_X1 U24261 ( .A1(n16973), .A2(\xmem_data[84][2] ), .B1(n3231), .B2(
        \xmem_data[85][2] ), .ZN(n20228) );
  AOI22_X1 U24262 ( .A1(n23813), .A2(\xmem_data[86][2] ), .B1(n3358), .B2(
        \xmem_data[87][2] ), .ZN(n20227) );
  NAND4_X1 U24263 ( .A1(n20230), .A2(n20229), .A3(n20228), .A4(n20227), .ZN(
        n20236) );
  AOI22_X1 U24264 ( .A1(n20730), .A2(\xmem_data[64][2] ), .B1(n24510), .B2(
        \xmem_data[65][2] ), .ZN(n20234) );
  AOI22_X1 U24265 ( .A1(n20731), .A2(\xmem_data[66][2] ), .B1(n25679), .B2(
        \xmem_data[67][2] ), .ZN(n20233) );
  AOI22_X1 U24266 ( .A1(n20732), .A2(\xmem_data[68][2] ), .B1(n24223), .B2(
        \xmem_data[69][2] ), .ZN(n20232) );
  AOI22_X1 U24267 ( .A1(n20734), .A2(\xmem_data[70][2] ), .B1(n20733), .B2(
        \xmem_data[71][2] ), .ZN(n20231) );
  NAND4_X1 U24268 ( .A1(n20234), .A2(n20233), .A3(n20232), .A4(n20231), .ZN(
        n20235) );
  OR3_X1 U24269 ( .A1(n20237), .A2(n20236), .A3(n20235), .ZN(n20238) );
  OAI21_X1 U24270 ( .B1(n20239), .B2(n20238), .A(n20833), .ZN(n20284) );
  AOI22_X1 U24271 ( .A1(n20826), .A2(\xmem_data[40][2] ), .B1(n24686), .B2(
        \xmem_data[41][2] ), .ZN(n20243) );
  AOI22_X1 U24272 ( .A1(n20827), .A2(\xmem_data[42][2] ), .B1(n20709), .B2(
        \xmem_data[43][2] ), .ZN(n20242) );
  AOI22_X1 U24273 ( .A1(n20828), .A2(\xmem_data[44][2] ), .B1(n27437), .B2(
        \xmem_data[45][2] ), .ZN(n20241) );
  AOI22_X1 U24274 ( .A1(n30592), .A2(\xmem_data[46][2] ), .B1(n3219), .B2(
        \xmem_data[47][2] ), .ZN(n20240) );
  NAND4_X1 U24275 ( .A1(n20243), .A2(n20242), .A3(n20241), .A4(n20240), .ZN(
        n20260) );
  AOI22_X1 U24276 ( .A1(n20799), .A2(\xmem_data[56][2] ), .B1(n24132), .B2(
        \xmem_data[57][2] ), .ZN(n20247) );
  AOI22_X1 U24277 ( .A1(n30514), .A2(\xmem_data[58][2] ), .B1(n20798), .B2(
        \xmem_data[59][2] ), .ZN(n20246) );
  AOI22_X1 U24278 ( .A1(n31354), .A2(\xmem_data[60][2] ), .B1(n27864), .B2(
        \xmem_data[61][2] ), .ZN(n20245) );
  AOI22_X1 U24279 ( .A1(n20800), .A2(\xmem_data[62][2] ), .B1(n25715), .B2(
        \xmem_data[63][2] ), .ZN(n20244) );
  NAND4_X1 U24280 ( .A1(n20247), .A2(n20246), .A3(n20245), .A4(n20244), .ZN(
        n20258) );
  AOI22_X1 U24281 ( .A1(n20805), .A2(\xmem_data[48][2] ), .B1(n20598), .B2(
        \xmem_data[49][2] ), .ZN(n20251) );
  AOI22_X1 U24282 ( .A1(n20807), .A2(\xmem_data[50][2] ), .B1(n20806), .B2(
        \xmem_data[51][2] ), .ZN(n20250) );
  AOI22_X1 U24283 ( .A1(n20808), .A2(\xmem_data[52][2] ), .B1(n25450), .B2(
        \xmem_data[53][2] ), .ZN(n20249) );
  AOI22_X1 U24284 ( .A1(n20809), .A2(\xmem_data[54][2] ), .B1(n29180), .B2(
        \xmem_data[55][2] ), .ZN(n20248) );
  NAND4_X1 U24285 ( .A1(n20251), .A2(n20250), .A3(n20249), .A4(n20248), .ZN(
        n20257) );
  AOI22_X1 U24286 ( .A1(n20815), .A2(\xmem_data[32][2] ), .B1(n20814), .B2(
        \xmem_data[33][2] ), .ZN(n20255) );
  AOI22_X1 U24287 ( .A1(n21010), .A2(\xmem_data[34][2] ), .B1(n20506), .B2(
        \xmem_data[35][2] ), .ZN(n20254) );
  AOI22_X1 U24288 ( .A1(n20817), .A2(\xmem_data[36][2] ), .B1(n24570), .B2(
        \xmem_data[37][2] ), .ZN(n20253) );
  AOI22_X1 U24289 ( .A1(n20818), .A2(\xmem_data[38][2] ), .B1(n29247), .B2(
        \xmem_data[39][2] ), .ZN(n20252) );
  NAND4_X1 U24290 ( .A1(n20255), .A2(n20254), .A3(n20253), .A4(n20252), .ZN(
        n20256) );
  OR3_X1 U24291 ( .A1(n20258), .A2(n20257), .A3(n20256), .ZN(n20259) );
  OAI21_X1 U24292 ( .B1(n20260), .B2(n20259), .A(n20765), .ZN(n20283) );
  AOI22_X1 U24293 ( .A1(n20708), .A2(\xmem_data[104][2] ), .B1(n20707), .B2(
        \xmem_data[105][2] ), .ZN(n20264) );
  AOI22_X1 U24294 ( .A1(n20710), .A2(\xmem_data[106][2] ), .B1(n20709), .B2(
        \xmem_data[107][2] ), .ZN(n20263) );
  AOI22_X1 U24295 ( .A1(n3348), .A2(\xmem_data[108][2] ), .B1(n20711), .B2(
        \xmem_data[109][2] ), .ZN(n20262) );
  AOI22_X1 U24296 ( .A1(n30962), .A2(\xmem_data[110][2] ), .B1(n3221), .B2(
        \xmem_data[111][2] ), .ZN(n20261) );
  NAND4_X1 U24297 ( .A1(n20264), .A2(n20263), .A3(n20262), .A4(n20261), .ZN(
        n20281) );
  AOI22_X1 U24298 ( .A1(n20716), .A2(\xmem_data[120][2] ), .B1(n27535), .B2(
        \xmem_data[121][2] ), .ZN(n20268) );
  AOI22_X1 U24299 ( .A1(n28334), .A2(\xmem_data[122][2] ), .B1(n20717), .B2(
        \xmem_data[123][2] ), .ZN(n20267) );
  AOI22_X1 U24300 ( .A1(n3158), .A2(\xmem_data[124][2] ), .B1(n24134), .B2(
        \xmem_data[125][2] ), .ZN(n20266) );
  AOI22_X1 U24301 ( .A1(n13149), .A2(\xmem_data[126][2] ), .B1(n25398), .B2(
        \xmem_data[127][2] ), .ZN(n20265) );
  NAND4_X1 U24302 ( .A1(n20268), .A2(n20267), .A3(n20266), .A4(n20265), .ZN(
        n20279) );
  AOI22_X1 U24303 ( .A1(n20724), .A2(\xmem_data[112][2] ), .B1(n20723), .B2(
        \xmem_data[113][2] ), .ZN(n20272) );
  AOI22_X1 U24304 ( .A1(n20725), .A2(\xmem_data[114][2] ), .B1(n20806), .B2(
        \xmem_data[115][2] ), .ZN(n20271) );
  AOI22_X1 U24305 ( .A1(n21074), .A2(\xmem_data[116][2] ), .B1(n28307), .B2(
        \xmem_data[117][2] ), .ZN(n20270) );
  AOI22_X1 U24306 ( .A1(n31321), .A2(\xmem_data[118][2] ), .B1(n28415), .B2(
        \xmem_data[119][2] ), .ZN(n20269) );
  NAND4_X1 U24307 ( .A1(n20272), .A2(n20271), .A3(n20270), .A4(n20269), .ZN(
        n20278) );
  AOI22_X1 U24308 ( .A1(n20730), .A2(\xmem_data[96][2] ), .B1(n25435), .B2(
        \xmem_data[97][2] ), .ZN(n20276) );
  AOI22_X1 U24309 ( .A1(n20731), .A2(\xmem_data[98][2] ), .B1(n25581), .B2(
        \xmem_data[99][2] ), .ZN(n20275) );
  AOI22_X1 U24310 ( .A1(n20732), .A2(\xmem_data[100][2] ), .B1(n24167), .B2(
        \xmem_data[101][2] ), .ZN(n20274) );
  AOI22_X1 U24311 ( .A1(n20734), .A2(\xmem_data[102][2] ), .B1(n20733), .B2(
        \xmem_data[103][2] ), .ZN(n20273) );
  NAND4_X1 U24312 ( .A1(n20276), .A2(n20275), .A3(n20274), .A4(n20273), .ZN(
        n20277) );
  OR3_X1 U24313 ( .A1(n20279), .A2(n20278), .A3(n20277), .ZN(n20280) );
  OAI21_X1 U24314 ( .B1(n20281), .B2(n20280), .A(n20742), .ZN(n20282) );
  XNOR2_X1 U24315 ( .A(n33573), .B(\fmem_data[28][5] ), .ZN(n30980) );
  OAI22_X1 U24316 ( .A1(n32755), .A2(n33828), .B1(n30980), .B2(n33827), .ZN(
        n23188) );
  XNOR2_X1 U24317 ( .A(n31899), .B(\fmem_data[20][5] ), .ZN(n31987) );
  XNOR2_X1 U24318 ( .A(n32127), .B(\fmem_data[20][5] ), .ZN(n32522) );
  NOR2_X1 U24319 ( .A1(n23173), .A2(n23174), .ZN(n20287) );
  NAND2_X1 U24320 ( .A1(n23174), .A2(n23173), .ZN(n20286) );
  OAI21_X1 U24321 ( .B1(n20288), .B2(n20287), .A(n20286), .ZN(n23184) );
  FA_X1 U24322 ( .A(n20291), .B(n20290), .CI(n20289), .CO(n12718), .S(n23183)
         );
  XNOR2_X1 U24323 ( .A(n32064), .B(\fmem_data[0][5] ), .ZN(n33184) );
  AOI22_X1 U24324 ( .A1(n20939), .A2(\xmem_data[32][2] ), .B1(n20938), .B2(
        \xmem_data[33][2] ), .ZN(n20295) );
  AOI22_X1 U24325 ( .A1(n24214), .A2(\xmem_data[34][2] ), .B1(n20940), .B2(
        \xmem_data[35][2] ), .ZN(n20294) );
  AOI22_X1 U24326 ( .A1(n20942), .A2(\xmem_data[36][2] ), .B1(n20941), .B2(
        \xmem_data[37][2] ), .ZN(n20293) );
  AOI22_X1 U24327 ( .A1(n24190), .A2(\xmem_data[38][2] ), .B1(n20943), .B2(
        \xmem_data[39][2] ), .ZN(n20292) );
  NAND4_X1 U24328 ( .A1(n20295), .A2(n20294), .A3(n20293), .A4(n20292), .ZN(
        n20301) );
  AOI22_X1 U24329 ( .A1(n20962), .A2(\xmem_data[56][2] ), .B1(n27446), .B2(
        \xmem_data[57][2] ), .ZN(n20299) );
  AOI22_X1 U24330 ( .A1(n20961), .A2(\xmem_data[58][2] ), .B1(n24158), .B2(
        \xmem_data[59][2] ), .ZN(n20298) );
  AOI22_X1 U24331 ( .A1(n24157), .A2(\xmem_data[60][2] ), .B1(n20958), .B2(
        \xmem_data[61][2] ), .ZN(n20297) );
  AOI22_X1 U24332 ( .A1(n20959), .A2(\xmem_data[62][2] ), .B1(n24160), .B2(
        \xmem_data[63][2] ), .ZN(n20296) );
  NAND4_X1 U24333 ( .A1(n20299), .A2(n20298), .A3(n20297), .A4(n20296), .ZN(
        n20300) );
  NOR2_X1 U24334 ( .A1(n20301), .A2(n20300), .ZN(n20304) );
  AOI22_X1 U24335 ( .A1(n20953), .A2(\xmem_data[46][2] ), .B1(n30861), .B2(
        \xmem_data[47][2] ), .ZN(n20303) );
  AOI22_X1 U24336 ( .A1(n27439), .A2(\xmem_data[50][2] ), .B1(n3217), .B2(
        \xmem_data[51][2] ), .ZN(n20302) );
  NAND3_X1 U24337 ( .A1(n20304), .A2(n20303), .A3(n20302), .ZN(n20313) );
  AOI22_X1 U24338 ( .A1(n20969), .A2(\xmem_data[54][2] ), .B1(n28372), .B2(
        \xmem_data[55][2] ), .ZN(n20306) );
  AOI22_X1 U24339 ( .A1(n29026), .A2(\xmem_data[52][2] ), .B1(n23739), .B2(
        \xmem_data[53][2] ), .ZN(n20305) );
  AOI22_X1 U24340 ( .A1(n20952), .A2(\xmem_data[44][2] ), .B1(n20951), .B2(
        \xmem_data[45][2] ), .ZN(n20310) );
  AOI22_X1 U24341 ( .A1(n24467), .A2(\xmem_data[42][2] ), .B1(n25359), .B2(
        \xmem_data[43][2] ), .ZN(n20309) );
  AOI22_X1 U24342 ( .A1(n22728), .A2(\xmem_data[48][2] ), .B1(n29286), .B2(
        \xmem_data[49][2] ), .ZN(n20308) );
  AOI22_X1 U24343 ( .A1(n20950), .A2(\xmem_data[40][2] ), .B1(n20949), .B2(
        \xmem_data[41][2] ), .ZN(n20307) );
  NAND3_X1 U24344 ( .A1(n4010), .A2(n20310), .A3(n3557), .ZN(n20312) );
  AOI22_X1 U24345 ( .A1(n21048), .A2(\xmem_data[64][2] ), .B1(n20586), .B2(
        \xmem_data[65][2] ), .ZN(n20317) );
  AOI22_X1 U24346 ( .A1(n25573), .A2(\xmem_data[66][2] ), .B1(n29048), .B2(
        \xmem_data[67][2] ), .ZN(n20316) );
  AOI22_X1 U24347 ( .A1(n21050), .A2(\xmem_data[68][2] ), .B1(n21049), .B2(
        \xmem_data[69][2] ), .ZN(n20315) );
  AOI22_X1 U24348 ( .A1(n3326), .A2(\xmem_data[70][2] ), .B1(n25581), .B2(
        \xmem_data[71][2] ), .ZN(n20314) );
  NAND4_X1 U24349 ( .A1(n20317), .A2(n20316), .A3(n20315), .A4(n20314), .ZN(
        n20323) );
  AOI22_X1 U24350 ( .A1(n21074), .A2(\xmem_data[88][2] ), .B1(n25450), .B2(
        \xmem_data[89][2] ), .ZN(n20321) );
  AOI22_X1 U24351 ( .A1(n25422), .A2(\xmem_data[90][2] ), .B1(n24590), .B2(
        \xmem_data[91][2] ), .ZN(n20320) );
  AOI22_X1 U24352 ( .A1(n29451), .A2(\xmem_data[92][2] ), .B1(n21075), .B2(
        \xmem_data[93][2] ), .ZN(n20319) );
  AOI22_X1 U24353 ( .A1(n28298), .A2(\xmem_data[94][2] ), .B1(n21076), .B2(
        \xmem_data[95][2] ), .ZN(n20318) );
  NAND4_X1 U24354 ( .A1(n20321), .A2(n20320), .A3(n20319), .A4(n20318), .ZN(
        n20322) );
  NOR2_X1 U24355 ( .A1(n20323), .A2(n20322), .ZN(n20336) );
  AOI22_X1 U24356 ( .A1(n21061), .A2(\xmem_data[78][2] ), .B1(n30571), .B2(
        \xmem_data[79][2] ), .ZN(n20335) );
  AOI22_X1 U24357 ( .A1(n21069), .A2(\xmem_data[86][2] ), .B1(n21068), .B2(
        \xmem_data[87][2] ), .ZN(n20325) );
  AOI22_X1 U24358 ( .A1(n21067), .A2(\xmem_data[84][2] ), .B1(n30963), .B2(
        \xmem_data[85][2] ), .ZN(n20324) );
  NAND2_X1 U24359 ( .A1(n20325), .A2(n20324), .ZN(n20332) );
  AOI22_X1 U24360 ( .A1(n21058), .A2(\xmem_data[74][2] ), .B1(n21057), .B2(
        \xmem_data[75][2] ), .ZN(n20328) );
  AOI22_X1 U24361 ( .A1(n3144), .A2(\xmem_data[80][2] ), .B1(n28501), .B2(
        \xmem_data[81][2] ), .ZN(n20327) );
  AOI22_X1 U24362 ( .A1(n21056), .A2(\xmem_data[72][2] ), .B1(n28098), .B2(
        \xmem_data[73][2] ), .ZN(n20326) );
  AOI22_X1 U24363 ( .A1(n21060), .A2(\xmem_data[76][2] ), .B1(n21059), .B2(
        \xmem_data[77][2] ), .ZN(n20329) );
  INV_X1 U24364 ( .A(n20329), .ZN(n20330) );
  NOR3_X1 U24365 ( .A1(n20332), .A2(n20331), .A3(n20330), .ZN(n20334) );
  AOI22_X1 U24366 ( .A1(n21066), .A2(\xmem_data[82][2] ), .B1(n3221), .B2(
        \xmem_data[83][2] ), .ZN(n20333) );
  NAND4_X1 U24367 ( .A1(n20336), .A2(n20335), .A3(n20334), .A4(n20333), .ZN(
        n20337) );
  NAND2_X1 U24368 ( .A1(n20337), .A2(n21086), .ZN(n20390) );
  AOI22_X1 U24369 ( .A1(n21048), .A2(\xmem_data[96][2] ), .B1(n25574), .B2(
        \xmem_data[97][2] ), .ZN(n20341) );
  AOI22_X1 U24370 ( .A1(n24509), .A2(\xmem_data[98][2] ), .B1(n23796), .B2(
        \xmem_data[99][2] ), .ZN(n20340) );
  AOI22_X1 U24371 ( .A1(n21050), .A2(\xmem_data[100][2] ), .B1(n21049), .B2(
        \xmem_data[101][2] ), .ZN(n20339) );
  AOI22_X1 U24372 ( .A1(n28428), .A2(\xmem_data[102][2] ), .B1(n27856), .B2(
        \xmem_data[103][2] ), .ZN(n20338) );
  NAND4_X1 U24373 ( .A1(n20341), .A2(n20340), .A3(n20339), .A4(n20338), .ZN(
        n20347) );
  AOI22_X1 U24374 ( .A1(n21074), .A2(\xmem_data[120][2] ), .B1(n3231), .B2(
        \xmem_data[121][2] ), .ZN(n20345) );
  AOI22_X1 U24375 ( .A1(n16974), .A2(\xmem_data[122][2] ), .B1(n25456), .B2(
        \xmem_data[123][2] ), .ZN(n20344) );
  AOI22_X1 U24376 ( .A1(n30608), .A2(\xmem_data[124][2] ), .B1(n21075), .B2(
        \xmem_data[125][2] ), .ZN(n20343) );
  AOI22_X1 U24377 ( .A1(n20959), .A2(\xmem_data[126][2] ), .B1(n21076), .B2(
        \xmem_data[127][2] ), .ZN(n20342) );
  NAND4_X1 U24378 ( .A1(n20345), .A2(n20344), .A3(n20343), .A4(n20342), .ZN(
        n20346) );
  NOR2_X1 U24379 ( .A1(n20347), .A2(n20346), .ZN(n20360) );
  AOI22_X1 U24380 ( .A1(n21061), .A2(\xmem_data[110][2] ), .B1(n21309), .B2(
        \xmem_data[111][2] ), .ZN(n20359) );
  AOI22_X1 U24381 ( .A1(n21069), .A2(\xmem_data[118][2] ), .B1(n21068), .B2(
        \xmem_data[119][2] ), .ZN(n20349) );
  AOI22_X1 U24382 ( .A1(n21067), .A2(\xmem_data[116][2] ), .B1(n29255), .B2(
        \xmem_data[117][2] ), .ZN(n20348) );
  NAND2_X1 U24383 ( .A1(n20349), .A2(n20348), .ZN(n20356) );
  AOI22_X1 U24384 ( .A1(n21058), .A2(\xmem_data[106][2] ), .B1(n21057), .B2(
        \xmem_data[107][2] ), .ZN(n20352) );
  AOI22_X1 U24385 ( .A1(n3424), .A2(\xmem_data[112][2] ), .B1(n24439), .B2(
        \xmem_data[113][2] ), .ZN(n20351) );
  AOI22_X1 U24386 ( .A1(n21056), .A2(\xmem_data[104][2] ), .B1(n28098), .B2(
        \xmem_data[105][2] ), .ZN(n20350) );
  AOI22_X1 U24387 ( .A1(n21060), .A2(\xmem_data[108][2] ), .B1(n21059), .B2(
        \xmem_data[109][2] ), .ZN(n20353) );
  INV_X1 U24388 ( .A(n20353), .ZN(n20354) );
  NOR3_X1 U24389 ( .A1(n20356), .A2(n20355), .A3(n20354), .ZN(n20358) );
  AOI22_X1 U24390 ( .A1(n21066), .A2(\xmem_data[114][2] ), .B1(n3221), .B2(
        \xmem_data[115][2] ), .ZN(n20357) );
  NAND4_X1 U24391 ( .A1(n20360), .A2(n20359), .A3(n20358), .A4(n20357), .ZN(
        n20361) );
  NAND2_X1 U24392 ( .A1(n20361), .A2(n21088), .ZN(n20389) );
  AOI22_X1 U24393 ( .A1(n21005), .A2(\xmem_data[0][2] ), .B1(n22742), .B2(
        \xmem_data[1][2] ), .ZN(n20365) );
  AOI22_X1 U24394 ( .A1(n21007), .A2(\xmem_data[2][2] ), .B1(n21006), .B2(
        \xmem_data[3][2] ), .ZN(n20364) );
  AOI22_X1 U24395 ( .A1(n21008), .A2(\xmem_data[4][2] ), .B1(n29318), .B2(
        \xmem_data[5][2] ), .ZN(n20363) );
  AOI22_X1 U24396 ( .A1(n21010), .A2(\xmem_data[6][2] ), .B1(n25581), .B2(
        \xmem_data[7][2] ), .ZN(n20362) );
  NAND4_X1 U24397 ( .A1(n20365), .A2(n20364), .A3(n20363), .A4(n20362), .ZN(
        n20366) );
  AOI22_X1 U24398 ( .A1(n29591), .A2(\xmem_data[28][2] ), .B1(n21015), .B2(
        \xmem_data[29][2] ), .ZN(n20373) );
  AOI22_X1 U24399 ( .A1(n25459), .A2(\xmem_data[30][2] ), .B1(n25572), .B2(
        \xmem_data[31][2] ), .ZN(n20367) );
  INV_X1 U24400 ( .A(n20367), .ZN(n20371) );
  AOI22_X1 U24401 ( .A1(n25422), .A2(\xmem_data[26][2] ), .B1(n20982), .B2(
        \xmem_data[27][2] ), .ZN(n20369) );
  NAND2_X1 U24402 ( .A1(n25417), .A2(\xmem_data[24][2] ), .ZN(n20368) );
  NAND2_X1 U24403 ( .A1(n20369), .A2(n20368), .ZN(n20370) );
  NOR2_X1 U24404 ( .A1(n20371), .A2(n20370), .ZN(n20372) );
  NAND2_X1 U24405 ( .A1(n20373), .A2(n20372), .ZN(n20384) );
  AOI22_X1 U24406 ( .A1(n20984), .A2(\xmem_data[8][2] ), .B1(n20983), .B2(
        \xmem_data[9][2] ), .ZN(n20377) );
  AOI22_X1 U24407 ( .A1(n24166), .A2(\xmem_data[10][2] ), .B1(n29247), .B2(
        \xmem_data[11][2] ), .ZN(n20376) );
  AOI22_X1 U24408 ( .A1(n20985), .A2(\xmem_data[12][2] ), .B1(n31344), .B2(
        \xmem_data[13][2] ), .ZN(n20375) );
  AOI22_X1 U24409 ( .A1(n20986), .A2(\xmem_data[14][2] ), .B1(n29118), .B2(
        \xmem_data[15][2] ), .ZN(n20374) );
  NAND4_X1 U24410 ( .A1(n20377), .A2(n20376), .A3(n20375), .A4(n20374), .ZN(
        n20383) );
  AOI22_X1 U24411 ( .A1(n3332), .A2(\xmem_data[16][2] ), .B1(n27501), .B2(
        \xmem_data[17][2] ), .ZN(n20381) );
  AOI22_X1 U24412 ( .A1(n20991), .A2(\xmem_data[18][2] ), .B1(n3217), .B2(
        \xmem_data[19][2] ), .ZN(n20380) );
  AOI22_X1 U24413 ( .A1(n29065), .A2(\xmem_data[20][2] ), .B1(n20992), .B2(
        \xmem_data[21][2] ), .ZN(n20379) );
  AOI22_X1 U24414 ( .A1(n20994), .A2(\xmem_data[22][2] ), .B1(n20993), .B2(
        \xmem_data[23][2] ), .ZN(n20378) );
  NAND4_X1 U24415 ( .A1(n20381), .A2(n20380), .A3(n20379), .A4(n20378), .ZN(
        n20382) );
  NAND2_X1 U24416 ( .A1(n20387), .A2(n20980), .ZN(n20388) );
  AOI22_X1 U24417 ( .A1(n20488), .A2(\xmem_data[0][1] ), .B1(n25407), .B2(
        \xmem_data[1][1] ), .ZN(n20396) );
  AOI22_X1 U24418 ( .A1(n24686), .A2(\xmem_data[2][1] ), .B1(n28354), .B2(
        \xmem_data[3][1] ), .ZN(n20395) );
  AOI22_X1 U24419 ( .A1(n20489), .A2(\xmem_data[4][1] ), .B1(n3335), .B2(
        \xmem_data[5][1] ), .ZN(n20394) );
  AND2_X1 U24420 ( .A1(n20568), .A2(\xmem_data[6][1] ), .ZN(n20392) );
  AOI21_X1 U24421 ( .B1(n20518), .B2(\xmem_data[7][1] ), .A(n20392), .ZN(
        n20393) );
  NAND4_X1 U24422 ( .A1(n20396), .A2(n20395), .A3(n20394), .A4(n20393), .ZN(
        n20416) );
  AOI22_X1 U24423 ( .A1(n3221), .A2(\xmem_data[8][1] ), .B1(n27708), .B2(
        \xmem_data[9][1] ), .ZN(n20403) );
  AOI22_X1 U24424 ( .A1(n25616), .A2(\xmem_data[12][1] ), .B1(n25732), .B2(
        \xmem_data[13][1] ), .ZN(n20397) );
  INV_X1 U24425 ( .A(n20397), .ZN(n20401) );
  AOI22_X1 U24426 ( .A1(n20500), .A2(\xmem_data[10][1] ), .B1(n24141), .B2(
        \xmem_data[11][1] ), .ZN(n20399) );
  NAND2_X1 U24427 ( .A1(n23813), .A2(\xmem_data[15][1] ), .ZN(n20398) );
  NAND2_X1 U24428 ( .A1(n20399), .A2(n20398), .ZN(n20400) );
  NOR2_X1 U24429 ( .A1(n20401), .A2(n20400), .ZN(n20402) );
  NAND2_X1 U24430 ( .A1(n20403), .A2(n20402), .ZN(n20414) );
  AOI22_X1 U24431 ( .A1(n20505), .A2(\xmem_data[24][1] ), .B1(n27825), .B2(
        \xmem_data[25][1] ), .ZN(n20407) );
  AOI22_X1 U24432 ( .A1(n13481), .A2(\xmem_data[26][1] ), .B1(n21010), .B2(
        \xmem_data[27][1] ), .ZN(n20406) );
  AOI22_X1 U24433 ( .A1(n21009), .A2(\xmem_data[28][1] ), .B1(n3308), .B2(
        \xmem_data[29][1] ), .ZN(n20405) );
  AOI22_X1 U24434 ( .A1(n20507), .A2(\xmem_data[30][1] ), .B1(n24606), .B2(
        \xmem_data[31][1] ), .ZN(n20404) );
  NAND4_X1 U24435 ( .A1(n20407), .A2(n20406), .A3(n20405), .A4(n20404), .ZN(
        n20413) );
  AOI22_X1 U24436 ( .A1(n30884), .A2(\xmem_data[16][1] ), .B1(n20587), .B2(
        \xmem_data[17][1] ), .ZN(n20411) );
  AOI22_X1 U24437 ( .A1(n24448), .A2(\xmem_data[18][1] ), .B1(n28980), .B2(
        \xmem_data[19][1] ), .ZN(n20410) );
  AOI22_X1 U24438 ( .A1(n25458), .A2(\xmem_data[20][1] ), .B1(n27455), .B2(
        \xmem_data[21][1] ), .ZN(n20409) );
  AOI22_X1 U24439 ( .A1(n20938), .A2(\xmem_data[22][1] ), .B1(n24509), .B2(
        \xmem_data[23][1] ), .ZN(n20408) );
  NAND4_X1 U24440 ( .A1(n20411), .A2(n20410), .A3(n20409), .A4(n20408), .ZN(
        n20412) );
  OR3_X1 U24441 ( .A1(n20414), .A2(n20413), .A3(n20412), .ZN(n20415) );
  NOR2_X1 U24442 ( .A1(n20416), .A2(n20415), .ZN(n20417) );
  AOI22_X1 U24443 ( .A1(n30496), .A2(\xmem_data[32][1] ), .B1(n20577), .B2(
        \xmem_data[33][1] ), .ZN(n20421) );
  AOI22_X1 U24444 ( .A1(n20579), .A2(\xmem_data[34][1] ), .B1(n27959), .B2(
        \xmem_data[35][1] ), .ZN(n20420) );
  AOI22_X1 U24445 ( .A1(n20578), .A2(\xmem_data[36][1] ), .B1(n28677), .B2(
        \xmem_data[37][1] ), .ZN(n20419) );
  AOI22_X1 U24446 ( .A1(n31347), .A2(\xmem_data[38][1] ), .B1(n20576), .B2(
        \xmem_data[39][1] ), .ZN(n20418) );
  NAND4_X1 U24447 ( .A1(n20421), .A2(n20420), .A3(n20419), .A4(n20418), .ZN(
        n20437) );
  AOI22_X1 U24448 ( .A1(n3217), .A2(\xmem_data[40][1] ), .B1(n27831), .B2(
        \xmem_data[41][1] ), .ZN(n20425) );
  AOI22_X1 U24449 ( .A1(n20598), .A2(\xmem_data[42][1] ), .B1(n3341), .B2(
        \xmem_data[43][1] ), .ZN(n20424) );
  AOI22_X1 U24450 ( .A1(n29104), .A2(\xmem_data[44][1] ), .B1(n25377), .B2(
        \xmem_data[45][1] ), .ZN(n20423) );
  AOI22_X1 U24451 ( .A1(n29045), .A2(\xmem_data[46][1] ), .B1(n27551), .B2(
        \xmem_data[47][1] ), .ZN(n20422) );
  NAND4_X1 U24452 ( .A1(n20425), .A2(n20424), .A3(n20423), .A4(n20422), .ZN(
        n20436) );
  AOI22_X1 U24453 ( .A1(n20588), .A2(\xmem_data[48][1] ), .B1(n20587), .B2(
        \xmem_data[49][1] ), .ZN(n20429) );
  AOI22_X1 U24454 ( .A1(n25605), .A2(\xmem_data[50][1] ), .B1(n27537), .B2(
        \xmem_data[51][1] ), .ZN(n20428) );
  AOI22_X1 U24455 ( .A1(n20584), .A2(\xmem_data[52][1] ), .B1(n3121), .B2(
        \xmem_data[53][1] ), .ZN(n20427) );
  AOI22_X1 U24456 ( .A1(n20586), .A2(\xmem_data[54][1] ), .B1(n20585), .B2(
        \xmem_data[55][1] ), .ZN(n20426) );
  NAND4_X1 U24457 ( .A1(n20429), .A2(n20428), .A3(n20427), .A4(n20426), .ZN(
        n20435) );
  AOI22_X1 U24458 ( .A1(n25715), .A2(\xmem_data[56][1] ), .B1(n17021), .B2(
        \xmem_data[57][1] ), .ZN(n20433) );
  AOI22_X1 U24459 ( .A1(n25399), .A2(\xmem_data[58][1] ), .B1(n29100), .B2(
        \xmem_data[59][1] ), .ZN(n20432) );
  AOI22_X1 U24460 ( .A1(n24117), .A2(\xmem_data[60][1] ), .B1(n24522), .B2(
        \xmem_data[61][1] ), .ZN(n20431) );
  AOI22_X1 U24461 ( .A1(n30599), .A2(\xmem_data[62][1] ), .B1(n30497), .B2(
        \xmem_data[63][1] ), .ZN(n20430) );
  NAND4_X1 U24462 ( .A1(n20433), .A2(n20432), .A3(n20431), .A4(n20430), .ZN(
        n20434) );
  OR4_X1 U24463 ( .A1(n20437), .A2(n20436), .A3(n20435), .A4(n20434), .ZN(
        n20438) );
  NAND2_X1 U24464 ( .A1(n20438), .A2(n20606), .ZN(n20486) );
  AOI22_X1 U24465 ( .A1(n25520), .A2(\xmem_data[88][1] ), .B1(n29319), .B2(
        \xmem_data[89][1] ), .ZN(n20442) );
  AOI22_X1 U24466 ( .A1(n24709), .A2(\xmem_data[90][1] ), .B1(n28493), .B2(
        \xmem_data[91][1] ), .ZN(n20441) );
  AOI22_X1 U24467 ( .A1(n20551), .A2(\xmem_data[92][1] ), .B1(n3269), .B2(
        \xmem_data[93][1] ), .ZN(n20440) );
  AOI22_X1 U24468 ( .A1(n20553), .A2(\xmem_data[94][1] ), .B1(n20552), .B2(
        \xmem_data[95][1] ), .ZN(n20439) );
  NAND4_X1 U24469 ( .A1(n20442), .A2(n20441), .A3(n20440), .A4(n20439), .ZN(
        n20448) );
  AOI22_X1 U24470 ( .A1(n20546), .A2(\xmem_data[80][1] ), .B1(n20545), .B2(
        \xmem_data[81][1] ), .ZN(n20446) );
  AOI22_X1 U24471 ( .A1(n30552), .A2(\xmem_data[82][1] ), .B1(n20495), .B2(
        \xmem_data[83][1] ), .ZN(n20445) );
  AOI22_X1 U24472 ( .A1(n20544), .A2(\xmem_data[84][1] ), .B1(n17018), .B2(
        \xmem_data[85][1] ), .ZN(n20444) );
  AOI22_X1 U24473 ( .A1(n20543), .A2(\xmem_data[86][1] ), .B1(n20542), .B2(
        \xmem_data[87][1] ), .ZN(n20443) );
  NAND4_X1 U24474 ( .A1(n20446), .A2(n20445), .A3(n20444), .A4(n20443), .ZN(
        n20447) );
  NOR2_X1 U24475 ( .A1(n20448), .A2(n20447), .ZN(n20460) );
  AOI22_X1 U24476 ( .A1(n20568), .A2(\xmem_data[70][1] ), .B1(n20576), .B2(
        \xmem_data[71][1] ), .ZN(n20459) );
  AOI22_X1 U24477 ( .A1(n28500), .A2(\xmem_data[64][1] ), .B1(n20567), .B2(
        \xmem_data[65][1] ), .ZN(n20458) );
  AOI22_X1 U24478 ( .A1(n3220), .A2(\xmem_data[72][1] ), .B1(n29431), .B2(
        \xmem_data[73][1] ), .ZN(n20452) );
  AOI22_X1 U24479 ( .A1(n20558), .A2(\xmem_data[74][1] ), .B1(n25449), .B2(
        \xmem_data[75][1] ), .ZN(n20451) );
  AOI22_X1 U24480 ( .A1(n20559), .A2(\xmem_data[76][1] ), .B1(n16973), .B2(
        \xmem_data[77][1] ), .ZN(n20450) );
  AOI22_X1 U24481 ( .A1(n3231), .A2(\xmem_data[78][1] ), .B1(n27551), .B2(
        \xmem_data[79][1] ), .ZN(n20449) );
  NAND4_X1 U24482 ( .A1(n20452), .A2(n20451), .A3(n20450), .A4(n20449), .ZN(
        n20456) );
  AOI22_X1 U24483 ( .A1(n30861), .A2(\xmem_data[68][1] ), .B1(n20828), .B2(
        \xmem_data[69][1] ), .ZN(n20454) );
  AOI22_X1 U24484 ( .A1(n13487), .A2(\xmem_data[66][1] ), .B1(n3380), .B2(
        \xmem_data[67][1] ), .ZN(n20453) );
  NAND2_X1 U24485 ( .A1(n20454), .A2(n20453), .ZN(n20455) );
  NOR2_X1 U24486 ( .A1(n20456), .A2(n20455), .ZN(n20457) );
  NAND4_X1 U24487 ( .A1(n20460), .A2(n20459), .A3(n20458), .A4(n20457), .ZN(
        n20462) );
  NOR2_X1 U24488 ( .A1(n3232), .A2(n39015), .ZN(n20461) );
  AOI21_X1 U24489 ( .B1(n20462), .B2(n20573), .A(n3892), .ZN(n20485) );
  AOI22_X1 U24490 ( .A1(n30544), .A2(\xmem_data[120][1] ), .B1(n28781), .B2(
        \xmem_data[121][1] ), .ZN(n20466) );
  AOI22_X1 U24491 ( .A1(n27460), .A2(\xmem_data[122][1] ), .B1(n27462), .B2(
        \xmem_data[123][1] ), .ZN(n20465) );
  AOI22_X1 U24492 ( .A1(n20551), .A2(\xmem_data[124][1] ), .B1(n17004), .B2(
        \xmem_data[125][1] ), .ZN(n20464) );
  AOI22_X1 U24493 ( .A1(n20553), .A2(\xmem_data[126][1] ), .B1(n20552), .B2(
        \xmem_data[127][1] ), .ZN(n20463) );
  NAND4_X1 U24494 ( .A1(n20466), .A2(n20465), .A3(n20464), .A4(n20463), .ZN(
        n20475) );
  AOI22_X1 U24495 ( .A1(n3221), .A2(\xmem_data[104][1] ), .B1(n24632), .B2(
        \xmem_data[105][1] ), .ZN(n20470) );
  AOI22_X1 U24496 ( .A1(n20558), .A2(\xmem_data[106][1] ), .B1(n20807), .B2(
        \xmem_data[107][1] ), .ZN(n20469) );
  AOI22_X1 U24497 ( .A1(n20559), .A2(\xmem_data[108][1] ), .B1(n16973), .B2(
        \xmem_data[109][1] ), .ZN(n20468) );
  AOI22_X1 U24498 ( .A1(n24553), .A2(\xmem_data[110][1] ), .B1(n31321), .B2(
        \xmem_data[111][1] ), .ZN(n20467) );
  NAND4_X1 U24499 ( .A1(n20470), .A2(n20469), .A3(n20468), .A4(n20467), .ZN(
        n20474) );
  AOI22_X1 U24500 ( .A1(n31346), .A2(\xmem_data[100][1] ), .B1(n27813), .B2(
        \xmem_data[101][1] ), .ZN(n20472) );
  AOI22_X1 U24501 ( .A1(n27435), .A2(\xmem_data[98][1] ), .B1(n30588), .B2(
        \xmem_data[99][1] ), .ZN(n20471) );
  NAND2_X1 U24502 ( .A1(n20472), .A2(n20471), .ZN(n20473) );
  NOR3_X1 U24503 ( .A1(n20475), .A2(n20474), .A3(n20473), .ZN(n20482) );
  AOI22_X1 U24504 ( .A1(n28468), .A2(\xmem_data[96][1] ), .B1(n20567), .B2(
        \xmem_data[97][1] ), .ZN(n20481) );
  AOI22_X1 U24505 ( .A1(n20568), .A2(\xmem_data[102][1] ), .B1(n30592), .B2(
        \xmem_data[103][1] ), .ZN(n20480) );
  AOI22_X1 U24506 ( .A1(n20546), .A2(\xmem_data[112][1] ), .B1(n20545), .B2(
        \xmem_data[113][1] ), .ZN(n20479) );
  AOI22_X1 U24507 ( .A1(n14998), .A2(\xmem_data[114][1] ), .B1(n29023), .B2(
        \xmem_data[115][1] ), .ZN(n20478) );
  AOI22_X1 U24508 ( .A1(n20544), .A2(\xmem_data[116][1] ), .B1(n16988), .B2(
        \xmem_data[117][1] ), .ZN(n20477) );
  AOI22_X1 U24509 ( .A1(n20543), .A2(\xmem_data[118][1] ), .B1(n20542), .B2(
        \xmem_data[119][1] ), .ZN(n20476) );
  NAND4_X1 U24510 ( .A1(n20482), .A2(n20481), .A3(n20480), .A4(n3767), .ZN(
        n20483) );
  NAND2_X1 U24511 ( .A1(n20483), .A2(n20538), .ZN(n20484) );
  AOI22_X1 U24512 ( .A1(n20488), .A2(\xmem_data[0][0] ), .B1(n28192), .B2(
        \xmem_data[1][0] ), .ZN(n20494) );
  AOI22_X1 U24513 ( .A1(n27435), .A2(\xmem_data[2][0] ), .B1(n27436), .B2(
        \xmem_data[3][0] ), .ZN(n20493) );
  AOI22_X1 U24514 ( .A1(n20489), .A2(\xmem_data[4][0] ), .B1(n28164), .B2(
        \xmem_data[5][0] ), .ZN(n20492) );
  AND2_X1 U24515 ( .A1(n25485), .A2(\xmem_data[6][0] ), .ZN(n20490) );
  AOI21_X1 U24516 ( .B1(n20576), .B2(\xmem_data[7][0] ), .A(n20490), .ZN(
        n20491) );
  NAND4_X1 U24517 ( .A1(n20494), .A2(n20493), .A3(n20492), .A4(n20491), .ZN(
        n20517) );
  AOI22_X1 U24518 ( .A1(n24212), .A2(\xmem_data[18][0] ), .B1(n27537), .B2(
        \xmem_data[19][0] ), .ZN(n20499) );
  AOI22_X1 U24519 ( .A1(n28517), .A2(\xmem_data[20][0] ), .B1(n30543), .B2(
        \xmem_data[21][0] ), .ZN(n20498) );
  AOI22_X1 U24520 ( .A1(n3212), .A2(\xmem_data[22][0] ), .B1(n28059), .B2(
        \xmem_data[23][0] ), .ZN(n20497) );
  AOI22_X1 U24521 ( .A1(n24158), .A2(\xmem_data[16][0] ), .B1(n30886), .B2(
        \xmem_data[17][0] ), .ZN(n20496) );
  NAND4_X1 U24522 ( .A1(n20499), .A2(n20498), .A3(n20497), .A4(n20496), .ZN(
        n20514) );
  AOI22_X1 U24523 ( .A1(n3222), .A2(\xmem_data[8][0] ), .B1(n23770), .B2(
        \xmem_data[9][0] ), .ZN(n20504) );
  AOI22_X1 U24524 ( .A1(n20500), .A2(\xmem_data[10][0] ), .B1(n25617), .B2(
        \xmem_data[11][0] ), .ZN(n20503) );
  AOI22_X1 U24525 ( .A1(n22711), .A2(\xmem_data[12][0] ), .B1(n25377), .B2(
        \xmem_data[13][0] ), .ZN(n20502) );
  AOI22_X1 U24526 ( .A1(n25450), .A2(\xmem_data[14][0] ), .B1(n27447), .B2(
        \xmem_data[15][0] ), .ZN(n20501) );
  NAND4_X1 U24527 ( .A1(n20504), .A2(n20503), .A3(n20502), .A4(n20501), .ZN(
        n20513) );
  AOI22_X1 U24528 ( .A1(n20505), .A2(\xmem_data[24][0] ), .B1(n27855), .B2(
        \xmem_data[25][0] ), .ZN(n20511) );
  AOI22_X1 U24529 ( .A1(n13481), .A2(\xmem_data[26][0] ), .B1(n28385), .B2(
        \xmem_data[27][0] ), .ZN(n20510) );
  AOI22_X1 U24530 ( .A1(n3372), .A2(\xmem_data[28][0] ), .B1(n29324), .B2(
        \xmem_data[29][0] ), .ZN(n20509) );
  AOI22_X1 U24531 ( .A1(n20507), .A2(\xmem_data[30][0] ), .B1(n24166), .B2(
        \xmem_data[31][0] ), .ZN(n20508) );
  NAND4_X1 U24532 ( .A1(n20511), .A2(n20510), .A3(n20509), .A4(n20508), .ZN(
        n20512) );
  OAI21_X1 U24533 ( .B1(n20517), .B2(n20516), .A(n20515), .ZN(n20612) );
  AOI22_X1 U24534 ( .A1(n22751), .A2(\xmem_data[96][0] ), .B1(n20567), .B2(
        \xmem_data[97][0] ), .ZN(n20522) );
  AOI22_X1 U24535 ( .A1(n29248), .A2(\xmem_data[98][0] ), .B1(n25358), .B2(
        \xmem_data[99][0] ), .ZN(n20521) );
  AOI22_X1 U24536 ( .A1(n25357), .A2(\xmem_data[100][0] ), .B1(n28245), .B2(
        \xmem_data[101][0] ), .ZN(n20520) );
  AOI22_X1 U24537 ( .A1(n20568), .A2(\xmem_data[102][0] ), .B1(n20518), .B2(
        \xmem_data[103][0] ), .ZN(n20519) );
  NAND4_X1 U24538 ( .A1(n20522), .A2(n20521), .A3(n20520), .A4(n20519), .ZN(
        n20540) );
  AOI22_X1 U24539 ( .A1(n22740), .A2(\xmem_data[114][0] ), .B1(n20495), .B2(
        \xmem_data[115][0] ), .ZN(n20526) );
  AOI22_X1 U24540 ( .A1(n20544), .A2(\xmem_data[116][0] ), .B1(n31354), .B2(
        \xmem_data[117][0] ), .ZN(n20525) );
  AOI22_X1 U24541 ( .A1(n20543), .A2(\xmem_data[118][0] ), .B1(n20542), .B2(
        \xmem_data[119][0] ), .ZN(n20524) );
  AOI22_X1 U24542 ( .A1(n20546), .A2(\xmem_data[112][0] ), .B1(n20545), .B2(
        \xmem_data[113][0] ), .ZN(n20523) );
  NAND4_X1 U24543 ( .A1(n20526), .A2(n20525), .A3(n20524), .A4(n20523), .ZN(
        n20537) );
  AOI22_X1 U24544 ( .A1(n22718), .A2(\xmem_data[120][0] ), .B1(n21050), .B2(
        \xmem_data[121][0] ), .ZN(n20530) );
  AOI22_X1 U24545 ( .A1(n29238), .A2(\xmem_data[122][0] ), .B1(n3325), .B2(
        \xmem_data[123][0] ), .ZN(n20529) );
  AOI22_X1 U24546 ( .A1(n20551), .A2(\xmem_data[124][0] ), .B1(n29246), .B2(
        \xmem_data[125][0] ), .ZN(n20528) );
  AOI22_X1 U24547 ( .A1(n20553), .A2(\xmem_data[126][0] ), .B1(n20552), .B2(
        \xmem_data[127][0] ), .ZN(n20527) );
  NAND4_X1 U24548 ( .A1(n20530), .A2(n20529), .A3(n20528), .A4(n20527), .ZN(
        n20536) );
  AOI22_X1 U24549 ( .A1(n3222), .A2(\xmem_data[104][0] ), .B1(n17033), .B2(
        \xmem_data[105][0] ), .ZN(n20534) );
  AOI22_X1 U24550 ( .A1(n20558), .A2(\xmem_data[106][0] ), .B1(n29289), .B2(
        \xmem_data[107][0] ), .ZN(n20533) );
  AOI22_X1 U24551 ( .A1(n20559), .A2(\xmem_data[108][0] ), .B1(n27396), .B2(
        \xmem_data[109][0] ), .ZN(n20532) );
  AOI22_X1 U24552 ( .A1(n29306), .A2(\xmem_data[110][0] ), .B1(n20809), .B2(
        \xmem_data[111][0] ), .ZN(n20531) );
  NAND4_X1 U24553 ( .A1(n20534), .A2(n20533), .A3(n20532), .A4(n20531), .ZN(
        n20535) );
  OAI21_X1 U24554 ( .B1(n20540), .B2(n20539), .A(n20538), .ZN(n20611) );
  AOI22_X1 U24555 ( .A1(n24132), .A2(\xmem_data[82][0] ), .B1(n20495), .B2(
        \xmem_data[83][0] ), .ZN(n20550) );
  AOI22_X1 U24556 ( .A1(n20543), .A2(\xmem_data[86][0] ), .B1(n20542), .B2(
        \xmem_data[87][0] ), .ZN(n20549) );
  AOI22_X1 U24557 ( .A1(n20544), .A2(\xmem_data[84][0] ), .B1(n28091), .B2(
        \xmem_data[85][0] ), .ZN(n20548) );
  AOI22_X1 U24558 ( .A1(n20546), .A2(\xmem_data[80][0] ), .B1(n20545), .B2(
        \xmem_data[81][0] ), .ZN(n20547) );
  NAND4_X1 U24559 ( .A1(n20550), .A2(n20549), .A3(n20548), .A4(n20547), .ZN(
        n20566) );
  AOI22_X1 U24560 ( .A1(n25398), .A2(\xmem_data[88][0] ), .B1(n29012), .B2(
        \xmem_data[89][0] ), .ZN(n20557) );
  AOI22_X1 U24561 ( .A1(n24460), .A2(\xmem_data[90][0] ), .B1(n3325), .B2(
        \xmem_data[91][0] ), .ZN(n20556) );
  AOI22_X1 U24562 ( .A1(n20551), .A2(\xmem_data[92][0] ), .B1(n25718), .B2(
        \xmem_data[93][0] ), .ZN(n20555) );
  AOI22_X1 U24563 ( .A1(n20553), .A2(\xmem_data[94][0] ), .B1(n20552), .B2(
        \xmem_data[95][0] ), .ZN(n20554) );
  NAND4_X1 U24564 ( .A1(n20557), .A2(n20556), .A3(n20555), .A4(n20554), .ZN(
        n20565) );
  AOI22_X1 U24565 ( .A1(n3219), .A2(\xmem_data[72][0] ), .B1(n22708), .B2(
        \xmem_data[73][0] ), .ZN(n20563) );
  AOI22_X1 U24566 ( .A1(n20558), .A2(\xmem_data[74][0] ), .B1(n23812), .B2(
        \xmem_data[75][0] ), .ZN(n20562) );
  AOI22_X1 U24567 ( .A1(n20559), .A2(\xmem_data[76][0] ), .B1(n29157), .B2(
        \xmem_data[77][0] ), .ZN(n20561) );
  AOI22_X1 U24568 ( .A1(n24657), .A2(\xmem_data[78][0] ), .B1(n25422), .B2(
        \xmem_data[79][0] ), .ZN(n20560) );
  NAND4_X1 U24569 ( .A1(n20563), .A2(n20562), .A3(n20561), .A4(n20560), .ZN(
        n20564) );
  AOI22_X1 U24570 ( .A1(n28500), .A2(\xmem_data[64][0] ), .B1(n20567), .B2(
        \xmem_data[65][0] ), .ZN(n20572) );
  AOI22_X1 U24571 ( .A1(n16999), .A2(\xmem_data[66][0] ), .B1(n24526), .B2(
        \xmem_data[67][0] ), .ZN(n20571) );
  AOI22_X1 U24572 ( .A1(n22729), .A2(\xmem_data[68][0] ), .B1(n23732), .B2(
        \xmem_data[69][0] ), .ZN(n20570) );
  AOI22_X1 U24573 ( .A1(n20568), .A2(\xmem_data[70][0] ), .B1(n24443), .B2(
        \xmem_data[71][0] ), .ZN(n20569) );
  NAND4_X1 U24574 ( .A1(n20572), .A2(n20571), .A3(n20570), .A4(n20569), .ZN(
        n20574) );
  OAI21_X1 U24575 ( .B1(n20575), .B2(n20574), .A(n20573), .ZN(n20610) );
  AOI22_X1 U24576 ( .A1(n31347), .A2(\xmem_data[38][0] ), .B1(n20576), .B2(
        \xmem_data[39][0] ), .ZN(n20583) );
  AOI22_X1 U24577 ( .A1(n28328), .A2(\xmem_data[32][0] ), .B1(n20577), .B2(
        \xmem_data[33][0] ), .ZN(n20582) );
  AOI22_X1 U24578 ( .A1(n20578), .A2(\xmem_data[36][0] ), .B1(n3142), .B2(
        \xmem_data[37][0] ), .ZN(n20581) );
  AOI22_X1 U24579 ( .A1(n20579), .A2(\xmem_data[34][0] ), .B1(n25724), .B2(
        \xmem_data[35][0] ), .ZN(n20580) );
  NAND4_X1 U24580 ( .A1(n20583), .A2(n20582), .A3(n20581), .A4(n20580), .ZN(
        n20608) );
  AOI22_X1 U24581 ( .A1(n20584), .A2(\xmem_data[52][0] ), .B1(n27945), .B2(
        \xmem_data[53][0] ), .ZN(n20592) );
  AOI22_X1 U24582 ( .A1(n29232), .A2(\xmem_data[50][0] ), .B1(n28980), .B2(
        \xmem_data[51][0] ), .ZN(n20591) );
  AOI22_X1 U24583 ( .A1(n20586), .A2(\xmem_data[54][0] ), .B1(n20585), .B2(
        \xmem_data[55][0] ), .ZN(n20590) );
  AOI22_X1 U24584 ( .A1(n20588), .A2(\xmem_data[48][0] ), .B1(n20587), .B2(
        \xmem_data[49][0] ), .ZN(n20589) );
  NAND4_X1 U24585 ( .A1(n20592), .A2(n20591), .A3(n20590), .A4(n20589), .ZN(
        n20605) );
  AOI22_X1 U24586 ( .A1(n24459), .A2(\xmem_data[56][0] ), .B1(n27855), .B2(
        \xmem_data[57][0] ), .ZN(n20597) );
  AOI22_X1 U24587 ( .A1(n27523), .A2(\xmem_data[58][0] ), .B1(n20593), .B2(
        \xmem_data[59][0] ), .ZN(n20596) );
  AOI22_X1 U24588 ( .A1(n23778), .A2(\xmem_data[60][0] ), .B1(n20950), .B2(
        \xmem_data[61][0] ), .ZN(n20595) );
  AOI22_X1 U24589 ( .A1(n14975), .A2(\xmem_data[62][0] ), .B1(n20552), .B2(
        \xmem_data[63][0] ), .ZN(n20594) );
  NAND4_X1 U24590 ( .A1(n20597), .A2(n20596), .A3(n20595), .A4(n20594), .ZN(
        n20604) );
  AOI22_X1 U24591 ( .A1(n3222), .A2(\xmem_data[40][0] ), .B1(n29065), .B2(
        \xmem_data[41][0] ), .ZN(n20602) );
  AOI22_X1 U24592 ( .A1(n20598), .A2(\xmem_data[42][0] ), .B1(n29289), .B2(
        \xmem_data[43][0] ), .ZN(n20601) );
  AOI22_X1 U24593 ( .A1(n27550), .A2(\xmem_data[44][0] ), .B1(n22668), .B2(
        \xmem_data[45][0] ), .ZN(n20600) );
  AOI22_X1 U24594 ( .A1(n3231), .A2(\xmem_data[46][0] ), .B1(n25604), .B2(
        \xmem_data[47][0] ), .ZN(n20599) );
  NAND4_X1 U24595 ( .A1(n20602), .A2(n20601), .A3(n20600), .A4(n20599), .ZN(
        n20603) );
  OAI21_X1 U24596 ( .B1(n20608), .B2(n20607), .A(n20606), .ZN(n20609) );
  XNOR2_X1 U24597 ( .A(n35120), .B(\fmem_data[6][1] ), .ZN(n31955) );
  AOI22_X1 U24598 ( .A1(n25707), .A2(\xmem_data[32][6] ), .B1(n3358), .B2(
        \xmem_data[33][6] ), .ZN(n20617) );
  AOI22_X1 U24599 ( .A1(n25708), .A2(\xmem_data[34][6] ), .B1(n22702), .B2(
        \xmem_data[35][6] ), .ZN(n20616) );
  AOI22_X1 U24600 ( .A1(n28980), .A2(\xmem_data[36][6] ), .B1(n25709), .B2(
        \xmem_data[37][6] ), .ZN(n20615) );
  AOI22_X1 U24601 ( .A1(n24545), .A2(\xmem_data[38][6] ), .B1(n31269), .B2(
        \xmem_data[39][6] ), .ZN(n20614) );
  NAND4_X1 U24602 ( .A1(n20617), .A2(n20616), .A3(n20615), .A4(n20614), .ZN(
        n20633) );
  AOI22_X1 U24603 ( .A1(n24509), .A2(\xmem_data[40][6] ), .B1(n25715), .B2(
        \xmem_data[41][6] ), .ZN(n20621) );
  AOI22_X1 U24604 ( .A1(n20815), .A2(\xmem_data[42][6] ), .B1(n25435), .B2(
        \xmem_data[43][6] ), .ZN(n20620) );
  AOI22_X1 U24605 ( .A1(n3325), .A2(\xmem_data[44][6] ), .B1(n3372), .B2(
        \xmem_data[45][6] ), .ZN(n20619) );
  AOI22_X1 U24606 ( .A1(n25718), .A2(\xmem_data[46][6] ), .B1(n20507), .B2(
        \xmem_data[47][6] ), .ZN(n20618) );
  NAND4_X1 U24607 ( .A1(n20621), .A2(n20620), .A3(n20619), .A4(n20618), .ZN(
        n20632) );
  AOI22_X1 U24608 ( .A1(n20782), .A2(\xmem_data[48][6] ), .B1(n25723), .B2(
        \xmem_data[49][6] ), .ZN(n20625) );
  AOI22_X1 U24609 ( .A1(n27568), .A2(\xmem_data[50][6] ), .B1(n31261), .B2(
        \xmem_data[51][6] ), .ZN(n20624) );
  AOI22_X1 U24610 ( .A1(n25724), .A2(\xmem_data[52][6] ), .B1(n24470), .B2(
        \xmem_data[53][6] ), .ZN(n20623) );
  AOI22_X1 U24611 ( .A1(n25725), .A2(\xmem_data[54][6] ), .B1(n20568), .B2(
        \xmem_data[55][6] ), .ZN(n20622) );
  NAND4_X1 U24612 ( .A1(n20625), .A2(n20624), .A3(n20623), .A4(n20622), .ZN(
        n20631) );
  AOI22_X1 U24613 ( .A1(n25730), .A2(\xmem_data[56][6] ), .B1(n3222), .B2(
        \xmem_data[57][6] ), .ZN(n20629) );
  AOI22_X1 U24614 ( .A1(n25731), .A2(\xmem_data[58][6] ), .B1(n20723), .B2(
        \xmem_data[59][6] ), .ZN(n20628) );
  AOI22_X1 U24615 ( .A1(n29174), .A2(\xmem_data[60][6] ), .B1(n25486), .B2(
        \xmem_data[61][6] ), .ZN(n20627) );
  AOI22_X1 U24616 ( .A1(n25732), .A2(\xmem_data[62][6] ), .B1(n3231), .B2(
        \xmem_data[63][6] ), .ZN(n20626) );
  NAND4_X1 U24617 ( .A1(n20629), .A2(n20628), .A3(n20627), .A4(n20626), .ZN(
        n20630) );
  OR4_X1 U24618 ( .A1(n20633), .A2(n20632), .A3(n20631), .A4(n20630), .ZN(
        n20661) );
  AOI22_X1 U24619 ( .A1(n28318), .A2(\xmem_data[24][6] ), .B1(n3217), .B2(
        \xmem_data[25][6] ), .ZN(n20640) );
  AOI22_X1 U24620 ( .A1(n25617), .A2(\xmem_data[28][6] ), .B1(n25616), .B2(
        \xmem_data[29][6] ), .ZN(n20634) );
  INV_X1 U24621 ( .A(n20634), .ZN(n20638) );
  AOI22_X1 U24622 ( .A1(n25612), .A2(\xmem_data[26][6] ), .B1(n29255), .B2(
        \xmem_data[27][6] ), .ZN(n20636) );
  NAND2_X1 U24623 ( .A1(n3281), .A2(\xmem_data[30][6] ), .ZN(n20635) );
  NAND2_X1 U24624 ( .A1(n20636), .A2(n20635), .ZN(n20637) );
  NOR2_X1 U24625 ( .A1(n20638), .A2(n20637), .ZN(n20639) );
  NAND2_X1 U24626 ( .A1(n20640), .A2(n20639), .ZN(n20648) );
  AOI22_X1 U24627 ( .A1(n25628), .A2(\xmem_data[18][6] ), .B1(n22727), .B2(
        \xmem_data[19][6] ), .ZN(n20646) );
  AND2_X1 U24628 ( .A1(n25630), .A2(\xmem_data[20][6] ), .ZN(n20644) );
  AOI22_X1 U24629 ( .A1(n27847), .A2(\xmem_data[16][6] ), .B1(n27526), .B2(
        \xmem_data[17][6] ), .ZN(n20642) );
  AOI22_X1 U24630 ( .A1(n25624), .A2(\xmem_data[22][6] ), .B1(n30589), .B2(
        \xmem_data[23][6] ), .ZN(n20641) );
  NAND2_X1 U24631 ( .A1(n20642), .A2(n20641), .ZN(n20643) );
  AOI211_X1 U24632 ( .C1(n25629), .C2(\xmem_data[21][6] ), .A(n20644), .B(
        n20643), .ZN(n20645) );
  NAND2_X1 U24633 ( .A1(n20646), .A2(n20645), .ZN(n20647) );
  NOR2_X1 U24634 ( .A1(n20648), .A2(n20647), .ZN(n20659) );
  AOI22_X1 U24635 ( .A1(n25604), .A2(\xmem_data[0][6] ), .B1(n25456), .B2(
        \xmem_data[1][6] ), .ZN(n20652) );
  AOI22_X1 U24636 ( .A1(n29403), .A2(\xmem_data[2][6] ), .B1(n25605), .B2(
        \xmem_data[3][6] ), .ZN(n20651) );
  AOI22_X1 U24637 ( .A1(n17041), .A2(\xmem_data[4][6] ), .B1(n25606), .B2(
        \xmem_data[5][6] ), .ZN(n20650) );
  AOI22_X1 U24638 ( .A1(n28516), .A2(\xmem_data[6][6] ), .B1(n29162), .B2(
        \xmem_data[7][6] ), .ZN(n20649) );
  NAND4_X1 U24639 ( .A1(n20652), .A2(n20651), .A3(n20650), .A4(n20649), .ZN(
        n20658) );
  AOI22_X1 U24640 ( .A1(n25635), .A2(\xmem_data[8][6] ), .B1(n29316), .B2(
        \xmem_data[9][6] ), .ZN(n20656) );
  AOI22_X1 U24641 ( .A1(n25400), .A2(\xmem_data[10][6] ), .B1(n29049), .B2(
        \xmem_data[11][6] ), .ZN(n20655) );
  AOI22_X1 U24642 ( .A1(n25632), .A2(\xmem_data[12][6] ), .B1(n27951), .B2(
        \xmem_data[13][6] ), .ZN(n20654) );
  AOI22_X1 U24643 ( .A1(n25636), .A2(\xmem_data[14][6] ), .B1(n31362), .B2(
        \xmem_data[15][6] ), .ZN(n20653) );
  NAND4_X1 U24644 ( .A1(n20656), .A2(n20655), .A3(n20654), .A4(n20653), .ZN(
        n20657) );
  AOI21_X1 U24645 ( .B1(n20659), .B2(n3549), .A(n25647), .ZN(n20660) );
  AOI21_X1 U24646 ( .B1(n20661), .B2(n25741), .A(n20660), .ZN(n20706) );
  AOI22_X1 U24647 ( .A1(n25670), .A2(\xmem_data[96][6] ), .B1(n24130), .B2(
        \xmem_data[97][6] ), .ZN(n20665) );
  AOI22_X1 U24648 ( .A1(n27911), .A2(\xmem_data[98][6] ), .B1(n25605), .B2(
        \xmem_data[99][6] ), .ZN(n20664) );
  AOI22_X1 U24649 ( .A1(n16986), .A2(\xmem_data[100][6] ), .B1(n25671), .B2(
        \xmem_data[101][6] ), .ZN(n20663) );
  AOI22_X1 U24650 ( .A1(n25672), .A2(\xmem_data[102][6] ), .B1(n28993), .B2(
        \xmem_data[103][6] ), .ZN(n20662) );
  NAND4_X1 U24651 ( .A1(n20665), .A2(n20664), .A3(n20663), .A4(n20662), .ZN(
        n20681) );
  AOI22_X1 U24652 ( .A1(n14937), .A2(\xmem_data[104][6] ), .B1(n25677), .B2(
        \xmem_data[105][6] ), .ZN(n20669) );
  AOI22_X1 U24653 ( .A1(n25678), .A2(\xmem_data[106][6] ), .B1(n29101), .B2(
        \xmem_data[107][6] ), .ZN(n20668) );
  AOI22_X1 U24654 ( .A1(n25521), .A2(\xmem_data[108][6] ), .B1(n28429), .B2(
        \xmem_data[109][6] ), .ZN(n20667) );
  AOI22_X1 U24655 ( .A1(n3151), .A2(\xmem_data[110][6] ), .B1(n31362), .B2(
        \xmem_data[111][6] ), .ZN(n20666) );
  NAND4_X1 U24656 ( .A1(n20669), .A2(n20668), .A3(n20667), .A4(n20666), .ZN(
        n20680) );
  AOI22_X1 U24657 ( .A1(n28293), .A2(\xmem_data[112][6] ), .B1(n29086), .B2(
        \xmem_data[113][6] ), .ZN(n20673) );
  AOI22_X1 U24658 ( .A1(n25684), .A2(\xmem_data[114][6] ), .B1(n27435), .B2(
        \xmem_data[115][6] ), .ZN(n20672) );
  AOI22_X1 U24659 ( .A1(n25686), .A2(\xmem_data[116][6] ), .B1(n25685), .B2(
        \xmem_data[117][6] ), .ZN(n20671) );
  AOI22_X1 U24660 ( .A1(n22728), .A2(\xmem_data[118][6] ), .B1(n25687), .B2(
        \xmem_data[119][6] ), .ZN(n20670) );
  NAND4_X1 U24661 ( .A1(n20673), .A2(n20672), .A3(n20671), .A4(n20670), .ZN(
        n20679) );
  AOI22_X1 U24662 ( .A1(n25692), .A2(\xmem_data[120][6] ), .B1(n3218), .B2(
        \xmem_data[121][6] ), .ZN(n20677) );
  AOI22_X1 U24663 ( .A1(n25693), .A2(\xmem_data[122][6] ), .B1(n25562), .B2(
        \xmem_data[123][6] ), .ZN(n20676) );
  AOI22_X1 U24664 ( .A1(n25694), .A2(\xmem_data[124][6] ), .B1(n27550), .B2(
        \xmem_data[125][6] ), .ZN(n20675) );
  AOI22_X1 U24665 ( .A1(n3134), .A2(\xmem_data[126][6] ), .B1(n28510), .B2(
        \xmem_data[127][6] ), .ZN(n20674) );
  NAND4_X1 U24666 ( .A1(n20677), .A2(n20676), .A3(n20675), .A4(n20674), .ZN(
        n20678) );
  OR4_X1 U24667 ( .A1(n20681), .A2(n20680), .A3(n20679), .A4(n20678), .ZN(
        n20704) );
  AOI22_X1 U24668 ( .A1(n25707), .A2(\xmem_data[64][6] ), .B1(n3357), .B2(
        \xmem_data[65][6] ), .ZN(n20686) );
  AOI22_X1 U24669 ( .A1(n25708), .A2(n20682), .B1(n25605), .B2(
        \xmem_data[67][6] ), .ZN(n20685) );
  AOI22_X1 U24670 ( .A1(n29023), .A2(\xmem_data[68][6] ), .B1(n25709), .B2(
        \xmem_data[69][6] ), .ZN(n20684) );
  AOI22_X1 U24671 ( .A1(n28752), .A2(\xmem_data[70][6] ), .B1(n28299), .B2(
        \xmem_data[71][6] ), .ZN(n20683) );
  NAND4_X1 U24672 ( .A1(n20686), .A2(n20685), .A3(n20684), .A4(n20683), .ZN(
        n20702) );
  AOI22_X1 U24673 ( .A1(n25635), .A2(\xmem_data[72][6] ), .B1(n25715), .B2(
        \xmem_data[73][6] ), .ZN(n20690) );
  AOI22_X1 U24674 ( .A1(n22682), .A2(\xmem_data[74][6] ), .B1(n25576), .B2(
        \xmem_data[75][6] ), .ZN(n20689) );
  AOI22_X1 U24675 ( .A1(n25717), .A2(\xmem_data[76][6] ), .B1(n30598), .B2(
        \xmem_data[77][6] ), .ZN(n20688) );
  AOI22_X1 U24676 ( .A1(n25718), .A2(\xmem_data[78][6] ), .B1(n24167), .B2(
        \xmem_data[79][6] ), .ZN(n20687) );
  NAND4_X1 U24677 ( .A1(n20690), .A2(n20689), .A3(n20688), .A4(n20687), .ZN(
        n20701) );
  AOI22_X1 U24678 ( .A1(n29325), .A2(\xmem_data[80][6] ), .B1(n25723), .B2(
        \xmem_data[81][6] ), .ZN(n20694) );
  AOI22_X1 U24679 ( .A1(n23730), .A2(\xmem_data[82][6] ), .B1(n25388), .B2(
        \xmem_data[83][6] ), .ZN(n20693) );
  AOI22_X1 U24680 ( .A1(n25724), .A2(\xmem_data[84][6] ), .B1(n29328), .B2(
        \xmem_data[85][6] ), .ZN(n20692) );
  AOI22_X1 U24681 ( .A1(n25725), .A2(\xmem_data[86][6] ), .B1(n27437), .B2(
        \xmem_data[87][6] ), .ZN(n20691) );
  NAND4_X1 U24682 ( .A1(n20694), .A2(n20693), .A3(n20692), .A4(n20691), .ZN(
        n20700) );
  AOI22_X1 U24683 ( .A1(n25730), .A2(\xmem_data[88][6] ), .B1(n3222), .B2(
        \xmem_data[89][6] ), .ZN(n20698) );
  AOI22_X1 U24684 ( .A1(n25731), .A2(\xmem_data[90][6] ), .B1(n23769), .B2(
        \xmem_data[91][6] ), .ZN(n20697) );
  AOI22_X1 U24685 ( .A1(n21069), .A2(\xmem_data[92][6] ), .B1(n3255), .B2(
        \xmem_data[93][6] ), .ZN(n20696) );
  AOI22_X1 U24686 ( .A1(n25732), .A2(\xmem_data[94][6] ), .B1(n27547), .B2(
        \xmem_data[95][6] ), .ZN(n20695) );
  NAND4_X1 U24687 ( .A1(n20698), .A2(n20697), .A3(n20696), .A4(n20695), .ZN(
        n20699) );
  OR4_X1 U24688 ( .A1(n20702), .A2(n20701), .A3(n20700), .A4(n20699), .ZN(
        n20703) );
  AOI22_X1 U24689 ( .A1(n25706), .A2(n20704), .B1(n25704), .B2(n20703), .ZN(
        n20705) );
  XNOR2_X1 U24690 ( .A(n31656), .B(\fmem_data[28][3] ), .ZN(n32644) );
  AOI22_X1 U24691 ( .A1(n20708), .A2(\xmem_data[104][4] ), .B1(n20707), .B2(
        \xmem_data[105][4] ), .ZN(n20715) );
  AOI22_X1 U24692 ( .A1(n20710), .A2(\xmem_data[106][4] ), .B1(n20709), .B2(
        \xmem_data[107][4] ), .ZN(n20714) );
  AOI22_X1 U24693 ( .A1(n3245), .A2(\xmem_data[108][4] ), .B1(n20711), .B2(
        \xmem_data[109][4] ), .ZN(n20713) );
  AOI22_X1 U24694 ( .A1(n21066), .A2(\xmem_data[110][4] ), .B1(n3220), .B2(
        \xmem_data[111][4] ), .ZN(n20712) );
  NAND4_X1 U24695 ( .A1(n20715), .A2(n20714), .A3(n20713), .A4(n20712), .ZN(
        n20744) );
  AOI22_X1 U24696 ( .A1(n20716), .A2(\xmem_data[120][4] ), .B1(n28416), .B2(
        \xmem_data[121][4] ), .ZN(n20722) );
  AOI22_X1 U24697 ( .A1(n30614), .A2(\xmem_data[122][4] ), .B1(n20717), .B2(
        \xmem_data[123][4] ), .ZN(n20721) );
  AOI22_X1 U24698 ( .A1(n29605), .A2(\xmem_data[124][4] ), .B1(n3212), .B2(
        \xmem_data[125][4] ), .ZN(n20720) );
  AOI22_X1 U24699 ( .A1(n23764), .A2(\xmem_data[126][4] ), .B1(n17043), .B2(
        \xmem_data[127][4] ), .ZN(n20719) );
  NAND4_X1 U24700 ( .A1(n20722), .A2(n20721), .A3(n20720), .A4(n20719), .ZN(
        n20741) );
  AOI22_X1 U24701 ( .A1(n20724), .A2(\xmem_data[112][4] ), .B1(n20723), .B2(
        \xmem_data[113][4] ), .ZN(n20729) );
  AOI22_X1 U24702 ( .A1(n20725), .A2(\xmem_data[114][4] ), .B1(n13444), .B2(
        \xmem_data[115][4] ), .ZN(n20728) );
  AOI22_X1 U24703 ( .A1(n20808), .A2(\xmem_data[116][4] ), .B1(n25514), .B2(
        \xmem_data[117][4] ), .ZN(n20727) );
  AOI22_X1 U24704 ( .A1(n30551), .A2(\xmem_data[118][4] ), .B1(n29180), .B2(
        \xmem_data[119][4] ), .ZN(n20726) );
  NAND4_X1 U24705 ( .A1(n20729), .A2(n20728), .A3(n20727), .A4(n20726), .ZN(
        n20740) );
  AOI22_X1 U24706 ( .A1(n20730), .A2(\xmem_data[96][4] ), .B1(n25435), .B2(
        \xmem_data[97][4] ), .ZN(n20738) );
  AOI22_X1 U24707 ( .A1(n20731), .A2(\xmem_data[98][4] ), .B1(n21009), .B2(
        \xmem_data[99][4] ), .ZN(n20737) );
  AOI22_X1 U24708 ( .A1(n20732), .A2(\xmem_data[100][4] ), .B1(n24622), .B2(
        \xmem_data[101][4] ), .ZN(n20736) );
  AOI22_X1 U24709 ( .A1(n20734), .A2(\xmem_data[102][4] ), .B1(n20733), .B2(
        \xmem_data[103][4] ), .ZN(n20735) );
  NAND4_X1 U24710 ( .A1(n20738), .A2(n20737), .A3(n20736), .A4(n20735), .ZN(
        n20739) );
  AOI22_X1 U24711 ( .A1(n20826), .A2(\xmem_data[40][4] ), .B1(n30524), .B2(
        \xmem_data[41][4] ), .ZN(n20749) );
  AOI22_X1 U24712 ( .A1(n20827), .A2(\xmem_data[42][4] ), .B1(n20578), .B2(
        \xmem_data[43][4] ), .ZN(n20748) );
  AOI22_X1 U24713 ( .A1(n20828), .A2(\xmem_data[44][4] ), .B1(n22753), .B2(
        \xmem_data[45][4] ), .ZN(n20747) );
  AND2_X1 U24714 ( .A1(n3221), .A2(\xmem_data[47][4] ), .ZN(n20745) );
  AOI21_X1 U24715 ( .B1(n28044), .B2(\xmem_data[46][4] ), .A(n20745), .ZN(
        n20746) );
  NAND4_X1 U24716 ( .A1(n20749), .A2(n20748), .A3(n20747), .A4(n20746), .ZN(
        n20767) );
  AOI22_X1 U24717 ( .A1(n29310), .A2(\xmem_data[58][4] ), .B1(n20798), .B2(
        \xmem_data[59][4] ), .ZN(n20753) );
  AOI22_X1 U24718 ( .A1(n20799), .A2(\xmem_data[56][4] ), .B1(n22702), .B2(
        \xmem_data[57][4] ), .ZN(n20752) );
  AOI22_X1 U24719 ( .A1(n20800), .A2(\xmem_data[62][4] ), .B1(n21006), .B2(
        \xmem_data[63][4] ), .ZN(n20751) );
  AOI22_X1 U24720 ( .A1(n28335), .A2(\xmem_data[61][4] ), .B1(
        \xmem_data[60][4] ), .B2(n20776), .ZN(n20750) );
  NAND4_X1 U24721 ( .A1(n20753), .A2(n20752), .A3(n20751), .A4(n20750), .ZN(
        n20764) );
  AOI22_X1 U24722 ( .A1(n20805), .A2(\xmem_data[48][4] ), .B1(n27507), .B2(
        \xmem_data[49][4] ), .ZN(n20757) );
  AOI22_X1 U24723 ( .A1(n20807), .A2(\xmem_data[50][4] ), .B1(n20806), .B2(
        \xmem_data[51][4] ), .ZN(n20756) );
  AOI22_X1 U24724 ( .A1(n20808), .A2(\xmem_data[52][4] ), .B1(n29103), .B2(
        \xmem_data[53][4] ), .ZN(n20755) );
  AOI22_X1 U24725 ( .A1(n20809), .A2(\xmem_data[54][4] ), .B1(n28415), .B2(
        \xmem_data[55][4] ), .ZN(n20754) );
  NAND4_X1 U24726 ( .A1(n20757), .A2(n20756), .A3(n20755), .A4(n20754), .ZN(
        n20763) );
  AOI22_X1 U24727 ( .A1(n20815), .A2(\xmem_data[32][4] ), .B1(n20814), .B2(
        \xmem_data[33][4] ), .ZN(n20761) );
  AOI22_X1 U24728 ( .A1(n3325), .A2(\xmem_data[34][4] ), .B1(n3372), .B2(
        \xmem_data[35][4] ), .ZN(n20760) );
  AOI22_X1 U24729 ( .A1(n20817), .A2(\xmem_data[36][4] ), .B1(n28098), .B2(
        \xmem_data[37][4] ), .ZN(n20759) );
  AOI22_X1 U24730 ( .A1(n20818), .A2(\xmem_data[38][4] ), .B1(n25527), .B2(
        \xmem_data[39][4] ), .ZN(n20758) );
  NAND4_X1 U24731 ( .A1(n20761), .A2(n20760), .A3(n20759), .A4(n20758), .ZN(
        n20762) );
  AOI22_X1 U24732 ( .A1(n30295), .A2(\xmem_data[20][4] ), .B1(n24553), .B2(
        \xmem_data[21][4] ), .ZN(n20768) );
  INV_X1 U24733 ( .A(n20768), .ZN(n20797) );
  AOI22_X1 U24734 ( .A1(n20770), .A2(\xmem_data[8][4] ), .B1(n20769), .B2(
        \xmem_data[9][4] ), .ZN(n20774) );
  AOI22_X1 U24735 ( .A1(n27925), .A2(\xmem_data[10][4] ), .B1(n29118), .B2(
        \xmem_data[11][4] ), .ZN(n20773) );
  AOI22_X1 U24736 ( .A1(n3305), .A2(\xmem_data[12][4] ), .B1(n25687), .B2(
        \xmem_data[13][4] ), .ZN(n20772) );
  AOI22_X1 U24737 ( .A1(n24562), .A2(\xmem_data[14][4] ), .B1(n3221), .B2(
        \xmem_data[15][4] ), .ZN(n20771) );
  NAND4_X1 U24738 ( .A1(n20774), .A2(n20773), .A3(n20772), .A4(n20771), .ZN(
        n20794) );
  AOI22_X1 U24739 ( .A1(n30608), .A2(\xmem_data[24][4] ), .B1(n20775), .B2(
        \xmem_data[25][4] ), .ZN(n20780) );
  AOI22_X1 U24740 ( .A1(n29023), .A2(\xmem_data[26][4] ), .B1(n25572), .B2(
        \xmem_data[27][4] ), .ZN(n20779) );
  AOI22_X1 U24741 ( .A1(n27517), .A2(\xmem_data[28][4] ), .B1(n27454), .B2(
        \xmem_data[29][4] ), .ZN(n20778) );
  AOI22_X1 U24742 ( .A1(n25635), .A2(\xmem_data[30][4] ), .B1(n20940), .B2(
        \xmem_data[31][4] ), .ZN(n20777) );
  NAND4_X1 U24743 ( .A1(n20780), .A2(n20779), .A3(n20778), .A4(n20777), .ZN(
        n20793) );
  AOI22_X1 U24744 ( .A1(n23802), .A2(\xmem_data[0][4] ), .B1(n28380), .B2(
        \xmem_data[1][4] ), .ZN(n20786) );
  AOI22_X1 U24745 ( .A1(n14881), .A2(\xmem_data[2][4] ), .B1(n29281), .B2(
        \xmem_data[3][4] ), .ZN(n20785) );
  AOI22_X1 U24746 ( .A1(n25636), .A2(\xmem_data[4][4] ), .B1(n20781), .B2(
        \xmem_data[5][4] ), .ZN(n20784) );
  AOI22_X1 U24747 ( .A1(n20782), .A2(\xmem_data[6][4] ), .B1(n11008), .B2(
        \xmem_data[7][4] ), .ZN(n20783) );
  NAND4_X1 U24748 ( .A1(n20786), .A2(n20785), .A3(n20784), .A4(n20783), .ZN(
        n20792) );
  AOI22_X1 U24749 ( .A1(n25617), .A2(\xmem_data[18][4] ), .B1(n13444), .B2(
        \xmem_data[19][4] ), .ZN(n20790) );
  AOI22_X1 U24750 ( .A1(n27447), .A2(\xmem_data[22][4] ), .B1(n24590), .B2(
        \xmem_data[23][4] ), .ZN(n20789) );
  AOI22_X1 U24751 ( .A1(n29698), .A2(\xmem_data[16][4] ), .B1(n20787), .B2(
        \xmem_data[17][4] ), .ZN(n20788) );
  NAND3_X1 U24752 ( .A1(n20790), .A2(n20789), .A3(n20788), .ZN(n20791) );
  OR4_X1 U24753 ( .A1(n20794), .A2(n20793), .A3(n20792), .A4(n20791), .ZN(
        n20796) );
  OAI21_X1 U24754 ( .B1(n20797), .B2(n20796), .A(n20795), .ZN(n20837) );
  AOI22_X1 U24755 ( .A1(n27515), .A2(\xmem_data[90][4] ), .B1(n20798), .B2(
        \xmem_data[91][4] ), .ZN(n20804) );
  AOI22_X1 U24756 ( .A1(n20799), .A2(\xmem_data[88][4] ), .B1(n22740), .B2(
        \xmem_data[89][4] ), .ZN(n20803) );
  AOI22_X1 U24757 ( .A1(n20800), .A2(\xmem_data[94][4] ), .B1(n25715), .B2(
        \xmem_data[95][4] ), .ZN(n20802) );
  AOI22_X1 U24758 ( .A1(n24134), .A2(\xmem_data[93][4] ), .B1(
        \xmem_data[92][4] ), .B2(n3158), .ZN(n20801) );
  NAND4_X1 U24759 ( .A1(n20804), .A2(n20803), .A3(n20802), .A4(n20801), .ZN(
        n20825) );
  AOI22_X1 U24760 ( .A1(n20805), .A2(\xmem_data[80][4] ), .B1(n20723), .B2(
        \xmem_data[81][4] ), .ZN(n20813) );
  AOI22_X1 U24761 ( .A1(n20807), .A2(\xmem_data[82][4] ), .B1(n20806), .B2(
        \xmem_data[83][4] ), .ZN(n20812) );
  AOI22_X1 U24762 ( .A1(n20808), .A2(\xmem_data[84][4] ), .B1(n25450), .B2(
        \xmem_data[85][4] ), .ZN(n20811) );
  AOI22_X1 U24763 ( .A1(n20809), .A2(\xmem_data[86][4] ), .B1(n3358), .B2(
        \xmem_data[87][4] ), .ZN(n20810) );
  NAND4_X1 U24764 ( .A1(n20813), .A2(n20812), .A3(n20811), .A4(n20810), .ZN(
        n20824) );
  AOI22_X1 U24765 ( .A1(n20815), .A2(\xmem_data[64][4] ), .B1(n20814), .B2(
        \xmem_data[65][4] ), .ZN(n20822) );
  AOI22_X1 U24766 ( .A1(n28061), .A2(\xmem_data[66][4] ), .B1(n25581), .B2(
        \xmem_data[67][4] ), .ZN(n20821) );
  AOI22_X1 U24767 ( .A1(n20817), .A2(\xmem_data[68][4] ), .B1(n20949), .B2(
        \xmem_data[69][4] ), .ZN(n20820) );
  AOI22_X1 U24768 ( .A1(n20818), .A2(\xmem_data[70][4] ), .B1(n29247), .B2(
        \xmem_data[71][4] ), .ZN(n20819) );
  NAND4_X1 U24769 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20823) );
  AOI22_X1 U24770 ( .A1(n20826), .A2(\xmem_data[72][4] ), .B1(n25528), .B2(
        \xmem_data[73][4] ), .ZN(n20832) );
  AOI22_X1 U24771 ( .A1(n20827), .A2(\xmem_data[74][4] ), .B1(n25357), .B2(
        \xmem_data[75][4] ), .ZN(n20831) );
  AOI22_X1 U24772 ( .A1(n20828), .A2(\xmem_data[76][4] ), .B1(n25442), .B2(
        \xmem_data[77][4] ), .ZN(n20830) );
  AOI22_X1 U24773 ( .A1(n30906), .A2(\xmem_data[78][4] ), .B1(n3221), .B2(
        \xmem_data[79][4] ), .ZN(n20829) );
  NAND4_X1 U24774 ( .A1(n20832), .A2(n20831), .A3(n20830), .A4(n20829), .ZN(
        n20834) );
  XNOR2_X1 U24775 ( .A(n30156), .B(\fmem_data[28][3] ), .ZN(n31898) );
  OAI22_X1 U24776 ( .A1(n32644), .A2(n33855), .B1(n31898), .B2(n33853), .ZN(
        n26381) );
  XNOR2_X1 U24777 ( .A(n31221), .B(\fmem_data[2][3] ), .ZN(n32166) );
  XNOR2_X1 U24778 ( .A(n3359), .B(\fmem_data[2][3] ), .ZN(n32641) );
  OAI22_X1 U24779 ( .A1(n32166), .A2(n33796), .B1(n33797), .B2(n32641), .ZN(
        n26380) );
  INV_X1 U24780 ( .A(n35581), .ZN(n20840) );
  INV_X1 U24781 ( .A(n35730), .ZN(n20841) );
  AOI22_X1 U24782 ( .A1(n23730), .A2(\xmem_data[112][0] ), .B1(n28035), .B2(
        \xmem_data[113][0] ), .ZN(n20845) );
  AOI22_X1 U24783 ( .A1(n20986), .A2(\xmem_data[114][0] ), .B1(n12471), .B2(
        \xmem_data[115][0] ), .ZN(n20844) );
  AOI22_X1 U24784 ( .A1(n23732), .A2(\xmem_data[116][0] ), .B1(n23731), .B2(
        \xmem_data[117][0] ), .ZN(n20843) );
  AOI22_X1 U24785 ( .A1(n23734), .A2(\xmem_data[118][0] ), .B1(n3219), .B2(
        \xmem_data[119][0] ), .ZN(n20842) );
  NAND4_X1 U24786 ( .A1(n20845), .A2(n20844), .A3(n20843), .A4(n20842), .ZN(
        n20862) );
  AOI22_X1 U24787 ( .A1(n29308), .A2(\xmem_data[96][0] ), .B1(n24448), .B2(
        \xmem_data[97][0] ), .ZN(n20849) );
  AOI22_X1 U24788 ( .A1(n28298), .A2(\xmem_data[98][0] ), .B1(n23715), .B2(
        \xmem_data[99][0] ), .ZN(n20848) );
  AOI22_X1 U24789 ( .A1(n30892), .A2(\xmem_data[100][0] ), .B1(n23716), .B2(
        \xmem_data[101][0] ), .ZN(n20847) );
  AOI22_X1 U24790 ( .A1(n23717), .A2(\xmem_data[102][0] ), .B1(n23796), .B2(
        \xmem_data[103][0] ), .ZN(n20846) );
  NAND4_X1 U24791 ( .A1(n20849), .A2(n20848), .A3(n20847), .A4(n20846), .ZN(
        n20860) );
  AOI22_X1 U24792 ( .A1(n23740), .A2(\xmem_data[120][0] ), .B1(n23739), .B2(
        \xmem_data[121][0] ), .ZN(n20853) );
  AOI22_X1 U24793 ( .A1(n23741), .A2(\xmem_data[122][0] ), .B1(n13444), .B2(
        \xmem_data[123][0] ), .ZN(n20852) );
  AOI22_X1 U24794 ( .A1(n23742), .A2(\xmem_data[124][0] ), .B1(n25450), .B2(
        \xmem_data[125][0] ), .ZN(n20851) );
  AOI22_X1 U24795 ( .A1(n27447), .A2(\xmem_data[126][0] ), .B1(n3358), .B2(
        \xmem_data[127][0] ), .ZN(n20850) );
  NAND4_X1 U24796 ( .A1(n20853), .A2(n20852), .A3(n20851), .A4(n20850), .ZN(
        n20859) );
  AOI22_X1 U24797 ( .A1(n23722), .A2(\xmem_data[104][0] ), .B1(n29318), .B2(
        \xmem_data[105][0] ), .ZN(n20857) );
  AOI22_X1 U24798 ( .A1(n17002), .A2(\xmem_data[106][0] ), .B1(n17001), .B2(
        \xmem_data[107][0] ), .ZN(n20856) );
  AOI22_X1 U24799 ( .A1(n23724), .A2(\xmem_data[108][0] ), .B1(n23723), .B2(
        \xmem_data[109][0] ), .ZN(n20855) );
  AOI22_X1 U24800 ( .A1(n24685), .A2(\xmem_data[110][0] ), .B1(n23725), .B2(
        \xmem_data[111][0] ), .ZN(n20854) );
  NAND4_X1 U24801 ( .A1(n20857), .A2(n20856), .A3(n20855), .A4(n20854), .ZN(
        n20858) );
  OAI21_X1 U24802 ( .B1(n20862), .B2(n20861), .A(n23751), .ZN(n20886) );
  AOI22_X1 U24803 ( .A1(n23730), .A2(\xmem_data[80][0] ), .B1(n27435), .B2(
        \xmem_data[81][0] ), .ZN(n20867) );
  AOI22_X1 U24804 ( .A1(n25686), .A2(\xmem_data[82][0] ), .B1(n20578), .B2(
        \xmem_data[83][0] ), .ZN(n20866) );
  AOI22_X1 U24805 ( .A1(n23732), .A2(\xmem_data[84][0] ), .B1(n23731), .B2(
        \xmem_data[85][0] ), .ZN(n20865) );
  AND2_X1 U24806 ( .A1(n3220), .A2(\xmem_data[87][0] ), .ZN(n20863) );
  AOI21_X1 U24807 ( .B1(n23734), .B2(\xmem_data[86][0] ), .A(n20863), .ZN(
        n20864) );
  NAND4_X1 U24808 ( .A1(n20867), .A2(n20866), .A3(n20865), .A4(n20864), .ZN(
        n20884) );
  AOI22_X1 U24809 ( .A1(n30886), .A2(\xmem_data[64][0] ), .B1(n24212), .B2(
        \xmem_data[65][0] ), .ZN(n20871) );
  AOI22_X1 U24810 ( .A1(n28334), .A2(\xmem_data[66][0] ), .B1(n23715), .B2(
        \xmem_data[67][0] ), .ZN(n20870) );
  AOI22_X1 U24811 ( .A1(n28516), .A2(\xmem_data[68][0] ), .B1(n23716), .B2(
        \xmem_data[69][0] ), .ZN(n20869) );
  AOI22_X1 U24812 ( .A1(n23717), .A2(\xmem_data[70][0] ), .B1(n30544), .B2(
        \xmem_data[71][0] ), .ZN(n20868) );
  NAND4_X1 U24813 ( .A1(n20871), .A2(n20870), .A3(n20869), .A4(n20868), .ZN(
        n20882) );
  AOI22_X1 U24814 ( .A1(n23740), .A2(\xmem_data[88][0] ), .B1(n23739), .B2(
        \xmem_data[89][0] ), .ZN(n20875) );
  AOI22_X1 U24815 ( .A1(n23741), .A2(\xmem_data[90][0] ), .B1(n3256), .B2(
        \xmem_data[91][0] ), .ZN(n20874) );
  AOI22_X1 U24816 ( .A1(n23742), .A2(\xmem_data[92][0] ), .B1(n25492), .B2(
        \xmem_data[93][0] ), .ZN(n20873) );
  AOI22_X1 U24817 ( .A1(n27447), .A2(\xmem_data[94][0] ), .B1(n20546), .B2(
        \xmem_data[95][0] ), .ZN(n20872) );
  NAND4_X1 U24818 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20881) );
  AOI22_X1 U24819 ( .A1(n23722), .A2(\xmem_data[72][0] ), .B1(n25367), .B2(
        \xmem_data[73][0] ), .ZN(n20879) );
  AOI22_X1 U24820 ( .A1(n3325), .A2(\xmem_data[74][0] ), .B1(n17001), .B2(
        \xmem_data[75][0] ), .ZN(n20878) );
  AOI22_X1 U24821 ( .A1(n23724), .A2(\xmem_data[76][0] ), .B1(n23723), .B2(
        \xmem_data[77][0] ), .ZN(n20877) );
  AOI22_X1 U24822 ( .A1(n20734), .A2(\xmem_data[78][0] ), .B1(n23725), .B2(
        \xmem_data[79][0] ), .ZN(n20876) );
  NAND4_X1 U24823 ( .A1(n20879), .A2(n20878), .A3(n20877), .A4(n20876), .ZN(
        n20880) );
  OAI21_X1 U24824 ( .B1(n20884), .B2(n20883), .A(n23713), .ZN(n20885) );
  AND2_X1 U24825 ( .A1(n20886), .A2(n20885), .ZN(n33465) );
  AOI22_X1 U24826 ( .A1(n30901), .A2(\xmem_data[16][0] ), .B1(n25388), .B2(
        \xmem_data[17][0] ), .ZN(n20890) );
  AOI22_X1 U24827 ( .A1(n24526), .A2(\xmem_data[18][0] ), .B1(n25629), .B2(
        \xmem_data[19][0] ), .ZN(n20889) );
  AOI22_X1 U24828 ( .A1(n29661), .A2(\xmem_data[20][0] ), .B1(n22753), .B2(
        \xmem_data[21][0] ), .ZN(n20888) );
  AOI22_X1 U24829 ( .A1(n25354), .A2(\xmem_data[22][0] ), .B1(n3218), .B2(
        \xmem_data[23][0] ), .ZN(n20887) );
  NAND4_X1 U24830 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n20896) );
  AOI22_X1 U24831 ( .A1(n23792), .A2(\xmem_data[0][0] ), .B1(n27535), .B2(
        \xmem_data[1][0] ), .ZN(n20894) );
  AOI22_X1 U24832 ( .A1(n28298), .A2(\xmem_data[2][0] ), .B1(n23793), .B2(
        \xmem_data[3][0] ), .ZN(n20893) );
  AOI22_X1 U24833 ( .A1(n28091), .A2(\xmem_data[4][0] ), .B1(n3208), .B2(
        \xmem_data[5][0] ), .ZN(n20892) );
  AOI22_X1 U24834 ( .A1(n24708), .A2(\xmem_data[6][0] ), .B1(n23796), .B2(
        \xmem_data[7][0] ), .ZN(n20891) );
  NAND4_X1 U24835 ( .A1(n20894), .A2(n20893), .A3(n20892), .A4(n20891), .ZN(
        n20895) );
  AOI22_X1 U24836 ( .A1(n23802), .A2(\xmem_data[8][0] ), .B1(n23801), .B2(
        \xmem_data[9][0] ), .ZN(n20900) );
  AOI22_X1 U24837 ( .A1(n28428), .A2(\xmem_data[10][0] ), .B1(n25716), .B2(
        \xmem_data[11][0] ), .ZN(n20899) );
  AOI22_X1 U24838 ( .A1(n3269), .A2(\xmem_data[12][0] ), .B1(n23723), .B2(
        \xmem_data[13][0] ), .ZN(n20898) );
  AOI22_X1 U24839 ( .A1(n24685), .A2(\xmem_data[14][0] ), .B1(n22751), .B2(
        \xmem_data[15][0] ), .ZN(n20897) );
  NAND4_X1 U24840 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20901) );
  OR2_X1 U24841 ( .A1(n20901), .A2(n4002), .ZN(n20910) );
  AOI22_X1 U24842 ( .A1(n23812), .A2(\xmem_data[26][0] ), .B1(n23811), .B2(
        \xmem_data[27][0] ), .ZN(n20908) );
  AOI22_X1 U24843 ( .A1(n25731), .A2(\xmem_data[24][0] ), .B1(n20992), .B2(
        \xmem_data[25][0] ), .ZN(n20902) );
  INV_X1 U24844 ( .A(n20902), .ZN(n20906) );
  AND2_X1 U24845 ( .A1(n3282), .A2(\xmem_data[28][0] ), .ZN(n20905) );
  AOI22_X1 U24846 ( .A1(n23813), .A2(\xmem_data[30][0] ), .B1(n13475), .B2(
        \xmem_data[31][0] ), .ZN(n20903) );
  INV_X1 U24847 ( .A(n20903), .ZN(n20904) );
  NOR3_X1 U24848 ( .A1(n20906), .A2(n20905), .A3(n20904), .ZN(n20907) );
  NAND2_X1 U24849 ( .A1(n20908), .A2(n20907), .ZN(n20909) );
  OR2_X1 U24850 ( .A1(n20910), .A2(n20909), .ZN(n20911) );
  OAI21_X1 U24851 ( .B1(n20912), .B2(n20911), .A(n23822), .ZN(n20936) );
  AOI22_X1 U24852 ( .A1(n23753), .A2(\xmem_data[48][0] ), .B1(n28329), .B2(
        \xmem_data[49][0] ), .ZN(n20917) );
  AOI22_X1 U24853 ( .A1(n21061), .A2(\xmem_data[50][0] ), .B1(n30861), .B2(
        \xmem_data[51][0] ), .ZN(n20916) );
  AOI22_X1 U24854 ( .A1(n23754), .A2(\xmem_data[52][0] ), .B1(n28501), .B2(
        \xmem_data[53][0] ), .ZN(n20915) );
  AND2_X1 U24855 ( .A1(n3219), .A2(\xmem_data[55][0] ), .ZN(n20913) );
  AOI21_X1 U24856 ( .B1(n23756), .B2(\xmem_data[54][0] ), .A(n20913), .ZN(
        n20914) );
  NAND4_X1 U24857 ( .A1(n20917), .A2(n20916), .A3(n20915), .A4(n20914), .ZN(
        n20934) );
  AOI22_X1 U24858 ( .A1(n23777), .A2(\xmem_data[40][0] ), .B1(n23776), .B2(
        \xmem_data[41][0] ), .ZN(n20921) );
  AOI22_X1 U24859 ( .A1(n28385), .A2(\xmem_data[42][0] ), .B1(n23778), .B2(
        \xmem_data[43][0] ), .ZN(n20920) );
  AOI22_X1 U24860 ( .A1(n23780), .A2(\xmem_data[44][0] ), .B1(n23779), .B2(
        \xmem_data[45][0] ), .ZN(n20919) );
  AOI22_X1 U24861 ( .A1(n20782), .A2(\xmem_data[46][0] ), .B1(n23781), .B2(
        \xmem_data[47][0] ), .ZN(n20918) );
  NAND4_X1 U24862 ( .A1(n20921), .A2(n20920), .A3(n20919), .A4(n20918), .ZN(
        n20932) );
  AOI22_X1 U24863 ( .A1(n23770), .A2(\xmem_data[56][0] ), .B1(n23769), .B2(
        \xmem_data[57][0] ), .ZN(n20925) );
  AOI22_X1 U24864 ( .A1(n22666), .A2(\xmem_data[58][0] ), .B1(n22711), .B2(
        \xmem_data[59][0] ), .ZN(n20924) );
  AOI22_X1 U24865 ( .A1(n21074), .A2(\xmem_data[60][0] ), .B1(n28510), .B2(
        \xmem_data[61][0] ), .ZN(n20923) );
  AOI22_X1 U24866 ( .A1(n27447), .A2(\xmem_data[62][0] ), .B1(n27943), .B2(
        \xmem_data[63][0] ), .ZN(n20922) );
  NAND4_X1 U24867 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        n20931) );
  AOI22_X1 U24868 ( .A1(n23762), .A2(\xmem_data[32][0] ), .B1(n23761), .B2(
        \xmem_data[33][0] ), .ZN(n20929) );
  AOI22_X1 U24869 ( .A1(n23763), .A2(\xmem_data[34][0] ), .B1(n30513), .B2(
        \xmem_data[35][0] ), .ZN(n20928) );
  AOI22_X1 U24870 ( .A1(n20718), .A2(\xmem_data[36][0] ), .B1(n27516), .B2(
        \xmem_data[37][0] ), .ZN(n20927) );
  AOI22_X1 U24871 ( .A1(n23764), .A2(\xmem_data[38][0] ), .B1(n29048), .B2(
        \xmem_data[39][0] ), .ZN(n20926) );
  NAND4_X1 U24872 ( .A1(n20929), .A2(n20928), .A3(n20927), .A4(n20926), .ZN(
        n20930) );
  OR3_X1 U24873 ( .A1(n20932), .A2(n20931), .A3(n20930), .ZN(n20933) );
  OAI21_X1 U24874 ( .B1(n20934), .B2(n20933), .A(n23790), .ZN(n20935) );
  AND2_X1 U24875 ( .A1(n20936), .A2(n20935), .ZN(n33466) );
  INV_X1 U24876 ( .A(n35749), .ZN(n20937) );
  AOI22_X1 U24877 ( .A1(n20939), .A2(\xmem_data[32][1] ), .B1(n20938), .B2(
        \xmem_data[33][1] ), .ZN(n20947) );
  AOI22_X1 U24878 ( .A1(n17020), .A2(\xmem_data[34][1] ), .B1(n20940), .B2(
        \xmem_data[35][1] ), .ZN(n20946) );
  AOI22_X1 U24879 ( .A1(n20942), .A2(\xmem_data[36][1] ), .B1(n20941), .B2(
        \xmem_data[37][1] ), .ZN(n20945) );
  AOI22_X1 U24880 ( .A1(n3206), .A2(\xmem_data[38][1] ), .B1(n20943), .B2(
        \xmem_data[39][1] ), .ZN(n20944) );
  NAND4_X1 U24881 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20948) );
  AOI22_X1 U24882 ( .A1(n20950), .A2(\xmem_data[40][1] ), .B1(n20949), .B2(
        \xmem_data[41][1] ), .ZN(n20957) );
  AOI22_X1 U24883 ( .A1(n22719), .A2(\xmem_data[42][1] ), .B1(n27463), .B2(
        \xmem_data[43][1] ), .ZN(n20956) );
  AOI22_X1 U24884 ( .A1(n20952), .A2(\xmem_data[44][1] ), .B1(n20951), .B2(
        \xmem_data[45][1] ), .ZN(n20955) );
  AOI22_X1 U24885 ( .A1(n20953), .A2(\xmem_data[46][1] ), .B1(n28317), .B2(
        \xmem_data[47][1] ), .ZN(n20954) );
  NAND4_X1 U24886 ( .A1(n20957), .A2(n20956), .A3(n20955), .A4(n20954), .ZN(
        n20976) );
  AOI22_X1 U24887 ( .A1(n28051), .A2(\xmem_data[60][1] ), .B1(n20958), .B2(
        \xmem_data[61][1] ), .ZN(n20968) );
  AOI22_X1 U24888 ( .A1(n20959), .A2(\xmem_data[62][1] ), .B1(n28090), .B2(
        \xmem_data[63][1] ), .ZN(n20960) );
  INV_X1 U24889 ( .A(n20960), .ZN(n20966) );
  AOI22_X1 U24890 ( .A1(n20961), .A2(\xmem_data[58][1] ), .B1(n20982), .B2(
        \xmem_data[59][1] ), .ZN(n20964) );
  NAND2_X1 U24891 ( .A1(n20962), .A2(\xmem_data[56][1] ), .ZN(n20963) );
  NAND2_X1 U24892 ( .A1(n20964), .A2(n20963), .ZN(n20965) );
  NOR2_X1 U24893 ( .A1(n20966), .A2(n20965), .ZN(n20967) );
  NAND2_X1 U24894 ( .A1(n20968), .A2(n20967), .ZN(n20975) );
  AOI22_X1 U24895 ( .A1(n3334), .A2(\xmem_data[48][1] ), .B1(n29253), .B2(
        \xmem_data[49][1] ), .ZN(n20973) );
  AOI22_X1 U24896 ( .A1(n27902), .A2(\xmem_data[50][1] ), .B1(n3217), .B2(
        \xmem_data[51][1] ), .ZN(n20972) );
  AOI22_X1 U24897 ( .A1(n24533), .A2(\xmem_data[52][1] ), .B1(n22710), .B2(
        \xmem_data[53][1] ), .ZN(n20971) );
  AOI22_X1 U24898 ( .A1(n20969), .A2(\xmem_data[54][1] ), .B1(n14890), .B2(
        \xmem_data[55][1] ), .ZN(n20970) );
  NAND4_X1 U24899 ( .A1(n20973), .A2(n20972), .A3(n20971), .A4(n20970), .ZN(
        n20974) );
  OR4_X1 U24900 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n20979) );
  NAND2_X1 U24901 ( .A1(n20979), .A2(n20311), .ZN(n21025) );
  INV_X1 U24902 ( .A(n21025), .ZN(n20981) );
  OR2_X1 U24903 ( .A1(n20981), .A2(n20980), .ZN(n21027) );
  NAND2_X1 U24904 ( .A1(n20982), .A2(\xmem_data[27][1] ), .ZN(n21004) );
  AOI22_X1 U24905 ( .A1(n20984), .A2(\xmem_data[8][1] ), .B1(n20983), .B2(
        \xmem_data[9][1] ), .ZN(n20990) );
  AOI22_X1 U24906 ( .A1(n29151), .A2(\xmem_data[10][1] ), .B1(n31256), .B2(
        \xmem_data[11][1] ), .ZN(n20989) );
  AOI22_X1 U24907 ( .A1(n20985), .A2(\xmem_data[12][1] ), .B1(n29248), .B2(
        \xmem_data[13][1] ), .ZN(n20988) );
  AOI22_X1 U24908 ( .A1(n20986), .A2(\xmem_data[14][1] ), .B1(n29118), .B2(
        \xmem_data[15][1] ), .ZN(n20987) );
  NAND4_X1 U24909 ( .A1(n20990), .A2(n20989), .A3(n20988), .A4(n20987), .ZN(
        n21002) );
  AOI22_X1 U24910 ( .A1(n3332), .A2(\xmem_data[16][1] ), .B1(n20711), .B2(
        \xmem_data[17][1] ), .ZN(n20998) );
  AOI22_X1 U24911 ( .A1(n20991), .A2(\xmem_data[18][1] ), .B1(n3220), .B2(
        \xmem_data[19][1] ), .ZN(n20997) );
  AOI22_X1 U24912 ( .A1(n30278), .A2(\xmem_data[20][1] ), .B1(n20992), .B2(
        \xmem_data[21][1] ), .ZN(n20996) );
  AOI22_X1 U24913 ( .A1(n20994), .A2(\xmem_data[22][1] ), .B1(n20993), .B2(
        \xmem_data[23][1] ), .ZN(n20995) );
  NAND4_X1 U24914 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n21001) );
  AND2_X1 U24915 ( .A1(n30663), .A2(\xmem_data[28][1] ), .ZN(n21000) );
  AND2_X1 U24916 ( .A1(n24160), .A2(\xmem_data[31][1] ), .ZN(n20999) );
  NOR4_X1 U24917 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  AND2_X1 U24918 ( .A1(n21004), .A2(n21003), .ZN(n21024) );
  AOI22_X1 U24919 ( .A1(n21005), .A2(\xmem_data[0][1] ), .B1(n3208), .B2(
        \xmem_data[1][1] ), .ZN(n21014) );
  AOI22_X1 U24920 ( .A1(n21007), .A2(\xmem_data[2][1] ), .B1(n21006), .B2(
        \xmem_data[3][1] ), .ZN(n21013) );
  AOI22_X1 U24921 ( .A1(n21008), .A2(\xmem_data[4][1] ), .B1(n30515), .B2(
        \xmem_data[5][1] ), .ZN(n21012) );
  AOI22_X1 U24922 ( .A1(n21010), .A2(\xmem_data[6][1] ), .B1(n25581), .B2(
        \xmem_data[7][1] ), .ZN(n21011) );
  NAND4_X1 U24923 ( .A1(n21014), .A2(n21013), .A3(n21012), .A4(n21011), .ZN(
        n21021) );
  AOI22_X1 U24924 ( .A1(n20495), .A2(\xmem_data[30][1] ), .B1(n21015), .B2(
        \xmem_data[29][1] ), .ZN(n21019) );
  AND2_X1 U24925 ( .A1(n25670), .A2(\xmem_data[26][1] ), .ZN(n21017) );
  AND2_X1 U24926 ( .A1(n30295), .A2(\xmem_data[24][1] ), .ZN(n21016) );
  NOR2_X1 U24927 ( .A1(n21017), .A2(n21016), .ZN(n21018) );
  NAND2_X1 U24928 ( .A1(n21019), .A2(n21018), .ZN(n21020) );
  NOR2_X1 U24929 ( .A1(n21021), .A2(n21020), .ZN(n21023) );
  NAND2_X1 U24930 ( .A1(n29103), .A2(\xmem_data[25][1] ), .ZN(n21022) );
  NAND4_X1 U24931 ( .A1(n21025), .A2(n21024), .A3(n21023), .A4(n21022), .ZN(
        n21026) );
  NAND2_X1 U24932 ( .A1(n21027), .A2(n21026), .ZN(n21090) );
  AOI22_X1 U24933 ( .A1(n21048), .A2(\xmem_data[96][1] ), .B1(n27864), .B2(
        \xmem_data[97][1] ), .ZN(n21031) );
  AOI22_X1 U24934 ( .A1(n25573), .A2(\xmem_data[98][1] ), .B1(n25715), .B2(
        \xmem_data[99][1] ), .ZN(n21030) );
  AOI22_X1 U24935 ( .A1(n21050), .A2(\xmem_data[100][1] ), .B1(n21049), .B2(
        \xmem_data[101][1] ), .ZN(n21029) );
  AOI22_X1 U24936 ( .A1(n3178), .A2(\xmem_data[102][1] ), .B1(n25581), .B2(
        \xmem_data[103][1] ), .ZN(n21028) );
  NAND4_X1 U24937 ( .A1(n21031), .A2(n21030), .A3(n21029), .A4(n21028), .ZN(
        n21047) );
  AOI22_X1 U24938 ( .A1(n21056), .A2(\xmem_data[104][1] ), .B1(n20507), .B2(
        \xmem_data[105][1] ), .ZN(n21035) );
  AOI22_X1 U24939 ( .A1(n21058), .A2(\xmem_data[106][1] ), .B1(n21057), .B2(
        \xmem_data[107][1] ), .ZN(n21034) );
  AOI22_X1 U24940 ( .A1(n21060), .A2(\xmem_data[108][1] ), .B1(n21059), .B2(
        \xmem_data[109][1] ), .ZN(n21033) );
  AOI22_X1 U24941 ( .A1(n21061), .A2(\xmem_data[110][1] ), .B1(n24525), .B2(
        \xmem_data[111][1] ), .ZN(n21032) );
  NAND4_X1 U24942 ( .A1(n21035), .A2(n21034), .A3(n21033), .A4(n21032), .ZN(
        n21046) );
  AOI22_X1 U24943 ( .A1(n3424), .A2(\xmem_data[112][1] ), .B1(n3247), .B2(
        \xmem_data[113][1] ), .ZN(n21039) );
  AOI22_X1 U24944 ( .A1(n21066), .A2(\xmem_data[114][1] ), .B1(n3221), .B2(
        \xmem_data[115][1] ), .ZN(n21038) );
  AOI22_X1 U24945 ( .A1(n21067), .A2(\xmem_data[116][1] ), .B1(n20723), .B2(
        \xmem_data[117][1] ), .ZN(n21037) );
  AOI22_X1 U24946 ( .A1(n21069), .A2(\xmem_data[118][1] ), .B1(n21068), .B2(
        \xmem_data[119][1] ), .ZN(n21036) );
  NAND4_X1 U24947 ( .A1(n21039), .A2(n21038), .A3(n21037), .A4(n21036), .ZN(
        n21045) );
  AOI22_X1 U24948 ( .A1(n21074), .A2(\xmem_data[120][1] ), .B1(n30877), .B2(
        \xmem_data[121][1] ), .ZN(n21043) );
  AOI22_X1 U24949 ( .A1(n25670), .A2(\xmem_data[122][1] ), .B1(n28415), .B2(
        \xmem_data[123][1] ), .ZN(n21042) );
  AOI22_X1 U24950 ( .A1(n30083), .A2(\xmem_data[124][1] ), .B1(n21075), .B2(
        \xmem_data[125][1] ), .ZN(n21041) );
  AOI22_X1 U24951 ( .A1(n17041), .A2(\xmem_data[126][1] ), .B1(n21076), .B2(
        \xmem_data[127][1] ), .ZN(n21040) );
  NAND4_X1 U24952 ( .A1(n21043), .A2(n21042), .A3(n21041), .A4(n21040), .ZN(
        n21044) );
  OR4_X1 U24953 ( .A1(n21047), .A2(n21046), .A3(n21045), .A4(n21044), .ZN(
        n21087) );
  AOI22_X1 U24954 ( .A1(n21048), .A2(\xmem_data[64][1] ), .B1(n20938), .B2(
        \xmem_data[65][1] ), .ZN(n21055) );
  AOI22_X1 U24955 ( .A1(n13149), .A2(\xmem_data[66][1] ), .B1(n30544), .B2(
        \xmem_data[67][1] ), .ZN(n21054) );
  AOI22_X1 U24956 ( .A1(n21050), .A2(\xmem_data[68][1] ), .B1(n21049), .B2(
        \xmem_data[69][1] ), .ZN(n21053) );
  AOI22_X1 U24957 ( .A1(n3325), .A2(\xmem_data[70][1] ), .B1(n21051), .B2(
        \xmem_data[71][1] ), .ZN(n21052) );
  NAND4_X1 U24958 ( .A1(n21055), .A2(n21054), .A3(n21053), .A4(n21052), .ZN(
        n21084) );
  AOI22_X1 U24959 ( .A1(n21056), .A2(\xmem_data[72][1] ), .B1(n24622), .B2(
        \xmem_data[73][1] ), .ZN(n21065) );
  AOI22_X1 U24960 ( .A1(n21058), .A2(\xmem_data[74][1] ), .B1(n21057), .B2(
        \xmem_data[75][1] ), .ZN(n21064) );
  AOI22_X1 U24961 ( .A1(n21060), .A2(\xmem_data[76][1] ), .B1(n21059), .B2(
        \xmem_data[77][1] ), .ZN(n21063) );
  AOI22_X1 U24962 ( .A1(n21061), .A2(\xmem_data[78][1] ), .B1(n28317), .B2(
        \xmem_data[79][1] ), .ZN(n21062) );
  NAND4_X1 U24963 ( .A1(n21065), .A2(n21064), .A3(n21063), .A4(n21062), .ZN(
        n21083) );
  AOI22_X1 U24964 ( .A1(n3384), .A2(\xmem_data[80][1] ), .B1(n31347), .B2(
        \xmem_data[81][1] ), .ZN(n21073) );
  AOI22_X1 U24965 ( .A1(n21066), .A2(\xmem_data[82][1] ), .B1(n3219), .B2(
        \xmem_data[83][1] ), .ZN(n21072) );
  AOI22_X1 U24966 ( .A1(n21067), .A2(\xmem_data[84][1] ), .B1(n29028), .B2(
        \xmem_data[85][1] ), .ZN(n21071) );
  AOI22_X1 U24967 ( .A1(n21069), .A2(\xmem_data[86][1] ), .B1(n21068), .B2(
        \xmem_data[87][1] ), .ZN(n21070) );
  NAND4_X1 U24968 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21082) );
  AOI22_X1 U24969 ( .A1(n21074), .A2(\xmem_data[88][1] ), .B1(n24657), .B2(
        \xmem_data[89][1] ), .ZN(n21080) );
  AOI22_X1 U24970 ( .A1(n27447), .A2(\xmem_data[90][1] ), .B1(n3358), .B2(
        \xmem_data[91][1] ), .ZN(n21079) );
  AOI22_X1 U24971 ( .A1(n20799), .A2(\xmem_data[92][1] ), .B1(n21075), .B2(
        \xmem_data[93][1] ), .ZN(n21078) );
  AOI22_X1 U24972 ( .A1(n3176), .A2(\xmem_data[94][1] ), .B1(n21076), .B2(
        \xmem_data[95][1] ), .ZN(n21077) );
  NAND4_X1 U24973 ( .A1(n21080), .A2(n21079), .A3(n21078), .A4(n21077), .ZN(
        n21081) );
  OR4_X1 U24974 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n21081), .ZN(
        n21085) );
  AOI22_X1 U24975 ( .A1(n21088), .A2(n21087), .B1(n21086), .B2(n21085), .ZN(
        n21089) );
  NOR2_X1 U24976 ( .A1(n26376), .A2(n26375), .ZN(n21092) );
  OAI21_X1 U24977 ( .B1(n21093), .B2(n21092), .A(n21091), .ZN(n23182) );
  AOI22_X1 U24978 ( .A1(n3220), .A2(\xmem_data[96][4] ), .B1(n29256), .B2(
        \xmem_data[97][4] ), .ZN(n21097) );
  AOI22_X1 U24979 ( .A1(n31367), .A2(\xmem_data[98][4] ), .B1(n28083), .B2(
        \xmem_data[99][4] ), .ZN(n21096) );
  AOI22_X1 U24980 ( .A1(n30882), .A2(\xmem_data[100][4] ), .B1(n23742), .B2(
        \xmem_data[101][4] ), .ZN(n21095) );
  AOI22_X1 U24981 ( .A1(n28007), .A2(\xmem_data[102][4] ), .B1(n28374), .B2(
        \xmem_data[103][4] ), .ZN(n21094) );
  NAND4_X1 U24982 ( .A1(n21097), .A2(n21096), .A3(n21095), .A4(n21094), .ZN(
        n21114) );
  AOI22_X1 U24983 ( .A1(n24158), .A2(\xmem_data[104][4] ), .B1(n24157), .B2(
        \xmem_data[105][4] ), .ZN(n21101) );
  AOI22_X1 U24984 ( .A1(n24159), .A2(\xmem_data[106][4] ), .B1(n13436), .B2(
        \xmem_data[107][4] ), .ZN(n21100) );
  AOI22_X1 U24985 ( .A1(n24160), .A2(\xmem_data[108][4] ), .B1(n27755), .B2(
        \xmem_data[109][4] ), .ZN(n21099) );
  AOI22_X1 U24986 ( .A1(n24134), .A2(\xmem_data[110][4] ), .B1(n23717), .B2(
        \xmem_data[111][4] ), .ZN(n21098) );
  NAND4_X1 U24987 ( .A1(n21101), .A2(n21100), .A3(n21099), .A4(n21098), .ZN(
        n21113) );
  AOI22_X1 U24988 ( .A1(n22718), .A2(\xmem_data[112][4] ), .B1(n29439), .B2(
        \xmem_data[113][4] ), .ZN(n21105) );
  AOI22_X1 U24989 ( .A1(n24165), .A2(\xmem_data[114][4] ), .B1(n24548), .B2(
        \xmem_data[115][4] ), .ZN(n21104) );
  AOI22_X1 U24990 ( .A1(n20816), .A2(\xmem_data[116][4] ), .B1(n28226), .B2(
        \xmem_data[117][4] ), .ZN(n21103) );
  AOI22_X1 U24991 ( .A1(n24167), .A2(\xmem_data[118][4] ), .B1(n24166), .B2(
        \xmem_data[119][4] ), .ZN(n21102) );
  NAND4_X1 U24992 ( .A1(n21105), .A2(n21104), .A3(n21103), .A4(n21102), .ZN(
        n21112) );
  AOI22_X1 U24993 ( .A1(n27463), .A2(\xmem_data[120][4] ), .B1(n20567), .B2(
        \xmem_data[121][4] ), .ZN(n21110) );
  AOI22_X1 U24994 ( .A1(n28329), .A2(\xmem_data[122][4] ), .B1(n24688), .B2(
        \xmem_data[123][4] ), .ZN(n21109) );
  AOI22_X1 U24995 ( .A1(n31262), .A2(\xmem_data[124][4] ), .B1(n23732), .B2(
        \xmem_data[125][4] ), .ZN(n21108) );
  AND2_X1 U24996 ( .A1(n24172), .A2(\xmem_data[126][4] ), .ZN(n21106) );
  AOI21_X1 U24997 ( .B1(n23756), .B2(\xmem_data[127][4] ), .A(n21106), .ZN(
        n21107) );
  NAND4_X1 U24998 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21111) );
  OR4_X1 U24999 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21137) );
  AOI22_X1 U25000 ( .A1(n11008), .A2(\xmem_data[88][4] ), .B1(n29327), .B2(
        \xmem_data[89][4] ), .ZN(n21119) );
  AOI22_X1 U25001 ( .A1(n20951), .A2(\xmem_data[90][4] ), .B1(n25358), .B2(
        \xmem_data[91][4] ), .ZN(n21118) );
  AOI22_X1 U25002 ( .A1(n24625), .A2(\xmem_data[92][4] ), .B1(n3334), .B2(
        \xmem_data[93][4] ), .ZN(n21117) );
  AND2_X1 U25003 ( .A1(n20711), .A2(\xmem_data[94][4] ), .ZN(n21115) );
  AOI21_X1 U25004 ( .B1(n24694), .B2(\xmem_data[95][4] ), .A(n21115), .ZN(
        n21116) );
  NAND4_X1 U25005 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21135) );
  AOI22_X1 U25006 ( .A1(n3358), .A2(\xmem_data[72][4] ), .B1(n29308), .B2(
        \xmem_data[73][4] ), .ZN(n21123) );
  AOI22_X1 U25007 ( .A1(n24212), .A2(\xmem_data[74][4] ), .B1(n28298), .B2(
        \xmem_data[75][4] ), .ZN(n21122) );
  AOI22_X1 U25008 ( .A1(n24597), .A2(\xmem_data[76][4] ), .B1(n30892), .B2(
        \xmem_data[77][4] ), .ZN(n21121) );
  AOI22_X1 U25009 ( .A1(n29279), .A2(\xmem_data[78][4] ), .B1(n24214), .B2(
        \xmem_data[79][4] ), .ZN(n21120) );
  NAND4_X1 U25010 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21134) );
  AOI22_X1 U25011 ( .A1(n24219), .A2(\xmem_data[80][4] ), .B1(n16990), .B2(
        \xmem_data[81][4] ), .ZN(n21127) );
  AOI22_X1 U25012 ( .A1(n24221), .A2(\xmem_data[82][4] ), .B1(n25632), .B2(
        \xmem_data[83][4] ), .ZN(n21126) );
  AOI22_X1 U25013 ( .A1(n24222), .A2(\xmem_data[84][4] ), .B1(n20732), .B2(
        \xmem_data[85][4] ), .ZN(n21125) );
  AOI22_X1 U25014 ( .A1(n24223), .A2(\xmem_data[86][4] ), .B1(n29325), .B2(
        \xmem_data[87][4] ), .ZN(n21124) );
  NAND4_X1 U25015 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21133) );
  AOI22_X1 U25016 ( .A1(n3220), .A2(\xmem_data[64][4] ), .B1(n28367), .B2(
        \xmem_data[65][4] ), .ZN(n21131) );
  AOI22_X1 U25017 ( .A1(n24207), .A2(\xmem_data[66][4] ), .B1(n22709), .B2(
        \xmem_data[67][4] ), .ZN(n21130) );
  AOI22_X1 U25018 ( .A1(n28342), .A2(\xmem_data[68][4] ), .B1(n23742), .B2(
        \xmem_data[69][4] ), .ZN(n21129) );
  AOI22_X1 U25019 ( .A1(n28510), .A2(\xmem_data[70][4] ), .B1(n25604), .B2(
        \xmem_data[71][4] ), .ZN(n21128) );
  NAND4_X1 U25020 ( .A1(n21131), .A2(n21130), .A3(n21129), .A4(n21128), .ZN(
        n21132) );
  OR4_X1 U25021 ( .A1(n21135), .A2(n21134), .A3(n21133), .A4(n21132), .ZN(
        n21136) );
  AOI22_X1 U25022 ( .A1(n21137), .A2(n24205), .B1(n24204), .B2(n21136), .ZN(
        n21189) );
  AOI22_X1 U25023 ( .A1(n3220), .A2(\xmem_data[32][4] ), .B1(n20805), .B2(
        \xmem_data[33][4] ), .ZN(n21141) );
  AOI22_X1 U25024 ( .A1(n24207), .A2(\xmem_data[34][4] ), .B1(n24565), .B2(
        \xmem_data[35][4] ), .ZN(n21140) );
  AOI22_X1 U25025 ( .A1(n25415), .A2(\xmem_data[36][4] ), .B1(n25417), .B2(
        \xmem_data[37][4] ), .ZN(n21139) );
  AOI22_X1 U25026 ( .A1(n24657), .A2(\xmem_data[38][4] ), .B1(n25604), .B2(
        \xmem_data[39][4] ), .ZN(n21138) );
  NAND4_X1 U25027 ( .A1(n21141), .A2(n21140), .A3(n21139), .A4(n21138), .ZN(
        n21157) );
  AOI22_X1 U25028 ( .A1(n22701), .A2(\xmem_data[40][4] ), .B1(n31353), .B2(
        \xmem_data[41][4] ), .ZN(n21145) );
  AOI22_X1 U25029 ( .A1(n24212), .A2(\xmem_data[42][4] ), .B1(n16986), .B2(
        \xmem_data[43][4] ), .ZN(n21144) );
  AOI22_X1 U25030 ( .A1(n29271), .A2(\xmem_data[44][4] ), .B1(n20776), .B2(
        \xmem_data[45][4] ), .ZN(n21143) );
  AOI22_X1 U25031 ( .A1(n23716), .A2(\xmem_data[46][4] ), .B1(n24214), .B2(
        \xmem_data[47][4] ), .ZN(n21142) );
  NAND4_X1 U25032 ( .A1(n21145), .A2(n21144), .A3(n21143), .A4(n21142), .ZN(
        n21156) );
  AOI22_X1 U25033 ( .A1(n24219), .A2(\xmem_data[48][4] ), .B1(n30872), .B2(
        \xmem_data[49][4] ), .ZN(n21149) );
  AOI22_X1 U25034 ( .A1(n24221), .A2(\xmem_data[50][4] ), .B1(n20731), .B2(
        \xmem_data[51][4] ), .ZN(n21148) );
  AOI22_X1 U25035 ( .A1(n24222), .A2(\xmem_data[52][4] ), .B1(n3338), .B2(
        \xmem_data[53][4] ), .ZN(n21147) );
  AOI22_X1 U25036 ( .A1(n24223), .A2(\xmem_data[54][4] ), .B1(n29325), .B2(
        \xmem_data[55][4] ), .ZN(n21146) );
  NAND4_X1 U25037 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21155) );
  AOI22_X1 U25038 ( .A1(n27526), .A2(\xmem_data[56][4] ), .B1(n29298), .B2(
        \xmem_data[57][4] ), .ZN(n21153) );
  AOI22_X1 U25039 ( .A1(n28035), .A2(\xmem_data[58][4] ), .B1(n24607), .B2(
        \xmem_data[59][4] ), .ZN(n21152) );
  AOI22_X1 U25040 ( .A1(n30908), .A2(\xmem_data[60][4] ), .B1(n3383), .B2(
        \xmem_data[61][4] ), .ZN(n21151) );
  AOI22_X1 U25041 ( .A1(n25485), .A2(\xmem_data[62][4] ), .B1(n24562), .B2(
        \xmem_data[63][4] ), .ZN(n21150) );
  NAND4_X1 U25042 ( .A1(n21153), .A2(n21152), .A3(n21151), .A4(n21150), .ZN(
        n21154) );
  OR4_X1 U25043 ( .A1(n21157), .A2(n21156), .A3(n21155), .A4(n21154), .ZN(
        n21187) );
  AOI22_X1 U25044 ( .A1(n25723), .A2(\xmem_data[24][4] ), .B1(n30754), .B2(
        \xmem_data[25][4] ), .ZN(n21162) );
  AOI22_X1 U25045 ( .A1(n24122), .A2(\xmem_data[26][4] ), .B1(n25358), .B2(
        \xmem_data[27][4] ), .ZN(n21161) );
  AOI22_X1 U25046 ( .A1(n29328), .A2(\xmem_data[28][4] ), .B1(n28039), .B2(
        \xmem_data[29][4] ), .ZN(n21160) );
  AND2_X1 U25047 ( .A1(n30589), .A2(\xmem_data[30][4] ), .ZN(n21158) );
  AOI21_X1 U25048 ( .B1(n20518), .B2(\xmem_data[31][4] ), .A(n21158), .ZN(
        n21159) );
  NAND4_X1 U25049 ( .A1(n21162), .A2(n21161), .A3(n21160), .A4(n21159), .ZN(
        n21182) );
  AOI22_X1 U25050 ( .A1(n29048), .A2(\xmem_data[16][4] ), .B1(n24115), .B2(
        \xmem_data[17][4] ), .ZN(n21166) );
  AOI22_X1 U25051 ( .A1(n24116), .A2(\xmem_data[18][4] ), .B1(n3326), .B2(
        \xmem_data[19][4] ), .ZN(n21165) );
  AOI22_X1 U25052 ( .A1(n24117), .A2(\xmem_data[20][4] ), .B1(n30686), .B2(
        \xmem_data[21][4] ), .ZN(n21164) );
  AOI22_X1 U25053 ( .A1(n28983), .A2(\xmem_data[22][4] ), .B1(n24572), .B2(
        \xmem_data[23][4] ), .ZN(n21163) );
  NAND4_X1 U25054 ( .A1(n21166), .A2(n21165), .A3(n21164), .A4(n21163), .ZN(
        n21181) );
  AOI22_X1 U25055 ( .A1(n24130), .A2(\xmem_data[8][4] ), .B1(n23792), .B2(
        \xmem_data[9][4] ), .ZN(n21170) );
  AOI22_X1 U25056 ( .A1(n24132), .A2(\xmem_data[10][4] ), .B1(n28980), .B2(
        \xmem_data[11][4] ), .ZN(n21169) );
  AOI22_X1 U25057 ( .A1(n22741), .A2(\xmem_data[12][4] ), .B1(n29605), .B2(
        \xmem_data[13][4] ), .ZN(n21168) );
  AOI22_X1 U25058 ( .A1(n24134), .A2(\xmem_data[14][4] ), .B1(n24133), .B2(
        \xmem_data[15][4] ), .ZN(n21167) );
  NAND4_X1 U25059 ( .A1(n21170), .A2(n21169), .A3(n21168), .A4(n21167), .ZN(
        n21180) );
  AOI22_X1 U25060 ( .A1(n24140), .A2(\xmem_data[4][4] ), .B1(n3140), .B2(
        \xmem_data[5][4] ), .ZN(n21178) );
  NAND2_X1 U25061 ( .A1(n3217), .A2(\xmem_data[0][4] ), .ZN(n21172) );
  NAND2_X1 U25062 ( .A1(n24139), .A2(\xmem_data[1][4] ), .ZN(n21171) );
  NAND2_X1 U25063 ( .A1(n21172), .A2(n21171), .ZN(n21176) );
  AOI22_X1 U25064 ( .A1(n14989), .A2(\xmem_data[2][4] ), .B1(n24141), .B2(
        \xmem_data[3][4] ), .ZN(n21173) );
  INV_X1 U25065 ( .A(n21173), .ZN(n21175) );
  AND2_X1 U25066 ( .A1(n23813), .A2(\xmem_data[7][4] ), .ZN(n21174) );
  NOR3_X1 U25067 ( .A1(n21176), .A2(n21175), .A3(n21174), .ZN(n21177) );
  NAND2_X1 U25068 ( .A1(n21178), .A2(n21177), .ZN(n21179) );
  NOR4_X1 U25069 ( .A1(n21182), .A2(n21181), .A3(n21180), .A4(n21179), .ZN(
        n21185) );
  NOR2_X1 U25070 ( .A1(n24151), .A2(n39032), .ZN(n21183) );
  NAND2_X1 U25071 ( .A1(n13474), .A2(n21183), .ZN(n21184) );
  OAI21_X1 U25072 ( .B1(n21185), .B2(n24151), .A(n21184), .ZN(n21186) );
  AOI21_X1 U25073 ( .B1(n21187), .B2(n24236), .A(n21186), .ZN(n21188) );
  XNOR2_X1 U25074 ( .A(n28539), .B(\fmem_data[13][3] ), .ZN(n30847) );
  XNOR2_X1 U25075 ( .A(n31668), .B(\fmem_data[13][3] ), .ZN(n31965) );
  OAI22_X1 U25076 ( .A1(n30847), .A2(n33570), .B1(n33568), .B2(n31965), .ZN(
        n34005) );
  AOI22_X1 U25077 ( .A1(n24693), .A2(\xmem_data[72][0] ), .B1(n28501), .B2(
        \xmem_data[73][0] ), .ZN(n21195) );
  AND2_X1 U25078 ( .A1(n3217), .A2(\xmem_data[75][0] ), .ZN(n21191) );
  AOI21_X1 U25079 ( .B1(n24694), .B2(\xmem_data[74][0] ), .A(n21191), .ZN(
        n21194) );
  AOI22_X1 U25080 ( .A1(n24696), .A2(\xmem_data[76][0] ), .B1(n24695), .B2(
        \xmem_data[77][0] ), .ZN(n21193) );
  AOI22_X1 U25081 ( .A1(n24697), .A2(\xmem_data[78][0] ), .B1(n31275), .B2(
        \xmem_data[79][0] ), .ZN(n21192) );
  NAND4_X1 U25082 ( .A1(n21195), .A2(n21194), .A3(n21193), .A4(n21192), .ZN(
        n21211) );
  AOI22_X1 U25083 ( .A1(n20984), .A2(\xmem_data[64][0] ), .B1(n24622), .B2(
        \xmem_data[65][0] ), .ZN(n21199) );
  AOI22_X1 U25084 ( .A1(n24685), .A2(\xmem_data[66][0] ), .B1(n27526), .B2(
        \xmem_data[67][0] ), .ZN(n21198) );
  AOI22_X1 U25085 ( .A1(n24687), .A2(\xmem_data[68][0] ), .B1(n24686), .B2(
        \xmem_data[69][0] ), .ZN(n21197) );
  AOI22_X1 U25086 ( .A1(n24688), .A2(\xmem_data[70][0] ), .B1(n29328), .B2(
        \xmem_data[71][0] ), .ZN(n21196) );
  NAND4_X1 U25087 ( .A1(n21199), .A2(n21198), .A3(n21197), .A4(n21196), .ZN(
        n21210) );
  AOI22_X1 U25088 ( .A1(n24702), .A2(\xmem_data[80][0] ), .B1(n29103), .B2(
        \xmem_data[81][0] ), .ZN(n21203) );
  AOI22_X1 U25089 ( .A1(n22712), .A2(\xmem_data[82][0] ), .B1(n24158), .B2(
        \xmem_data[83][0] ), .ZN(n21202) );
  AOI22_X1 U25090 ( .A1(n28309), .A2(\xmem_data[84][0] ), .B1(n13168), .B2(
        \xmem_data[85][0] ), .ZN(n21201) );
  AOI22_X1 U25091 ( .A1(n25459), .A2(\xmem_data[86][0] ), .B1(n20544), .B2(
        \xmem_data[87][0] ), .ZN(n21200) );
  NAND4_X1 U25092 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21209) );
  AOI22_X1 U25093 ( .A1(n27945), .A2(\xmem_data[88][0] ), .B1(n27864), .B2(
        \xmem_data[89][0] ), .ZN(n21207) );
  AOI22_X1 U25094 ( .A1(n24708), .A2(\xmem_data[90][0] ), .B1(n24707), .B2(
        \xmem_data[91][0] ), .ZN(n21206) );
  AOI22_X1 U25095 ( .A1(n24710), .A2(\xmem_data[92][0] ), .B1(n24709), .B2(
        \xmem_data[93][0] ), .ZN(n21205) );
  AOI22_X1 U25096 ( .A1(n28061), .A2(\xmem_data[94][0] ), .B1(n20551), .B2(
        \xmem_data[95][0] ), .ZN(n21204) );
  NAND4_X1 U25097 ( .A1(n21207), .A2(n21206), .A3(n21205), .A4(n21204), .ZN(
        n21208) );
  OR4_X1 U25098 ( .A1(n21211), .A2(n21210), .A3(n21209), .A4(n21208), .ZN(
        n21212) );
  NAND2_X1 U25099 ( .A1(n21212), .A2(n24720), .ZN(n21283) );
  AOI22_X1 U25100 ( .A1(n24693), .A2(\xmem_data[104][0] ), .B1(n30863), .B2(
        \xmem_data[105][0] ), .ZN(n21217) );
  AND2_X1 U25101 ( .A1(n3220), .A2(\xmem_data[107][0] ), .ZN(n21213) );
  AOI21_X1 U25102 ( .B1(n24694), .B2(\xmem_data[106][0] ), .A(n21213), .ZN(
        n21216) );
  AOI22_X1 U25103 ( .A1(n24696), .A2(\xmem_data[108][0] ), .B1(n24695), .B2(
        \xmem_data[109][0] ), .ZN(n21215) );
  AOI22_X1 U25104 ( .A1(n24697), .A2(\xmem_data[110][0] ), .B1(n24140), .B2(
        \xmem_data[111][0] ), .ZN(n21214) );
  NAND4_X1 U25105 ( .A1(n21217), .A2(n21216), .A3(n21215), .A4(n21214), .ZN(
        n21233) );
  AOI22_X1 U25106 ( .A1(n23724), .A2(\xmem_data[96][0] ), .B1(n31314), .B2(
        \xmem_data[97][0] ), .ZN(n21221) );
  AOI22_X1 U25107 ( .A1(n24685), .A2(\xmem_data[98][0] ), .B1(n28500), .B2(
        \xmem_data[99][0] ), .ZN(n21220) );
  AOI22_X1 U25108 ( .A1(n24687), .A2(\xmem_data[100][0] ), .B1(n24686), .B2(
        \xmem_data[101][0] ), .ZN(n21219) );
  AOI22_X1 U25109 ( .A1(n24688), .A2(\xmem_data[102][0] ), .B1(n29118), .B2(
        \xmem_data[103][0] ), .ZN(n21218) );
  NAND4_X1 U25110 ( .A1(n21221), .A2(n21220), .A3(n21219), .A4(n21218), .ZN(
        n21232) );
  AOI22_X1 U25111 ( .A1(n24702), .A2(\xmem_data[112][0] ), .B1(n29103), .B2(
        \xmem_data[113][0] ), .ZN(n21225) );
  AOI22_X1 U25112 ( .A1(n25422), .A2(\xmem_data[114][0] ), .B1(n25456), .B2(
        \xmem_data[115][0] ), .ZN(n21224) );
  AOI22_X1 U25113 ( .A1(n23762), .A2(\xmem_data[116][0] ), .B1(n13168), .B2(
        \xmem_data[117][0] ), .ZN(n21223) );
  AOI22_X1 U25114 ( .A1(n28298), .A2(\xmem_data[118][0] ), .B1(n30541), .B2(
        \xmem_data[119][0] ), .ZN(n21222) );
  NAND4_X1 U25115 ( .A1(n21225), .A2(n21224), .A3(n21223), .A4(n21222), .ZN(
        n21231) );
  AOI22_X1 U25116 ( .A1(n25607), .A2(\xmem_data[120][0] ), .B1(n29279), .B2(
        \xmem_data[121][0] ), .ZN(n21229) );
  AOI22_X1 U25117 ( .A1(n24708), .A2(\xmem_data[122][0] ), .B1(n24707), .B2(
        \xmem_data[123][0] ), .ZN(n21228) );
  AOI22_X1 U25118 ( .A1(n24710), .A2(\xmem_data[124][0] ), .B1(n24709), .B2(
        \xmem_data[125][0] ), .ZN(n21227) );
  AOI22_X1 U25119 ( .A1(n28385), .A2(\xmem_data[126][0] ), .B1(n24117), .B2(
        \xmem_data[127][0] ), .ZN(n21226) );
  NAND4_X1 U25120 ( .A1(n21229), .A2(n21228), .A3(n21227), .A4(n21226), .ZN(
        n21230) );
  OR4_X1 U25121 ( .A1(n21233), .A2(n21232), .A3(n21231), .A4(n21230), .ZN(
        n21234) );
  NAND2_X1 U25122 ( .A1(n21234), .A2(n24722), .ZN(n21282) );
  AOI22_X1 U25123 ( .A1(n24630), .A2(\xmem_data[40][0] ), .B1(n3247), .B2(
        \xmem_data[41][0] ), .ZN(n21239) );
  AND2_X1 U25124 ( .A1(n3218), .A2(\xmem_data[43][0] ), .ZN(n21235) );
  AOI21_X1 U25125 ( .B1(n24631), .B2(\xmem_data[42][0] ), .A(n21235), .ZN(
        n21238) );
  AOI22_X1 U25126 ( .A1(n24632), .A2(\xmem_data[44][0] ), .B1(n25491), .B2(
        \xmem_data[45][0] ), .ZN(n21237) );
  AOI22_X1 U25127 ( .A1(n3342), .A2(\xmem_data[46][0] ), .B1(n24633), .B2(
        \xmem_data[47][0] ), .ZN(n21236) );
  NAND4_X1 U25128 ( .A1(n21239), .A2(n21238), .A3(n21237), .A4(n21236), .ZN(
        n21256) );
  AOI22_X1 U25129 ( .A1(n24623), .A2(\xmem_data[32][0] ), .B1(n24622), .B2(
        \xmem_data[33][0] ), .ZN(n21244) );
  AOI22_X1 U25130 ( .A1(n24685), .A2(\xmem_data[34][0] ), .B1(n11008), .B2(
        \xmem_data[35][0] ), .ZN(n21243) );
  AND2_X1 U25131 ( .A1(n24624), .A2(\xmem_data[37][0] ), .ZN(n21240) );
  AOI21_X1 U25132 ( .B1(n29298), .B2(\xmem_data[36][0] ), .A(n21240), .ZN(
        n21242) );
  AOI22_X1 U25133 ( .A1(n24688), .A2(\xmem_data[38][0] ), .B1(n24625), .B2(
        \xmem_data[39][0] ), .ZN(n21241) );
  NAND4_X1 U25134 ( .A1(n21244), .A2(n21243), .A3(n21242), .A4(n21241), .ZN(
        n21255) );
  AOI22_X1 U25135 ( .A1(n3282), .A2(\xmem_data[48][0] ), .B1(n30877), .B2(
        \xmem_data[49][0] ), .ZN(n21248) );
  AOI22_X1 U25136 ( .A1(n24638), .A2(\xmem_data[50][0] ), .B1(n28373), .B2(
        \xmem_data[51][0] ), .ZN(n21247) );
  AOI22_X1 U25137 ( .A1(n24640), .A2(\xmem_data[52][0] ), .B1(n24639), .B2(
        \xmem_data[53][0] ), .ZN(n21246) );
  AOI22_X1 U25138 ( .A1(n30614), .A2(\xmem_data[54][0] ), .B1(n29271), .B2(
        \xmem_data[55][0] ), .ZN(n21245) );
  NAND4_X1 U25139 ( .A1(n21248), .A2(n21247), .A3(n21246), .A4(n21245), .ZN(
        n21254) );
  AOI22_X1 U25140 ( .A1(n3157), .A2(\xmem_data[56][0] ), .B1(n30542), .B2(
        \xmem_data[57][0] ), .ZN(n21252) );
  AOI22_X1 U25141 ( .A1(n20542), .A2(\xmem_data[58][0] ), .B1(n24645), .B2(
        \xmem_data[59][0] ), .ZN(n21251) );
  AOI22_X1 U25142 ( .A1(n23777), .A2(\xmem_data[60][0] ), .B1(n24646), .B2(
        \xmem_data[61][0] ), .ZN(n21250) );
  AOI22_X1 U25143 ( .A1(n24647), .A2(\xmem_data[62][0] ), .B1(n29055), .B2(
        \xmem_data[63][0] ), .ZN(n21249) );
  NAND4_X1 U25144 ( .A1(n21252), .A2(n21251), .A3(n21250), .A4(n21249), .ZN(
        n21253) );
  OR4_X1 U25145 ( .A1(n21256), .A2(n21255), .A3(n21254), .A4(n21253), .ZN(
        n21257) );
  NAND2_X1 U25146 ( .A1(n21257), .A2(n24659), .ZN(n21281) );
  AOI22_X1 U25147 ( .A1(n25401), .A2(\xmem_data[0][0] ), .B1(n28983), .B2(
        \xmem_data[1][0] ), .ZN(n21261) );
  AOI22_X1 U25148 ( .A1(n24606), .A2(\xmem_data[2][0] ), .B1(n27981), .B2(
        \xmem_data[3][0] ), .ZN(n21260) );
  AOI22_X1 U25149 ( .A1(n14982), .A2(\xmem_data[4][0] ), .B1(n27567), .B2(
        \xmem_data[5][0] ), .ZN(n21259) );
  AOI22_X1 U25150 ( .A1(n24607), .A2(\xmem_data[6][0] ), .B1(n24470), .B2(
        \xmem_data[7][0] ), .ZN(n21258) );
  NAND4_X1 U25151 ( .A1(n21261), .A2(n21260), .A3(n21259), .A4(n21258), .ZN(
        n21277) );
  AOI22_X1 U25152 ( .A1(n23732), .A2(\xmem_data[8][0] ), .B1(n3247), .B2(
        \xmem_data[9][0] ), .ZN(n21265) );
  AOI22_X1 U25153 ( .A1(n23734), .A2(\xmem_data[10][0] ), .B1(n3219), .B2(
        \xmem_data[11][0] ), .ZN(n21264) );
  AOI22_X1 U25154 ( .A1(n31368), .A2(\xmem_data[12][0] ), .B1(n20723), .B2(
        \xmem_data[13][0] ), .ZN(n21263) );
  AOI22_X1 U25155 ( .A1(n24141), .A2(\xmem_data[14][0] ), .B1(n17061), .B2(
        \xmem_data[15][0] ), .ZN(n21262) );
  NAND4_X1 U25156 ( .A1(n21265), .A2(n21264), .A3(n21263), .A4(n21262), .ZN(
        n21276) );
  AOI22_X1 U25157 ( .A1(n29762), .A2(\xmem_data[16][0] ), .B1(n24657), .B2(
        \xmem_data[17][0] ), .ZN(n21269) );
  AOI22_X1 U25158 ( .A1(n24554), .A2(\xmem_data[18][0] ), .B1(n24590), .B2(
        \xmem_data[19][0] ), .ZN(n21268) );
  AOI22_X1 U25159 ( .A1(n30508), .A2(\xmem_data[20][0] ), .B1(n13168), .B2(
        \xmem_data[21][0] ), .ZN(n21267) );
  AOI22_X1 U25160 ( .A1(n30614), .A2(\xmem_data[22][0] ), .B1(n24597), .B2(
        \xmem_data[23][0] ), .ZN(n21266) );
  NAND4_X1 U25161 ( .A1(n21269), .A2(n21268), .A3(n21267), .A4(n21266), .ZN(
        n21275) );
  AOI22_X1 U25162 ( .A1(n3157), .A2(\xmem_data[24][0] ), .B1(n28993), .B2(
        \xmem_data[25][0] ), .ZN(n21273) );
  AOI22_X1 U25163 ( .A1(n24593), .A2(\xmem_data[26][0] ), .B1(n24219), .B2(
        \xmem_data[27][0] ), .ZN(n21272) );
  AOI22_X1 U25164 ( .A1(n31255), .A2(\xmem_data[28][0] ), .B1(n24592), .B2(
        \xmem_data[29][0] ), .ZN(n21271) );
  AOI22_X1 U25165 ( .A1(n3326), .A2(\xmem_data[30][0] ), .B1(n3372), .B2(
        \xmem_data[31][0] ), .ZN(n21270) );
  NAND4_X1 U25166 ( .A1(n21273), .A2(n21272), .A3(n21271), .A4(n21270), .ZN(
        n21274) );
  OR4_X1 U25167 ( .A1(n21277), .A2(n21276), .A3(n21275), .A4(n21274), .ZN(
        n21279) );
  INV_X1 U25168 ( .A(n35490), .ZN(n21284) );
  AOI22_X1 U25169 ( .A1(n16999), .A2(\xmem_data[118][0] ), .B1(n27500), .B2(
        \xmem_data[119][0] ), .ZN(n21286) );
  AOI22_X1 U25170 ( .A1(n29028), .A2(\xmem_data[126][0] ), .B1(n29027), .B2(
        \xmem_data[127][0] ), .ZN(n21285) );
  AOI22_X1 U25171 ( .A1(n29281), .A2(\xmem_data[112][0] ), .B1(n28955), .B2(
        \xmem_data[113][0] ), .ZN(n21289) );
  AOI22_X1 U25172 ( .A1(n28062), .A2(\xmem_data[114][0] ), .B1(n3172), .B2(
        \xmem_data[115][0] ), .ZN(n21288) );
  AOI22_X1 U25173 ( .A1(n28974), .A2(\xmem_data[120][0] ), .B1(n21308), .B2(
        \xmem_data[121][0] ), .ZN(n21287) );
  AOI22_X1 U25174 ( .A1(n29017), .A2(\xmem_data[116][0] ), .B1(n28241), .B2(
        \xmem_data[117][0] ), .ZN(n21290) );
  NAND2_X1 U25175 ( .A1(n3903), .A2(n21290), .ZN(n21291) );
  AND2_X1 U25176 ( .A1(n20568), .A2(\xmem_data[122][0] ), .ZN(n21293) );
  AOI21_X1 U25177 ( .B1(n28470), .B2(\xmem_data[123][0] ), .A(n21293), .ZN(
        n21294) );
  INV_X1 U25178 ( .A(n21294), .ZN(n21297) );
  AOI22_X1 U25179 ( .A1(n3219), .A2(\xmem_data[124][0] ), .B1(n29026), .B2(
        \xmem_data[125][0] ), .ZN(n21295) );
  NOR2_X1 U25180 ( .A1(n21297), .A2(n21296), .ZN(n21306) );
  AOI22_X1 U25181 ( .A1(n29009), .A2(\xmem_data[104][0] ), .B1(n29008), .B2(
        \xmem_data[105][0] ), .ZN(n21301) );
  AOI22_X1 U25182 ( .A1(n3213), .A2(\xmem_data[106][0] ), .B1(n29010), .B2(
        \xmem_data[107][0] ), .ZN(n21300) );
  AOI22_X1 U25183 ( .A1(n24459), .A2(\xmem_data[108][0] ), .B1(n29012), .B2(
        \xmem_data[109][0] ), .ZN(n21299) );
  AOI22_X1 U25184 ( .A1(n30871), .A2(\xmem_data[110][0] ), .B1(n28061), .B2(
        \xmem_data[111][0] ), .ZN(n21298) );
  AOI22_X1 U25185 ( .A1(n25415), .A2(\xmem_data[96][0] ), .B1(n29231), .B2(
        \xmem_data[97][0] ), .ZN(n21305) );
  AOI22_X1 U25186 ( .A1(n29103), .A2(\xmem_data[98][0] ), .B1(n28972), .B2(
        \xmem_data[99][0] ), .ZN(n21304) );
  AOI22_X1 U25187 ( .A1(n29180), .A2(\xmem_data[100][0] ), .B1(n17013), .B2(
        \xmem_data[101][0] ), .ZN(n21303) );
  AOI22_X1 U25188 ( .A1(n23761), .A2(\xmem_data[102][0] ), .B1(n28980), .B2(
        \xmem_data[103][0] ), .ZN(n21302) );
  NAND3_X1 U25189 ( .A1(n21306), .A2(n3531), .A3(n3904), .ZN(n21307) );
  OAI21_X1 U25190 ( .B1(n3985), .B2(n21307), .A(n28968), .ZN(n21393) );
  AOI22_X1 U25191 ( .A1(n21309), .A2(\xmem_data[88][0] ), .B1(n21308), .B2(
        \xmem_data[89][0] ), .ZN(n21310) );
  NAND2_X1 U25192 ( .A1(n30257), .A2(\xmem_data[85][0] ), .ZN(n21312) );
  NAND2_X1 U25193 ( .A1(n29017), .A2(\xmem_data[84][0] ), .ZN(n21311) );
  NAND2_X1 U25194 ( .A1(n21312), .A2(n21311), .ZN(n21316) );
  AOI22_X1 U25195 ( .A1(n21059), .A2(\xmem_data[86][0] ), .B1(n29057), .B2(
        \xmem_data[87][0] ), .ZN(n21314) );
  AOI22_X1 U25196 ( .A1(n29028), .A2(\xmem_data[94][0] ), .B1(n29027), .B2(
        \xmem_data[95][0] ), .ZN(n21313) );
  NOR3_X1 U25197 ( .A1(n21317), .A2(n21316), .A3(n21315), .ZN(n21327) );
  AOI22_X1 U25198 ( .A1(n30882), .A2(\xmem_data[64][0] ), .B1(n3375), .B2(
        \xmem_data[65][0] ), .ZN(n21321) );
  AOI22_X1 U25199 ( .A1(n29045), .A2(\xmem_data[66][0] ), .B1(n24450), .B2(
        \xmem_data[67][0] ), .ZN(n21320) );
  AOI22_X1 U25200 ( .A1(n30854), .A2(\xmem_data[68][0] ), .B1(n25457), .B2(
        \xmem_data[69][0] ), .ZN(n21319) );
  AOI22_X1 U25201 ( .A1(n28375), .A2(\xmem_data[70][0] ), .B1(n20541), .B2(
        \xmem_data[71][0] ), .ZN(n21318) );
  AOI22_X1 U25202 ( .A1(n24134), .A2(\xmem_data[74][0] ), .B1(n29010), .B2(
        \xmem_data[75][0] ), .ZN(n21325) );
  AOI22_X1 U25203 ( .A1(n29009), .A2(\xmem_data[72][0] ), .B1(n29008), .B2(
        \xmem_data[73][0] ), .ZN(n21324) );
  AOI22_X1 U25204 ( .A1(n29048), .A2(\xmem_data[76][0] ), .B1(n29012), .B2(
        \xmem_data[77][0] ), .ZN(n21323) );
  AOI22_X1 U25205 ( .A1(n29238), .A2(\xmem_data[78][0] ), .B1(n30849), .B2(
        \xmem_data[79][0] ), .ZN(n21322) );
  NAND3_X1 U25206 ( .A1(n21327), .A2(n3788), .A3(n21326), .ZN(n21337) );
  AOI22_X1 U25207 ( .A1(n20816), .A2(\xmem_data[80][0] ), .B1(n28955), .B2(
        \xmem_data[81][0] ), .ZN(n21328) );
  INV_X1 U25208 ( .A(n21328), .ZN(n21332) );
  AOI22_X1 U25209 ( .A1(n3218), .A2(\xmem_data[92][0] ), .B1(n29026), .B2(
        \xmem_data[93][0] ), .ZN(n21330) );
  AOI22_X1 U25210 ( .A1(n14975), .A2(\xmem_data[82][0] ), .B1(n13486), .B2(
        \xmem_data[83][0] ), .ZN(n21329) );
  NAND2_X1 U25211 ( .A1(n21330), .A2(n21329), .ZN(n21331) );
  NAND2_X1 U25212 ( .A1(n28082), .A2(\xmem_data[91][0] ), .ZN(n21334) );
  NAND2_X1 U25213 ( .A1(n30589), .A2(\xmem_data[90][0] ), .ZN(n21333) );
  NAND2_X1 U25214 ( .A1(n21334), .A2(n21333), .ZN(n21335) );
  OAI21_X1 U25215 ( .B1(n21337), .B2(n21336), .A(n29041), .ZN(n21392) );
  AND2_X1 U25216 ( .A1(n25442), .A2(\xmem_data[58][0] ), .ZN(n21338) );
  AOI21_X1 U25217 ( .B1(n20518), .B2(\xmem_data[59][0] ), .A(n21338), .ZN(
        n21345) );
  AOI22_X1 U25218 ( .A1(n23739), .A2(\xmem_data[62][0] ), .B1(n25694), .B2(
        \xmem_data[63][0] ), .ZN(n21339) );
  INV_X1 U25219 ( .A(n21339), .ZN(n21343) );
  AOI22_X1 U25220 ( .A1(n3222), .A2(\xmem_data[60][0] ), .B1(n29065), .B2(
        \xmem_data[61][0] ), .ZN(n21341) );
  AOI22_X1 U25221 ( .A1(n31262), .A2(\xmem_data[56][0] ), .B1(n21308), .B2(
        \xmem_data[57][0] ), .ZN(n21340) );
  NAND2_X1 U25222 ( .A1(n21340), .A2(n21341), .ZN(n21342) );
  NOR2_X1 U25223 ( .A1(n21343), .A2(n21342), .ZN(n21344) );
  NAND2_X1 U25224 ( .A1(n21345), .A2(n21344), .ZN(n21352) );
  AOI22_X1 U25225 ( .A1(n29055), .A2(\xmem_data[48][0] ), .B1(n29054), .B2(
        \xmem_data[49][0] ), .ZN(n21350) );
  AOI22_X1 U25226 ( .A1(n29245), .A2(\xmem_data[50][0] ), .B1(n22684), .B2(
        \xmem_data[51][0] ), .ZN(n21349) );
  AND2_X1 U25227 ( .A1(n20733), .A2(\xmem_data[52][0] ), .ZN(n21346) );
  AOI21_X1 U25228 ( .B1(n27568), .B2(\xmem_data[53][0] ), .A(n21346), .ZN(
        n21348) );
  AOI22_X1 U25229 ( .A1(n27957), .A2(\xmem_data[54][0] ), .B1(n29057), .B2(
        \xmem_data[55][0] ), .ZN(n21347) );
  NAND4_X1 U25230 ( .A1(n21350), .A2(n21349), .A3(n21348), .A4(n21347), .ZN(
        n21351) );
  AOI22_X1 U25231 ( .A1(n29046), .A2(\xmem_data[40][0] ), .B1(n25607), .B2(
        \xmem_data[41][0] ), .ZN(n21356) );
  AOI22_X1 U25232 ( .A1(n13188), .A2(\xmem_data[42][0] ), .B1(n31330), .B2(
        \xmem_data[43][0] ), .ZN(n21355) );
  AOI22_X1 U25233 ( .A1(n29048), .A2(\xmem_data[44][0] ), .B1(n29047), .B2(
        \xmem_data[45][0] ), .ZN(n21354) );
  AOI22_X1 U25234 ( .A1(n29049), .A2(\xmem_data[46][0] ), .B1(n3178), .B2(
        \xmem_data[47][0] ), .ZN(n21353) );
  NAND4_X1 U25235 ( .A1(n21356), .A2(n21355), .A3(n21354), .A4(n21353), .ZN(
        n21362) );
  AOI22_X1 U25236 ( .A1(n28509), .A2(\xmem_data[32][0] ), .B1(n28952), .B2(
        \xmem_data[33][0] ), .ZN(n21360) );
  AOI22_X1 U25237 ( .A1(n29103), .A2(\xmem_data[34][0] ), .B1(n25422), .B2(
        \xmem_data[35][0] ), .ZN(n21359) );
  AOI22_X1 U25238 ( .A1(n28373), .A2(\xmem_data[36][0] ), .B1(n23792), .B2(
        \xmem_data[37][0] ), .ZN(n21358) );
  AOI22_X1 U25239 ( .A1(n24212), .A2(\xmem_data[38][0] ), .B1(n16986), .B2(
        \xmem_data[39][0] ), .ZN(n21357) );
  NAND4_X1 U25240 ( .A1(n21360), .A2(n21359), .A3(n21358), .A4(n21357), .ZN(
        n21361) );
  OAI21_X1 U25241 ( .B1(n21364), .B2(n21363), .A(n29078), .ZN(n21391) );
  AND2_X1 U25242 ( .A1(n28979), .A2(\xmem_data[20][0] ), .ZN(n21365) );
  AOI21_X1 U25243 ( .B1(n29657), .B2(\xmem_data[21][0] ), .A(n21365), .ZN(
        n21366) );
  INV_X1 U25244 ( .A(n21366), .ZN(n21371) );
  AOI22_X1 U25245 ( .A1(n28429), .A2(\xmem_data[16][0] ), .B1(n28955), .B2(
        \xmem_data[17][0] ), .ZN(n21369) );
  AOI22_X1 U25246 ( .A1(n29125), .A2(\xmem_data[22][0] ), .B1(n20953), .B2(
        \xmem_data[23][0] ), .ZN(n21368) );
  AOI22_X1 U25247 ( .A1(n28983), .A2(\xmem_data[18][0] ), .B1(n3172), .B2(
        \xmem_data[19][0] ), .ZN(n21367) );
  NOR2_X1 U25248 ( .A1(n21371), .A2(n21370), .ZN(n21382) );
  AOI22_X1 U25249 ( .A1(n29309), .A2(\xmem_data[8][0] ), .B1(n31328), .B2(
        \xmem_data[9][0] ), .ZN(n21375) );
  AOI22_X1 U25250 ( .A1(n28993), .A2(\xmem_data[10][0] ), .B1(n21007), .B2(
        \xmem_data[11][0] ), .ZN(n21374) );
  AOI22_X1 U25251 ( .A1(n29048), .A2(\xmem_data[12][0] ), .B1(n28994), .B2(
        \xmem_data[13][0] ), .ZN(n21373) );
  AOI22_X1 U25252 ( .A1(n23776), .A2(\xmem_data[14][0] ), .B1(n3326), .B2(
        \xmem_data[15][0] ), .ZN(n21372) );
  NAND4_X1 U25253 ( .A1(n21375), .A2(n21374), .A3(n21373), .A4(n21372), .ZN(
        n21380) );
  AOI22_X1 U25254 ( .A1(n25629), .A2(\xmem_data[24][0] ), .B1(n25443), .B2(
        \xmem_data[25][0] ), .ZN(n21378) );
  AOI22_X1 U25255 ( .A1(n23739), .A2(\xmem_data[30][0] ), .B1(n20994), .B2(
        \xmem_data[31][0] ), .ZN(n21377) );
  AOI22_X1 U25256 ( .A1(n3221), .A2(\xmem_data[28][0] ), .B1(n27445), .B2(
        \xmem_data[29][0] ), .ZN(n21376) );
  NAND3_X1 U25257 ( .A1(n21378), .A2(n21377), .A3(n21376), .ZN(n21379) );
  NOR2_X1 U25258 ( .A1(n21380), .A2(n21379), .ZN(n21381) );
  NAND2_X1 U25259 ( .A1(n21382), .A2(n21381), .ZN(n21389) );
  AOI22_X1 U25260 ( .A1(n28509), .A2(\xmem_data[0][0] ), .B1(n28952), .B2(
        \xmem_data[1][0] ), .ZN(n21386) );
  AOI22_X1 U25261 ( .A1(n29103), .A2(\xmem_data[2][0] ), .B1(n25422), .B2(
        \xmem_data[3][0] ), .ZN(n21385) );
  AOI22_X1 U25262 ( .A1(n30884), .A2(\xmem_data[4][0] ), .B1(n27453), .B2(
        \xmem_data[5][0] ), .ZN(n21384) );
  AOI22_X1 U25263 ( .A1(n24212), .A2(\xmem_data[6][0] ), .B1(n28980), .B2(
        \xmem_data[7][0] ), .ZN(n21383) );
  AOI22_X1 U25264 ( .A1(n29286), .A2(\xmem_data[26][0] ), .B1(n30503), .B2(
        \xmem_data[27][0] ), .ZN(n21387) );
  NAND2_X1 U25265 ( .A1(n3909), .A2(n21387), .ZN(n21388) );
  OAI21_X1 U25266 ( .B1(n21389), .B2(n21388), .A(n29002), .ZN(n21390) );
  INV_X1 U25267 ( .A(n35726), .ZN(n21394) );
  INV_X1 U25268 ( .A(n35592), .ZN(n21395) );
  XNOR2_X1 U25269 ( .A(n31798), .B(\fmem_data[14][3] ), .ZN(n31945) );
  AOI22_X1 U25270 ( .A1(n30949), .A2(\xmem_data[16][4] ), .B1(n25398), .B2(
        \xmem_data[17][4] ), .ZN(n21401) );
  AOI22_X1 U25271 ( .A1(n27855), .A2(\xmem_data[18][4] ), .B1(n29049), .B2(
        \xmem_data[19][4] ), .ZN(n21400) );
  AOI22_X1 U25272 ( .A1(n25575), .A2(\xmem_data[20][4] ), .B1(n3372), .B2(
        \xmem_data[21][4] ), .ZN(n21399) );
  AOI22_X1 U25273 ( .A1(n29816), .A2(\xmem_data[22][4] ), .B1(n31362), .B2(
        \xmem_data[23][4] ), .ZN(n21398) );
  NAND4_X1 U25274 ( .A1(n21401), .A2(n21400), .A3(n21399), .A4(n21398), .ZN(
        n21407) );
  AOI22_X1 U25275 ( .A1(n27847), .A2(\xmem_data[24][4] ), .B1(n29017), .B2(
        \xmem_data[25][4] ), .ZN(n21405) );
  AOI22_X1 U25276 ( .A1(n27852), .A2(\xmem_data[26][4] ), .B1(n22727), .B2(
        \xmem_data[27][4] ), .ZN(n21404) );
  AOI22_X1 U25277 ( .A1(n27436), .A2(\xmem_data[28][4] ), .B1(n29118), .B2(
        \xmem_data[29][4] ), .ZN(n21403) );
  AOI22_X1 U25278 ( .A1(n3317), .A2(\xmem_data[30][4] ), .B1(n28501), .B2(
        \xmem_data[31][4] ), .ZN(n21402) );
  NAND4_X1 U25279 ( .A1(n21405), .A2(n21404), .A3(n21403), .A4(n21402), .ZN(
        n21406) );
  OR2_X1 U25280 ( .A1(n21407), .A2(n21406), .ZN(n21421) );
  AOI22_X1 U25281 ( .A1(n24631), .A2(\xmem_data[0][4] ), .B1(n3217), .B2(
        \xmem_data[1][4] ), .ZN(n21408) );
  INV_X1 U25282 ( .A(n21408), .ZN(n21419) );
  AOI22_X1 U25283 ( .A1(n25707), .A2(\xmem_data[8][4] ), .B1(n27863), .B2(
        \xmem_data[9][4] ), .ZN(n21412) );
  AOI22_X1 U25284 ( .A1(n29308), .A2(\xmem_data[10][4] ), .B1(n13168), .B2(
        \xmem_data[11][4] ), .ZN(n21411) );
  AOI22_X1 U25285 ( .A1(n27515), .A2(\xmem_data[12][4] ), .B1(n25572), .B2(
        \xmem_data[13][4] ), .ZN(n21410) );
  AOI22_X1 U25286 ( .A1(n29008), .A2(\xmem_data[14][4] ), .B1(n27864), .B2(
        \xmem_data[15][4] ), .ZN(n21409) );
  NAND4_X1 U25287 ( .A1(n21412), .A2(n21411), .A3(n21410), .A4(n21409), .ZN(
        n21418) );
  AOI22_X1 U25288 ( .A1(n20807), .A2(\xmem_data[4][4] ), .B1(n17061), .B2(
        \xmem_data[5][4] ), .ZN(n21414) );
  NAND2_X1 U25289 ( .A1(n29706), .A2(\xmem_data[6][4] ), .ZN(n21413) );
  NAND2_X1 U25290 ( .A1(n21414), .A2(n21413), .ZN(n21417) );
  AOI22_X1 U25291 ( .A1(n31368), .A2(\xmem_data[2][4] ), .B1(n27869), .B2(
        \xmem_data[3][4] ), .ZN(n21415) );
  NOR2_X1 U25292 ( .A1(n21421), .A2(n21420), .ZN(n21422) );
  NOR2_X1 U25293 ( .A1(n21422), .A2(n27877), .ZN(n21445) );
  AOI22_X1 U25294 ( .A1(n28503), .A2(\xmem_data[32][4] ), .B1(n3221), .B2(
        \xmem_data[33][4] ), .ZN(n21426) );
  AOI22_X1 U25295 ( .A1(n28367), .A2(\xmem_data[34][4] ), .B1(n27444), .B2(
        \xmem_data[35][4] ), .ZN(n21425) );
  AOI22_X1 U25296 ( .A1(n27938), .A2(\xmem_data[36][4] ), .B1(n24633), .B2(
        \xmem_data[37][4] ), .ZN(n21424) );
  AOI22_X1 U25297 ( .A1(n3375), .A2(\xmem_data[38][4] ), .B1(n29306), .B2(
        \xmem_data[39][4] ), .ZN(n21423) );
  NAND4_X1 U25298 ( .A1(n21426), .A2(n21425), .A3(n21424), .A4(n21423), .ZN(
        n21442) );
  AOI22_X1 U25299 ( .A1(n25422), .A2(\xmem_data[40][4] ), .B1(n3358), .B2(
        \xmem_data[41][4] ), .ZN(n21430) );
  AOI22_X1 U25300 ( .A1(n27944), .A2(\xmem_data[42][4] ), .B1(n24212), .B2(
        \xmem_data[43][4] ), .ZN(n21429) );
  AOI22_X1 U25301 ( .A1(n31268), .A2(\xmem_data[44][4] ), .B1(n27536), .B2(
        \xmem_data[45][4] ), .ZN(n21428) );
  AOI22_X1 U25302 ( .A1(n23795), .A2(\xmem_data[46][4] ), .B1(n27516), .B2(
        \xmem_data[47][4] ), .ZN(n21427) );
  NAND4_X1 U25303 ( .A1(n21430), .A2(n21429), .A3(n21428), .A4(n21427), .ZN(
        n21441) );
  AOI22_X1 U25304 ( .A1(n21007), .A2(\xmem_data[48][4] ), .B1(n29048), .B2(
        \xmem_data[49][4] ), .ZN(n21434) );
  AOI22_X1 U25305 ( .A1(n22717), .A2(\xmem_data[50][4] ), .B1(n27950), .B2(
        \xmem_data[51][4] ), .ZN(n21433) );
  AOI22_X1 U25306 ( .A1(n27952), .A2(\xmem_data[52][4] ), .B1(n27951), .B2(
        \xmem_data[53][4] ), .ZN(n21432) );
  AOI22_X1 U25307 ( .A1(n3270), .A2(\xmem_data[54][4] ), .B1(n20553), .B2(
        \xmem_data[55][4] ), .ZN(n21431) );
  NAND4_X1 U25308 ( .A1(n21434), .A2(n21433), .A3(n21432), .A4(n21431), .ZN(
        n21440) );
  AOI22_X1 U25309 ( .A1(n25582), .A2(\xmem_data[56][4] ), .B1(n25359), .B2(
        \xmem_data[57][4] ), .ZN(n21438) );
  AOI22_X1 U25310 ( .A1(n20770), .A2(\xmem_data[58][4] ), .B1(n27957), .B2(
        \xmem_data[59][4] ), .ZN(n21437) );
  AOI22_X1 U25311 ( .A1(n27959), .A2(\xmem_data[60][4] ), .B1(n27958), .B2(
        \xmem_data[61][4] ), .ZN(n21436) );
  AOI22_X1 U25312 ( .A1(n3228), .A2(\xmem_data[62][4] ), .B1(n30863), .B2(
        \xmem_data[63][4] ), .ZN(n21435) );
  NAND4_X1 U25313 ( .A1(n21438), .A2(n21437), .A3(n21436), .A4(n21435), .ZN(
        n21439) );
  OR4_X1 U25314 ( .A1(n21442), .A2(n21441), .A3(n21440), .A4(n21439), .ZN(
        n21443) );
  AND2_X1 U25315 ( .A1(n21443), .A2(n27968), .ZN(n21444) );
  NOR2_X1 U25316 ( .A1(n21445), .A2(n21444), .ZN(n21491) );
  NOR2_X1 U25317 ( .A1(n27877), .A2(n39039), .ZN(n21446) );
  NAND2_X1 U25318 ( .A1(n30877), .A2(n21446), .ZN(n21490) );
  AOI22_X1 U25319 ( .A1(n27902), .A2(\xmem_data[96][4] ), .B1(n3221), .B2(
        \xmem_data[97][4] ), .ZN(n21450) );
  AOI22_X1 U25320 ( .A1(n29288), .A2(\xmem_data[98][4] ), .B1(n31367), .B2(
        \xmem_data[99][4] ), .ZN(n21449) );
  AOI22_X1 U25321 ( .A1(n27904), .A2(\xmem_data[100][4] ), .B1(n27903), .B2(
        \xmem_data[101][4] ), .ZN(n21448) );
  AOI22_X1 U25322 ( .A1(n27905), .A2(\xmem_data[102][4] ), .B1(n29306), .B2(
        \xmem_data[103][4] ), .ZN(n21447) );
  NAND4_X1 U25323 ( .A1(n21450), .A2(n21449), .A3(n21448), .A4(n21447), .ZN(
        n21466) );
  AOI22_X1 U25324 ( .A1(n27910), .A2(\xmem_data[104][4] ), .B1(n29180), .B2(
        \xmem_data[105][4] ), .ZN(n21454) );
  AOI22_X1 U25325 ( .A1(n27911), .A2(\xmem_data[106][4] ), .B1(n28515), .B2(
        \xmem_data[107][4] ), .ZN(n21453) );
  AOI22_X1 U25326 ( .A1(n3176), .A2(\xmem_data[108][4] ), .B1(n27912), .B2(
        \xmem_data[109][4] ), .ZN(n21452) );
  AOI22_X1 U25327 ( .A1(n28091), .A2(\xmem_data[110][4] ), .B1(n23716), .B2(
        \xmem_data[111][4] ), .ZN(n21451) );
  NAND4_X1 U25328 ( .A1(n21454), .A2(n21453), .A3(n21452), .A4(n21451), .ZN(
        n21465) );
  AOI22_X1 U25329 ( .A1(n27919), .A2(\xmem_data[112][4] ), .B1(n27918), .B2(
        \xmem_data[113][4] ), .ZN(n21458) );
  AOI22_X1 U25330 ( .A1(n22682), .A2(\xmem_data[114][4] ), .B1(n27920), .B2(
        \xmem_data[115][4] ), .ZN(n21457) );
  AOI22_X1 U25331 ( .A1(n3325), .A2(\xmem_data[116][4] ), .B1(n28429), .B2(
        \xmem_data[117][4] ), .ZN(n21456) );
  AOI22_X1 U25332 ( .A1(n30686), .A2(\xmem_data[118][4] ), .B1(n30599), .B2(
        \xmem_data[119][4] ), .ZN(n21455) );
  NAND4_X1 U25333 ( .A1(n21458), .A2(n21457), .A3(n21456), .A4(n21455), .ZN(
        n21464) );
  AOI22_X1 U25334 ( .A1(n22719), .A2(\xmem_data[120][4] ), .B1(n11008), .B2(
        \xmem_data[121][4] ), .ZN(n21462) );
  AOI22_X1 U25335 ( .A1(n29298), .A2(\xmem_data[122][4] ), .B1(n24624), .B2(
        \xmem_data[123][4] ), .ZN(n21461) );
  AOI22_X1 U25336 ( .A1(n27925), .A2(\xmem_data[124][4] ), .B1(n27563), .B2(
        \xmem_data[125][4] ), .ZN(n21460) );
  AOI22_X1 U25337 ( .A1(n29661), .A2(\xmem_data[126][4] ), .B1(n25442), .B2(
        \xmem_data[127][4] ), .ZN(n21459) );
  NAND4_X1 U25338 ( .A1(n21462), .A2(n21461), .A3(n21460), .A4(n21459), .ZN(
        n21463) );
  OR4_X1 U25339 ( .A1(n21466), .A2(n21465), .A3(n21464), .A4(n21463), .ZN(
        n21488) );
  AOI22_X1 U25340 ( .A1(n25730), .A2(\xmem_data[64][4] ), .B1(n3218), .B2(
        \xmem_data[65][4] ), .ZN(n21470) );
  AOI22_X1 U25341 ( .A1(n29288), .A2(\xmem_data[66][4] ), .B1(n30963), .B2(
        \xmem_data[67][4] ), .ZN(n21469) );
  AOI22_X1 U25342 ( .A1(n27938), .A2(\xmem_data[68][4] ), .B1(n29104), .B2(
        \xmem_data[69][4] ), .ZN(n21468) );
  AOI22_X1 U25343 ( .A1(n27905), .A2(\xmem_data[70][4] ), .B1(n23771), .B2(
        \xmem_data[71][4] ), .ZN(n21467) );
  NAND4_X1 U25344 ( .A1(n21470), .A2(n21469), .A3(n21468), .A4(n21467), .ZN(
        n21486) );
  AOI22_X1 U25345 ( .A1(n27508), .A2(\xmem_data[72][4] ), .B1(n3357), .B2(
        \xmem_data[73][4] ), .ZN(n21474) );
  AOI22_X1 U25346 ( .A1(n27944), .A2(\xmem_data[74][4] ), .B1(n24212), .B2(
        \xmem_data[75][4] ), .ZN(n21473) );
  AOI22_X1 U25347 ( .A1(n31268), .A2(\xmem_data[76][4] ), .B1(n28052), .B2(
        \xmem_data[77][4] ), .ZN(n21472) );
  AOI22_X1 U25348 ( .A1(n29396), .A2(\xmem_data[78][4] ), .B1(n27516), .B2(
        \xmem_data[79][4] ), .ZN(n21471) );
  NAND4_X1 U25349 ( .A1(n21474), .A2(n21473), .A3(n21472), .A4(n21471), .ZN(
        n21485) );
  AOI22_X1 U25350 ( .A1(n20542), .A2(\xmem_data[80][4] ), .B1(n25398), .B2(
        \xmem_data[81][4] ), .ZN(n21478) );
  AOI22_X1 U25351 ( .A1(n21008), .A2(\xmem_data[82][4] ), .B1(n27950), .B2(
        \xmem_data[83][4] ), .ZN(n21477) );
  AOI22_X1 U25352 ( .A1(n27952), .A2(\xmem_data[84][4] ), .B1(n27951), .B2(
        \xmem_data[85][4] ), .ZN(n21476) );
  AOI22_X1 U25353 ( .A1(n25401), .A2(\xmem_data[86][4] ), .B1(n24622), .B2(
        \xmem_data[87][4] ), .ZN(n21475) );
  NAND4_X1 U25354 ( .A1(n21478), .A2(n21477), .A3(n21476), .A4(n21475), .ZN(
        n21484) );
  AOI22_X1 U25355 ( .A1(n25582), .A2(\xmem_data[88][4] ), .B1(n23781), .B2(
        \xmem_data[89][4] ), .ZN(n21482) );
  AOI22_X1 U25356 ( .A1(n30674), .A2(\xmem_data[90][4] ), .B1(n27957), .B2(
        \xmem_data[91][4] ), .ZN(n21481) );
  AOI22_X1 U25357 ( .A1(n27959), .A2(\xmem_data[92][4] ), .B1(n27958), .B2(
        \xmem_data[93][4] ), .ZN(n21480) );
  AOI22_X1 U25358 ( .A1(n3229), .A2(\xmem_data[94][4] ), .B1(n24439), .B2(
        \xmem_data[95][4] ), .ZN(n21479) );
  NAND4_X1 U25359 ( .A1(n21482), .A2(n21481), .A3(n21480), .A4(n21479), .ZN(
        n21483) );
  OR4_X1 U25360 ( .A1(n21486), .A2(n21485), .A3(n21484), .A4(n21483), .ZN(
        n21487) );
  AOI22_X1 U25361 ( .A1(n27937), .A2(n21488), .B1(n27935), .B2(n21487), .ZN(
        n21489) );
  OAI22_X1 U25362 ( .A1(n31945), .A2(n33741), .B1(n26271), .B2(n33603), .ZN(
        n34003) );
  AOI22_X1 U25363 ( .A1(n27902), .A2(\xmem_data[96][0] ), .B1(n3221), .B2(
        \xmem_data[97][0] ), .ZN(n21495) );
  AOI22_X1 U25364 ( .A1(n29065), .A2(\xmem_data[98][0] ), .B1(n24695), .B2(
        \xmem_data[99][0] ), .ZN(n21494) );
  AOI22_X1 U25365 ( .A1(n27904), .A2(\xmem_data[100][0] ), .B1(n27903), .B2(
        \xmem_data[101][0] ), .ZN(n21493) );
  AOI22_X1 U25366 ( .A1(n27905), .A2(\xmem_data[102][0] ), .B1(n25514), .B2(
        \xmem_data[103][0] ), .ZN(n21492) );
  NAND4_X1 U25367 ( .A1(n21495), .A2(n21494), .A3(n21493), .A4(n21492), .ZN(
        n21511) );
  AOI22_X1 U25368 ( .A1(n27910), .A2(\xmem_data[104][0] ), .B1(n29307), .B2(
        \xmem_data[105][0] ), .ZN(n21499) );
  AOI22_X1 U25369 ( .A1(n27911), .A2(\xmem_data[106][0] ), .B1(n25605), .B2(
        \xmem_data[107][0] ), .ZN(n21498) );
  AOI22_X1 U25370 ( .A1(n3176), .A2(\xmem_data[108][0] ), .B1(n27912), .B2(
        \xmem_data[109][0] ), .ZN(n21497) );
  AOI22_X1 U25371 ( .A1(n27455), .A2(\xmem_data[110][0] ), .B1(n25460), .B2(
        \xmem_data[111][0] ), .ZN(n21496) );
  NAND4_X1 U25372 ( .A1(n21499), .A2(n21498), .A3(n21497), .A4(n21496), .ZN(
        n21510) );
  AOI22_X1 U25373 ( .A1(n27919), .A2(\xmem_data[112][0] ), .B1(n27918), .B2(
        \xmem_data[113][0] ), .ZN(n21503) );
  AOI22_X1 U25374 ( .A1(n23722), .A2(\xmem_data[114][0] ), .B1(n27920), .B2(
        \xmem_data[115][0] ), .ZN(n21502) );
  AOI22_X1 U25375 ( .A1(n28493), .A2(\xmem_data[116][0] ), .B1(n30898), .B2(
        \xmem_data[117][0] ), .ZN(n21501) );
  AOI22_X1 U25376 ( .A1(n25718), .A2(\xmem_data[118][0] ), .B1(n24521), .B2(
        \xmem_data[119][0] ), .ZN(n21500) );
  NAND4_X1 U25377 ( .A1(n21503), .A2(n21502), .A3(n21501), .A4(n21500), .ZN(
        n21509) );
  AOI22_X1 U25378 ( .A1(n14976), .A2(\xmem_data[120][0] ), .B1(n27463), .B2(
        \xmem_data[121][0] ), .ZN(n21507) );
  AOI22_X1 U25379 ( .A1(n30901), .A2(\xmem_data[122][0] ), .B1(n30524), .B2(
        \xmem_data[123][0] ), .ZN(n21506) );
  AOI22_X1 U25380 ( .A1(n27925), .A2(\xmem_data[124][0] ), .B1(n31262), .B2(
        \xmem_data[125][0] ), .ZN(n21505) );
  AOI22_X1 U25381 ( .A1(n3388), .A2(\xmem_data[126][0] ), .B1(n25485), .B2(
        \xmem_data[127][0] ), .ZN(n21504) );
  NAND4_X1 U25382 ( .A1(n21507), .A2(n21506), .A3(n21505), .A4(n21504), .ZN(
        n21508) );
  OR4_X1 U25383 ( .A1(n21511), .A2(n21510), .A3(n21509), .A4(n21508), .ZN(
        n21533) );
  AOI22_X1 U25384 ( .A1(n27902), .A2(\xmem_data[64][0] ), .B1(n3218), .B2(
        \xmem_data[65][0] ), .ZN(n21515) );
  AOI22_X1 U25385 ( .A1(n25414), .A2(\xmem_data[66][0] ), .B1(n27444), .B2(
        \xmem_data[67][0] ), .ZN(n21514) );
  AOI22_X1 U25386 ( .A1(n27904), .A2(\xmem_data[68][0] ), .B1(n27903), .B2(
        \xmem_data[69][0] ), .ZN(n21513) );
  AOI22_X1 U25387 ( .A1(n27905), .A2(\xmem_data[70][0] ), .B1(n28007), .B2(
        \xmem_data[71][0] ), .ZN(n21512) );
  NAND4_X1 U25388 ( .A1(n21515), .A2(n21514), .A3(n21513), .A4(n21512), .ZN(
        n21531) );
  AOI22_X1 U25389 ( .A1(n29325), .A2(\xmem_data[88][0] ), .B1(n27981), .B2(
        \xmem_data[89][0] ), .ZN(n21519) );
  AOI22_X1 U25390 ( .A1(n28241), .A2(\xmem_data[90][0] ), .B1(n16999), .B2(
        \xmem_data[91][0] ), .ZN(n21518) );
  AOI22_X1 U25391 ( .A1(n27925), .A2(\xmem_data[92][0] ), .B1(n30908), .B2(
        \xmem_data[93][0] ), .ZN(n21517) );
  AOI22_X1 U25392 ( .A1(n25443), .A2(\xmem_data[94][0] ), .B1(n25485), .B2(
        \xmem_data[95][0] ), .ZN(n21516) );
  NAND4_X1 U25393 ( .A1(n21519), .A2(n21518), .A3(n21517), .A4(n21516), .ZN(
        n21530) );
  AOI22_X1 U25394 ( .A1(n27919), .A2(\xmem_data[80][0] ), .B1(n27918), .B2(
        \xmem_data[81][0] ), .ZN(n21523) );
  AOI22_X1 U25395 ( .A1(n16990), .A2(\xmem_data[82][0] ), .B1(n27920), .B2(
        \xmem_data[83][0] ), .ZN(n21522) );
  AOI22_X1 U25396 ( .A1(n28061), .A2(\xmem_data[84][0] ), .B1(n30495), .B2(
        \xmem_data[85][0] ), .ZN(n21521) );
  AOI22_X1 U25397 ( .A1(n3269), .A2(\xmem_data[86][0] ), .B1(n24521), .B2(
        \xmem_data[87][0] ), .ZN(n21520) );
  NAND4_X1 U25398 ( .A1(n21523), .A2(n21522), .A3(n21521), .A4(n21520), .ZN(
        n21529) );
  AOI22_X1 U25399 ( .A1(n27910), .A2(\xmem_data[72][0] ), .B1(n28415), .B2(
        \xmem_data[73][0] ), .ZN(n21527) );
  AOI22_X1 U25400 ( .A1(n27911), .A2(\xmem_data[74][0] ), .B1(n24212), .B2(
        \xmem_data[75][0] ), .ZN(n21526) );
  AOI22_X1 U25401 ( .A1(n3176), .A2(\xmem_data[76][0] ), .B1(n27912), .B2(
        \xmem_data[77][0] ), .ZN(n21525) );
  AOI22_X1 U25402 ( .A1(n31328), .A2(\xmem_data[78][0] ), .B1(n25383), .B2(
        \xmem_data[79][0] ), .ZN(n21524) );
  NAND4_X1 U25403 ( .A1(n21527), .A2(n21526), .A3(n21525), .A4(n21524), .ZN(
        n21528) );
  OR4_X1 U25404 ( .A1(n21531), .A2(n21530), .A3(n21529), .A4(n21528), .ZN(
        n21532) );
  AOI22_X1 U25405 ( .A1(n21533), .A2(n27937), .B1(n27935), .B2(n21532), .ZN(
        n21582) );
  AOI22_X1 U25406 ( .A1(n25422), .A2(\xmem_data[8][0] ), .B1(n27863), .B2(
        \xmem_data[9][0] ), .ZN(n21537) );
  AOI22_X1 U25407 ( .A1(n28152), .A2(\xmem_data[10][0] ), .B1(n13168), .B2(
        \xmem_data[11][0] ), .ZN(n21536) );
  AOI22_X1 U25408 ( .A1(n17041), .A2(\xmem_data[12][0] ), .B1(n25671), .B2(
        \xmem_data[13][0] ), .ZN(n21535) );
  AOI22_X1 U25409 ( .A1(n27818), .A2(\xmem_data[14][0] ), .B1(n27864), .B2(
        \xmem_data[15][0] ), .ZN(n21534) );
  NAND4_X1 U25410 ( .A1(n21537), .A2(n21536), .A3(n21535), .A4(n21534), .ZN(
        n21545) );
  AOI22_X1 U25411 ( .A1(n24562), .A2(\xmem_data[0][0] ), .B1(n3222), .B2(
        \xmem_data[1][0] ), .ZN(n21538) );
  INV_X1 U25412 ( .A(n21538), .ZN(n21544) );
  AOI22_X1 U25413 ( .A1(n23741), .A2(\xmem_data[4][0] ), .B1(n25415), .B2(
        \xmem_data[5][0] ), .ZN(n21539) );
  INV_X1 U25414 ( .A(n21539), .ZN(n21543) );
  AOI22_X1 U25415 ( .A1(n29494), .A2(\xmem_data[2][0] ), .B1(n27869), .B2(
        \xmem_data[3][0] ), .ZN(n21541) );
  NAND2_X1 U25416 ( .A1(n3375), .A2(\xmem_data[6][0] ), .ZN(n21540) );
  NAND2_X1 U25417 ( .A1(n21541), .A2(n21540), .ZN(n21542) );
  NOR3_X1 U25418 ( .A1(n21545), .A2(n21544), .A3(n3994), .ZN(n21551) );
  AOI22_X1 U25419 ( .A1(n27847), .A2(\xmem_data[24][0] ), .B1(n17049), .B2(
        \xmem_data[25][0] ), .ZN(n21549) );
  AOI22_X1 U25420 ( .A1(n27852), .A2(\xmem_data[26][0] ), .B1(n20951), .B2(
        \xmem_data[27][0] ), .ZN(n21548) );
  AOI22_X1 U25421 ( .A1(n29057), .A2(\xmem_data[28][0] ), .B1(n27563), .B2(
        \xmem_data[29][0] ), .ZN(n21547) );
  AOI22_X1 U25422 ( .A1(n3412), .A2(\xmem_data[30][0] ), .B1(n31347), .B2(
        \xmem_data[31][0] ), .ZN(n21546) );
  AND4_X1 U25423 ( .A1(n21549), .A2(n21548), .A3(n21547), .A4(n21546), .ZN(
        n21550) );
  NAND2_X1 U25424 ( .A1(n21551), .A2(n21550), .ZN(n21558) );
  AOI22_X1 U25425 ( .A1(n27919), .A2(\xmem_data[16][0] ), .B1(n16989), .B2(
        \xmem_data[17][0] ), .ZN(n21555) );
  AOI22_X1 U25426 ( .A1(n27855), .A2(\xmem_data[18][0] ), .B1(n30515), .B2(
        \xmem_data[19][0] ), .ZN(n21554) );
  AOI22_X1 U25427 ( .A1(n17002), .A2(\xmem_data[20][0] ), .B1(n25716), .B2(
        \xmem_data[21][0] ), .ZN(n21553) );
  AOI22_X1 U25428 ( .A1(n29297), .A2(\xmem_data[22][0] ), .B1(n28495), .B2(
        \xmem_data[23][0] ), .ZN(n21552) );
  NAND4_X1 U25429 ( .A1(n21555), .A2(n21554), .A3(n21553), .A4(n21552), .ZN(
        n21556) );
  AOI22_X1 U25430 ( .A1(n29254), .A2(\xmem_data[32][0] ), .B1(n3219), .B2(
        \xmem_data[33][0] ), .ZN(n21562) );
  AOI22_X1 U25431 ( .A1(n24533), .A2(\xmem_data[34][0] ), .B1(n23739), .B2(
        \xmem_data[35][0] ), .ZN(n21561) );
  AOI22_X1 U25432 ( .A1(n27938), .A2(\xmem_data[36][0] ), .B1(n28342), .B2(
        \xmem_data[37][0] ), .ZN(n21560) );
  AOI22_X1 U25433 ( .A1(n25451), .A2(\xmem_data[38][0] ), .B1(n31252), .B2(
        \xmem_data[39][0] ), .ZN(n21559) );
  NAND4_X1 U25434 ( .A1(n21562), .A2(n21561), .A3(n21560), .A4(n21559), .ZN(
        n21578) );
  AOI22_X1 U25435 ( .A1(n27447), .A2(\xmem_data[40][0] ), .B1(n28373), .B2(
        \xmem_data[41][0] ), .ZN(n21566) );
  AOI22_X1 U25436 ( .A1(n27944), .A2(\xmem_data[42][0] ), .B1(n24212), .B2(
        \xmem_data[43][0] ), .ZN(n21565) );
  AOI22_X1 U25437 ( .A1(n23763), .A2(\xmem_data[44][0] ), .B1(n29046), .B2(
        \xmem_data[45][0] ), .ZN(n21564) );
  AOI22_X1 U25438 ( .A1(n29605), .A2(\xmem_data[46][0] ), .B1(n20543), .B2(
        \xmem_data[47][0] ), .ZN(n21563) );
  NAND4_X1 U25439 ( .A1(n21566), .A2(n21565), .A3(n21564), .A4(n21563), .ZN(
        n21577) );
  AOI22_X1 U25440 ( .A1(n21007), .A2(\xmem_data[48][0] ), .B1(n20505), .B2(
        \xmem_data[49][0] ), .ZN(n21570) );
  AOI22_X1 U25441 ( .A1(n30617), .A2(\xmem_data[50][0] ), .B1(n27950), .B2(
        \xmem_data[51][0] ), .ZN(n21569) );
  AOI22_X1 U25442 ( .A1(n27952), .A2(\xmem_data[52][0] ), .B1(n27951), .B2(
        \xmem_data[53][0] ), .ZN(n21568) );
  AOI22_X1 U25443 ( .A1(n20817), .A2(\xmem_data[54][0] ), .B1(n25583), .B2(
        \xmem_data[55][0] ), .ZN(n21567) );
  NAND4_X1 U25444 ( .A1(n21570), .A2(n21569), .A3(n21568), .A4(n21567), .ZN(
        n21576) );
  AOI22_X1 U25445 ( .A1(n29151), .A2(\xmem_data[56][0] ), .B1(n20488), .B2(
        \xmem_data[57][0] ), .ZN(n21574) );
  AOI22_X1 U25446 ( .A1(n21060), .A2(\xmem_data[58][0] ), .B1(n27957), .B2(
        \xmem_data[59][0] ), .ZN(n21573) );
  AOI22_X1 U25447 ( .A1(n27959), .A2(\xmem_data[60][0] ), .B1(n27958), .B2(
        \xmem_data[61][0] ), .ZN(n21572) );
  AOI22_X1 U25448 ( .A1(n3153), .A2(\xmem_data[62][0] ), .B1(n3247), .B2(
        \xmem_data[63][0] ), .ZN(n21571) );
  NAND4_X1 U25449 ( .A1(n21574), .A2(n21573), .A3(n21572), .A4(n21571), .ZN(
        n21575) );
  OR4_X1 U25450 ( .A1(n21578), .A2(n21577), .A3(n21576), .A4(n21575), .ZN(
        n21579) );
  NAND3_X2 U25451 ( .A1(n21582), .A2(n21581), .A3(n21580), .ZN(n36244) );
  AOI22_X1 U25452 ( .A1(n25434), .A2(\xmem_data[32][0] ), .B1(n25677), .B2(
        \xmem_data[33][0] ), .ZN(n21587) );
  AOI22_X1 U25453 ( .A1(n14971), .A2(\xmem_data[34][0] ), .B1(n25435), .B2(
        \xmem_data[35][0] ), .ZN(n21586) );
  AOI22_X1 U25454 ( .A1(n28428), .A2(\xmem_data[36][0] ), .B1(n20551), .B2(
        \xmem_data[37][0] ), .ZN(n21585) );
  AOI22_X1 U25455 ( .A1(n3308), .A2(\xmem_data[38][0] ), .B1(n27525), .B2(
        \xmem_data[39][0] ), .ZN(n21584) );
  NAND4_X1 U25456 ( .A1(n21587), .A2(n21586), .A3(n21585), .A4(n21584), .ZN(
        n21603) );
  AOI22_X1 U25457 ( .A1(n25526), .A2(\xmem_data[40][0] ), .B1(n25406), .B2(
        \xmem_data[41][0] ), .ZN(n21591) );
  AOI22_X1 U25458 ( .A1(n30674), .A2(\xmem_data[42][0] ), .B1(n25440), .B2(
        \xmem_data[43][0] ), .ZN(n21590) );
  AOI22_X1 U25459 ( .A1(n25441), .A2(\xmem_data[44][0] ), .B1(n12471), .B2(
        \xmem_data[45][0] ), .ZN(n21589) );
  AOI22_X1 U25460 ( .A1(n25443), .A2(\xmem_data[46][0] ), .B1(n25442), .B2(
        \xmem_data[47][0] ), .ZN(n21588) );
  NAND4_X1 U25461 ( .A1(n21591), .A2(n21590), .A3(n21589), .A4(n21588), .ZN(
        n21602) );
  AOI22_X1 U25462 ( .A1(n27439), .A2(\xmem_data[48][0] ), .B1(n3221), .B2(
        \xmem_data[49][0] ), .ZN(n21595) );
  AOI22_X1 U25463 ( .A1(n25448), .A2(\xmem_data[50][0] ), .B1(n23739), .B2(
        \xmem_data[51][0] ), .ZN(n21594) );
  AOI22_X1 U25464 ( .A1(n25449), .A2(\xmem_data[52][0] ), .B1(n20993), .B2(
        \xmem_data[53][0] ), .ZN(n21593) );
  AOI22_X1 U25465 ( .A1(n25451), .A2(\xmem_data[54][0] ), .B1(n23771), .B2(
        \xmem_data[55][0] ), .ZN(n21592) );
  NAND4_X1 U25466 ( .A1(n21595), .A2(n21594), .A3(n21593), .A4(n21592), .ZN(
        n21601) );
  AOI22_X1 U25467 ( .A1(n25422), .A2(\xmem_data[56][0] ), .B1(n22739), .B2(
        \xmem_data[57][0] ), .ZN(n21599) );
  AOI22_X1 U25468 ( .A1(n25457), .A2(\xmem_data[58][0] ), .B1(n30552), .B2(
        \xmem_data[59][0] ), .ZN(n21598) );
  AOI22_X1 U25469 ( .A1(n25459), .A2(\xmem_data[60][0] ), .B1(n25458), .B2(
        \xmem_data[61][0] ), .ZN(n21597) );
  AOI22_X1 U25470 ( .A1(n29437), .A2(\xmem_data[62][0] ), .B1(n25460), .B2(
        \xmem_data[63][0] ), .ZN(n21596) );
  NAND4_X1 U25471 ( .A1(n21599), .A2(n21598), .A3(n21597), .A4(n21596), .ZN(
        n21600) );
  OR4_X1 U25472 ( .A1(n21603), .A2(n21602), .A3(n21601), .A4(n21600), .ZN(
        n21628) );
  AOI22_X1 U25473 ( .A1(n30497), .A2(\xmem_data[8][0] ), .B1(n25359), .B2(
        \xmem_data[9][0] ), .ZN(n21607) );
  AOI22_X1 U25474 ( .A1(n30674), .A2(\xmem_data[10][0] ), .B1(n25388), .B2(
        \xmem_data[11][0] ), .ZN(n21606) );
  AOI22_X1 U25475 ( .A1(n25358), .A2(\xmem_data[12][0] ), .B1(n25357), .B2(
        \xmem_data[13][0] ), .ZN(n21605) );
  AOI22_X1 U25476 ( .A1(n24693), .A2(\xmem_data[14][0] ), .B1(n25360), .B2(
        \xmem_data[15][0] ), .ZN(n21604) );
  AND4_X1 U25477 ( .A1(n21607), .A2(n21606), .A3(n21605), .A4(n21604), .ZN(
        n21615) );
  AOI22_X1 U25478 ( .A1(n25354), .A2(\xmem_data[16][0] ), .B1(n3217), .B2(
        \xmem_data[17][0] ), .ZN(n21614) );
  AOI22_X1 U25479 ( .A1(n3342), .A2(\xmem_data[20][0] ), .B1(n24140), .B2(
        \xmem_data[21][0] ), .ZN(n21608) );
  INV_X1 U25480 ( .A(n21608), .ZN(n21612) );
  AOI22_X1 U25481 ( .A1(n30593), .A2(\xmem_data[18][0] ), .B1(n24695), .B2(
        \xmem_data[19][0] ), .ZN(n21610) );
  NAND2_X1 U25482 ( .A1(n25377), .A2(\xmem_data[22][0] ), .ZN(n21609) );
  NAND2_X1 U25483 ( .A1(n21610), .A2(n21609), .ZN(n21611) );
  NOR2_X1 U25484 ( .A1(n21612), .A2(n21611), .ZN(n21613) );
  NAND3_X1 U25485 ( .A1(n21615), .A2(n21614), .A3(n21613), .ZN(n21626) );
  AOI22_X1 U25486 ( .A1(n27551), .A2(\xmem_data[24][0] ), .B1(n22701), .B2(
        \xmem_data[25][0] ), .ZN(n21619) );
  AOI22_X1 U25487 ( .A1(n29591), .A2(\xmem_data[26][0] ), .B1(n28515), .B2(
        \xmem_data[27][0] ), .ZN(n21618) );
  AOI22_X1 U25488 ( .A1(n29109), .A2(\xmem_data[28][0] ), .B1(n25382), .B2(
        \xmem_data[29][0] ), .ZN(n21617) );
  AOI22_X1 U25489 ( .A1(n29807), .A2(\xmem_data[30][0] ), .B1(n25383), .B2(
        \xmem_data[31][0] ), .ZN(n21616) );
  NAND4_X1 U25490 ( .A1(n21619), .A2(n21618), .A3(n21617), .A4(n21616), .ZN(
        n21625) );
  AOI22_X1 U25491 ( .A1(n25573), .A2(\xmem_data[0][0] ), .B1(n31329), .B2(
        \xmem_data[1][0] ), .ZN(n21623) );
  AOI22_X1 U25492 ( .A1(n28754), .A2(\xmem_data[2][0] ), .B1(n25367), .B2(
        \xmem_data[3][0] ), .ZN(n21622) );
  AOI22_X1 U25493 ( .A1(n3177), .A2(\xmem_data[4][0] ), .B1(n25364), .B2(
        \xmem_data[5][0] ), .ZN(n21621) );
  AOI22_X1 U25494 ( .A1(n30686), .A2(\xmem_data[6][0] ), .B1(n28495), .B2(
        \xmem_data[7][0] ), .ZN(n21620) );
  NAND4_X1 U25495 ( .A1(n21623), .A2(n21622), .A3(n21621), .A4(n21620), .ZN(
        n21624) );
  AOI22_X1 U25496 ( .A1(n23764), .A2(\xmem_data[96][0] ), .B1(n25398), .B2(
        \xmem_data[97][0] ), .ZN(n21632) );
  AOI22_X1 U25497 ( .A1(n25400), .A2(\xmem_data[98][0] ), .B1(n25399), .B2(
        \xmem_data[99][0] ), .ZN(n21631) );
  AOI22_X1 U25498 ( .A1(n27974), .A2(\xmem_data[100][0] ), .B1(n17001), .B2(
        \xmem_data[101][0] ), .ZN(n21630) );
  AOI22_X1 U25499 ( .A1(n25401), .A2(\xmem_data[102][0] ), .B1(n14975), .B2(
        \xmem_data[103][0] ), .ZN(n21629) );
  NAND4_X1 U25500 ( .A1(n21632), .A2(n21631), .A3(n21630), .A4(n21629), .ZN(
        n21648) );
  AOI22_X1 U25501 ( .A1(n3209), .A2(\xmem_data[104][0] ), .B1(n25406), .B2(
        \xmem_data[105][0] ), .ZN(n21636) );
  AOI22_X1 U25502 ( .A1(n25407), .A2(\xmem_data[106][0] ), .B1(n21059), .B2(
        \xmem_data[107][0] ), .ZN(n21635) );
  AOI22_X1 U25503 ( .A1(n25408), .A2(\xmem_data[108][0] ), .B1(n30861), .B2(
        \xmem_data[109][0] ), .ZN(n21634) );
  AOI22_X1 U25504 ( .A1(n3318), .A2(\xmem_data[110][0] ), .B1(n28501), .B2(
        \xmem_data[111][0] ), .ZN(n21633) );
  NAND4_X1 U25505 ( .A1(n21636), .A2(n21635), .A3(n21634), .A4(n21633), .ZN(
        n21647) );
  AOI22_X1 U25506 ( .A1(n25413), .A2(\xmem_data[112][0] ), .B1(n3220), .B2(
        \xmem_data[113][0] ), .ZN(n21640) );
  AOI22_X1 U25507 ( .A1(n25414), .A2(\xmem_data[114][0] ), .B1(n29028), .B2(
        \xmem_data[115][0] ), .ZN(n21639) );
  AOI22_X1 U25508 ( .A1(n25416), .A2(\xmem_data[116][0] ), .B1(n25415), .B2(
        \xmem_data[117][0] ), .ZN(n21638) );
  AOI22_X1 U25509 ( .A1(n25417), .A2(\xmem_data[118][0] ), .B1(n28045), .B2(
        \xmem_data[119][0] ), .ZN(n21637) );
  NAND4_X1 U25510 ( .A1(n21640), .A2(n21639), .A3(n21638), .A4(n21637), .ZN(
        n21646) );
  AOI22_X1 U25511 ( .A1(n25422), .A2(\xmem_data[120][0] ), .B1(n22739), .B2(
        \xmem_data[121][0] ), .ZN(n21644) );
  AOI22_X1 U25512 ( .A1(n25424), .A2(\xmem_data[122][0] ), .B1(n25423), .B2(
        \xmem_data[123][0] ), .ZN(n21643) );
  AOI22_X1 U25513 ( .A1(n25425), .A2(\xmem_data[124][0] ), .B1(n29046), .B2(
        \xmem_data[125][0] ), .ZN(n21642) );
  AOI22_X1 U25514 ( .A1(n29807), .A2(\xmem_data[126][0] ), .B1(n3213), .B2(
        \xmem_data[127][0] ), .ZN(n21641) );
  NAND4_X1 U25515 ( .A1(n21644), .A2(n21643), .A3(n21642), .A4(n21641), .ZN(
        n21645) );
  OR4_X1 U25516 ( .A1(n21648), .A2(n21647), .A3(n21646), .A4(n21645), .ZN(
        n21670) );
  AOI22_X1 U25517 ( .A1(n30949), .A2(\xmem_data[64][0] ), .B1(n25398), .B2(
        \xmem_data[65][0] ), .ZN(n21652) );
  AOI22_X1 U25518 ( .A1(n25400), .A2(\xmem_data[66][0] ), .B1(n25399), .B2(
        \xmem_data[67][0] ), .ZN(n21651) );
  AOI22_X1 U25519 ( .A1(n25521), .A2(\xmem_data[68][0] ), .B1(n27856), .B2(
        \xmem_data[69][0] ), .ZN(n21650) );
  AOI22_X1 U25520 ( .A1(n25401), .A2(\xmem_data[70][0] ), .B1(n14975), .B2(
        \xmem_data[71][0] ), .ZN(n21649) );
  NAND4_X1 U25521 ( .A1(n21652), .A2(n21651), .A3(n21650), .A4(n21649), .ZN(
        n21668) );
  AOI22_X1 U25522 ( .A1(n24572), .A2(\xmem_data[72][0] ), .B1(n25406), .B2(
        \xmem_data[73][0] ), .ZN(n21656) );
  AOI22_X1 U25523 ( .A1(n25407), .A2(\xmem_data[74][0] ), .B1(n21059), .B2(
        \xmem_data[75][0] ), .ZN(n21655) );
  AOI22_X1 U25524 ( .A1(n25408), .A2(\xmem_data[76][0] ), .B1(n28317), .B2(
        \xmem_data[77][0] ), .ZN(n21654) );
  AOI22_X1 U25525 ( .A1(n3318), .A2(\xmem_data[78][0] ), .B1(n25687), .B2(
        \xmem_data[79][0] ), .ZN(n21653) );
  NAND4_X1 U25526 ( .A1(n21656), .A2(n21655), .A3(n21654), .A4(n21653), .ZN(
        n21667) );
  AOI22_X1 U25527 ( .A1(n25413), .A2(\xmem_data[80][0] ), .B1(n3221), .B2(
        \xmem_data[81][0] ), .ZN(n21660) );
  AOI22_X1 U25528 ( .A1(n25414), .A2(\xmem_data[82][0] ), .B1(n20992), .B2(
        \xmem_data[83][0] ), .ZN(n21659) );
  AOI22_X1 U25529 ( .A1(n25416), .A2(\xmem_data[84][0] ), .B1(n25415), .B2(
        \xmem_data[85][0] ), .ZN(n21658) );
  AOI22_X1 U25530 ( .A1(n25417), .A2(\xmem_data[86][0] ), .B1(n30877), .B2(
        \xmem_data[87][0] ), .ZN(n21657) );
  NAND4_X1 U25531 ( .A1(n21660), .A2(n21659), .A3(n21658), .A4(n21657), .ZN(
        n21666) );
  AOI22_X1 U25532 ( .A1(n25422), .A2(\xmem_data[88][0] ), .B1(n30854), .B2(
        \xmem_data[89][0] ), .ZN(n21664) );
  AOI22_X1 U25533 ( .A1(n25424), .A2(\xmem_data[90][0] ), .B1(n25423), .B2(
        \xmem_data[91][0] ), .ZN(n21663) );
  AOI22_X1 U25534 ( .A1(n25425), .A2(\xmem_data[92][0] ), .B1(n20584), .B2(
        \xmem_data[93][0] ), .ZN(n21662) );
  AOI22_X1 U25535 ( .A1(n29008), .A2(\xmem_data[94][0] ), .B1(n24134), .B2(
        \xmem_data[95][0] ), .ZN(n21661) );
  NAND4_X1 U25536 ( .A1(n21664), .A2(n21663), .A3(n21662), .A4(n21661), .ZN(
        n21665) );
  OR4_X1 U25537 ( .A1(n21668), .A2(n21667), .A3(n21666), .A4(n21665), .ZN(
        n21669) );
  AOI22_X1 U25538 ( .A1(n25473), .A2(n21670), .B1(n25471), .B2(n21669), .ZN(
        n21671) );
  XOR2_X1 U25539 ( .A(\fmem_data[30][6] ), .B(\fmem_data[30][7] ), .Z(n21673)
         );
  AOI22_X1 U25540 ( .A1(n30525), .A2(\xmem_data[96][0] ), .B1(n28292), .B2(
        \xmem_data[97][0] ), .ZN(n21678) );
  AOI22_X1 U25541 ( .A1(n28036), .A2(\xmem_data[98][0] ), .B1(n28035), .B2(
        \xmem_data[99][0] ), .ZN(n21677) );
  AOI22_X1 U25542 ( .A1(n28038), .A2(\xmem_data[100][0] ), .B1(n28037), .B2(
        \xmem_data[101][0] ), .ZN(n21676) );
  AOI22_X1 U25543 ( .A1(n28039), .A2(\xmem_data[102][0] ), .B1(n24439), .B2(
        \xmem_data[103][0] ), .ZN(n21675) );
  NAND4_X1 U25544 ( .A1(n21678), .A2(n21677), .A3(n21676), .A4(n21675), .ZN(
        n21694) );
  AOI22_X1 U25545 ( .A1(n28044), .A2(\xmem_data[104][0] ), .B1(n3217), .B2(
        \xmem_data[105][0] ), .ZN(n21682) );
  AOI22_X1 U25546 ( .A1(n24632), .A2(\xmem_data[106][0] ), .B1(n20723), .B2(
        \xmem_data[107][0] ), .ZN(n21681) );
  AOI22_X1 U25547 ( .A1(n24697), .A2(\xmem_data[108][0] ), .B1(n22759), .B2(
        \xmem_data[109][0] ), .ZN(n21680) );
  AOI22_X1 U25548 ( .A1(n20962), .A2(\xmem_data[110][0] ), .B1(n25450), .B2(
        \xmem_data[111][0] ), .ZN(n21679) );
  NAND4_X1 U25549 ( .A1(n21682), .A2(n21681), .A3(n21680), .A4(n21679), .ZN(
        n21693) );
  AOI22_X1 U25550 ( .A1(n28050), .A2(\xmem_data[112][0] ), .B1(n27863), .B2(
        \xmem_data[113][0] ), .ZN(n21686) );
  AOI22_X1 U25551 ( .A1(n28051), .A2(\xmem_data[114][0] ), .B1(n24132), .B2(
        \xmem_data[115][0] ), .ZN(n21685) );
  AOI22_X1 U25552 ( .A1(n28980), .A2(\xmem_data[116][0] ), .B1(n28052), .B2(
        \xmem_data[117][0] ), .ZN(n21684) );
  AOI22_X1 U25553 ( .A1(n30948), .A2(\xmem_data[118][0] ), .B1(n24457), .B2(
        \xmem_data[119][0] ), .ZN(n21683) );
  NAND4_X1 U25554 ( .A1(n21686), .A2(n21685), .A3(n21684), .A4(n21683), .ZN(
        n21692) );
  AOI22_X1 U25555 ( .A1(n28059), .A2(\xmem_data[120][0] ), .B1(n28058), .B2(
        \xmem_data[121][0] ), .ZN(n21690) );
  AOI22_X1 U25556 ( .A1(n16990), .A2(\xmem_data[122][0] ), .B1(n25399), .B2(
        \xmem_data[123][0] ), .ZN(n21689) );
  AOI22_X1 U25557 ( .A1(n28061), .A2(\xmem_data[124][0] ), .B1(n28060), .B2(
        \xmem_data[125][0] ), .ZN(n21688) );
  AOI22_X1 U25558 ( .A1(n30645), .A2(\xmem_data[126][0] ), .B1(n28062), .B2(
        \xmem_data[127][0] ), .ZN(n21687) );
  NAND4_X1 U25559 ( .A1(n21690), .A2(n21689), .A3(n21688), .A4(n21687), .ZN(
        n21691) );
  OR4_X1 U25560 ( .A1(n21694), .A2(n21693), .A3(n21692), .A4(n21691), .ZN(
        n21716) );
  AOI22_X1 U25561 ( .A1(n24166), .A2(\xmem_data[64][0] ), .B1(n28500), .B2(
        \xmem_data[65][0] ), .ZN(n21698) );
  AOI22_X1 U25562 ( .A1(n28036), .A2(\xmem_data[66][0] ), .B1(n28035), .B2(
        \xmem_data[67][0] ), .ZN(n21697) );
  AOI22_X1 U25563 ( .A1(n28038), .A2(\xmem_data[68][0] ), .B1(n28037), .B2(
        \xmem_data[69][0] ), .ZN(n21696) );
  AOI22_X1 U25564 ( .A1(n28039), .A2(\xmem_data[70][0] ), .B1(n28501), .B2(
        \xmem_data[71][0] ), .ZN(n21695) );
  NAND4_X1 U25565 ( .A1(n21698), .A2(n21697), .A3(n21696), .A4(n21695), .ZN(
        n21714) );
  AOI22_X1 U25566 ( .A1(n28044), .A2(\xmem_data[72][0] ), .B1(n3217), .B2(
        \xmem_data[73][0] ), .ZN(n21702) );
  AOI22_X1 U25567 ( .A1(n25448), .A2(\xmem_data[74][0] ), .B1(n22667), .B2(
        \xmem_data[75][0] ), .ZN(n21701) );
  AOI22_X1 U25568 ( .A1(n25449), .A2(\xmem_data[76][0] ), .B1(n30882), .B2(
        \xmem_data[77][0] ), .ZN(n21700) );
  AOI22_X1 U25569 ( .A1(n29762), .A2(\xmem_data[78][0] ), .B1(n25450), .B2(
        \xmem_data[79][0] ), .ZN(n21699) );
  NAND4_X1 U25570 ( .A1(n21702), .A2(n21701), .A3(n21700), .A4(n21699), .ZN(
        n21713) );
  AOI22_X1 U25571 ( .A1(n28050), .A2(\xmem_data[80][0] ), .B1(n27943), .B2(
        \xmem_data[81][0] ), .ZN(n21706) );
  AOI22_X1 U25572 ( .A1(n28051), .A2(\xmem_data[82][0] ), .B1(n31326), .B2(
        \xmem_data[83][0] ), .ZN(n21705) );
  AOI22_X1 U25573 ( .A1(n25425), .A2(\xmem_data[84][0] ), .B1(n28052), .B2(
        \xmem_data[85][0] ), .ZN(n21704) );
  AOI22_X1 U25574 ( .A1(n28752), .A2(\xmem_data[86][0] ), .B1(n3207), .B2(
        \xmem_data[87][0] ), .ZN(n21703) );
  NAND4_X1 U25575 ( .A1(n21706), .A2(n21705), .A3(n21704), .A4(n21703), .ZN(
        n21712) );
  AOI22_X1 U25576 ( .A1(n28059), .A2(\xmem_data[88][0] ), .B1(n28058), .B2(
        \xmem_data[89][0] ), .ZN(n21710) );
  AOI22_X1 U25577 ( .A1(n28781), .A2(\xmem_data[90][0] ), .B1(n25576), .B2(
        \xmem_data[91][0] ), .ZN(n21709) );
  AOI22_X1 U25578 ( .A1(n28061), .A2(\xmem_data[92][0] ), .B1(n28060), .B2(
        \xmem_data[93][0] ), .ZN(n21708) );
  AOI22_X1 U25579 ( .A1(n3307), .A2(\xmem_data[94][0] ), .B1(n28062), .B2(
        \xmem_data[95][0] ), .ZN(n21707) );
  NAND4_X1 U25580 ( .A1(n21710), .A2(n21709), .A3(n21708), .A4(n21707), .ZN(
        n21711) );
  OR4_X1 U25581 ( .A1(n21714), .A2(n21713), .A3(n21712), .A4(n21711), .ZN(
        n21715) );
  AOI22_X1 U25582 ( .A1(n28071), .A2(n21716), .B1(n28033), .B2(n21715), .ZN(
        n21765) );
  AOI22_X1 U25583 ( .A1(n20734), .A2(\xmem_data[32][0] ), .B1(n20488), .B2(
        \xmem_data[33][0] ), .ZN(n21720) );
  AOI22_X1 U25584 ( .A1(n27568), .A2(\xmem_data[34][0] ), .B1(n17050), .B2(
        \xmem_data[35][0] ), .ZN(n21719) );
  AOI22_X1 U25585 ( .A1(n28076), .A2(\xmem_data[36][0] ), .B1(n28075), .B2(
        \xmem_data[37][0] ), .ZN(n21718) );
  AOI22_X1 U25586 ( .A1(n3434), .A2(\xmem_data[38][0] ), .B1(n3247), .B2(
        \xmem_data[39][0] ), .ZN(n21717) );
  NAND4_X1 U25587 ( .A1(n21720), .A2(n21719), .A3(n21718), .A4(n21717), .ZN(
        n21736) );
  AOI22_X1 U25588 ( .A1(n28082), .A2(\xmem_data[40][0] ), .B1(n3220), .B2(
        \xmem_data[41][0] ), .ZN(n21724) );
  AOI22_X1 U25589 ( .A1(n29256), .A2(\xmem_data[42][0] ), .B1(n27869), .B2(
        \xmem_data[43][0] ), .ZN(n21723) );
  AOI22_X1 U25590 ( .A1(n28083), .A2(\xmem_data[44][0] ), .B1(n24564), .B2(
        \xmem_data[45][0] ), .ZN(n21722) );
  AOI22_X1 U25591 ( .A1(n28084), .A2(\xmem_data[46][0] ), .B1(n28007), .B2(
        \xmem_data[47][0] ), .ZN(n21721) );
  NAND4_X1 U25592 ( .A1(n21724), .A2(n21723), .A3(n21722), .A4(n21721), .ZN(
        n21735) );
  AOI22_X1 U25593 ( .A1(n27551), .A2(\xmem_data[48][0] ), .B1(n13475), .B2(
        \xmem_data[49][0] ), .ZN(n21728) );
  AOI22_X1 U25594 ( .A1(n28089), .A2(\xmem_data[50][0] ), .B1(n24212), .B2(
        \xmem_data[51][0] ), .ZN(n21727) );
  AOI22_X1 U25595 ( .A1(n28334), .A2(\xmem_data[52][0] ), .B1(n28090), .B2(
        \xmem_data[53][0] ), .ZN(n21726) );
  AOI22_X1 U25596 ( .A1(n28231), .A2(\xmem_data[54][0] ), .B1(n27989), .B2(
        \xmem_data[55][0] ), .ZN(n21725) );
  NAND4_X1 U25597 ( .A1(n21728), .A2(n21727), .A3(n21726), .A4(n21725), .ZN(
        n21734) );
  AOI22_X1 U25598 ( .A1(n28096), .A2(\xmem_data[56][0] ), .B1(n25398), .B2(
        \xmem_data[57][0] ), .ZN(n21732) );
  AOI22_X1 U25599 ( .A1(n20815), .A2(\xmem_data[58][0] ), .B1(n28097), .B2(
        \xmem_data[59][0] ), .ZN(n21731) );
  AOI22_X1 U25600 ( .A1(n28428), .A2(\xmem_data[60][0] ), .B1(n3372), .B2(
        \xmem_data[61][0] ), .ZN(n21730) );
  AOI22_X1 U25601 ( .A1(n28202), .A2(\xmem_data[62][0] ), .B1(n28098), .B2(
        \xmem_data[63][0] ), .ZN(n21729) );
  NAND4_X1 U25602 ( .A1(n21732), .A2(n21731), .A3(n21730), .A4(n21729), .ZN(
        n21733) );
  OR4_X1 U25603 ( .A1(n21736), .A2(n21735), .A3(n21734), .A4(n21733), .ZN(
        n21737) );
  AOI22_X1 U25604 ( .A1(n25422), .A2(\xmem_data[16][0] ), .B1(n27988), .B2(
        \xmem_data[17][0] ), .ZN(n21741) );
  AOI22_X1 U25605 ( .A1(n17064), .A2(\xmem_data[18][0] ), .B1(n13168), .B2(
        \xmem_data[19][0] ), .ZN(n21740) );
  AOI22_X1 U25606 ( .A1(n16986), .A2(\xmem_data[20][0] ), .B1(n25709), .B2(
        \xmem_data[21][0] ), .ZN(n21739) );
  AOI22_X1 U25607 ( .A1(n30948), .A2(\xmem_data[22][0] ), .B1(n27989), .B2(
        \xmem_data[23][0] ), .ZN(n21738) );
  NAND4_X1 U25608 ( .A1(n21741), .A2(n21740), .A3(n21739), .A4(n21738), .ZN(
        n21755) );
  AOI22_X1 U25609 ( .A1(n20552), .A2(\xmem_data[0][0] ), .B1(n27981), .B2(
        \xmem_data[1][0] ), .ZN(n21745) );
  AOI22_X1 U25610 ( .A1(n29820), .A2(\xmem_data[2][0] ), .B1(n20769), .B2(
        \xmem_data[3][0] ), .ZN(n21744) );
  AOI22_X1 U25611 ( .A1(n25408), .A2(\xmem_data[4][0] ), .B1(n27563), .B2(
        \xmem_data[5][0] ), .ZN(n21743) );
  AOI22_X1 U25612 ( .A1(n3449), .A2(\xmem_data[6][0] ), .B1(n3247), .B2(
        \xmem_data[7][0] ), .ZN(n21742) );
  AND4_X1 U25613 ( .A1(n21745), .A2(n21744), .A3(n21743), .A4(n21742), .ZN(
        n21753) );
  AOI22_X1 U25614 ( .A1(n28355), .A2(\xmem_data[8][0] ), .B1(n3222), .B2(
        \xmem_data[9][0] ), .ZN(n21752) );
  AOI22_X1 U25615 ( .A1(n30883), .A2(\xmem_data[12][0] ), .B1(n27994), .B2(
        \xmem_data[13][0] ), .ZN(n21746) );
  INV_X1 U25616 ( .A(n21746), .ZN(n21750) );
  AOI22_X1 U25617 ( .A1(n29431), .A2(\xmem_data[10][0] ), .B1(n24695), .B2(
        \xmem_data[11][0] ), .ZN(n21748) );
  NAND2_X1 U25618 ( .A1(n30295), .A2(\xmem_data[14][0] ), .ZN(n21747) );
  NAND2_X1 U25619 ( .A1(n21748), .A2(n21747), .ZN(n21749) );
  NOR2_X1 U25620 ( .A1(n21750), .A2(n21749), .ZN(n21751) );
  NAND3_X1 U25621 ( .A1(n21753), .A2(n21752), .A3(n21751), .ZN(n21754) );
  OR2_X1 U25622 ( .A1(n21755), .A2(n21754), .ZN(n21762) );
  AOI22_X1 U25623 ( .A1(n20585), .A2(\xmem_data[24][0] ), .B1(n28492), .B2(
        \xmem_data[25][0] ), .ZN(n21759) );
  AOI22_X1 U25624 ( .A1(n29047), .A2(\xmem_data[26][0] ), .B1(n25367), .B2(
        \xmem_data[27][0] ), .ZN(n21758) );
  AOI22_X1 U25625 ( .A1(n27974), .A2(\xmem_data[28][0] ), .B1(n28429), .B2(
        \xmem_data[29][0] ), .ZN(n21757) );
  AOI22_X1 U25626 ( .A1(n3329), .A2(\xmem_data[30][0] ), .B1(n27975), .B2(
        \xmem_data[31][0] ), .ZN(n21756) );
  NAND4_X1 U25627 ( .A1(n21759), .A2(n21758), .A3(n21757), .A4(n21756), .ZN(
        n21760) );
  OAI21_X1 U25628 ( .B1(n21762), .B2(n21761), .A(n25287), .ZN(n21763) );
  NAND3_X2 U25629 ( .A1(n21765), .A2(n21764), .A3(n21763), .ZN(n36243) );
  AOI22_X1 U25630 ( .A1(n30849), .A2(\xmem_data[120][3] ), .B1(n28291), .B2(
        \xmem_data[121][3] ), .ZN(n21770) );
  AOI22_X1 U25631 ( .A1(n29246), .A2(\xmem_data[122][3] ), .B1(n24622), .B2(
        \xmem_data[123][3] ), .ZN(n21769) );
  AOI22_X1 U25632 ( .A1(n28293), .A2(\xmem_data[124][3] ), .B1(n28292), .B2(
        \xmem_data[125][3] ), .ZN(n21768) );
  AOI22_X1 U25633 ( .A1(n28241), .A2(\xmem_data[126][3] ), .B1(n27567), .B2(
        \xmem_data[127][3] ), .ZN(n21767) );
  NAND4_X1 U25634 ( .A1(n21770), .A2(n21769), .A3(n21768), .A4(n21767), .ZN(
        n21781) );
  AOI22_X1 U25635 ( .A1(n28298), .A2(\xmem_data[112][3] ), .B1(n28517), .B2(
        \xmem_data[113][3] ), .ZN(n21774) );
  AOI22_X1 U25636 ( .A1(n28053), .A2(\xmem_data[114][3] ), .B1(n28299), .B2(
        \xmem_data[115][3] ), .ZN(n21773) );
  AOI22_X1 U25637 ( .A1(n20585), .A2(\xmem_data[116][3] ), .B1(n29048), .B2(
        \xmem_data[117][3] ), .ZN(n21772) );
  AOI22_X1 U25638 ( .A1(n28302), .A2(\xmem_data[118][3] ), .B1(n28301), .B2(
        \xmem_data[119][3] ), .ZN(n21771) );
  NAND4_X1 U25639 ( .A1(n21774), .A2(n21773), .A3(n21772), .A4(n21771), .ZN(
        n21780) );
  AOI22_X1 U25640 ( .A1(n27938), .A2(\xmem_data[104][3] ), .B1(n25415), .B2(
        \xmem_data[105][3] ), .ZN(n21778) );
  AOI22_X1 U25641 ( .A1(n28308), .A2(\xmem_data[106][3] ), .B1(n28307), .B2(
        \xmem_data[107][3] ), .ZN(n21777) );
  AOI22_X1 U25642 ( .A1(n24554), .A2(\xmem_data[108][3] ), .B1(n20982), .B2(
        \xmem_data[109][3] ), .ZN(n21776) );
  AOI22_X1 U25643 ( .A1(n28309), .A2(\xmem_data[110][3] ), .B1(n25605), .B2(
        \xmem_data[111][3] ), .ZN(n21775) );
  NAND4_X1 U25644 ( .A1(n21778), .A2(n21777), .A3(n21776), .A4(n21775), .ZN(
        n21779) );
  OR3_X1 U25645 ( .A1(n21781), .A2(n21780), .A3(n21779), .ZN(n21788) );
  AND2_X1 U25646 ( .A1(n3220), .A2(\xmem_data[101][3] ), .ZN(n21782) );
  AOI21_X1 U25647 ( .B1(n28318), .B2(\xmem_data[100][3] ), .A(n21782), .ZN(
        n21786) );
  AOI22_X1 U25648 ( .A1(n3424), .A2(\xmem_data[98][3] ), .B1(n30589), .B2(
        \xmem_data[99][3] ), .ZN(n21785) );
  AOI22_X1 U25649 ( .A1(n25724), .A2(\xmem_data[96][3] ), .B1(n28317), .B2(
        \xmem_data[97][3] ), .ZN(n21784) );
  AOI22_X1 U25650 ( .A1(n30593), .A2(\xmem_data[102][3] ), .B1(n28319), .B2(
        \xmem_data[103][3] ), .ZN(n21783) );
  NAND4_X1 U25651 ( .A1(n21786), .A2(n21785), .A3(n21784), .A4(n21783), .ZN(
        n21787) );
  OAI21_X1 U25652 ( .B1(n21788), .B2(n21787), .A(n28288), .ZN(n21860) );
  AOI22_X1 U25653 ( .A1(n3325), .A2(\xmem_data[56][3] ), .B1(n25679), .B2(
        \xmem_data[57][3] ), .ZN(n21792) );
  AOI22_X1 U25654 ( .A1(n20732), .A2(\xmem_data[58][3] ), .B1(n25583), .B2(
        \xmem_data[59][3] ), .ZN(n21791) );
  AOI22_X1 U25655 ( .A1(n3179), .A2(\xmem_data[60][3] ), .B1(n28328), .B2(
        \xmem_data[61][3] ), .ZN(n21790) );
  AOI22_X1 U25656 ( .A1(n20985), .A2(\xmem_data[62][3] ), .B1(n28329), .B2(
        \xmem_data[63][3] ), .ZN(n21789) );
  NAND4_X1 U25657 ( .A1(n21792), .A2(n21791), .A3(n21790), .A4(n21789), .ZN(
        n21803) );
  AOI22_X1 U25658 ( .A1(n28334), .A2(\xmem_data[48][3] ), .B1(n20584), .B2(
        \xmem_data[49][3] ), .ZN(n21796) );
  AOI22_X1 U25659 ( .A1(n28336), .A2(\xmem_data[50][3] ), .B1(n28335), .B2(
        \xmem_data[51][3] ), .ZN(n21795) );
  AOI22_X1 U25660 ( .A1(n28337), .A2(\xmem_data[52][3] ), .B1(n28492), .B2(
        \xmem_data[53][3] ), .ZN(n21794) );
  AOI22_X1 U25661 ( .A1(n23722), .A2(\xmem_data[54][3] ), .B1(n24221), .B2(
        \xmem_data[55][3] ), .ZN(n21793) );
  NAND4_X1 U25662 ( .A1(n21796), .A2(n21795), .A3(n21794), .A4(n21793), .ZN(
        n21802) );
  AOI22_X1 U25663 ( .A1(n24438), .A2(\xmem_data[40][3] ), .B1(n28342), .B2(
        \xmem_data[41][3] ), .ZN(n21800) );
  AOI22_X1 U25664 ( .A1(n28344), .A2(\xmem_data[42][3] ), .B1(n25450), .B2(
        \xmem_data[43][3] ), .ZN(n21799) );
  AOI22_X1 U25665 ( .A1(n25422), .A2(\xmem_data[44][3] ), .B1(n27863), .B2(
        \xmem_data[45][3] ), .ZN(n21798) );
  AOI22_X1 U25666 ( .A1(n28346), .A2(\xmem_data[46][3] ), .B1(n28345), .B2(
        \xmem_data[47][3] ), .ZN(n21797) );
  NAND4_X1 U25667 ( .A1(n21800), .A2(n21799), .A3(n21798), .A4(n21797), .ZN(
        n21801) );
  OR3_X1 U25668 ( .A1(n21803), .A2(n21802), .A3(n21801), .ZN(n21810) );
  AND2_X1 U25669 ( .A1(n3220), .A2(\xmem_data[37][3] ), .ZN(n21804) );
  AOI21_X1 U25670 ( .B1(n28355), .B2(\xmem_data[36][3] ), .A(n21804), .ZN(
        n21808) );
  AOI22_X1 U25671 ( .A1(n30864), .A2(\xmem_data[34][3] ), .B1(n3247), .B2(
        \xmem_data[35][3] ), .ZN(n21807) );
  AOI22_X1 U25672 ( .A1(n28354), .A2(\xmem_data[32][3] ), .B1(n28075), .B2(
        \xmem_data[33][3] ), .ZN(n21806) );
  AOI22_X1 U25673 ( .A1(n24533), .A2(\xmem_data[38][3] ), .B1(n28356), .B2(
        \xmem_data[39][3] ), .ZN(n21805) );
  NAND4_X1 U25674 ( .A1(n21808), .A2(n21807), .A3(n21806), .A4(n21805), .ZN(
        n21809) );
  OAI21_X1 U25675 ( .B1(n21810), .B2(n21809), .A(n28361), .ZN(n21859) );
  AND2_X1 U25676 ( .A1(n3218), .A2(\xmem_data[69][3] ), .ZN(n21811) );
  AOI21_X1 U25677 ( .B1(n28318), .B2(\xmem_data[68][3] ), .A(n21811), .ZN(
        n21818) );
  AOI22_X1 U25678 ( .A1(n17030), .A2(\xmem_data[64][3] ), .B1(n28317), .B2(
        \xmem_data[65][3] ), .ZN(n21817) );
  AOI22_X1 U25679 ( .A1(n21067), .A2(\xmem_data[70][3] ), .B1(n28319), .B2(
        \xmem_data[71][3] ), .ZN(n21812) );
  INV_X1 U25680 ( .A(n21812), .ZN(n21815) );
  AOI22_X1 U25681 ( .A1(n3245), .A2(\xmem_data[66][3] ), .B1(n28501), .B2(
        \xmem_data[67][3] ), .ZN(n21813) );
  INV_X1 U25682 ( .A(n21813), .ZN(n21814) );
  NOR2_X1 U25683 ( .A1(n21815), .A2(n21814), .ZN(n21816) );
  NAND3_X1 U25684 ( .A1(n21818), .A2(n21817), .A3(n21816), .ZN(n21834) );
  AOI22_X1 U25685 ( .A1(n28298), .A2(\xmem_data[80][3] ), .B1(n29046), .B2(
        \xmem_data[81][3] ), .ZN(n21822) );
  AOI22_X1 U25686 ( .A1(n20939), .A2(\xmem_data[82][3] ), .B1(n28299), .B2(
        \xmem_data[83][3] ), .ZN(n21821) );
  AOI22_X1 U25687 ( .A1(n21007), .A2(\xmem_data[84][3] ), .B1(n25398), .B2(
        \xmem_data[85][3] ), .ZN(n21820) );
  AOI22_X1 U25688 ( .A1(n28302), .A2(\xmem_data[86][3] ), .B1(n28301), .B2(
        \xmem_data[87][3] ), .ZN(n21819) );
  NAND4_X1 U25689 ( .A1(n21822), .A2(n21821), .A3(n21820), .A4(n21819), .ZN(
        n21833) );
  AOI22_X1 U25690 ( .A1(n25617), .A2(\xmem_data[72][3] ), .B1(n20806), .B2(
        \xmem_data[73][3] ), .ZN(n21826) );
  AOI22_X1 U25691 ( .A1(n28308), .A2(\xmem_data[74][3] ), .B1(n28307), .B2(
        \xmem_data[75][3] ), .ZN(n21825) );
  AOI22_X1 U25692 ( .A1(n20809), .A2(\xmem_data[76][3] ), .B1(n24590), .B2(
        \xmem_data[77][3] ), .ZN(n21824) );
  AOI22_X1 U25693 ( .A1(n28309), .A2(\xmem_data[78][3] ), .B1(n28416), .B2(
        \xmem_data[79][3] ), .ZN(n21823) );
  NAND4_X1 U25694 ( .A1(n21826), .A2(n21825), .A3(n21824), .A4(n21823), .ZN(
        n21832) );
  AOI22_X1 U25695 ( .A1(n25632), .A2(\xmem_data[88][3] ), .B1(n28291), .B2(
        \xmem_data[89][3] ), .ZN(n21830) );
  AOI22_X1 U25696 ( .A1(n23724), .A2(\xmem_data[90][3] ), .B1(n27525), .B2(
        \xmem_data[91][3] ), .ZN(n21829) );
  AOI22_X1 U25697 ( .A1(n28293), .A2(\xmem_data[92][3] ), .B1(n28292), .B2(
        \xmem_data[93][3] ), .ZN(n21828) );
  AOI22_X1 U25698 ( .A1(n17051), .A2(\xmem_data[94][3] ), .B1(n24122), .B2(
        \xmem_data[95][3] ), .ZN(n21827) );
  NAND4_X1 U25699 ( .A1(n21830), .A2(n21829), .A3(n21828), .A4(n21827), .ZN(
        n21831) );
  OR4_X1 U25700 ( .A1(n21834), .A2(n21833), .A3(n21832), .A4(n21831), .ZN(
        n21835) );
  NAND2_X1 U25701 ( .A1(n21835), .A2(n28324), .ZN(n21858) );
  AOI22_X1 U25702 ( .A1(n3380), .A2(\xmem_data[0][3] ), .B1(n28366), .B2(
        \xmem_data[1][3] ), .ZN(n21839) );
  AOI22_X1 U25703 ( .A1(n3306), .A2(\xmem_data[2][3] ), .B1(n30589), .B2(
        \xmem_data[3][3] ), .ZN(n21838) );
  AOI22_X1 U25704 ( .A1(n28364), .A2(\xmem_data[4][3] ), .B1(n3219), .B2(
        \xmem_data[5][3] ), .ZN(n21837) );
  AOI22_X1 U25705 ( .A1(n28367), .A2(\xmem_data[6][3] ), .B1(n31367), .B2(
        \xmem_data[7][3] ), .ZN(n21836) );
  NAND4_X1 U25706 ( .A1(n21839), .A2(n21838), .A3(n21837), .A4(n21836), .ZN(
        n21855) );
  AOI22_X1 U25707 ( .A1(n28385), .A2(\xmem_data[24][3] ), .B1(n30598), .B2(
        \xmem_data[25][3] ), .ZN(n21843) );
  AOI22_X1 U25708 ( .A1(n30686), .A2(\xmem_data[26][3] ), .B1(n29245), .B2(
        \xmem_data[27][3] ), .ZN(n21842) );
  AOI22_X1 U25709 ( .A1(n24685), .A2(\xmem_data[28][3] ), .B1(n28468), .B2(
        \xmem_data[29][3] ), .ZN(n21841) );
  AOI22_X1 U25710 ( .A1(n30901), .A2(\xmem_data[30][3] ), .B1(n29248), .B2(
        \xmem_data[31][3] ), .ZN(n21840) );
  NAND4_X1 U25711 ( .A1(n21843), .A2(n21842), .A3(n21841), .A4(n21840), .ZN(
        n21854) );
  AOI22_X1 U25712 ( .A1(n28980), .A2(\xmem_data[16][3] ), .B1(n27912), .B2(
        \xmem_data[17][3] ), .ZN(n21847) );
  AOI22_X1 U25713 ( .A1(n25672), .A2(\xmem_data[18][3] ), .B1(n20586), .B2(
        \xmem_data[19][3] ), .ZN(n21846) );
  AOI22_X1 U25714 ( .A1(n28059), .A2(\xmem_data[20][3] ), .B1(n27518), .B2(
        \xmem_data[21][3] ), .ZN(n21845) );
  AOI22_X1 U25715 ( .A1(n20730), .A2(\xmem_data[22][3] ), .B1(n28380), .B2(
        \xmem_data[23][3] ), .ZN(n21844) );
  NAND4_X1 U25716 ( .A1(n21847), .A2(n21846), .A3(n21845), .A4(n21844), .ZN(
        n21853) );
  AOI22_X1 U25717 ( .A1(n29257), .A2(\xmem_data[8][3] ), .B1(n28372), .B2(
        \xmem_data[9][3] ), .ZN(n21851) );
  AOI22_X1 U25718 ( .A1(n3280), .A2(\xmem_data[10][3] ), .B1(n30877), .B2(
        \xmem_data[11][3] ), .ZN(n21850) );
  AOI22_X1 U25719 ( .A1(n28374), .A2(\xmem_data[12][3] ), .B1(n20546), .B2(
        \xmem_data[13][3] ), .ZN(n21849) );
  AOI22_X1 U25720 ( .A1(n25424), .A2(\xmem_data[14][3] ), .B1(n28375), .B2(
        \xmem_data[15][3] ), .ZN(n21848) );
  NAND4_X1 U25721 ( .A1(n21851), .A2(n21850), .A3(n21849), .A4(n21848), .ZN(
        n21852) );
  OR4_X1 U25722 ( .A1(n21855), .A2(n21854), .A3(n21853), .A4(n21852), .ZN(
        n21856) );
  NAND2_X1 U25723 ( .A1(n21856), .A2(n28395), .ZN(n21857) );
  NAND4_X1 U25724 ( .A1(n21860), .A2(n21859), .A3(n21858), .A4(n21857), .ZN(
        n32283) );
  XNOR2_X1 U25725 ( .A(n32283), .B(\fmem_data[18][5] ), .ZN(n27327) );
  AOI22_X1 U25726 ( .A1(n28355), .A2(\xmem_data[36][4] ), .B1(n3217), .B2(
        \xmem_data[37][4] ), .ZN(n21864) );
  AOI22_X1 U25727 ( .A1(n3318), .A2(\xmem_data[34][4] ), .B1(n22753), .B2(
        \xmem_data[35][4] ), .ZN(n21863) );
  AOI22_X1 U25728 ( .A1(n28354), .A2(\xmem_data[32][4] ), .B1(n20489), .B2(
        \xmem_data[33][4] ), .ZN(n21862) );
  AOI22_X1 U25729 ( .A1(n25693), .A2(\xmem_data[38][4] ), .B1(n28356), .B2(
        \xmem_data[39][4] ), .ZN(n21861) );
  NAND4_X1 U25730 ( .A1(n21864), .A2(n21863), .A3(n21862), .A4(n21861), .ZN(
        n21881) );
  AOI22_X1 U25731 ( .A1(n25632), .A2(\xmem_data[56][4] ), .B1(n21051), .B2(
        \xmem_data[57][4] ), .ZN(n21868) );
  AOI22_X1 U25732 ( .A1(n17004), .A2(\xmem_data[58][4] ), .B1(n24223), .B2(
        \xmem_data[59][4] ), .ZN(n21867) );
  AOI22_X1 U25733 ( .A1(n3179), .A2(\xmem_data[60][4] ), .B1(n28328), .B2(
        \xmem_data[61][4] ), .ZN(n21866) );
  AOI22_X1 U25734 ( .A1(n30901), .A2(\xmem_data[62][4] ), .B1(n28329), .B2(
        \xmem_data[63][4] ), .ZN(n21865) );
  NAND4_X1 U25735 ( .A1(n21868), .A2(n21867), .A3(n21866), .A4(n21865), .ZN(
        n21879) );
  AOI22_X1 U25736 ( .A1(n28334), .A2(\xmem_data[48][4] ), .B1(n14999), .B2(
        \xmem_data[49][4] ), .ZN(n21872) );
  AOI22_X1 U25737 ( .A1(n28336), .A2(\xmem_data[50][4] ), .B1(n28335), .B2(
        \xmem_data[51][4] ), .ZN(n21871) );
  AOI22_X1 U25738 ( .A1(n28337), .A2(\xmem_data[52][4] ), .B1(n29316), .B2(
        \xmem_data[53][4] ), .ZN(n21870) );
  AOI22_X1 U25739 ( .A1(n22717), .A2(\xmem_data[54][4] ), .B1(n27523), .B2(
        \xmem_data[55][4] ), .ZN(n21869) );
  NAND4_X1 U25740 ( .A1(n21872), .A2(n21871), .A3(n21870), .A4(n21869), .ZN(
        n21878) );
  AOI22_X1 U25741 ( .A1(n17010), .A2(\xmem_data[40][4] ), .B1(n28342), .B2(
        \xmem_data[41][4] ), .ZN(n21876) );
  AOI22_X1 U25742 ( .A1(n28344), .A2(\xmem_data[42][4] ), .B1(n28007), .B2(
        \xmem_data[43][4] ), .ZN(n21875) );
  AOI22_X1 U25743 ( .A1(n24554), .A2(\xmem_data[44][4] ), .B1(n24158), .B2(
        \xmem_data[45][4] ), .ZN(n21874) );
  AOI22_X1 U25744 ( .A1(n28346), .A2(\xmem_data[46][4] ), .B1(n28345), .B2(
        \xmem_data[47][4] ), .ZN(n21873) );
  NAND4_X1 U25745 ( .A1(n21876), .A2(n21875), .A3(n21874), .A4(n21873), .ZN(
        n21877) );
  OR3_X1 U25746 ( .A1(n21879), .A2(n21878), .A3(n21877), .ZN(n21880) );
  OAI21_X1 U25747 ( .B1(n21881), .B2(n21880), .A(n28361), .ZN(n21952) );
  AOI22_X1 U25748 ( .A1(n28318), .A2(\xmem_data[100][4] ), .B1(n3218), .B2(
        \xmem_data[101][4] ), .ZN(n21885) );
  AOI22_X1 U25749 ( .A1(n3424), .A2(\xmem_data[98][4] ), .B1(n27437), .B2(
        \xmem_data[99][4] ), .ZN(n21884) );
  AOI22_X1 U25750 ( .A1(n27925), .A2(\xmem_data[96][4] ), .B1(n28317), .B2(
        \xmem_data[97][4] ), .ZN(n21883) );
  AOI22_X1 U25751 ( .A1(n23740), .A2(\xmem_data[102][4] ), .B1(n28319), .B2(
        \xmem_data[103][4] ), .ZN(n21882) );
  NAND4_X1 U25752 ( .A1(n21885), .A2(n21884), .A3(n21883), .A4(n21882), .ZN(
        n21902) );
  AOI22_X1 U25753 ( .A1(n3326), .A2(\xmem_data[120][4] ), .B1(n28291), .B2(
        \xmem_data[121][4] ), .ZN(n21889) );
  AOI22_X1 U25754 ( .A1(n31315), .A2(\xmem_data[122][4] ), .B1(n31314), .B2(
        \xmem_data[123][4] ), .ZN(n21888) );
  AOI22_X1 U25755 ( .A1(n28293), .A2(\xmem_data[124][4] ), .B1(n28292), .B2(
        \xmem_data[125][4] ), .ZN(n21887) );
  AOI22_X1 U25756 ( .A1(n29383), .A2(\xmem_data[126][4] ), .B1(n24524), .B2(
        \xmem_data[127][4] ), .ZN(n21886) );
  NAND4_X1 U25757 ( .A1(n21889), .A2(n21888), .A3(n21887), .A4(n21886), .ZN(
        n21900) );
  AOI22_X1 U25758 ( .A1(n28298), .A2(\xmem_data[112][4] ), .B1(n28517), .B2(
        \xmem_data[113][4] ), .ZN(n21893) );
  AOI22_X1 U25759 ( .A1(n29008), .A2(\xmem_data[114][4] ), .B1(n28299), .B2(
        \xmem_data[115][4] ), .ZN(n21892) );
  AOI22_X1 U25760 ( .A1(n23717), .A2(\xmem_data[116][4] ), .B1(n29316), .B2(
        \xmem_data[117][4] ), .ZN(n21891) );
  AOI22_X1 U25761 ( .A1(n28302), .A2(\xmem_data[118][4] ), .B1(n28301), .B2(
        \xmem_data[119][4] ), .ZN(n21890) );
  NAND4_X1 U25762 ( .A1(n21893), .A2(n21892), .A3(n21891), .A4(n21890), .ZN(
        n21899) );
  AOI22_X1 U25763 ( .A1(n28083), .A2(\xmem_data[104][4] ), .B1(n27550), .B2(
        \xmem_data[105][4] ), .ZN(n21897) );
  AOI22_X1 U25764 ( .A1(n28308), .A2(\xmem_data[106][4] ), .B1(n28307), .B2(
        \xmem_data[107][4] ), .ZN(n21896) );
  AOI22_X1 U25765 ( .A1(n27447), .A2(\xmem_data[108][4] ), .B1(n29180), .B2(
        \xmem_data[109][4] ), .ZN(n21895) );
  AOI22_X1 U25766 ( .A1(n28309), .A2(\xmem_data[110][4] ), .B1(n28416), .B2(
        \xmem_data[111][4] ), .ZN(n21894) );
  NAND4_X1 U25767 ( .A1(n21897), .A2(n21896), .A3(n21895), .A4(n21894), .ZN(
        n21898) );
  OR3_X1 U25768 ( .A1(n21900), .A2(n21899), .A3(n21898), .ZN(n21901) );
  OAI21_X1 U25769 ( .B1(n21902), .B2(n21901), .A(n28288), .ZN(n21951) );
  AOI22_X1 U25770 ( .A1(n3178), .A2(\xmem_data[88][4] ), .B1(n3372), .B2(
        \xmem_data[89][4] ), .ZN(n21906) );
  AOI22_X1 U25771 ( .A1(n20732), .A2(\xmem_data[90][4] ), .B1(n31362), .B2(
        \xmem_data[91][4] ), .ZN(n21905) );
  AOI22_X1 U25772 ( .A1(n3179), .A2(\xmem_data[92][4] ), .B1(n28328), .B2(
        \xmem_data[93][4] ), .ZN(n21904) );
  AOI22_X1 U25773 ( .A1(n27498), .A2(\xmem_data[94][4] ), .B1(n28329), .B2(
        \xmem_data[95][4] ), .ZN(n21903) );
  NAND4_X1 U25774 ( .A1(n21903), .A2(n21905), .A3(n21904), .A4(n21906), .ZN(
        n21917) );
  AOI22_X1 U25775 ( .A1(n28334), .A2(\xmem_data[80][4] ), .B1(n25709), .B2(
        \xmem_data[81][4] ), .ZN(n21910) );
  AOI22_X1 U25776 ( .A1(n28336), .A2(\xmem_data[82][4] ), .B1(n28335), .B2(
        \xmem_data[83][4] ), .ZN(n21909) );
  AOI22_X1 U25777 ( .A1(n28337), .A2(\xmem_data[84][4] ), .B1(n31270), .B2(
        \xmem_data[85][4] ), .ZN(n21908) );
  AOI22_X1 U25778 ( .A1(n25678), .A2(\xmem_data[86][4] ), .B1(n29318), .B2(
        \xmem_data[87][4] ), .ZN(n21907) );
  NAND4_X1 U25779 ( .A1(n21910), .A2(n21909), .A3(n21908), .A4(n21907), .ZN(
        n21916) );
  AOI22_X1 U25780 ( .A1(n20994), .A2(\xmem_data[72][4] ), .B1(n28342), .B2(
        \xmem_data[73][4] ), .ZN(n21914) );
  AOI22_X1 U25781 ( .A1(n28344), .A2(\xmem_data[74][4] ), .B1(n27547), .B2(
        \xmem_data[75][4] ), .ZN(n21913) );
  AOI22_X1 U25782 ( .A1(n27447), .A2(\xmem_data[76][4] ), .B1(n28373), .B2(
        \xmem_data[77][4] ), .ZN(n21912) );
  AOI22_X1 U25783 ( .A1(n28346), .A2(\xmem_data[78][4] ), .B1(n28345), .B2(
        \xmem_data[79][4] ), .ZN(n21911) );
  NAND4_X1 U25784 ( .A1(n21914), .A2(n21913), .A3(n21912), .A4(n21911), .ZN(
        n21915) );
  OR3_X1 U25785 ( .A1(n21917), .A2(n21916), .A3(n21915), .ZN(n21927) );
  AND2_X1 U25786 ( .A1(n3220), .A2(\xmem_data[69][4] ), .ZN(n21918) );
  AOI21_X1 U25787 ( .B1(n28355), .B2(\xmem_data[68][4] ), .A(n21918), .ZN(
        n21925) );
  AOI22_X1 U25788 ( .A1(n28354), .A2(\xmem_data[64][4] ), .B1(n30571), .B2(
        \xmem_data[65][4] ), .ZN(n21924) );
  AOI22_X1 U25789 ( .A1(n25612), .A2(\xmem_data[70][4] ), .B1(n28356), .B2(
        \xmem_data[71][4] ), .ZN(n21919) );
  INV_X1 U25790 ( .A(n21919), .ZN(n21922) );
  AOI22_X1 U25791 ( .A1(n16980), .A2(\xmem_data[66][4] ), .B1(n29286), .B2(
        \xmem_data[67][4] ), .ZN(n21920) );
  INV_X1 U25792 ( .A(n21920), .ZN(n21921) );
  NOR2_X1 U25793 ( .A1(n21922), .A2(n21921), .ZN(n21923) );
  NAND3_X1 U25794 ( .A1(n21925), .A2(n21924), .A3(n21923), .ZN(n21926) );
  OAI21_X1 U25795 ( .B1(n21927), .B2(n21926), .A(n28324), .ZN(n21950) );
  AOI22_X1 U25796 ( .A1(n28364), .A2(\xmem_data[4][4] ), .B1(n3218), .B2(
        \xmem_data[5][4] ), .ZN(n21931) );
  AOI22_X1 U25797 ( .A1(n3306), .A2(\xmem_data[2][4] ), .B1(n24439), .B2(
        \xmem_data[3][4] ), .ZN(n21930) );
  AOI22_X1 U25798 ( .A1(n27500), .A2(\xmem_data[0][4] ), .B1(n28366), .B2(
        \xmem_data[1][4] ), .ZN(n21929) );
  AOI22_X1 U25799 ( .A1(n28367), .A2(\xmem_data[6][4] ), .B1(n29255), .B2(
        \xmem_data[7][4] ), .ZN(n21928) );
  NAND4_X1 U25800 ( .A1(n21931), .A2(n21930), .A3(n21929), .A4(n21928), .ZN(
        n21947) );
  AOI22_X1 U25801 ( .A1(n28385), .A2(\xmem_data[24][4] ), .B1(n20506), .B2(
        \xmem_data[25][4] ), .ZN(n21935) );
  AOI22_X1 U25802 ( .A1(n29324), .A2(\xmem_data[26][4] ), .B1(n24622), .B2(
        \xmem_data[27][4] ), .ZN(n21934) );
  AOI22_X1 U25803 ( .A1(n24467), .A2(\xmem_data[28][4] ), .B1(n11008), .B2(
        \xmem_data[29][4] ), .ZN(n21933) );
  AOI22_X1 U25804 ( .A1(n30901), .A2(\xmem_data[30][4] ), .B1(n24122), .B2(
        \xmem_data[31][4] ), .ZN(n21932) );
  NAND4_X1 U25805 ( .A1(n21935), .A2(n21934), .A3(n21933), .A4(n21932), .ZN(
        n21946) );
  AOI22_X1 U25806 ( .A1(n20541), .A2(\xmem_data[16][4] ), .B1(n25458), .B2(
        \xmem_data[17][4] ), .ZN(n21939) );
  AOI22_X1 U25807 ( .A1(n3465), .A2(\xmem_data[18][4] ), .B1(n28299), .B2(
        \xmem_data[19][4] ), .ZN(n21938) );
  AOI22_X1 U25808 ( .A1(n24708), .A2(\xmem_data[20][4] ), .B1(n25677), .B2(
        \xmem_data[21][4] ), .ZN(n21937) );
  AOI22_X1 U25809 ( .A1(n30872), .A2(\xmem_data[22][4] ), .B1(n28380), .B2(
        \xmem_data[23][4] ), .ZN(n21936) );
  NAND4_X1 U25810 ( .A1(n21939), .A2(n21938), .A3(n21937), .A4(n21936), .ZN(
        n21945) );
  AOI22_X1 U25811 ( .A1(n20994), .A2(\xmem_data[8][4] ), .B1(n28372), .B2(
        \xmem_data[9][4] ), .ZN(n21943) );
  AOI22_X1 U25812 ( .A1(n25451), .A2(\xmem_data[10][4] ), .B1(n28510), .B2(
        \xmem_data[11][4] ), .ZN(n21942) );
  AOI22_X1 U25813 ( .A1(n28374), .A2(\xmem_data[12][4] ), .B1(n25456), .B2(
        \xmem_data[13][4] ), .ZN(n21941) );
  AOI22_X1 U25814 ( .A1(n20587), .A2(\xmem_data[14][4] ), .B1(n28375), .B2(
        \xmem_data[15][4] ), .ZN(n21940) );
  NAND4_X1 U25815 ( .A1(n21943), .A2(n21942), .A3(n21941), .A4(n21940), .ZN(
        n21944) );
  OR4_X1 U25816 ( .A1(n21947), .A2(n21946), .A3(n21945), .A4(n21944), .ZN(
        n21948) );
  NAND2_X1 U25817 ( .A1(n21948), .A2(n28395), .ZN(n21949) );
  XNOR2_X1 U25818 ( .A(n31383), .B(\fmem_data[18][5] ), .ZN(n33033) );
  XNOR2_X1 U25819 ( .A(n32163), .B(\fmem_data[26][3] ), .ZN(n26151) );
  XNOR2_X1 U25820 ( .A(n31670), .B(\fmem_data[26][3] ), .ZN(n32020) );
  OAI22_X1 U25821 ( .A1(n26151), .A2(n32779), .B1(n32020), .B2(n32780), .ZN(
        n34237) );
  AOI22_X1 U25822 ( .A1(n28427), .A2(\xmem_data[104][1] ), .B1(n22682), .B2(
        \xmem_data[105][1] ), .ZN(n21957) );
  AOI22_X1 U25823 ( .A1(n27950), .A2(\xmem_data[106][1] ), .B1(n22683), .B2(
        \xmem_data[107][1] ), .ZN(n21956) );
  AOI22_X1 U25824 ( .A1(n25581), .A2(\xmem_data[108][1] ), .B1(n3302), .B2(
        \xmem_data[109][1] ), .ZN(n21955) );
  AOI22_X1 U25825 ( .A1(n22685), .A2(\xmem_data[110][1] ), .B1(n22684), .B2(
        \xmem_data[111][1] ), .ZN(n21954) );
  NAND4_X1 U25826 ( .A1(n21957), .A2(n21956), .A3(n21955), .A4(n21954), .ZN(
        n21961) );
  AND2_X1 U25827 ( .A1(n14983), .A2(\xmem_data[118][1] ), .ZN(n21958) );
  AOI21_X1 U25828 ( .B1(n28364), .B2(\xmem_data[119][1] ), .A(n21958), .ZN(
        n21959) );
  INV_X1 U25829 ( .A(n21959), .ZN(n21960) );
  NOR2_X1 U25830 ( .A1(n21961), .A2(n21960), .ZN(n21979) );
  AOI22_X1 U25831 ( .A1(n23781), .A2(\xmem_data[112][1] ), .B1(n25684), .B2(
        \xmem_data[113][1] ), .ZN(n21978) );
  AOI22_X1 U25832 ( .A1(n28415), .A2(\xmem_data[96][1] ), .B1(n27453), .B2(
        \xmem_data[97][1] ), .ZN(n21965) );
  AOI22_X1 U25833 ( .A1(n22675), .A2(\xmem_data[98][1] ), .B1(n28334), .B2(
        \xmem_data[99][1] ), .ZN(n21964) );
  AOI22_X1 U25834 ( .A1(n22674), .A2(\xmem_data[100][1] ), .B1(n29605), .B2(
        \xmem_data[101][1] ), .ZN(n21963) );
  AOI22_X1 U25835 ( .A1(n22677), .A2(\xmem_data[102][1] ), .B1(n22676), .B2(
        \xmem_data[103][1] ), .ZN(n21962) );
  NAND4_X1 U25836 ( .A1(n21965), .A2(n21964), .A3(n21963), .A4(n21962), .ZN(
        n21968) );
  AOI22_X1 U25837 ( .A1(n28317), .A2(\xmem_data[116][1] ), .B1(n3424), .B2(
        \xmem_data[117][1] ), .ZN(n21966) );
  INV_X1 U25838 ( .A(n21966), .ZN(n21967) );
  NOR2_X1 U25839 ( .A1(n21968), .A2(n21967), .ZN(n21977) );
  AOI22_X1 U25840 ( .A1(n3219), .A2(\xmem_data[120][1] ), .B1(n28137), .B2(
        \xmem_data[121][1] ), .ZN(n21972) );
  AOI22_X1 U25841 ( .A1(n22667), .A2(\xmem_data[122][1] ), .B1(n22666), .B2(
        \xmem_data[123][1] ), .ZN(n21971) );
  AOI22_X1 U25842 ( .A1(n22669), .A2(\xmem_data[124][1] ), .B1(n22668), .B2(
        \xmem_data[125][1] ), .ZN(n21970) );
  AOI22_X1 U25843 ( .A1(n29103), .A2(\xmem_data[126][1] ), .B1(n23813), .B2(
        \xmem_data[127][1] ), .ZN(n21969) );
  NAND4_X1 U25844 ( .A1(n21972), .A2(n21971), .A3(n21970), .A4(n21969), .ZN(
        n21975) );
  AOI22_X1 U25845 ( .A1(n29125), .A2(\xmem_data[114][1] ), .B1(n27564), .B2(
        \xmem_data[115][1] ), .ZN(n21973) );
  INV_X1 U25846 ( .A(n21973), .ZN(n21974) );
  NOR2_X1 U25847 ( .A1(n21975), .A2(n21974), .ZN(n21976) );
  NAND4_X1 U25848 ( .A1(n21979), .A2(n21978), .A3(n21977), .A4(n21976), .ZN(
        n21980) );
  NAND2_X1 U25849 ( .A1(n21980), .A2(n22698), .ZN(n22054) );
  AOI22_X1 U25850 ( .A1(n22718), .A2(\xmem_data[40][1] ), .B1(n22717), .B2(
        \xmem_data[41][1] ), .ZN(n21984) );
  AOI22_X1 U25851 ( .A1(n30545), .A2(\xmem_data[42][1] ), .B1(n28493), .B2(
        \xmem_data[43][1] ), .ZN(n21983) );
  AOI22_X1 U25852 ( .A1(n28060), .A2(\xmem_data[44][1] ), .B1(n3338), .B2(
        \xmem_data[45][1] ), .ZN(n21982) );
  AOI22_X1 U25853 ( .A1(n25583), .A2(\xmem_data[46][1] ), .B1(n22719), .B2(
        \xmem_data[47][1] ), .ZN(n21981) );
  AOI22_X1 U25854 ( .A1(n31256), .A2(\xmem_data[48][1] ), .B1(n29725), .B2(
        \xmem_data[49][1] ), .ZN(n21986) );
  AOI22_X1 U25855 ( .A1(n20711), .A2(\xmem_data[54][1] ), .B1(n30906), .B2(
        \xmem_data[55][1] ), .ZN(n21985) );
  AOI22_X1 U25856 ( .A1(n22701), .A2(\xmem_data[32][1] ), .B1(n29179), .B2(
        \xmem_data[33][1] ), .ZN(n21990) );
  AOI22_X1 U25857 ( .A1(n22702), .A2(\xmem_data[34][1] ), .B1(n16986), .B2(
        \xmem_data[35][1] ), .ZN(n21989) );
  AOI22_X1 U25858 ( .A1(n22703), .A2(\xmem_data[36][1] ), .B1(n29396), .B2(
        \xmem_data[37][1] ), .ZN(n21988) );
  AOI22_X1 U25859 ( .A1(n28993), .A2(\xmem_data[38][1] ), .B1(n28096), .B2(
        \xmem_data[39][1] ), .ZN(n21987) );
  AOI22_X1 U25860 ( .A1(n22727), .A2(\xmem_data[50][1] ), .B1(n28076), .B2(
        \xmem_data[51][1] ), .ZN(n21996) );
  AOI22_X1 U25861 ( .A1(n3222), .A2(\xmem_data[56][1] ), .B1(n22708), .B2(
        \xmem_data[57][1] ), .ZN(n21994) );
  AOI22_X1 U25862 ( .A1(n22710), .A2(\xmem_data[58][1] ), .B1(n22709), .B2(
        \xmem_data[59][1] ), .ZN(n21993) );
  AOI22_X1 U25863 ( .A1(n22711), .A2(\xmem_data[60][1] ), .B1(n27396), .B2(
        \xmem_data[61][1] ), .ZN(n21992) );
  AOI22_X1 U25864 ( .A1(n28045), .A2(\xmem_data[62][1] ), .B1(n22712), .B2(
        \xmem_data[63][1] ), .ZN(n21991) );
  AOI22_X1 U25865 ( .A1(n22729), .A2(\xmem_data[52][1] ), .B1(n22728), .B2(
        \xmem_data[53][1] ), .ZN(n21995) );
  NAND4_X1 U25866 ( .A1(n3862), .A2(n21996), .A3(n3532), .A4(n21995), .ZN(
        n21997) );
  OAI21_X1 U25867 ( .B1(n21998), .B2(n21997), .A(n22735), .ZN(n22053) );
  AOI22_X1 U25868 ( .A1(n22741), .A2(\xmem_data[4][1] ), .B1(n27818), .B2(
        \xmem_data[5][1] ), .ZN(n22002) );
  AOI22_X1 U25869 ( .A1(n22740), .A2(\xmem_data[2][1] ), .B1(n25425), .B2(
        \xmem_data[3][1] ), .ZN(n22001) );
  AOI22_X1 U25870 ( .A1(n22739), .A2(\xmem_data[0][1] ), .B1(n22738), .B2(
        \xmem_data[1][1] ), .ZN(n22000) );
  AOI22_X1 U25871 ( .A1(n22742), .A2(\xmem_data[6][1] ), .B1(n31330), .B2(
        \xmem_data[7][1] ), .ZN(n21999) );
  AND4_X1 U25872 ( .A1(n22002), .A2(n22001), .A3(n22000), .A4(n21999), .ZN(
        n22010) );
  AOI22_X1 U25873 ( .A1(n3219), .A2(\xmem_data[24][1] ), .B1(n28367), .B2(
        \xmem_data[25][1] ), .ZN(n22003) );
  INV_X1 U25874 ( .A(n22003), .ZN(n22008) );
  AOI22_X1 U25875 ( .A1(n22759), .A2(\xmem_data[28][1] ), .B1(n29567), .B2(
        \xmem_data[29][1] ), .ZN(n22006) );
  AOI22_X1 U25876 ( .A1(n22710), .A2(\xmem_data[26][1] ), .B1(n22758), .B2(
        \xmem_data[27][1] ), .ZN(n22005) );
  NAND2_X1 U25877 ( .A1(n27447), .A2(\xmem_data[31][1] ), .ZN(n22004) );
  NAND3_X1 U25878 ( .A1(n22006), .A2(n22005), .A3(n22004), .ZN(n22007) );
  NOR2_X1 U25879 ( .A1(n22008), .A2(n22007), .ZN(n22009) );
  NAND2_X1 U25880 ( .A1(n22010), .A2(n22009), .ZN(n22021) );
  AOI22_X1 U25881 ( .A1(n22751), .A2(\xmem_data[16][1] ), .B1(n28772), .B2(
        \xmem_data[17][1] ), .ZN(n22014) );
  AOI22_X1 U25882 ( .A1(n31261), .A2(\xmem_data[18][1] ), .B1(n28354), .B2(
        \xmem_data[19][1] ), .ZN(n22013) );
  AOI22_X1 U25883 ( .A1(n22752), .A2(\xmem_data[20][1] ), .B1(n3413), .B2(
        \xmem_data[21][1] ), .ZN(n22012) );
  AOI22_X1 U25884 ( .A1(n22753), .A2(\xmem_data[22][1] ), .B1(n29064), .B2(
        \xmem_data[23][1] ), .ZN(n22011) );
  NAND4_X1 U25885 ( .A1(n22014), .A2(n22013), .A3(n22012), .A4(n22011), .ZN(
        n22020) );
  AOI22_X1 U25886 ( .A1(n28058), .A2(\xmem_data[8][1] ), .B1(n29410), .B2(
        \xmem_data[9][1] ), .ZN(n22018) );
  AOI22_X1 U25887 ( .A1(n29238), .A2(\xmem_data[10][1] ), .B1(n28428), .B2(
        \xmem_data[11][1] ), .ZN(n22017) );
  AOI22_X1 U25888 ( .A1(n25581), .A2(\xmem_data[12][1] ), .B1(n31315), .B2(
        \xmem_data[13][1] ), .ZN(n22016) );
  AOI22_X1 U25889 ( .A1(n27975), .A2(\xmem_data[14][1] ), .B1(n20818), .B2(
        \xmem_data[15][1] ), .ZN(n22015) );
  NAND4_X1 U25890 ( .A1(n22018), .A2(n22017), .A3(n22016), .A4(n22015), .ZN(
        n22019) );
  NOR2_X1 U25891 ( .A1(n22022), .A2(n39014), .ZN(n22023) );
  AOI21_X1 U25892 ( .B1(n22024), .B2(n22768), .A(n3884), .ZN(n22052) );
  AOI22_X1 U25893 ( .A1(n3220), .A2(\xmem_data[88][1] ), .B1(n29789), .B2(
        \xmem_data[89][1] ), .ZN(n22028) );
  AOI22_X1 U25894 ( .A1(n22667), .A2(\xmem_data[90][1] ), .B1(n22666), .B2(
        \xmem_data[91][1] ), .ZN(n22027) );
  AOI22_X1 U25895 ( .A1(n22669), .A2(\xmem_data[92][1] ), .B1(n22668), .B2(
        \xmem_data[93][1] ), .ZN(n22026) );
  AOI22_X1 U25896 ( .A1(n25450), .A2(\xmem_data[94][1] ), .B1(n30551), .B2(
        \xmem_data[95][1] ), .ZN(n22025) );
  AOI22_X1 U25897 ( .A1(n30861), .A2(\xmem_data[84][1] ), .B1(n3229), .B2(
        \xmem_data[85][1] ), .ZN(n22045) );
  AOI22_X1 U25898 ( .A1(n31360), .A2(\xmem_data[74][1] ), .B1(n22683), .B2(
        \xmem_data[75][1] ), .ZN(n22029) );
  INV_X1 U25899 ( .A(n22029), .ZN(n22034) );
  AOI22_X1 U25900 ( .A1(n29089), .A2(\xmem_data[76][1] ), .B1(n3301), .B2(
        \xmem_data[77][1] ), .ZN(n22032) );
  AOI22_X1 U25901 ( .A1(n22685), .A2(\xmem_data[78][1] ), .B1(n22684), .B2(
        \xmem_data[79][1] ), .ZN(n22031) );
  AOI22_X1 U25902 ( .A1(n14970), .A2(\xmem_data[72][1] ), .B1(n22682), .B2(
        \xmem_data[73][1] ), .ZN(n22030) );
  NOR2_X1 U25903 ( .A1(n22034), .A2(n22033), .ZN(n22044) );
  AOI22_X1 U25904 ( .A1(n22675), .A2(\xmem_data[66][1] ), .B1(n16986), .B2(
        \xmem_data[67][1] ), .ZN(n22036) );
  AOI22_X1 U25905 ( .A1(n22674), .A2(\xmem_data[68][1] ), .B1(n16988), .B2(
        \xmem_data[69][1] ), .ZN(n22035) );
  NAND2_X1 U25906 ( .A1(n22036), .A2(n22035), .ZN(n22042) );
  AOI22_X1 U25907 ( .A1(n22677), .A2(\xmem_data[70][1] ), .B1(n22676), .B2(
        \xmem_data[71][1] ), .ZN(n22037) );
  INV_X1 U25908 ( .A(n22037), .ZN(n22041) );
  AOI22_X1 U25909 ( .A1(n28415), .A2(\xmem_data[64][1] ), .B1(n27911), .B2(
        \xmem_data[65][1] ), .ZN(n22039) );
  AOI22_X1 U25910 ( .A1(n20951), .A2(\xmem_data[82][1] ), .B1(n17056), .B2(
        \xmem_data[83][1] ), .ZN(n22038) );
  NAND2_X1 U25911 ( .A1(n22039), .A2(n22038), .ZN(n22040) );
  NOR3_X1 U25912 ( .A1(n22042), .A2(n22041), .A3(n22040), .ZN(n22043) );
  NAND4_X1 U25913 ( .A1(n3854), .A2(n22045), .A3(n22044), .A4(n22043), .ZN(
        n22050) );
  AOI22_X1 U25914 ( .A1(n27463), .A2(\xmem_data[80][1] ), .B1(n28036), .B2(
        \xmem_data[81][1] ), .ZN(n22048) );
  AND2_X1 U25915 ( .A1(n30863), .A2(\xmem_data[86][1] ), .ZN(n22046) );
  AOI21_X1 U25916 ( .B1(n30906), .B2(\xmem_data[87][1] ), .A(n22046), .ZN(
        n22047) );
  NAND2_X1 U25917 ( .A1(n22048), .A2(n22047), .ZN(n22049) );
  OAI21_X1 U25918 ( .B1(n22050), .B2(n22049), .A(n22663), .ZN(n22051) );
  AOI22_X1 U25919 ( .A1(n22701), .A2(\xmem_data[32][2] ), .B1(n29308), .B2(
        \xmem_data[33][2] ), .ZN(n22058) );
  AOI22_X1 U25920 ( .A1(n22702), .A2(\xmem_data[34][2] ), .B1(n28298), .B2(
        \xmem_data[35][2] ), .ZN(n22057) );
  AOI22_X1 U25921 ( .A1(n22703), .A2(\xmem_data[36][2] ), .B1(n29237), .B2(
        \xmem_data[37][2] ), .ZN(n22056) );
  AOI22_X1 U25922 ( .A1(n29279), .A2(\xmem_data[38][2] ), .B1(n17020), .B2(
        \xmem_data[39][2] ), .ZN(n22055) );
  NAND4_X1 U25923 ( .A1(n22058), .A2(n22057), .A3(n22056), .A4(n22055), .ZN(
        n22074) );
  AOI22_X1 U25924 ( .A1(n22718), .A2(\xmem_data[40][2] ), .B1(n22717), .B2(
        \xmem_data[41][2] ), .ZN(n22062) );
  AOI22_X1 U25925 ( .A1(n25435), .A2(\xmem_data[42][2] ), .B1(n3178), .B2(
        \xmem_data[43][2] ), .ZN(n22061) );
  AOI22_X1 U25926 ( .A1(n20816), .A2(\xmem_data[44][2] ), .B1(n3338), .B2(
        \xmem_data[45][2] ), .ZN(n22060) );
  AOI22_X1 U25927 ( .A1(n28098), .A2(\xmem_data[46][2] ), .B1(n22719), .B2(
        \xmem_data[47][2] ), .ZN(n22059) );
  NAND4_X1 U25928 ( .A1(n22062), .A2(n22061), .A3(n22060), .A4(n22059), .ZN(
        n22073) );
  AOI22_X1 U25929 ( .A1(n27526), .A2(\xmem_data[48][2] ), .B1(n30257), .B2(
        \xmem_data[49][2] ), .ZN(n22066) );
  AOI22_X1 U25930 ( .A1(n22727), .A2(\xmem_data[50][2] ), .B1(n24607), .B2(
        \xmem_data[51][2] ), .ZN(n22065) );
  AOI22_X1 U25931 ( .A1(n22729), .A2(\xmem_data[52][2] ), .B1(n22728), .B2(
        \xmem_data[53][2] ), .ZN(n22064) );
  AOI22_X1 U25932 ( .A1(n22753), .A2(\xmem_data[54][2] ), .B1(n25354), .B2(
        \xmem_data[55][2] ), .ZN(n22063) );
  NAND4_X1 U25933 ( .A1(n22066), .A2(n22065), .A3(n22064), .A4(n22063), .ZN(
        n22072) );
  AOI22_X1 U25934 ( .A1(n3218), .A2(\xmem_data[56][2] ), .B1(n22708), .B2(
        \xmem_data[57][2] ), .ZN(n22070) );
  AOI22_X1 U25935 ( .A1(n22710), .A2(\xmem_data[58][2] ), .B1(n22709), .B2(
        \xmem_data[59][2] ), .ZN(n22069) );
  AOI22_X1 U25936 ( .A1(n22711), .A2(\xmem_data[60][2] ), .B1(n28952), .B2(
        \xmem_data[61][2] ), .ZN(n22068) );
  AOI22_X1 U25937 ( .A1(n24657), .A2(\xmem_data[62][2] ), .B1(n22712), .B2(
        \xmem_data[63][2] ), .ZN(n22067) );
  NAND4_X1 U25938 ( .A1(n22070), .A2(n22069), .A3(n22068), .A4(n22067), .ZN(
        n22071) );
  OR4_X1 U25939 ( .A1(n22074), .A2(n22073), .A3(n22072), .A4(n22071), .ZN(
        n22104) );
  AOI22_X1 U25940 ( .A1(n3222), .A2(\xmem_data[24][2] ), .B1(n28733), .B2(
        \xmem_data[25][2] ), .ZN(n22081) );
  AOI22_X1 U25941 ( .A1(n22759), .A2(\xmem_data[28][2] ), .B1(n22668), .B2(
        \xmem_data[29][2] ), .ZN(n22075) );
  INV_X1 U25942 ( .A(n22075), .ZN(n22079) );
  AOI22_X1 U25943 ( .A1(n20992), .A2(\xmem_data[26][2] ), .B1(n22758), .B2(
        \xmem_data[27][2] ), .ZN(n22077) );
  NAND2_X1 U25944 ( .A1(n25422), .A2(\xmem_data[31][2] ), .ZN(n22076) );
  NAND2_X1 U25945 ( .A1(n22077), .A2(n22076), .ZN(n22078) );
  NOR2_X1 U25946 ( .A1(n22079), .A2(n22078), .ZN(n22080) );
  NAND2_X1 U25947 ( .A1(n22081), .A2(n22080), .ZN(n22087) );
  AOI22_X1 U25948 ( .A1(n22739), .A2(\xmem_data[0][2] ), .B1(n22738), .B2(
        \xmem_data[1][2] ), .ZN(n22085) );
  AOI22_X1 U25949 ( .A1(n22740), .A2(\xmem_data[2][2] ), .B1(n17041), .B2(
        \xmem_data[3][2] ), .ZN(n22084) );
  AOI22_X1 U25950 ( .A1(n22741), .A2(\xmem_data[4][2] ), .B1(n3158), .B2(
        \xmem_data[5][2] ), .ZN(n22083) );
  AOI22_X1 U25951 ( .A1(n22742), .A2(\xmem_data[6][2] ), .B1(n17020), .B2(
        \xmem_data[7][2] ), .ZN(n22082) );
  NAND4_X1 U25952 ( .A1(n22085), .A2(n22084), .A3(n22083), .A4(n22082), .ZN(
        n22086) );
  OR2_X1 U25953 ( .A1(n22087), .A2(n22086), .ZN(n22100) );
  AND2_X1 U25954 ( .A1(n22751), .A2(\xmem_data[16][2] ), .ZN(n22088) );
  AOI21_X1 U25955 ( .B1(n29657), .B2(\xmem_data[17][2] ), .A(n22088), .ZN(
        n22092) );
  AOI22_X1 U25956 ( .A1(n28035), .A2(\xmem_data[18][2] ), .B1(n27564), .B2(
        \xmem_data[19][2] ), .ZN(n22091) );
  AOI22_X1 U25957 ( .A1(n22752), .A2(\xmem_data[20][2] ), .B1(n3228), .B2(
        \xmem_data[21][2] ), .ZN(n22090) );
  AOI22_X1 U25958 ( .A1(n22753), .A2(\xmem_data[22][2] ), .B1(n29064), .B2(
        \xmem_data[23][2] ), .ZN(n22089) );
  NAND4_X1 U25959 ( .A1(n22092), .A2(n22091), .A3(n22090), .A4(n22089), .ZN(
        n22098) );
  AOI22_X1 U25960 ( .A1(n23796), .A2(\xmem_data[8][2] ), .B1(n23722), .B2(
        \xmem_data[9][2] ), .ZN(n22096) );
  AOI22_X1 U25961 ( .A1(n29190), .A2(\xmem_data[10][2] ), .B1(n28385), .B2(
        \xmem_data[11][2] ), .ZN(n22095) );
  AOI22_X1 U25962 ( .A1(n27856), .A2(\xmem_data[12][2] ), .B1(n3300), .B2(
        \xmem_data[13][2] ), .ZN(n22094) );
  AOI22_X1 U25963 ( .A1(n22685), .A2(\xmem_data[14][2] ), .B1(n3171), .B2(
        \xmem_data[15][2] ), .ZN(n22093) );
  NAND4_X1 U25964 ( .A1(n22096), .A2(n22095), .A3(n22094), .A4(n22093), .ZN(
        n22097) );
  OR2_X1 U25965 ( .A1(n22098), .A2(n22097), .ZN(n22099) );
  NOR2_X1 U25966 ( .A1(n22100), .A2(n22099), .ZN(n22102) );
  NAND2_X1 U25967 ( .A1(n23771), .A2(\xmem_data[30][2] ), .ZN(n22101) );
  AOI21_X1 U25968 ( .B1(n22102), .B2(n22101), .A(n22022), .ZN(n22103) );
  AOI21_X1 U25969 ( .B1(n22104), .B2(n22735), .A(n22103), .ZN(n22150) );
  AOI22_X1 U25970 ( .A1(n28415), .A2(\xmem_data[64][2] ), .B1(n27453), .B2(
        \xmem_data[65][2] ), .ZN(n22108) );
  AOI22_X1 U25971 ( .A1(n22675), .A2(\xmem_data[66][2] ), .B1(n28298), .B2(
        \xmem_data[67][2] ), .ZN(n22107) );
  AOI22_X1 U25972 ( .A1(n22674), .A2(\xmem_data[68][2] ), .B1(n29237), .B2(
        \xmem_data[69][2] ), .ZN(n22106) );
  AOI22_X1 U25973 ( .A1(n22677), .A2(\xmem_data[70][2] ), .B1(n22676), .B2(
        \xmem_data[71][2] ), .ZN(n22105) );
  NAND4_X1 U25974 ( .A1(n22108), .A2(n22107), .A3(n22106), .A4(n22105), .ZN(
        n22125) );
  AOI22_X1 U25975 ( .A1(n28058), .A2(\xmem_data[72][2] ), .B1(n22682), .B2(
        \xmem_data[73][2] ), .ZN(n22112) );
  AOI22_X1 U25976 ( .A1(n30545), .A2(\xmem_data[74][2] ), .B1(n22683), .B2(
        \xmem_data[75][2] ), .ZN(n22111) );
  AOI22_X1 U25977 ( .A1(n25581), .A2(\xmem_data[76][2] ), .B1(n17004), .B2(
        \xmem_data[77][2] ), .ZN(n22110) );
  AOI22_X1 U25978 ( .A1(n22685), .A2(\xmem_data[78][2] ), .B1(n22684), .B2(
        \xmem_data[79][2] ), .ZN(n22109) );
  NAND4_X1 U25979 ( .A1(n22112), .A2(n22111), .A3(n22110), .A4(n22109), .ZN(
        n22124) );
  AOI22_X1 U25980 ( .A1(n27526), .A2(\xmem_data[80][2] ), .B1(n30674), .B2(
        \xmem_data[81][2] ), .ZN(n22117) );
  AOI22_X1 U25981 ( .A1(n31344), .A2(\xmem_data[82][2] ), .B1(n20710), .B2(
        \xmem_data[83][2] ), .ZN(n22116) );
  AOI22_X1 U25982 ( .A1(n31309), .A2(\xmem_data[84][2] ), .B1(n3229), .B2(
        \xmem_data[85][2] ), .ZN(n22115) );
  AND2_X1 U25983 ( .A1(n25360), .A2(\xmem_data[86][2] ), .ZN(n22113) );
  AOI21_X1 U25984 ( .B1(n30503), .B2(\xmem_data[87][2] ), .A(n22113), .ZN(
        n22114) );
  NAND4_X1 U25985 ( .A1(n22117), .A2(n22116), .A3(n22115), .A4(n22114), .ZN(
        n22123) );
  AOI22_X1 U25986 ( .A1(n3219), .A2(\xmem_data[88][2] ), .B1(n24632), .B2(
        \xmem_data[89][2] ), .ZN(n22121) );
  AOI22_X1 U25987 ( .A1(n22667), .A2(\xmem_data[90][2] ), .B1(n22666), .B2(
        \xmem_data[91][2] ), .ZN(n22120) );
  AOI22_X1 U25988 ( .A1(n22669), .A2(\xmem_data[92][2] ), .B1(n22668), .B2(
        \xmem_data[93][2] ), .ZN(n22119) );
  AOI22_X1 U25989 ( .A1(n30877), .A2(\xmem_data[94][2] ), .B1(n28374), .B2(
        \xmem_data[95][2] ), .ZN(n22118) );
  NAND4_X1 U25990 ( .A1(n22121), .A2(n22120), .A3(n22119), .A4(n22118), .ZN(
        n22122) );
  OR4_X1 U25991 ( .A1(n22125), .A2(n22124), .A3(n22123), .A4(n22122), .ZN(
        n22148) );
  AOI22_X1 U25992 ( .A1(n3357), .A2(\xmem_data[96][2] ), .B1(n25457), .B2(
        \xmem_data[97][2] ), .ZN(n22129) );
  AOI22_X1 U25993 ( .A1(n22675), .A2(\xmem_data[98][2] ), .B1(n25425), .B2(
        \xmem_data[99][2] ), .ZN(n22128) );
  AOI22_X1 U25994 ( .A1(n22674), .A2(\xmem_data[100][2] ), .B1(n24213), .B2(
        \xmem_data[101][2] ), .ZN(n22127) );
  AOI22_X1 U25995 ( .A1(n22677), .A2(\xmem_data[102][2] ), .B1(n22676), .B2(
        \xmem_data[103][2] ), .ZN(n22126) );
  NAND4_X1 U25996 ( .A1(n22129), .A2(n22128), .A3(n22127), .A4(n22126), .ZN(
        n22146) );
  AOI22_X1 U25997 ( .A1(n24459), .A2(\xmem_data[104][2] ), .B1(n22682), .B2(
        \xmem_data[105][2] ), .ZN(n22133) );
  AOI22_X1 U25998 ( .A1(n29049), .A2(\xmem_data[106][2] ), .B1(n22683), .B2(
        \xmem_data[107][2] ), .ZN(n22132) );
  AOI22_X1 U25999 ( .A1(n28494), .A2(\xmem_data[108][2] ), .B1(n3329), .B2(
        \xmem_data[109][2] ), .ZN(n22131) );
  AOI22_X1 U26000 ( .A1(n22685), .A2(\xmem_data[110][2] ), .B1(n22684), .B2(
        \xmem_data[111][2] ), .ZN(n22130) );
  NAND4_X1 U26001 ( .A1(n22133), .A2(n22132), .A3(n22131), .A4(n22130), .ZN(
        n22145) );
  AOI22_X1 U26002 ( .A1(n25406), .A2(\xmem_data[112][2] ), .B1(n17051), .B2(
        \xmem_data[113][2] ), .ZN(n22138) );
  AOI22_X1 U26003 ( .A1(n29125), .A2(\xmem_data[114][2] ), .B1(n25441), .B2(
        \xmem_data[115][2] ), .ZN(n22137) );
  AOI22_X1 U26004 ( .A1(n30908), .A2(\xmem_data[116][2] ), .B1(n3350), .B2(
        \xmem_data[117][2] ), .ZN(n22136) );
  AND2_X1 U26005 ( .A1(n14983), .A2(\xmem_data[118][2] ), .ZN(n22134) );
  AOI21_X1 U26006 ( .B1(n23734), .B2(\xmem_data[119][2] ), .A(n22134), .ZN(
        n22135) );
  NAND4_X1 U26007 ( .A1(n22138), .A2(n22137), .A3(n22136), .A4(n22135), .ZN(
        n22144) );
  AOI22_X1 U26008 ( .A1(n3217), .A2(\xmem_data[120][2] ), .B1(n22708), .B2(
        \xmem_data[121][2] ), .ZN(n22142) );
  AOI22_X1 U26009 ( .A1(n22667), .A2(\xmem_data[122][2] ), .B1(n22666), .B2(
        \xmem_data[123][2] ), .ZN(n22141) );
  AOI22_X1 U26010 ( .A1(n22669), .A2(\xmem_data[124][2] ), .B1(n22668), .B2(
        \xmem_data[125][2] ), .ZN(n22140) );
  AOI22_X1 U26011 ( .A1(n29306), .A2(\xmem_data[126][2] ), .B1(n28374), .B2(
        \xmem_data[127][2] ), .ZN(n22139) );
  NAND4_X1 U26012 ( .A1(n22142), .A2(n22141), .A3(n22140), .A4(n22139), .ZN(
        n22143) );
  OR4_X1 U26013 ( .A1(n22146), .A2(n22145), .A3(n22144), .A4(n22143), .ZN(
        n22147) );
  AOI22_X1 U26014 ( .A1(n22148), .A2(n22663), .B1(n22147), .B2(n22698), .ZN(
        n22149) );
  XNOR2_X1 U26015 ( .A(n32419), .B(\fmem_data[5][7] ), .ZN(n30358) );
  OAI21_X1 U26016 ( .B1(n34030), .B2(n34029), .A(n34031), .ZN(n22152) );
  NAND2_X1 U26017 ( .A1(n34030), .A2(n34029), .ZN(n22151) );
  NAND2_X1 U26018 ( .A1(n22152), .A2(n22151), .ZN(n23181) );
  FA_X1 U26019 ( .A(n22154), .B(n22155), .CI(n22153), .CO(n26264), .S(n27316)
         );
  XNOR2_X1 U26020 ( .A(n31489), .B(\fmem_data[21][3] ), .ZN(n32116) );
  XNOR2_X1 U26021 ( .A(n31882), .B(\fmem_data[21][3] ), .ZN(n33159) );
  OAI22_X1 U26022 ( .A1(n32116), .A2(n34199), .B1(n34201), .B2(n33159), .ZN(
        n29529) );
  AOI22_X1 U26023 ( .A1(n24157), .A2(\xmem_data[12][5] ), .B1(n24448), .B2(
        \xmem_data[13][5] ), .ZN(n22162) );
  AOI22_X1 U26024 ( .A1(n30514), .A2(\xmem_data[14][5] ), .B1(n22741), .B2(
        \xmem_data[15][5] ), .ZN(n22156) );
  INV_X1 U26025 ( .A(n22156), .ZN(n22160) );
  AOI22_X1 U26026 ( .A1(n24450), .A2(\xmem_data[10][5] ), .B1(n29307), .B2(
        \xmem_data[11][5] ), .ZN(n22158) );
  NAND2_X1 U26027 ( .A1(n29706), .A2(\xmem_data[8][5] ), .ZN(n22157) );
  NAND2_X1 U26028 ( .A1(n22158), .A2(n22157), .ZN(n22159) );
  NOR2_X1 U26029 ( .A1(n22160), .A2(n22159), .ZN(n22161) );
  NAND2_X1 U26030 ( .A1(n22162), .A2(n22161), .ZN(n22178) );
  AOI22_X1 U26031 ( .A1(n3350), .A2(\xmem_data[0][5] ), .B1(n24439), .B2(
        \xmem_data[1][5] ), .ZN(n22166) );
  AOI22_X1 U26032 ( .A1(n24443), .A2(\xmem_data[2][5] ), .B1(n3221), .B2(
        \xmem_data[3][5] ), .ZN(n22165) );
  AOI22_X1 U26033 ( .A1(n28137), .A2(\xmem_data[4][5] ), .B1(n29095), .B2(
        \xmem_data[5][5] ), .ZN(n22164) );
  AOI22_X1 U26034 ( .A1(n24438), .A2(\xmem_data[6][5] ), .B1(n20806), .B2(
        \xmem_data[7][5] ), .ZN(n22163) );
  NAND4_X1 U26035 ( .A1(n22166), .A2(n22165), .A3(n22164), .A4(n22163), .ZN(
        n22177) );
  AOI22_X1 U26036 ( .A1(n3338), .A2(\xmem_data[24][5] ), .B1(n28983), .B2(
        \xmem_data[25][5] ), .ZN(n22170) );
  AOI22_X1 U26037 ( .A1(n24467), .A2(\xmem_data[26][5] ), .B1(n23781), .B2(
        \xmem_data[27][5] ), .ZN(n22169) );
  AOI22_X1 U26038 ( .A1(n29657), .A2(\xmem_data[28][5] ), .B1(n24468), .B2(
        \xmem_data[29][5] ), .ZN(n22168) );
  AOI22_X1 U26039 ( .A1(n25630), .A2(\xmem_data[30][5] ), .B1(n24470), .B2(
        \xmem_data[31][5] ), .ZN(n22167) );
  NAND4_X1 U26040 ( .A1(n22170), .A2(n22169), .A3(n22168), .A4(n22167), .ZN(
        n22176) );
  AOI22_X1 U26041 ( .A1(n24458), .A2(\xmem_data[16][5] ), .B1(n24457), .B2(
        \xmem_data[17][5] ), .ZN(n22174) );
  AOI22_X1 U26042 ( .A1(n24133), .A2(\xmem_data[18][5] ), .B1(n24459), .B2(
        \xmem_data[19][5] ), .ZN(n22173) );
  AOI22_X1 U26043 ( .A1(n16990), .A2(\xmem_data[20][5] ), .B1(n24460), .B2(
        \xmem_data[21][5] ), .ZN(n22172) );
  AOI22_X1 U26044 ( .A1(n3178), .A2(\xmem_data[22][5] ), .B1(n3372), .B2(
        \xmem_data[23][5] ), .ZN(n22171) );
  NAND4_X1 U26045 ( .A1(n22174), .A2(n22173), .A3(n22172), .A4(n22171), .ZN(
        n22175) );
  NOR2_X1 U26046 ( .A1(n22298), .A2(n39031), .ZN(n22179) );
  AOI22_X1 U26047 ( .A1(n24562), .A2(\xmem_data[66][5] ), .B1(n3220), .B2(
        \xmem_data[67][5] ), .ZN(n22188) );
  AOI22_X1 U26048 ( .A1(n24565), .A2(\xmem_data[70][5] ), .B1(n24564), .B2(
        \xmem_data[71][5] ), .ZN(n22182) );
  INV_X1 U26049 ( .A(n22182), .ZN(n22186) );
  AOI22_X1 U26050 ( .A1(n24563), .A2(\xmem_data[68][5] ), .B1(n24695), .B2(
        \xmem_data[69][5] ), .ZN(n22184) );
  AOI22_X1 U26051 ( .A1(n3245), .A2(\xmem_data[64][5] ), .B1(n31347), .B2(
        \xmem_data[65][5] ), .ZN(n22183) );
  NAND2_X1 U26052 ( .A1(n22184), .A2(n22183), .ZN(n22185) );
  NOR2_X1 U26053 ( .A1(n22186), .A2(n22185), .ZN(n22187) );
  NAND2_X1 U26054 ( .A1(n22188), .A2(n22187), .ZN(n22204) );
  AOI22_X1 U26055 ( .A1(n29231), .A2(\xmem_data[72][5] ), .B1(n24553), .B2(
        \xmem_data[73][5] ), .ZN(n22192) );
  AOI22_X1 U26056 ( .A1(n24554), .A2(\xmem_data[74][5] ), .B1(n28373), .B2(
        \xmem_data[75][5] ), .ZN(n22191) );
  AOI22_X1 U26057 ( .A1(n24556), .A2(\xmem_data[76][5] ), .B1(n24555), .B2(
        \xmem_data[77][5] ), .ZN(n22190) );
  AOI22_X1 U26058 ( .A1(n16986), .A2(\xmem_data[78][5] ), .B1(n25709), .B2(
        \xmem_data[79][5] ), .ZN(n22189) );
  NAND4_X1 U26059 ( .A1(n22192), .A2(n22191), .A3(n22190), .A4(n22189), .ZN(
        n22203) );
  AOI22_X1 U26060 ( .A1(n24545), .A2(\xmem_data[80][5] ), .B1(n31269), .B2(
        \xmem_data[81][5] ), .ZN(n22196) );
  AOI22_X1 U26061 ( .A1(n24547), .A2(\xmem_data[82][5] ), .B1(n24546), .B2(
        \xmem_data[83][5] ), .ZN(n22195) );
  AOI22_X1 U26062 ( .A1(n24115), .A2(\xmem_data[84][5] ), .B1(n31360), .B2(
        \xmem_data[85][5] ), .ZN(n22194) );
  AOI22_X1 U26063 ( .A1(n29100), .A2(\xmem_data[86][5] ), .B1(n25581), .B2(
        \xmem_data[87][5] ), .ZN(n22193) );
  NAND4_X1 U26064 ( .A1(n22196), .A2(n22195), .A3(n22194), .A4(n22193), .ZN(
        n22202) );
  AOI22_X1 U26065 ( .A1(n24571), .A2(\xmem_data[88][5] ), .B1(n24570), .B2(
        \xmem_data[89][5] ), .ZN(n22200) );
  AOI22_X1 U26066 ( .A1(n24572), .A2(\xmem_data[90][5] ), .B1(n28500), .B2(
        \xmem_data[91][5] ), .ZN(n22199) );
  AOI22_X1 U26067 ( .A1(n23753), .A2(\xmem_data[92][5] ), .B1(n30601), .B2(
        \xmem_data[93][5] ), .ZN(n22198) );
  AOI22_X1 U26068 ( .A1(n30909), .A2(\xmem_data[94][5] ), .B1(n24573), .B2(
        \xmem_data[95][5] ), .ZN(n22197) );
  NAND4_X1 U26069 ( .A1(n22200), .A2(n22199), .A3(n22198), .A4(n22197), .ZN(
        n22201) );
  OR4_X1 U26070 ( .A1(n22204), .A2(n22203), .A3(n22202), .A4(n22201), .ZN(
        n22205) );
  NAND2_X1 U26071 ( .A1(n22205), .A2(n24581), .ZN(n22250) );
  AOI22_X1 U26072 ( .A1(n3351), .A2(\xmem_data[32][5] ), .B1(n27437), .B2(
        \xmem_data[33][5] ), .ZN(n22209) );
  AOI22_X1 U26073 ( .A1(n24562), .A2(\xmem_data[34][5] ), .B1(n3222), .B2(
        \xmem_data[35][5] ), .ZN(n22208) );
  AOI22_X1 U26074 ( .A1(n24563), .A2(\xmem_data[36][5] ), .B1(n22710), .B2(
        \xmem_data[37][5] ), .ZN(n22207) );
  AOI22_X1 U26075 ( .A1(n24565), .A2(\xmem_data[38][5] ), .B1(n24564), .B2(
        \xmem_data[39][5] ), .ZN(n22206) );
  NAND4_X1 U26076 ( .A1(n22209), .A2(n22208), .A3(n22207), .A4(n22206), .ZN(
        n22225) );
  AOI22_X1 U26077 ( .A1(n16973), .A2(\xmem_data[40][5] ), .B1(n24553), .B2(
        \xmem_data[41][5] ), .ZN(n22213) );
  AOI22_X1 U26078 ( .A1(n24554), .A2(\xmem_data[42][5] ), .B1(n27943), .B2(
        \xmem_data[43][5] ), .ZN(n22212) );
  AOI22_X1 U26079 ( .A1(n24556), .A2(\xmem_data[44][5] ), .B1(n24555), .B2(
        \xmem_data[45][5] ), .ZN(n22211) );
  AOI22_X1 U26080 ( .A1(n28298), .A2(\xmem_data[46][5] ), .B1(n25382), .B2(
        \xmem_data[47][5] ), .ZN(n22210) );
  NAND4_X1 U26081 ( .A1(n22213), .A2(n22212), .A3(n22211), .A4(n22210), .ZN(
        n22224) );
  AOI22_X1 U26082 ( .A1(n24545), .A2(\xmem_data[48][5] ), .B1(n3207), .B2(
        \xmem_data[49][5] ), .ZN(n22217) );
  AOI22_X1 U26083 ( .A1(n24547), .A2(\xmem_data[50][5] ), .B1(n24546), .B2(
        \xmem_data[51][5] ), .ZN(n22216) );
  AOI22_X1 U26084 ( .A1(n28994), .A2(\xmem_data[52][5] ), .B1(n25435), .B2(
        \xmem_data[53][5] ), .ZN(n22215) );
  AOI22_X1 U26085 ( .A1(n3325), .A2(\xmem_data[54][5] ), .B1(n27856), .B2(
        \xmem_data[55][5] ), .ZN(n22214) );
  NAND4_X1 U26086 ( .A1(n22217), .A2(n22216), .A3(n22215), .A4(n22214), .ZN(
        n22223) );
  AOI22_X1 U26087 ( .A1(n24571), .A2(\xmem_data[56][5] ), .B1(n24570), .B2(
        \xmem_data[57][5] ), .ZN(n22221) );
  AOI22_X1 U26088 ( .A1(n24572), .A2(\xmem_data[58][5] ), .B1(n21057), .B2(
        \xmem_data[59][5] ), .ZN(n22220) );
  AOI22_X1 U26089 ( .A1(n21060), .A2(\xmem_data[60][5] ), .B1(n30900), .B2(
        \xmem_data[61][5] ), .ZN(n22219) );
  AOI22_X1 U26090 ( .A1(n25408), .A2(\xmem_data[62][5] ), .B1(n24573), .B2(
        \xmem_data[63][5] ), .ZN(n22218) );
  NAND4_X1 U26091 ( .A1(n22221), .A2(n22220), .A3(n22219), .A4(n22218), .ZN(
        n22222) );
  OR4_X1 U26092 ( .A1(n22225), .A2(n22224), .A3(n22223), .A4(n22222), .ZN(
        n22226) );
  NAND2_X1 U26093 ( .A1(n22226), .A2(n24508), .ZN(n22249) );
  AOI22_X1 U26094 ( .A1(n3424), .A2(\xmem_data[96][5] ), .B1(n24172), .B2(
        \xmem_data[97][5] ), .ZN(n22230) );
  AOI22_X1 U26095 ( .A1(n24532), .A2(\xmem_data[98][5] ), .B1(n3217), .B2(
        \xmem_data[99][5] ), .ZN(n22229) );
  AOI22_X1 U26096 ( .A1(n24533), .A2(\xmem_data[100][5] ), .B1(n13469), .B2(
        \xmem_data[101][5] ), .ZN(n22228) );
  AOI22_X1 U26097 ( .A1(n24534), .A2(\xmem_data[102][5] ), .B1(n31275), .B2(
        \xmem_data[103][5] ), .ZN(n22227) );
  NAND4_X1 U26098 ( .A1(n22230), .A2(n22229), .A3(n22228), .A4(n22227), .ZN(
        n22246) );
  AOI22_X1 U26099 ( .A1(n20962), .A2(\xmem_data[104][5] ), .B1(n25514), .B2(
        \xmem_data[105][5] ), .ZN(n22234) );
  AOI22_X1 U26100 ( .A1(n30551), .A2(\xmem_data[106][5] ), .B1(n24130), .B2(
        \xmem_data[107][5] ), .ZN(n22233) );
  AOI22_X1 U26101 ( .A1(n29403), .A2(\xmem_data[108][5] ), .B1(n24516), .B2(
        \xmem_data[109][5] ), .ZN(n22232) );
  AOI22_X1 U26102 ( .A1(n28334), .A2(\xmem_data[110][5] ), .B1(n27912), .B2(
        \xmem_data[111][5] ), .ZN(n22231) );
  NAND4_X1 U26103 ( .A1(n22234), .A2(n22233), .A3(n22232), .A4(n22231), .ZN(
        n22245) );
  AOI22_X1 U26104 ( .A1(n30892), .A2(\xmem_data[112][5] ), .B1(n24134), .B2(
        \xmem_data[113][5] ), .ZN(n22238) );
  AOI22_X1 U26105 ( .A1(n24509), .A2(\xmem_data[114][5] ), .B1(n27518), .B2(
        \xmem_data[115][5] ), .ZN(n22237) );
  AOI22_X1 U26106 ( .A1(n17044), .A2(\xmem_data[116][5] ), .B1(n24510), .B2(
        \xmem_data[117][5] ), .ZN(n22236) );
  AOI22_X1 U26107 ( .A1(n24511), .A2(\xmem_data[118][5] ), .B1(n23778), .B2(
        \xmem_data[119][5] ), .ZN(n22235) );
  NAND4_X1 U26108 ( .A1(n22238), .A2(n22237), .A3(n22236), .A4(n22235), .ZN(
        n22244) );
  AOI22_X1 U26109 ( .A1(n24522), .A2(\xmem_data[120][5] ), .B1(n24521), .B2(
        \xmem_data[121][5] ), .ZN(n22242) );
  AOI22_X1 U26110 ( .A1(n3209), .A2(\xmem_data[122][5] ), .B1(n28468), .B2(
        \xmem_data[123][5] ), .ZN(n22241) );
  AOI22_X1 U26111 ( .A1(n28467), .A2(\xmem_data[124][5] ), .B1(n24524), .B2(
        \xmem_data[125][5] ), .ZN(n22240) );
  AOI22_X1 U26112 ( .A1(n24526), .A2(\xmem_data[126][5] ), .B1(n24525), .B2(
        \xmem_data[127][5] ), .ZN(n22239) );
  NAND4_X1 U26113 ( .A1(n22242), .A2(n22241), .A3(n22240), .A4(n22239), .ZN(
        n22243) );
  OR4_X1 U26114 ( .A1(n22246), .A2(n22245), .A3(n22244), .A4(n22243), .ZN(
        n22247) );
  NAND2_X1 U26115 ( .A1(n22247), .A2(n24542), .ZN(n22248) );
  NAND4_X2 U26116 ( .A1(n22251), .A2(n22250), .A3(n22249), .A4(n22248), .ZN(
        n34862) );
  AOI22_X1 U26117 ( .A1(n3338), .A2(\xmem_data[24][4] ), .B1(n27525), .B2(
        \xmem_data[25][4] ), .ZN(n22255) );
  AOI22_X1 U26118 ( .A1(n24467), .A2(\xmem_data[26][4] ), .B1(n29136), .B2(
        \xmem_data[27][4] ), .ZN(n22254) );
  AOI22_X1 U26119 ( .A1(n21060), .A2(\xmem_data[28][4] ), .B1(n24468), .B2(
        \xmem_data[29][4] ), .ZN(n22253) );
  AOI22_X1 U26120 ( .A1(n30862), .A2(\xmem_data[30][4] ), .B1(n24470), .B2(
        \xmem_data[31][4] ), .ZN(n22252) );
  AOI22_X1 U26121 ( .A1(n24458), .A2(\xmem_data[16][4] ), .B1(n24457), .B2(
        \xmem_data[17][4] ), .ZN(n22259) );
  AOI22_X1 U26122 ( .A1(n24133), .A2(\xmem_data[18][4] ), .B1(n24459), .B2(
        \xmem_data[19][4] ), .ZN(n22258) );
  AOI22_X1 U26123 ( .A1(n22682), .A2(\xmem_data[20][4] ), .B1(n24460), .B2(
        \xmem_data[21][4] ), .ZN(n22257) );
  AOI22_X1 U26124 ( .A1(n3178), .A2(\xmem_data[22][4] ), .B1(n28494), .B2(
        \xmem_data[23][4] ), .ZN(n22256) );
  NAND4_X1 U26125 ( .A1(n22259), .A2(n22258), .A3(n22257), .A4(n22256), .ZN(
        n22260) );
  NOR2_X1 U26126 ( .A1(n22260), .A2(n3733), .ZN(n22275) );
  AOI22_X1 U26127 ( .A1(n3333), .A2(\xmem_data[0][4] ), .B1(n24439), .B2(
        \xmem_data[1][4] ), .ZN(n22261) );
  INV_X1 U26128 ( .A(n22261), .ZN(n22263) );
  AND2_X1 U26129 ( .A1(n3217), .A2(\xmem_data[3][4] ), .ZN(n22262) );
  AOI22_X1 U26130 ( .A1(n24438), .A2(\xmem_data[6][4] ), .B1(n30550), .B2(
        \xmem_data[7][4] ), .ZN(n22265) );
  AOI22_X1 U26131 ( .A1(n30292), .A2(\xmem_data[4][4] ), .B1(n23739), .B2(
        \xmem_data[5][4] ), .ZN(n22264) );
  NAND2_X1 U26132 ( .A1(n22265), .A2(n22264), .ZN(n22266) );
  NOR2_X1 U26133 ( .A1(n3981), .A2(n22266), .ZN(n22274) );
  AOI22_X1 U26134 ( .A1(n29403), .A2(\xmem_data[12][4] ), .B1(n24448), .B2(
        \xmem_data[13][4] ), .ZN(n22267) );
  INV_X1 U26135 ( .A(n22267), .ZN(n22273) );
  AOI22_X1 U26136 ( .A1(n24450), .A2(\xmem_data[10][4] ), .B1(n30854), .B2(
        \xmem_data[11][4] ), .ZN(n22269) );
  NAND2_X1 U26137 ( .A1(n27905), .A2(\xmem_data[8][4] ), .ZN(n22268) );
  NAND2_X1 U26138 ( .A1(n22269), .A2(n22268), .ZN(n22272) );
  AOI22_X1 U26139 ( .A1(n31268), .A2(\xmem_data[14][4] ), .B1(n20717), .B2(
        \xmem_data[15][4] ), .ZN(n22270) );
  INV_X1 U26140 ( .A(n22270), .ZN(n22271) );
  NAND4_X1 U26141 ( .A1(n3545), .A2(n22275), .A3(n22274), .A4(n3898), .ZN(
        n22276) );
  NAND2_X1 U26142 ( .A1(n22276), .A2(n22180), .ZN(n22357) );
  AOI22_X1 U26143 ( .A1(n25624), .A2(\xmem_data[64][4] ), .B1(n31347), .B2(
        \xmem_data[65][4] ), .ZN(n22280) );
  AOI22_X1 U26144 ( .A1(n24562), .A2(\xmem_data[66][4] ), .B1(n3217), .B2(
        \xmem_data[67][4] ), .ZN(n22279) );
  AOI22_X1 U26145 ( .A1(n24563), .A2(\xmem_data[68][4] ), .B1(n20598), .B2(
        \xmem_data[69][4] ), .ZN(n22278) );
  AOI22_X1 U26146 ( .A1(n24565), .A2(\xmem_data[70][4] ), .B1(n24564), .B2(
        \xmem_data[71][4] ), .ZN(n22277) );
  NAND4_X1 U26147 ( .A1(n22280), .A2(n22279), .A3(n22278), .A4(n22277), .ZN(
        n22297) );
  AOI22_X1 U26148 ( .A1(n24571), .A2(\xmem_data[88][4] ), .B1(n24570), .B2(
        \xmem_data[89][4] ), .ZN(n22285) );
  AOI22_X1 U26149 ( .A1(n24572), .A2(\xmem_data[90][4] ), .B1(n25723), .B2(
        \xmem_data[91][4] ), .ZN(n22284) );
  AOI22_X1 U26150 ( .A1(n23753), .A2(\xmem_data[92][4] ), .B1(n17050), .B2(
        \xmem_data[93][4] ), .ZN(n22283) );
  AND2_X1 U26151 ( .A1(n17056), .A2(\xmem_data[94][4] ), .ZN(n22281) );
  AOI21_X1 U26152 ( .B1(n24573), .B2(\xmem_data[95][4] ), .A(n22281), .ZN(
        n22282) );
  NAND4_X1 U26153 ( .A1(n22285), .A2(n22284), .A3(n22283), .A4(n22282), .ZN(
        n22296) );
  AOI22_X1 U26154 ( .A1(n24545), .A2(\xmem_data[80][4] ), .B1(n3207), .B2(
        \xmem_data[81][4] ), .ZN(n22289) );
  AOI22_X1 U26155 ( .A1(n24547), .A2(\xmem_data[82][4] ), .B1(n24546), .B2(
        \xmem_data[83][4] ), .ZN(n22288) );
  AOI22_X1 U26156 ( .A1(n24710), .A2(\xmem_data[84][4] ), .B1(n30616), .B2(
        \xmem_data[85][4] ), .ZN(n22287) );
  AOI22_X1 U26157 ( .A1(n24220), .A2(\xmem_data[86][4] ), .B1(n23778), .B2(
        \xmem_data[87][4] ), .ZN(n22286) );
  NAND4_X1 U26158 ( .A1(n22289), .A2(n22288), .A3(n22287), .A4(n22286), .ZN(
        n22295) );
  AOI22_X1 U26159 ( .A1(n30295), .A2(\xmem_data[72][4] ), .B1(n24553), .B2(
        \xmem_data[73][4] ), .ZN(n22293) );
  AOI22_X1 U26160 ( .A1(n24554), .A2(\xmem_data[74][4] ), .B1(n25456), .B2(
        \xmem_data[75][4] ), .ZN(n22292) );
  AOI22_X1 U26161 ( .A1(n24556), .A2(\xmem_data[76][4] ), .B1(n24555), .B2(
        \xmem_data[77][4] ), .ZN(n22291) );
  AOI22_X1 U26162 ( .A1(n28298), .A2(\xmem_data[78][4] ), .B1(n25382), .B2(
        \xmem_data[79][4] ), .ZN(n22290) );
  NAND4_X1 U26163 ( .A1(n22293), .A2(n22292), .A3(n22291), .A4(n22290), .ZN(
        n22294) );
  OR4_X1 U26164 ( .A1(n22297), .A2(n22296), .A3(n22295), .A4(n22294), .ZN(
        n22300) );
  NOR2_X1 U26165 ( .A1(n22298), .A2(n39038), .ZN(n22299) );
  AOI21_X1 U26166 ( .B1(n22300), .B2(n24581), .A(n3893), .ZN(n22356) );
  AOI22_X1 U26167 ( .A1(n24545), .A2(\xmem_data[48][4] ), .B1(n3207), .B2(
        \xmem_data[49][4] ), .ZN(n22304) );
  AOI22_X1 U26168 ( .A1(n24547), .A2(\xmem_data[50][4] ), .B1(n24546), .B2(
        \xmem_data[51][4] ), .ZN(n22303) );
  AOI22_X1 U26169 ( .A1(n14971), .A2(\xmem_data[52][4] ), .B1(n28380), .B2(
        \xmem_data[53][4] ), .ZN(n22302) );
  AOI22_X1 U26170 ( .A1(n24548), .A2(\xmem_data[54][4] ), .B1(n27856), .B2(
        \xmem_data[55][4] ), .ZN(n22301) );
  NAND4_X1 U26171 ( .A1(n22304), .A2(n22303), .A3(n22302), .A4(n22301), .ZN(
        n22308) );
  AND2_X1 U26172 ( .A1(n3222), .A2(\xmem_data[35][4] ), .ZN(n22305) );
  AOI21_X1 U26173 ( .B1(n24562), .B2(\xmem_data[34][4] ), .A(n22305), .ZN(
        n22306) );
  INV_X1 U26174 ( .A(n22306), .ZN(n22307) );
  NOR2_X1 U26175 ( .A1(n22308), .A2(n22307), .ZN(n22331) );
  AOI22_X1 U26176 ( .A1(n24565), .A2(\xmem_data[38][4] ), .B1(n24564), .B2(
        \xmem_data[39][4] ), .ZN(n22309) );
  INV_X1 U26177 ( .A(n22309), .ZN(n22313) );
  AOI22_X1 U26178 ( .A1(n24563), .A2(\xmem_data[36][4] ), .B1(n25562), .B2(
        \xmem_data[37][4] ), .ZN(n22311) );
  AOI22_X1 U26179 ( .A1(n25725), .A2(\xmem_data[32][4] ), .B1(n30863), .B2(
        \xmem_data[33][4] ), .ZN(n22310) );
  NAND2_X1 U26180 ( .A1(n22311), .A2(n22310), .ZN(n22312) );
  NOR2_X1 U26181 ( .A1(n22313), .A2(n22312), .ZN(n22330) );
  AND2_X1 U26182 ( .A1(n30588), .A2(\xmem_data[62][4] ), .ZN(n22314) );
  AOI21_X1 U26183 ( .B1(n24573), .B2(\xmem_data[63][4] ), .A(n22314), .ZN(
        n22315) );
  INV_X1 U26184 ( .A(n22315), .ZN(n22319) );
  AOI22_X1 U26185 ( .A1(n24572), .A2(\xmem_data[58][4] ), .B1(n29247), .B2(
        \xmem_data[59][4] ), .ZN(n22317) );
  AOI22_X1 U26186 ( .A1(n24571), .A2(\xmem_data[56][4] ), .B1(n24570), .B2(
        \xmem_data[57][4] ), .ZN(n22316) );
  NAND2_X1 U26187 ( .A1(n22317), .A2(n22316), .ZN(n22318) );
  NOR2_X1 U26188 ( .A1(n22319), .A2(n22318), .ZN(n22329) );
  AOI22_X1 U26189 ( .A1(n21074), .A2(\xmem_data[40][4] ), .B1(n24553), .B2(
        \xmem_data[41][4] ), .ZN(n22323) );
  AOI22_X1 U26190 ( .A1(n24554), .A2(\xmem_data[42][4] ), .B1(n29180), .B2(
        \xmem_data[43][4] ), .ZN(n22322) );
  AOI22_X1 U26191 ( .A1(n24556), .A2(\xmem_data[44][4] ), .B1(n24555), .B2(
        \xmem_data[45][4] ), .ZN(n22321) );
  AOI22_X1 U26192 ( .A1(n27515), .A2(\xmem_data[46][4] ), .B1(n24597), .B2(
        \xmem_data[47][4] ), .ZN(n22320) );
  NAND4_X1 U26193 ( .A1(n22323), .A2(n22322), .A3(n22321), .A4(n22320), .ZN(
        n22327) );
  NAND2_X1 U26194 ( .A1(n25684), .A2(\xmem_data[60][4] ), .ZN(n22325) );
  NAND2_X1 U26195 ( .A1(n25440), .A2(\xmem_data[61][4] ), .ZN(n22324) );
  NAND2_X1 U26196 ( .A1(n22325), .A2(n22324), .ZN(n22326) );
  NOR2_X1 U26197 ( .A1(n22327), .A2(n22326), .ZN(n22328) );
  NAND4_X1 U26198 ( .A1(n22331), .A2(n22330), .A3(n22329), .A4(n22328), .ZN(
        n22332) );
  NAND2_X1 U26199 ( .A1(n22332), .A2(n24508), .ZN(n22355) );
  AOI22_X1 U26200 ( .A1(n3383), .A2(\xmem_data[96][4] ), .B1(n23731), .B2(
        \xmem_data[97][4] ), .ZN(n22336) );
  AOI22_X1 U26201 ( .A1(n24532), .A2(\xmem_data[98][4] ), .B1(n3217), .B2(
        \xmem_data[99][4] ), .ZN(n22335) );
  AOI22_X1 U26202 ( .A1(n24533), .A2(\xmem_data[100][4] ), .B1(n20500), .B2(
        \xmem_data[101][4] ), .ZN(n22334) );
  AOI22_X1 U26203 ( .A1(n24534), .A2(\xmem_data[102][4] ), .B1(n28372), .B2(
        \xmem_data[103][4] ), .ZN(n22333) );
  NAND4_X1 U26204 ( .A1(n22336), .A2(n22335), .A3(n22334), .A4(n22333), .ZN(
        n22352) );
  AOI22_X1 U26205 ( .A1(n3282), .A2(\xmem_data[104][4] ), .B1(n25514), .B2(
        \xmem_data[105][4] ), .ZN(n22340) );
  AOI22_X1 U26206 ( .A1(n24638), .A2(\xmem_data[106][4] ), .B1(n28373), .B2(
        \xmem_data[107][4] ), .ZN(n22339) );
  AOI22_X1 U26207 ( .A1(n27763), .A2(\xmem_data[108][4] ), .B1(n24516), .B2(
        \xmem_data[109][4] ), .ZN(n22338) );
  AOI22_X1 U26208 ( .A1(n28334), .A2(\xmem_data[110][4] ), .B1(n24160), .B2(
        \xmem_data[111][4] ), .ZN(n22337) );
  NAND4_X1 U26209 ( .A1(n22340), .A2(n22339), .A3(n22338), .A4(n22337), .ZN(
        n22351) );
  AOI22_X1 U26210 ( .A1(n28752), .A2(\xmem_data[112][4] ), .B1(n3212), .B2(
        \xmem_data[113][4] ), .ZN(n22344) );
  AOI22_X1 U26211 ( .A1(n24509), .A2(\xmem_data[114][4] ), .B1(n21006), .B2(
        \xmem_data[115][4] ), .ZN(n22343) );
  AOI22_X1 U26212 ( .A1(n28302), .A2(\xmem_data[116][4] ), .B1(n24510), .B2(
        \xmem_data[117][4] ), .ZN(n22342) );
  AOI22_X1 U26213 ( .A1(n24511), .A2(\xmem_data[118][4] ), .B1(n28060), .B2(
        \xmem_data[119][4] ), .ZN(n22341) );
  NAND4_X1 U26214 ( .A1(n22344), .A2(n22343), .A3(n22342), .A4(n22341), .ZN(
        n22350) );
  AOI22_X1 U26215 ( .A1(n24522), .A2(\xmem_data[120][4] ), .B1(n24521), .B2(
        \xmem_data[121][4] ), .ZN(n22348) );
  AOI22_X1 U26216 ( .A1(n3209), .A2(\xmem_data[122][4] ), .B1(n25359), .B2(
        \xmem_data[123][4] ), .ZN(n22347) );
  AOI22_X1 U26217 ( .A1(n25628), .A2(\xmem_data[124][4] ), .B1(n24524), .B2(
        \xmem_data[125][4] ), .ZN(n22346) );
  AOI22_X1 U26218 ( .A1(n24526), .A2(\xmem_data[126][4] ), .B1(n24525), .B2(
        \xmem_data[127][4] ), .ZN(n22345) );
  NAND4_X1 U26219 ( .A1(n22348), .A2(n22347), .A3(n22346), .A4(n22345), .ZN(
        n22349) );
  OR4_X1 U26220 ( .A1(n22352), .A2(n22351), .A3(n22350), .A4(n22349), .ZN(
        n22353) );
  NAND2_X1 U26221 ( .A1(n22353), .A2(n24542), .ZN(n22354) );
  NAND4_X1 U26222 ( .A1(n22357), .A2(n22356), .A3(n22355), .A4(n22354), .ZN(
        n33225) );
  XNOR2_X1 U26223 ( .A(n33225), .B(\fmem_data[16][3] ), .ZN(n26270) );
  OAI22_X1 U26224 ( .A1(n34038), .A2(n34501), .B1(n26270), .B2(n34499), .ZN(
        n29528) );
  XNOR2_X1 U26225 ( .A(n35240), .B(\fmem_data[3][1] ), .ZN(n32189) );
  XNOR2_X1 U26226 ( .A(n35355), .B(\fmem_data[10][1] ), .ZN(n32730) );
  OAI21_X1 U26227 ( .B1(n29522), .B2(n29521), .A(n29520), .ZN(n22362) );
  NAND2_X1 U26228 ( .A1(n29522), .A2(n29521), .ZN(n22361) );
  NAND2_X1 U26229 ( .A1(n22362), .A2(n22361), .ZN(n24843) );
  AOI22_X1 U26230 ( .A1(n27713), .A2(\xmem_data[0][5] ), .B1(n29640), .B2(
        \xmem_data[1][5] ), .ZN(n22384) );
  AOI22_X1 U26231 ( .A1(n29726), .A2(\xmem_data[6][5] ), .B1(n30901), .B2(
        \xmem_data[7][5] ), .ZN(n22365) );
  AOI22_X1 U26232 ( .A1(n29382), .A2(\xmem_data[4][5] ), .B1(n28724), .B2(
        \xmem_data[5][5] ), .ZN(n22364) );
  AOI22_X1 U26233 ( .A1(n7446), .A2(\xmem_data[2][5] ), .B1(n28701), .B2(
        \xmem_data[3][5] ), .ZN(n22363) );
  NAND3_X1 U26234 ( .A1(n22365), .A2(n22364), .A3(n22363), .ZN(n22381) );
  AOI22_X1 U26235 ( .A1(n29769), .A2(\xmem_data[24][5] ), .B1(n30090), .B2(
        \xmem_data[25][5] ), .ZN(n22369) );
  AOI22_X1 U26236 ( .A1(n27756), .A2(\xmem_data[26][5] ), .B1(n25607), .B2(
        \xmem_data[27][5] ), .ZN(n22368) );
  AOI22_X1 U26237 ( .A1(n3167), .A2(\xmem_data[28][5] ), .B1(n3188), .B2(
        \xmem_data[29][5] ), .ZN(n22367) );
  AOI22_X1 U26238 ( .A1(n30684), .A2(\xmem_data[30][5] ), .B1(n27825), .B2(
        \xmem_data[31][5] ), .ZN(n22366) );
  NAND4_X1 U26239 ( .A1(n22369), .A2(n22368), .A3(n22367), .A4(n22366), .ZN(
        n22380) );
  AOI22_X1 U26240 ( .A1(n29419), .A2(\xmem_data[8][5] ), .B1(n27743), .B2(
        \xmem_data[9][5] ), .ZN(n22373) );
  AOI22_X1 U26241 ( .A1(n27742), .A2(\xmem_data[10][5] ), .B1(n3149), .B2(
        \xmem_data[11][5] ), .ZN(n22372) );
  AOI22_X1 U26242 ( .A1(n29421), .A2(\xmem_data[12][5] ), .B1(n27013), .B2(
        \xmem_data[13][5] ), .ZN(n22371) );
  AOI22_X1 U26243 ( .A1(n29628), .A2(\xmem_data[14][5] ), .B1(n30292), .B2(
        \xmem_data[15][5] ), .ZN(n22370) );
  NAND4_X1 U26244 ( .A1(n22373), .A2(n22372), .A3(n22371), .A4(n22370), .ZN(
        n22379) );
  AOI22_X1 U26245 ( .A1(n27771), .A2(\xmem_data[16][5] ), .B1(n29629), .B2(
        \xmem_data[17][5] ), .ZN(n22377) );
  AOI22_X1 U26246 ( .A1(n3223), .A2(\xmem_data[18][5] ), .B1(n3147), .B2(
        \xmem_data[19][5] ), .ZN(n22376) );
  AOI22_X1 U26247 ( .A1(n29647), .A2(\xmem_data[20][5] ), .B1(n30730), .B2(
        \xmem_data[21][5] ), .ZN(n22375) );
  AOI22_X1 U26248 ( .A1(n26879), .A2(\xmem_data[22][5] ), .B1(n27763), .B2(
        \xmem_data[23][5] ), .ZN(n22374) );
  NAND4_X1 U26249 ( .A1(n22377), .A2(n22376), .A3(n22375), .A4(n22374), .ZN(
        n22378) );
  NOR4_X1 U26250 ( .A1(n22379), .A2(n22380), .A3(n22381), .A4(n22378), .ZN(
        n22383) );
  INV_X1 U26251 ( .A(n27778), .ZN(n22382) );
  AOI21_X1 U26252 ( .B1(n22384), .B2(n22383), .A(n22382), .ZN(n22385) );
  INV_X1 U26253 ( .A(n22385), .ZN(n22452) );
  AOI22_X1 U26254 ( .A1(n30076), .A2(\xmem_data[96][5] ), .B1(n30765), .B2(
        \xmem_data[97][5] ), .ZN(n22389) );
  AOI22_X1 U26255 ( .A1(n27804), .A2(\xmem_data[98][5] ), .B1(n30686), .B2(
        \xmem_data[99][5] ), .ZN(n22388) );
  AOI22_X1 U26256 ( .A1(n28725), .A2(\xmem_data[100][5] ), .B1(n27805), .B2(
        \xmem_data[101][5] ), .ZN(n22387) );
  AOI22_X1 U26257 ( .A1(n27806), .A2(\xmem_data[102][5] ), .B1(n28241), .B2(
        \xmem_data[103][5] ), .ZN(n22386) );
  NAND4_X1 U26258 ( .A1(n22389), .A2(n22388), .A3(n22387), .A4(n22386), .ZN(
        n22405) );
  AOI22_X1 U26259 ( .A1(n7451), .A2(\xmem_data[104][5] ), .B1(n27812), .B2(
        \xmem_data[105][5] ), .ZN(n22393) );
  AOI22_X1 U26260 ( .A1(n27814), .A2(\xmem_data[106][5] ), .B1(n27813), .B2(
        \xmem_data[107][5] ), .ZN(n22392) );
  AOI22_X1 U26261 ( .A1(n29788), .A2(\xmem_data[108][5] ), .B1(n30222), .B2(
        \xmem_data[109][5] ), .ZN(n22391) );
  AOI22_X1 U26262 ( .A1(n3392), .A2(\xmem_data[110][5] ), .B1(n27831), .B2(
        \xmem_data[111][5] ), .ZN(n22390) );
  NAND4_X1 U26263 ( .A1(n22393), .A2(n22392), .A3(n22391), .A4(n22390), .ZN(
        n22404) );
  AOI22_X1 U26264 ( .A1(n27834), .A2(\xmem_data[112][5] ), .B1(n27833), .B2(
        \xmem_data[113][5] ), .ZN(n22397) );
  AOI22_X1 U26265 ( .A1(n3223), .A2(\xmem_data[114][5] ), .B1(n3140), .B2(
        \xmem_data[115][5] ), .ZN(n22396) );
  AOI22_X1 U26266 ( .A1(n3249), .A2(\xmem_data[116][5] ), .B1(n29646), .B2(
        \xmem_data[117][5] ), .ZN(n22395) );
  AOI22_X1 U26267 ( .A1(n29500), .A2(\xmem_data[118][5] ), .B1(n27763), .B2(
        \xmem_data[119][5] ), .ZN(n22394) );
  NAND4_X1 U26268 ( .A1(n22397), .A2(n22396), .A3(n22395), .A4(n22394), .ZN(
        n22403) );
  AOI22_X1 U26269 ( .A1(n30250), .A2(\xmem_data[120][5] ), .B1(n26884), .B2(
        \xmem_data[121][5] ), .ZN(n22401) );
  AOI22_X1 U26270 ( .A1(n27819), .A2(\xmem_data[122][5] ), .B1(n3465), .B2(
        \xmem_data[123][5] ), .ZN(n22400) );
  AOI22_X1 U26271 ( .A1(n3161), .A2(\xmem_data[124][5] ), .B1(n3184), .B2(
        \xmem_data[125][5] ), .ZN(n22399) );
  AOI22_X1 U26272 ( .A1(n30715), .A2(\xmem_data[126][5] ), .B1(n25678), .B2(
        \xmem_data[127][5] ), .ZN(n22398) );
  NAND4_X1 U26273 ( .A1(n22401), .A2(n22400), .A3(n22399), .A4(n22398), .ZN(
        n22402) );
  NAND2_X1 U26274 ( .A1(n22406), .A2(n27801), .ZN(n22451) );
  AOI22_X1 U26275 ( .A1(n27701), .A2(\xmem_data[80][5] ), .B1(n3170), .B2(
        \xmem_data[81][5] ), .ZN(n22410) );
  AOI22_X1 U26276 ( .A1(n27702), .A2(\xmem_data[82][5] ), .B1(n3140), .B2(
        \xmem_data[83][5] ), .ZN(n22409) );
  AOI22_X1 U26277 ( .A1(n30191), .A2(\xmem_data[84][5] ), .B1(n29646), .B2(
        \xmem_data[85][5] ), .ZN(n22408) );
  AOI22_X1 U26278 ( .A1(n29763), .A2(\xmem_data[86][5] ), .B1(n27763), .B2(
        \xmem_data[87][5] ), .ZN(n22407) );
  NAND4_X1 U26279 ( .A1(n22410), .A2(n22409), .A3(n22408), .A4(n22407), .ZN(
        n22426) );
  AOI22_X1 U26280 ( .A1(n29786), .A2(\xmem_data[72][5] ), .B1(n27723), .B2(
        \xmem_data[73][5] ), .ZN(n22414) );
  AOI22_X1 U26281 ( .A1(n27742), .A2(\xmem_data[74][5] ), .B1(n3149), .B2(
        \xmem_data[75][5] ), .ZN(n22413) );
  AOI22_X1 U26282 ( .A1(n27710), .A2(\xmem_data[76][5] ), .B1(n29753), .B2(
        \xmem_data[77][5] ), .ZN(n22412) );
  AOI22_X1 U26283 ( .A1(n28700), .A2(\xmem_data[78][5] ), .B1(n27708), .B2(
        \xmem_data[79][5] ), .ZN(n22411) );
  NAND4_X1 U26284 ( .A1(n22414), .A2(n22413), .A3(n22412), .A4(n22411), .ZN(
        n22425) );
  AOI22_X1 U26285 ( .A1(n29714), .A2(\xmem_data[88][5] ), .B1(n26884), .B2(
        \xmem_data[89][5] ), .ZN(n22418) );
  AOI22_X1 U26286 ( .A1(n27729), .A2(\xmem_data[90][5] ), .B1(n25607), .B2(
        \xmem_data[91][5] ), .ZN(n22417) );
  AOI22_X1 U26287 ( .A1(n3164), .A2(\xmem_data[92][5] ), .B1(n3186), .B2(
        \xmem_data[93][5] ), .ZN(n22416) );
  AOI22_X1 U26288 ( .A1(n29476), .A2(\xmem_data[94][5] ), .B1(n29410), .B2(
        \xmem_data[95][5] ), .ZN(n22415) );
  NAND4_X1 U26289 ( .A1(n22418), .A2(n22417), .A3(n22416), .A4(n22415), .ZN(
        n22424) );
  AOI22_X1 U26290 ( .A1(n29547), .A2(\xmem_data[64][5] ), .B1(n29721), .B2(
        \xmem_data[65][5] ), .ZN(n22422) );
  AOI22_X1 U26291 ( .A1(n27714), .A2(\xmem_data[66][5] ), .B1(n20817), .B2(
        \xmem_data[67][5] ), .ZN(n22421) );
  AOI22_X1 U26292 ( .A1(n27716), .A2(\xmem_data[68][5] ), .B1(n27715), .B2(
        \xmem_data[69][5] ), .ZN(n22420) );
  AOI22_X1 U26293 ( .A1(n27718), .A2(\xmem_data[70][5] ), .B1(n27717), .B2(
        \xmem_data[71][5] ), .ZN(n22419) );
  NAND4_X1 U26294 ( .A1(n22422), .A2(n22421), .A3(n22420), .A4(n22419), .ZN(
        n22423) );
  OR4_X1 U26295 ( .A1(n22426), .A2(n22425), .A3(n22424), .A4(n22423), .ZN(
        n22427) );
  NAND2_X1 U26296 ( .A1(n22427), .A2(n27839), .ZN(n22450) );
  AOI22_X1 U26297 ( .A1(n30766), .A2(\xmem_data[32][5] ), .B1(n30266), .B2(
        \xmem_data[33][5] ), .ZN(n22431) );
  AOI22_X1 U26298 ( .A1(n27714), .A2(\xmem_data[34][5] ), .B1(n29054), .B2(
        \xmem_data[35][5] ), .ZN(n22430) );
  AOI22_X1 U26299 ( .A1(n27716), .A2(\xmem_data[36][5] ), .B1(n27715), .B2(
        \xmem_data[37][5] ), .ZN(n22429) );
  AOI22_X1 U26300 ( .A1(n27718), .A2(\xmem_data[38][5] ), .B1(n27717), .B2(
        \xmem_data[39][5] ), .ZN(n22428) );
  NAND4_X1 U26301 ( .A1(n22431), .A2(n22430), .A3(n22429), .A4(n22428), .ZN(
        n22447) );
  AOI22_X1 U26302 ( .A1(n29786), .A2(\xmem_data[40][5] ), .B1(n27723), .B2(
        \xmem_data[41][5] ), .ZN(n22435) );
  AOI22_X1 U26303 ( .A1(n27742), .A2(\xmem_data[42][5] ), .B1(n3149), .B2(
        \xmem_data[43][5] ), .ZN(n22434) );
  AOI22_X1 U26304 ( .A1(n27710), .A2(\xmem_data[44][5] ), .B1(n27832), .B2(
        \xmem_data[45][5] ), .ZN(n22433) );
  AOI22_X1 U26305 ( .A1(n30215), .A2(\xmem_data[46][5] ), .B1(n27708), .B2(
        \xmem_data[47][5] ), .ZN(n22432) );
  NAND4_X1 U26306 ( .A1(n22432), .A2(n22434), .A3(n22433), .A4(n22435), .ZN(
        n22446) );
  AOI22_X1 U26307 ( .A1(n27701), .A2(\xmem_data[48][5] ), .B1(n30293), .B2(
        \xmem_data[49][5] ), .ZN(n22439) );
  AOI22_X1 U26308 ( .A1(n27702), .A2(\xmem_data[50][5] ), .B1(n3146), .B2(
        \xmem_data[51][5] ), .ZN(n22438) );
  AOI22_X1 U26309 ( .A1(n29705), .A2(\xmem_data[52][5] ), .B1(n29646), .B2(
        \xmem_data[53][5] ), .ZN(n22437) );
  AOI22_X1 U26310 ( .A1(n26879), .A2(\xmem_data[54][5] ), .B1(n27911), .B2(
        \xmem_data[55][5] ), .ZN(n22436) );
  NAND4_X1 U26311 ( .A1(n22439), .A2(n22438), .A3(n22437), .A4(n22436), .ZN(
        n22445) );
  AOI22_X1 U26312 ( .A1(n30665), .A2(\xmem_data[56][5] ), .B1(n30237), .B2(
        \xmem_data[57][5] ), .ZN(n22443) );
  AOI22_X1 U26313 ( .A1(n27729), .A2(\xmem_data[58][5] ), .B1(n30543), .B2(
        \xmem_data[59][5] ), .ZN(n22442) );
  AOI22_X1 U26314 ( .A1(n3168), .A2(\xmem_data[60][5] ), .B1(n3188), .B2(
        \xmem_data[61][5] ), .ZN(n22441) );
  AOI22_X1 U26315 ( .A1(n29610), .A2(\xmem_data[62][5] ), .B1(n29439), .B2(
        \xmem_data[63][5] ), .ZN(n22440) );
  NAND4_X1 U26316 ( .A1(n22443), .A2(n22442), .A3(n22441), .A4(n22440), .ZN(
        n22444) );
  OR4_X1 U26317 ( .A1(n22444), .A2(n22446), .A3(n22445), .A4(n22447), .ZN(
        n22448) );
  NAND2_X1 U26318 ( .A1(n22448), .A2(n27737), .ZN(n22449) );
  XNOR2_X1 U26319 ( .A(n31980), .B(\fmem_data[27][3] ), .ZN(n31894) );
  XNOR2_X1 U26320 ( .A(n3257), .B(\fmem_data[19][5] ), .ZN(n32183) );
  XNOR2_X1 U26321 ( .A(n35359), .B(\fmem_data[7][1] ), .ZN(n32181) );
  INV_X1 U26322 ( .A(n36218), .ZN(n22455) );
  NOR2_X1 U26323 ( .A1(n22455), .A2(\fmem_data[7][0] ), .ZN(n22456) );
  XNOR2_X1 U26324 ( .A(n24843), .B(n24842), .ZN(n22779) );
  AOI22_X1 U26325 ( .A1(n25708), .A2(\xmem_data[4][3] ), .B1(n24555), .B2(
        \xmem_data[5][3] ), .ZN(n22458) );
  AOI22_X1 U26326 ( .A1(n29271), .A2(\xmem_data[7][3] ), .B1(\xmem_data[3][3] ), .B2(n29180), .ZN(n22457) );
  NAND2_X1 U26327 ( .A1(n22458), .A2(n22457), .ZN(n22469) );
  AOI22_X1 U26328 ( .A1(n3335), .A2(\xmem_data[24][3] ), .B1(n29286), .B2(
        \xmem_data[25][3] ), .ZN(n22462) );
  AOI22_X1 U26329 ( .A1(n28318), .A2(\xmem_data[26][3] ), .B1(n3222), .B2(
        \xmem_data[27][3] ), .ZN(n22461) );
  AOI22_X1 U26330 ( .A1(n29288), .A2(\xmem_data[28][3] ), .B1(n27444), .B2(
        \xmem_data[29][3] ), .ZN(n22460) );
  AOI22_X1 U26331 ( .A1(n29289), .A2(\xmem_data[30][3] ), .B1(n27994), .B2(
        \xmem_data[31][3] ), .ZN(n22459) );
  NAND4_X1 U26332 ( .A1(n22462), .A2(n22461), .A3(n22460), .A4(n22459), .ZN(
        n22468) );
  AOI22_X1 U26333 ( .A1(n29297), .A2(\xmem_data[16][3] ), .B1(n25583), .B2(
        \xmem_data[17][3] ), .ZN(n22466) );
  AOI22_X1 U26334 ( .A1(n20552), .A2(\xmem_data[18][3] ), .B1(n28468), .B2(
        \xmem_data[19][3] ), .ZN(n22465) );
  AOI22_X1 U26335 ( .A1(n29298), .A2(\xmem_data[20][3] ), .B1(n17050), .B2(
        \xmem_data[21][3] ), .ZN(n22464) );
  AOI22_X1 U26336 ( .A1(n24526), .A2(\xmem_data[22][3] ), .B1(n28366), .B2(
        \xmem_data[23][3] ), .ZN(n22463) );
  NAND4_X1 U26337 ( .A1(n22466), .A2(n22465), .A3(n22464), .A4(n22463), .ZN(
        n22467) );
  OR3_X1 U26338 ( .A1(n22469), .A2(n22468), .A3(n22467), .ZN(n22481) );
  AOI22_X1 U26339 ( .A1(n25607), .A2(\xmem_data[8][3] ), .B1(n29279), .B2(
        \xmem_data[9][3] ), .ZN(n22473) );
  AOI22_X1 U26340 ( .A1(n23717), .A2(\xmem_data[10][3] ), .B1(n24645), .B2(
        \xmem_data[11][3] ), .ZN(n22472) );
  AOI22_X1 U26341 ( .A1(n27825), .A2(\xmem_data[12][3] ), .B1(n29280), .B2(
        \xmem_data[13][3] ), .ZN(n22471) );
  AOI22_X1 U26342 ( .A1(n3325), .A2(\xmem_data[14][3] ), .B1(n20506), .B2(
        \xmem_data[15][3] ), .ZN(n22470) );
  NAND4_X1 U26343 ( .A1(n22473), .A2(n22472), .A3(n22471), .A4(n22470), .ZN(
        n22477) );
  NAND2_X1 U26344 ( .A1(n28050), .A2(\xmem_data[2][3] ), .ZN(n22475) );
  NAND2_X1 U26345 ( .A1(n3146), .A2(\xmem_data[0][3] ), .ZN(n22474) );
  NAND2_X1 U26346 ( .A1(n22475), .A2(n22474), .ZN(n22476) );
  NOR2_X1 U26347 ( .A1(n22477), .A2(n22476), .ZN(n22479) );
  AOI21_X1 U26348 ( .B1(n3231), .B2(\xmem_data[1][3] ), .A(n22482), .ZN(n22548) );
  AOI22_X1 U26349 ( .A1(n29231), .A2(\xmem_data[96][3] ), .B1(n28007), .B2(
        \xmem_data[97][3] ), .ZN(n22486) );
  AOI22_X1 U26350 ( .A1(n27447), .A2(\xmem_data[98][3] ), .B1(n20546), .B2(
        \xmem_data[99][3] ), .ZN(n22485) );
  AOI22_X1 U26351 ( .A1(n28051), .A2(\xmem_data[100][3] ), .B1(n29232), .B2(
        \xmem_data[101][3] ), .ZN(n22484) );
  AOI22_X1 U26352 ( .A1(n25459), .A2(\xmem_data[102][3] ), .B1(n29271), .B2(
        \xmem_data[103][3] ), .ZN(n22483) );
  NAND4_X1 U26353 ( .A1(n22486), .A2(n22485), .A3(n22484), .A4(n22483), .ZN(
        n22502) );
  AOI22_X1 U26354 ( .A1(n3466), .A2(\xmem_data[104][3] ), .B1(n20543), .B2(
        \xmem_data[105][3] ), .ZN(n22490) );
  AOI22_X1 U26355 ( .A1(n13149), .A2(\xmem_data[106][3] ), .B1(n24219), .B2(
        \xmem_data[107][3] ), .ZN(n22489) );
  AOI22_X1 U26356 ( .A1(n29239), .A2(\xmem_data[108][3] ), .B1(n29238), .B2(
        \xmem_data[109][3] ), .ZN(n22488) );
  AOI22_X1 U26357 ( .A1(n29240), .A2(\xmem_data[110][3] ), .B1(n28327), .B2(
        \xmem_data[111][3] ), .ZN(n22487) );
  NAND4_X1 U26358 ( .A1(n22490), .A2(n22489), .A3(n22488), .A4(n22487), .ZN(
        n22501) );
  AOI22_X1 U26359 ( .A1(n29246), .A2(\xmem_data[112][3] ), .B1(n29245), .B2(
        \xmem_data[113][3] ), .ZN(n22494) );
  AOI22_X1 U26360 ( .A1(n27542), .A2(\xmem_data[114][3] ), .B1(n29247), .B2(
        \xmem_data[115][3] ), .ZN(n22493) );
  AOI22_X1 U26361 ( .A1(n28241), .A2(\xmem_data[116][3] ), .B1(n29248), .B2(
        \xmem_data[117][3] ), .ZN(n22492) );
  AOI22_X1 U26362 ( .A1(n20986), .A2(\xmem_data[118][3] ), .B1(n20709), .B2(
        \xmem_data[119][3] ), .ZN(n22491) );
  NAND4_X1 U26363 ( .A1(n22494), .A2(n22493), .A3(n22492), .A4(n22491), .ZN(
        n22500) );
  AOI22_X1 U26364 ( .A1(n3412), .A2(\xmem_data[120][3] ), .B1(n29253), .B2(
        \xmem_data[121][3] ), .ZN(n22498) );
  AOI22_X1 U26365 ( .A1(n29254), .A2(\xmem_data[122][3] ), .B1(n3218), .B2(
        \xmem_data[123][3] ), .ZN(n22497) );
  AOI22_X1 U26366 ( .A1(n29256), .A2(\xmem_data[124][3] ), .B1(n29255), .B2(
        \xmem_data[125][3] ), .ZN(n22496) );
  AOI22_X1 U26367 ( .A1(n29257), .A2(\xmem_data[126][3] ), .B1(n25486), .B2(
        \xmem_data[127][3] ), .ZN(n22495) );
  NAND4_X1 U26368 ( .A1(n22498), .A2(n22497), .A3(n22496), .A4(n22495), .ZN(
        n22499) );
  OR4_X1 U26369 ( .A1(n22502), .A2(n22501), .A3(n22500), .A4(n22499), .ZN(
        n22524) );
  AOI22_X1 U26370 ( .A1(n29231), .A2(\xmem_data[64][3] ), .B1(n25492), .B2(
        \xmem_data[65][3] ), .ZN(n22506) );
  AOI22_X1 U26371 ( .A1(n24554), .A2(\xmem_data[66][3] ), .B1(n27943), .B2(
        \xmem_data[67][3] ), .ZN(n22505) );
  AOI22_X1 U26372 ( .A1(n29179), .A2(\xmem_data[68][3] ), .B1(n29232), .B2(
        \xmem_data[69][3] ), .ZN(n22504) );
  AOI22_X1 U26373 ( .A1(n16986), .A2(\xmem_data[70][3] ), .B1(n20544), .B2(
        \xmem_data[71][3] ), .ZN(n22503) );
  NAND4_X1 U26374 ( .A1(n22506), .A2(n22505), .A3(n22504), .A4(n22503), .ZN(
        n22522) );
  AOI22_X1 U26375 ( .A1(n24213), .A2(\xmem_data[72][3] ), .B1(n27989), .B2(
        \xmem_data[73][3] ), .ZN(n22510) );
  AOI22_X1 U26376 ( .A1(n24509), .A2(\xmem_data[74][3] ), .B1(n28492), .B2(
        \xmem_data[75][3] ), .ZN(n22509) );
  AOI22_X1 U26377 ( .A1(n29239), .A2(\xmem_data[76][3] ), .B1(n29238), .B2(
        \xmem_data[77][3] ), .ZN(n22508) );
  AOI22_X1 U26378 ( .A1(n29240), .A2(\xmem_data[78][3] ), .B1(n3372), .B2(
        \xmem_data[79][3] ), .ZN(n22507) );
  NAND4_X1 U26379 ( .A1(n22510), .A2(n22509), .A3(n22508), .A4(n22507), .ZN(
        n22521) );
  AOI22_X1 U26380 ( .A1(n29246), .A2(\xmem_data[80][3] ), .B1(n29245), .B2(
        \xmem_data[81][3] ), .ZN(n22514) );
  AOI22_X1 U26381 ( .A1(n27542), .A2(\xmem_data[82][3] ), .B1(n29247), .B2(
        \xmem_data[83][3] ), .ZN(n22513) );
  AOI22_X1 U26382 ( .A1(n21060), .A2(\xmem_data[84][3] ), .B1(n29248), .B2(
        \xmem_data[85][3] ), .ZN(n22512) );
  AOI22_X1 U26383 ( .A1(n27925), .A2(\xmem_data[86][3] ), .B1(n29118), .B2(
        \xmem_data[87][3] ), .ZN(n22511) );
  NAND4_X1 U26384 ( .A1(n22514), .A2(n22513), .A3(n22512), .A4(n22511), .ZN(
        n22520) );
  AOI22_X1 U26385 ( .A1(n23754), .A2(\xmem_data[88][3] ), .B1(n29253), .B2(
        \xmem_data[89][3] ), .ZN(n22518) );
  AOI22_X1 U26386 ( .A1(n29254), .A2(\xmem_data[90][3] ), .B1(n3218), .B2(
        \xmem_data[91][3] ), .ZN(n22517) );
  AOI22_X1 U26387 ( .A1(n29256), .A2(\xmem_data[92][3] ), .B1(n29255), .B2(
        \xmem_data[93][3] ), .ZN(n22516) );
  AOI22_X1 U26388 ( .A1(n29257), .A2(\xmem_data[94][3] ), .B1(n22669), .B2(
        \xmem_data[95][3] ), .ZN(n22515) );
  NAND4_X1 U26389 ( .A1(n22518), .A2(n22517), .A3(n22516), .A4(n22515), .ZN(
        n22519) );
  OR4_X1 U26390 ( .A1(n22522), .A2(n22521), .A3(n22520), .A4(n22519), .ZN(
        n22523) );
  AOI22_X1 U26391 ( .A1(n29269), .A2(n22524), .B1(n29267), .B2(n22523), .ZN(
        n22547) );
  AOI22_X1 U26392 ( .A1(n3281), .A2(\xmem_data[32][3] ), .B1(n28045), .B2(
        \xmem_data[33][3] ), .ZN(n22528) );
  AOI22_X1 U26393 ( .A1(n25670), .A2(\xmem_data[34][3] ), .B1(n29307), .B2(
        \xmem_data[35][3] ), .ZN(n22527) );
  AOI22_X1 U26394 ( .A1(n29308), .A2(\xmem_data[36][3] ), .B1(n21015), .B2(
        \xmem_data[37][3] ), .ZN(n22526) );
  AOI22_X1 U26395 ( .A1(n29310), .A2(\xmem_data[38][3] ), .B1(n29309), .B2(
        \xmem_data[39][3] ), .ZN(n22525) );
  NAND4_X1 U26396 ( .A1(n22528), .A2(n22527), .A3(n22526), .A4(n22525), .ZN(
        n22544) );
  AOI22_X1 U26397 ( .A1(n3158), .A2(\xmem_data[40][3] ), .B1(n27989), .B2(
        \xmem_data[41][3] ), .ZN(n22532) );
  AOI22_X1 U26398 ( .A1(n29317), .A2(\xmem_data[42][3] ), .B1(n29316), .B2(
        \xmem_data[43][3] ), .ZN(n22531) );
  AOI22_X1 U26399 ( .A1(n29319), .A2(\xmem_data[44][3] ), .B1(n29318), .B2(
        \xmem_data[45][3] ), .ZN(n22530) );
  AOI22_X1 U26400 ( .A1(n25521), .A2(\xmem_data[46][3] ), .B1(n25581), .B2(
        \xmem_data[47][3] ), .ZN(n22529) );
  NAND4_X1 U26401 ( .A1(n22532), .A2(n22531), .A3(n22530), .A4(n22529), .ZN(
        n22543) );
  AOI22_X1 U26402 ( .A1(n29324), .A2(\xmem_data[48][3] ), .B1(n14975), .B2(
        \xmem_data[49][3] ), .ZN(n22536) );
  AOI22_X1 U26403 ( .A1(n29325), .A2(\xmem_data[50][3] ), .B1(n28468), .B2(
        \xmem_data[51][3] ), .ZN(n22535) );
  AOI22_X1 U26404 ( .A1(n29327), .A2(\xmem_data[52][3] ), .B1(n29326), .B2(
        \xmem_data[53][3] ), .ZN(n22534) );
  AOI22_X1 U26405 ( .A1(n27500), .A2(\xmem_data[54][3] ), .B1(n29328), .B2(
        \xmem_data[55][3] ), .ZN(n22533) );
  NAND4_X1 U26406 ( .A1(n22536), .A2(n22535), .A3(n22534), .A4(n22533), .ZN(
        n22542) );
  AOI22_X1 U26407 ( .A1(n3384), .A2(\xmem_data[56][3] ), .B1(n30863), .B2(
        \xmem_data[57][3] ), .ZN(n22540) );
  AOI22_X1 U26408 ( .A1(n24443), .A2(\xmem_data[58][3] ), .B1(n3221), .B2(
        \xmem_data[59][3] ), .ZN(n22539) );
  AOI22_X1 U26409 ( .A1(n25693), .A2(\xmem_data[60][3] ), .B1(n23739), .B2(
        \xmem_data[61][3] ), .ZN(n22538) );
  AOI22_X1 U26410 ( .A1(n30606), .A2(\xmem_data[62][3] ), .B1(n24140), .B2(
        \xmem_data[63][3] ), .ZN(n22537) );
  NAND4_X1 U26411 ( .A1(n22540), .A2(n22539), .A3(n22538), .A4(n22537), .ZN(
        n22541) );
  OR4_X1 U26412 ( .A1(n22544), .A2(n22543), .A3(n22542), .A4(n22541), .ZN(
        n22545) );
  NAND2_X1 U26413 ( .A1(n22545), .A2(n29343), .ZN(n22546) );
  AOI22_X1 U26414 ( .A1(n30295), .A2(\xmem_data[0][4] ), .B1(n28007), .B2(
        \xmem_data[1][4] ), .ZN(n22570) );
  AOI22_X1 U26415 ( .A1(n29451), .A2(\xmem_data[4][4] ), .B1(n20958), .B2(
        \xmem_data[5][4] ), .ZN(n22551) );
  AOI22_X1 U26416 ( .A1(n29272), .A2(\xmem_data[6][4] ), .B1(n29271), .B2(
        \xmem_data[7][4] ), .ZN(n22550) );
  AOI22_X1 U26417 ( .A1(n27447), .A2(\xmem_data[2][4] ), .B1(n25481), .B2(
        \xmem_data[3][4] ), .ZN(n22549) );
  NAND3_X1 U26418 ( .A1(n22551), .A2(n22550), .A3(n22549), .ZN(n22562) );
  AOI22_X1 U26419 ( .A1(n24213), .A2(\xmem_data[8][4] ), .B1(n29279), .B2(
        \xmem_data[9][4] ), .ZN(n22555) );
  AOI22_X1 U26420 ( .A1(n23717), .A2(\xmem_data[10][4] ), .B1(n29316), .B2(
        \xmem_data[11][4] ), .ZN(n22554) );
  AOI22_X1 U26421 ( .A1(n31255), .A2(\xmem_data[12][4] ), .B1(n29280), .B2(
        \xmem_data[13][4] ), .ZN(n22553) );
  AOI22_X1 U26422 ( .A1(n28061), .A2(\xmem_data[14][4] ), .B1(n25581), .B2(
        \xmem_data[15][4] ), .ZN(n22552) );
  NAND4_X1 U26423 ( .A1(n22555), .A2(n22554), .A3(n22553), .A4(n22552), .ZN(
        n22561) );
  AOI22_X1 U26424 ( .A1(n3334), .A2(\xmem_data[24][4] ), .B1(n29286), .B2(
        \xmem_data[25][4] ), .ZN(n22559) );
  AOI22_X1 U26425 ( .A1(n24443), .A2(\xmem_data[26][4] ), .B1(n3219), .B2(
        \xmem_data[27][4] ), .ZN(n22558) );
  AOI22_X1 U26426 ( .A1(n29288), .A2(\xmem_data[28][4] ), .B1(n24207), .B2(
        \xmem_data[29][4] ), .ZN(n22557) );
  AOI22_X1 U26427 ( .A1(n29289), .A2(\xmem_data[30][4] ), .B1(n27903), .B2(
        \xmem_data[31][4] ), .ZN(n22556) );
  NAND4_X1 U26428 ( .A1(n22559), .A2(n22558), .A3(n22557), .A4(n22556), .ZN(
        n22560) );
  OR3_X1 U26429 ( .A1(n22562), .A2(n22561), .A3(n22560), .ZN(n22568) );
  AOI22_X1 U26430 ( .A1(n29297), .A2(\xmem_data[16][4] ), .B1(n20983), .B2(
        \xmem_data[17][4] ), .ZN(n22566) );
  AOI22_X1 U26431 ( .A1(n29325), .A2(\xmem_data[18][4] ), .B1(n31256), .B2(
        \xmem_data[19][4] ), .ZN(n22565) );
  AOI22_X1 U26432 ( .A1(n29298), .A2(\xmem_data[20][4] ), .B1(n31261), .B2(
        \xmem_data[21][4] ), .ZN(n22564) );
  AOI22_X1 U26433 ( .A1(n29124), .A2(\xmem_data[22][4] ), .B1(n25629), .B2(
        \xmem_data[23][4] ), .ZN(n22563) );
  NAND4_X1 U26434 ( .A1(n22566), .A2(n22565), .A3(n22564), .A4(n22563), .ZN(
        n22567) );
  NOR2_X1 U26435 ( .A1(n22568), .A2(n22567), .ZN(n22569) );
  AOI21_X1 U26436 ( .B1(n22570), .B2(n22569), .A(n29341), .ZN(n22641) );
  AOI22_X1 U26437 ( .A1(n24630), .A2(\xmem_data[120][4] ), .B1(n29253), .B2(
        \xmem_data[121][4] ), .ZN(n22574) );
  AOI22_X1 U26438 ( .A1(n29254), .A2(\xmem_data[122][4] ), .B1(n3220), .B2(
        \xmem_data[123][4] ), .ZN(n22573) );
  AOI22_X1 U26439 ( .A1(n29256), .A2(\xmem_data[124][4] ), .B1(n29255), .B2(
        \xmem_data[125][4] ), .ZN(n22572) );
  AOI22_X1 U26440 ( .A1(n29257), .A2(\xmem_data[126][4] ), .B1(n22711), .B2(
        \xmem_data[127][4] ), .ZN(n22571) );
  NAND4_X1 U26441 ( .A1(n22574), .A2(n22573), .A3(n22572), .A4(n22571), .ZN(
        n22590) );
  AOI22_X1 U26442 ( .A1(n29246), .A2(\xmem_data[112][4] ), .B1(n29245), .B2(
        \xmem_data[113][4] ), .ZN(n22578) );
  AOI22_X1 U26443 ( .A1(n25582), .A2(\xmem_data[114][4] ), .B1(n29247), .B2(
        \xmem_data[115][4] ), .ZN(n22577) );
  AOI22_X1 U26444 ( .A1(n23753), .A2(\xmem_data[116][4] ), .B1(n29248), .B2(
        \xmem_data[117][4] ), .ZN(n22576) );
  AOI22_X1 U26445 ( .A1(n30909), .A2(\xmem_data[118][4] ), .B1(n29328), .B2(
        \xmem_data[119][4] ), .ZN(n22575) );
  NAND4_X1 U26446 ( .A1(n22578), .A2(n22577), .A3(n22576), .A4(n22575), .ZN(
        n22589) );
  AOI22_X1 U26447 ( .A1(n29231), .A2(\xmem_data[96][4] ), .B1(n30877), .B2(
        \xmem_data[97][4] ), .ZN(n22582) );
  AOI22_X1 U26448 ( .A1(n27447), .A2(\xmem_data[98][4] ), .B1(n3357), .B2(
        \xmem_data[99][4] ), .ZN(n22581) );
  AOI22_X1 U26449 ( .A1(n24556), .A2(\xmem_data[100][4] ), .B1(n29232), .B2(
        \xmem_data[101][4] ), .ZN(n22580) );
  AOI22_X1 U26450 ( .A1(n28334), .A2(\xmem_data[102][4] ), .B1(n14999), .B2(
        \xmem_data[103][4] ), .ZN(n22579) );
  NAND4_X1 U26451 ( .A1(n22582), .A2(n22581), .A3(n22580), .A4(n22579), .ZN(
        n22588) );
  AOI22_X1 U26452 ( .A1(n29396), .A2(\xmem_data[104][4] ), .B1(n23716), .B2(
        \xmem_data[105][4] ), .ZN(n22586) );
  AOI22_X1 U26453 ( .A1(n20585), .A2(\xmem_data[106][4] ), .B1(n29316), .B2(
        \xmem_data[107][4] ), .ZN(n22585) );
  AOI22_X1 U26454 ( .A1(n29239), .A2(\xmem_data[108][4] ), .B1(n29238), .B2(
        \xmem_data[109][4] ), .ZN(n22584) );
  AOI22_X1 U26455 ( .A1(n29240), .A2(\xmem_data[110][4] ), .B1(n28060), .B2(
        \xmem_data[111][4] ), .ZN(n22583) );
  NAND4_X1 U26456 ( .A1(n22586), .A2(n22585), .A3(n22584), .A4(n22583), .ZN(
        n22587) );
  OR4_X1 U26457 ( .A1(n22590), .A2(n22589), .A3(n22588), .A4(n22587), .ZN(
        n22591) );
  AND2_X1 U26458 ( .A1(n22591), .A2(n29269), .ZN(n22640) );
  AOI22_X1 U26459 ( .A1(n29324), .A2(\xmem_data[48][4] ), .B1(n28983), .B2(
        \xmem_data[49][4] ), .ZN(n22595) );
  AOI22_X1 U26460 ( .A1(n29325), .A2(\xmem_data[50][4] ), .B1(n28979), .B2(
        \xmem_data[51][4] ), .ZN(n22594) );
  AOI22_X1 U26461 ( .A1(n29327), .A2(\xmem_data[52][4] ), .B1(n29326), .B2(
        \xmem_data[53][4] ), .ZN(n22593) );
  AOI22_X1 U26462 ( .A1(n25358), .A2(\xmem_data[54][4] ), .B1(n29328), .B2(
        \xmem_data[55][4] ), .ZN(n22592) );
  NAND4_X1 U26463 ( .A1(n22595), .A2(n22594), .A3(n22593), .A4(n22592), .ZN(
        n22596) );
  NAND2_X1 U26464 ( .A1(n22596), .A2(n29343), .ZN(n22638) );
  AOI22_X1 U26465 ( .A1(n30543), .A2(\xmem_data[40][4] ), .B1(n24134), .B2(
        \xmem_data[41][4] ), .ZN(n22600) );
  AOI22_X1 U26466 ( .A1(n29317), .A2(\xmem_data[42][4] ), .B1(n29316), .B2(
        \xmem_data[43][4] ), .ZN(n22599) );
  AOI22_X1 U26467 ( .A1(n29319), .A2(\xmem_data[44][4] ), .B1(n29318), .B2(
        \xmem_data[45][4] ), .ZN(n22598) );
  AOI22_X1 U26468 ( .A1(n24220), .A2(\xmem_data[46][4] ), .B1(n24222), .B2(
        \xmem_data[47][4] ), .ZN(n22597) );
  NAND4_X1 U26469 ( .A1(n22600), .A2(n22599), .A3(n22598), .A4(n22597), .ZN(
        n22606) );
  AOI22_X1 U26470 ( .A1(n28344), .A2(\xmem_data[32][4] ), .B1(n25450), .B2(
        \xmem_data[33][4] ), .ZN(n22604) );
  AOI22_X1 U26471 ( .A1(n27551), .A2(\xmem_data[34][4] ), .B1(n29307), .B2(
        \xmem_data[35][4] ), .ZN(n22603) );
  AOI22_X1 U26472 ( .A1(n29308), .A2(\xmem_data[36][4] ), .B1(n14998), .B2(
        \xmem_data[37][4] ), .ZN(n22602) );
  AOI22_X1 U26473 ( .A1(n29310), .A2(\xmem_data[38][4] ), .B1(n29309), .B2(
        \xmem_data[39][4] ), .ZN(n22601) );
  NAND4_X1 U26474 ( .A1(n22604), .A2(n22603), .A3(n22602), .A4(n22601), .ZN(
        n22605) );
  OR2_X1 U26475 ( .A1(n22606), .A2(n22605), .ZN(n22612) );
  AOI22_X1 U26476 ( .A1(n3383), .A2(\xmem_data[56][4] ), .B1(n28501), .B2(
        \xmem_data[57][4] ), .ZN(n22610) );
  AOI22_X1 U26477 ( .A1(n27502), .A2(\xmem_data[58][4] ), .B1(n3218), .B2(
        \xmem_data[59][4] ), .ZN(n22609) );
  AOI22_X1 U26478 ( .A1(n25612), .A2(\xmem_data[60][4] ), .B1(n20723), .B2(
        \xmem_data[61][4] ), .ZN(n22608) );
  AOI22_X1 U26479 ( .A1(n30883), .A2(\xmem_data[62][4] ), .B1(n23811), .B2(
        \xmem_data[63][4] ), .ZN(n22607) );
  NAND4_X1 U26480 ( .A1(n22610), .A2(n22609), .A3(n22608), .A4(n22607), .ZN(
        n22611) );
  AOI22_X1 U26481 ( .A1(n3383), .A2(\xmem_data[88][4] ), .B1(n14875), .B2(
        \xmem_data[89][4] ), .ZN(n22616) );
  AOI22_X1 U26482 ( .A1(n28355), .A2(\xmem_data[90][4] ), .B1(n3219), .B2(
        \xmem_data[91][4] ), .ZN(n22615) );
  AOI22_X1 U26483 ( .A1(n25731), .A2(\xmem_data[92][4] ), .B1(n31367), .B2(
        \xmem_data[93][4] ), .ZN(n22614) );
  AOI22_X1 U26484 ( .A1(n27938), .A2(\xmem_data[94][4] ), .B1(n22759), .B2(
        \xmem_data[95][4] ), .ZN(n22613) );
  NAND4_X1 U26485 ( .A1(n22616), .A2(n22615), .A3(n22614), .A4(n22613), .ZN(
        n22628) );
  AOI22_X1 U26486 ( .A1(n29605), .A2(\xmem_data[72][4] ), .B1(n3213), .B2(
        \xmem_data[73][4] ), .ZN(n22620) );
  AOI22_X1 U26487 ( .A1(n29317), .A2(\xmem_data[74][4] ), .B1(n29316), .B2(
        \xmem_data[75][4] ), .ZN(n22619) );
  AOI22_X1 U26488 ( .A1(n29319), .A2(\xmem_data[76][4] ), .B1(n29318), .B2(
        \xmem_data[77][4] ), .ZN(n22618) );
  AOI22_X1 U26489 ( .A1(n3206), .A2(\xmem_data[78][4] ), .B1(n30955), .B2(
        \xmem_data[79][4] ), .ZN(n22617) );
  NAND4_X1 U26490 ( .A1(n22620), .A2(n22619), .A3(n22618), .A4(n22617), .ZN(
        n22626) );
  AOI22_X1 U26491 ( .A1(n16973), .A2(\xmem_data[64][4] ), .B1(n28343), .B2(
        \xmem_data[65][4] ), .ZN(n22624) );
  AOI22_X1 U26492 ( .A1(n25422), .A2(\xmem_data[66][4] ), .B1(n29307), .B2(
        \xmem_data[67][4] ), .ZN(n22623) );
  AOI22_X1 U26493 ( .A1(n29308), .A2(\xmem_data[68][4] ), .B1(n24132), .B2(
        \xmem_data[69][4] ), .ZN(n22622) );
  AOI22_X1 U26494 ( .A1(n29310), .A2(\xmem_data[70][4] ), .B1(n29309), .B2(
        \xmem_data[71][4] ), .ZN(n22621) );
  NAND4_X1 U26495 ( .A1(n22624), .A2(n22623), .A3(n22622), .A4(n22621), .ZN(
        n22625) );
  OAI21_X1 U26496 ( .B1(n22628), .B2(n22627), .A(n29267), .ZN(n22636) );
  AOI22_X1 U26497 ( .A1(n29324), .A2(\xmem_data[80][4] ), .B1(n31362), .B2(
        \xmem_data[81][4] ), .ZN(n22633) );
  AOI22_X1 U26498 ( .A1(n29325), .A2(\xmem_data[82][4] ), .B1(n28292), .B2(
        \xmem_data[83][4] ), .ZN(n22632) );
  AOI22_X1 U26499 ( .A1(n29327), .A2(\xmem_data[84][4] ), .B1(n29326), .B2(
        \xmem_data[85][4] ), .ZN(n22631) );
  AND2_X1 U26500 ( .A1(n28038), .A2(\xmem_data[86][4] ), .ZN(n22629) );
  AOI21_X1 U26501 ( .B1(n29328), .B2(\xmem_data[87][4] ), .A(n22629), .ZN(
        n22630) );
  NAND4_X1 U26502 ( .A1(n22633), .A2(n22632), .A3(n22631), .A4(n22630), .ZN(
        n22634) );
  NAND2_X1 U26503 ( .A1(n22634), .A2(n29267), .ZN(n22635) );
  NAND4_X1 U26504 ( .A1(n22638), .A2(n22637), .A3(n22636), .A4(n22635), .ZN(
        n22639) );
  XNOR2_X1 U26505 ( .A(n35238), .B(\fmem_data[11][1] ), .ZN(n32112) );
  INV_X1 U26506 ( .A(n22642), .ZN(n28911) );
  AOI22_X1 U26507 ( .A1(n28468), .A2(\xmem_data[80][0] ), .B1(n31308), .B2(
        \xmem_data[81][0] ), .ZN(n22646) );
  AOI22_X1 U26508 ( .A1(n24686), .A2(\xmem_data[82][0] ), .B1(n28354), .B2(
        \xmem_data[83][0] ), .ZN(n22645) );
  AOI22_X1 U26509 ( .A1(n29118), .A2(\xmem_data[84][0] ), .B1(n3434), .B2(
        \xmem_data[85][0] ), .ZN(n22644) );
  AOI22_X1 U26510 ( .A1(n30589), .A2(\xmem_data[86][0] ), .B1(n25508), .B2(
        \xmem_data[87][0] ), .ZN(n22643) );
  NAND4_X1 U26511 ( .A1(n22646), .A2(n22645), .A3(n22644), .A4(n22643), .ZN(
        n22665) );
  AOI22_X1 U26512 ( .A1(n25677), .A2(\xmem_data[72][0] ), .B1(n22682), .B2(
        \xmem_data[73][0] ), .ZN(n22650) );
  AOI22_X1 U26513 ( .A1(n29318), .A2(\xmem_data[74][0] ), .B1(n22683), .B2(
        \xmem_data[75][0] ), .ZN(n22649) );
  AOI22_X1 U26514 ( .A1(n30495), .A2(\xmem_data[76][0] ), .B1(n30269), .B2(
        \xmem_data[77][0] ), .ZN(n22648) );
  AOI22_X1 U26515 ( .A1(n22685), .A2(\xmem_data[78][0] ), .B1(n22684), .B2(
        \xmem_data[79][0] ), .ZN(n22647) );
  NAND4_X1 U26516 ( .A1(n22650), .A2(n22649), .A3(n22648), .A4(n22647), .ZN(
        n22662) );
  AOI22_X1 U26517 ( .A1(n22674), .A2(\xmem_data[68][0] ), .B1(n24458), .B2(
        \xmem_data[69][0] ), .ZN(n22655) );
  AOI22_X1 U26518 ( .A1(n22675), .A2(\xmem_data[66][0] ), .B1(n25425), .B2(
        \xmem_data[67][0] ), .ZN(n22654) );
  AOI22_X1 U26519 ( .A1(n28415), .A2(\xmem_data[64][0] ), .B1(n30608), .B2(
        \xmem_data[65][0] ), .ZN(n22653) );
  AND2_X1 U26520 ( .A1(n22676), .A2(\xmem_data[71][0] ), .ZN(n22651) );
  AOI21_X1 U26521 ( .B1(n22677), .B2(\xmem_data[70][0] ), .A(n22651), .ZN(
        n22652) );
  NAND4_X1 U26522 ( .A1(n22655), .A2(n22654), .A3(n22653), .A4(n22652), .ZN(
        n22661) );
  AOI22_X1 U26523 ( .A1(n3218), .A2(\xmem_data[88][0] ), .B1(n17033), .B2(
        \xmem_data[89][0] ), .ZN(n22659) );
  AOI22_X1 U26524 ( .A1(n22667), .A2(\xmem_data[90][0] ), .B1(n22666), .B2(
        \xmem_data[91][0] ), .ZN(n22658) );
  AOI22_X1 U26525 ( .A1(n22669), .A2(\xmem_data[92][0] ), .B1(n22668), .B2(
        \xmem_data[93][0] ), .ZN(n22657) );
  AOI22_X1 U26526 ( .A1(n25514), .A2(\xmem_data[94][0] ), .B1(n28374), .B2(
        \xmem_data[95][0] ), .ZN(n22656) );
  NAND4_X1 U26527 ( .A1(n22659), .A2(n22658), .A3(n22657), .A4(n22656), .ZN(
        n22660) );
  OR3_X1 U26528 ( .A1(n22662), .A2(n22661), .A3(n22660), .ZN(n22664) );
  OAI21_X1 U26529 ( .B1(n22665), .B2(n22664), .A(n22663), .ZN(n22773) );
  AOI22_X1 U26530 ( .A1(n3221), .A2(\xmem_data[120][0] ), .B1(n27445), .B2(
        \xmem_data[121][0] ), .ZN(n22673) );
  AOI22_X1 U26531 ( .A1(n22667), .A2(\xmem_data[122][0] ), .B1(n22666), .B2(
        \xmem_data[123][0] ), .ZN(n22672) );
  AOI22_X1 U26532 ( .A1(n22669), .A2(\xmem_data[124][0] ), .B1(n22668), .B2(
        \xmem_data[125][0] ), .ZN(n22671) );
  AOI22_X1 U26533 ( .A1(n23771), .A2(\xmem_data[126][0] ), .B1(n30551), .B2(
        \xmem_data[127][0] ), .ZN(n22670) );
  NAND4_X1 U26534 ( .A1(n22673), .A2(n22672), .A3(n22671), .A4(n22670), .ZN(
        n22692) );
  AOI22_X1 U26535 ( .A1(n3357), .A2(\xmem_data[96][0] ), .B1(n28309), .B2(
        \xmem_data[97][0] ), .ZN(n22681) );
  AOI22_X1 U26536 ( .A1(n22674), .A2(\xmem_data[100][0] ), .B1(n24213), .B2(
        \xmem_data[101][0] ), .ZN(n22680) );
  AOI22_X1 U26537 ( .A1(n22675), .A2(\xmem_data[98][0] ), .B1(n25425), .B2(
        \xmem_data[99][0] ), .ZN(n22679) );
  AOI22_X1 U26538 ( .A1(n22677), .A2(\xmem_data[102][0] ), .B1(n22676), .B2(
        \xmem_data[103][0] ), .ZN(n22678) );
  NAND4_X1 U26539 ( .A1(n22681), .A2(n22680), .A3(n22679), .A4(n22678), .ZN(
        n22691) );
  AOI22_X1 U26540 ( .A1(n24459), .A2(\xmem_data[104][0] ), .B1(n22682), .B2(
        \xmem_data[105][0] ), .ZN(n22689) );
  AOI22_X1 U26541 ( .A1(n29318), .A2(\xmem_data[106][0] ), .B1(n22683), .B2(
        \xmem_data[107][0] ), .ZN(n22688) );
  AOI22_X1 U26542 ( .A1(n25581), .A2(\xmem_data[108][0] ), .B1(n20817), .B2(
        \xmem_data[109][0] ), .ZN(n22687) );
  AOI22_X1 U26543 ( .A1(n22685), .A2(\xmem_data[110][0] ), .B1(n22684), .B2(
        \xmem_data[111][0] ), .ZN(n22686) );
  NAND4_X1 U26544 ( .A1(n22689), .A2(n22688), .A3(n22687), .A4(n22686), .ZN(
        n22690) );
  AOI22_X1 U26545 ( .A1(n30496), .A2(\xmem_data[112][0] ), .B1(n20567), .B2(
        \xmem_data[113][0] ), .ZN(n22697) );
  AOI22_X1 U26546 ( .A1(n27567), .A2(\xmem_data[114][0] ), .B1(n30862), .B2(
        \xmem_data[115][0] ), .ZN(n22696) );
  AOI22_X1 U26547 ( .A1(n20709), .A2(\xmem_data[116][0] ), .B1(n3352), .B2(
        \xmem_data[117][0] ), .ZN(n22695) );
  AND2_X1 U26548 ( .A1(n23731), .A2(\xmem_data[118][0] ), .ZN(n22693) );
  AOI21_X1 U26549 ( .B1(n30592), .B2(\xmem_data[119][0] ), .A(n22693), .ZN(
        n22694) );
  NAND4_X1 U26550 ( .A1(n22697), .A2(n22696), .A3(n22695), .A4(n22694), .ZN(
        n22699) );
  AOI22_X1 U26551 ( .A1(n22701), .A2(\xmem_data[32][0] ), .B1(n30608), .B2(
        \xmem_data[33][0] ), .ZN(n22707) );
  AOI22_X1 U26552 ( .A1(n22702), .A2(\xmem_data[34][0] ), .B1(n20495), .B2(
        \xmem_data[35][0] ), .ZN(n22706) );
  AOI22_X1 U26553 ( .A1(n22703), .A2(\xmem_data[36][0] ), .B1(n20718), .B2(
        \xmem_data[37][0] ), .ZN(n22705) );
  AOI22_X1 U26554 ( .A1(n3208), .A2(\xmem_data[38][0] ), .B1(n24214), .B2(
        \xmem_data[39][0] ), .ZN(n22704) );
  NAND4_X1 U26555 ( .A1(n22707), .A2(n22706), .A3(n22705), .A4(n22704), .ZN(
        n22726) );
  AOI22_X1 U26556 ( .A1(n3218), .A2(\xmem_data[56][0] ), .B1(n22708), .B2(
        \xmem_data[57][0] ), .ZN(n22716) );
  AOI22_X1 U26557 ( .A1(n22710), .A2(\xmem_data[58][0] ), .B1(n22709), .B2(
        \xmem_data[59][0] ), .ZN(n22715) );
  AOI22_X1 U26558 ( .A1(n22711), .A2(\xmem_data[60][0] ), .B1(n25417), .B2(
        \xmem_data[61][0] ), .ZN(n22714) );
  AOI22_X1 U26559 ( .A1(n28343), .A2(\xmem_data[62][0] ), .B1(n22712), .B2(
        \xmem_data[63][0] ), .ZN(n22713) );
  NAND4_X1 U26560 ( .A1(n22716), .A2(n22715), .A3(n22714), .A4(n22713), .ZN(
        n22725) );
  AOI22_X1 U26561 ( .A1(n24222), .A2(\xmem_data[44][0] ), .B1(n3328), .B2(
        \xmem_data[45][0] ), .ZN(n22723) );
  AOI22_X1 U26562 ( .A1(n22718), .A2(\xmem_data[40][0] ), .B1(n22717), .B2(
        \xmem_data[41][0] ), .ZN(n22722) );
  AOI22_X1 U26563 ( .A1(n24570), .A2(\xmem_data[46][0] ), .B1(n22719), .B2(
        \xmem_data[47][0] ), .ZN(n22721) );
  AOI22_X1 U26564 ( .A1(n20731), .A2(\xmem_data[43][0] ), .B1(
        \xmem_data[42][0] ), .B2(n13481), .ZN(n22720) );
  NAND4_X1 U26565 ( .A1(n22723), .A2(n22722), .A3(n22721), .A4(n22720), .ZN(
        n22724) );
  AOI22_X1 U26566 ( .A1(n27526), .A2(\xmem_data[48][0] ), .B1(n30674), .B2(
        \xmem_data[49][0] ), .ZN(n22734) );
  AOI22_X1 U26567 ( .A1(n22727), .A2(\xmem_data[50][0] ), .B1(n27436), .B2(
        \xmem_data[51][0] ), .ZN(n22733) );
  AOI22_X1 U26568 ( .A1(n22729), .A2(\xmem_data[52][0] ), .B1(n22728), .B2(
        \xmem_data[53][0] ), .ZN(n22732) );
  AND2_X1 U26569 ( .A1(n3247), .A2(\xmem_data[54][0] ), .ZN(n22730) );
  AOI21_X1 U26570 ( .B1(n27502), .B2(\xmem_data[55][0] ), .A(n22730), .ZN(
        n22731) );
  NAND4_X1 U26571 ( .A1(n22734), .A2(n22733), .A3(n22732), .A4(n22731), .ZN(
        n22736) );
  AOI22_X1 U26572 ( .A1(n22739), .A2(\xmem_data[0][0] ), .B1(n22738), .B2(
        \xmem_data[1][0] ), .ZN(n22746) );
  AOI22_X1 U26573 ( .A1(n22740), .A2(\xmem_data[2][0] ), .B1(n27537), .B2(
        \xmem_data[3][0] ), .ZN(n22745) );
  AOI22_X1 U26574 ( .A1(n22741), .A2(\xmem_data[4][0] ), .B1(n30746), .B2(
        \xmem_data[5][0] ), .ZN(n22744) );
  AOI22_X1 U26575 ( .A1(n22742), .A2(\xmem_data[6][0] ), .B1(n25573), .B2(
        \xmem_data[7][0] ), .ZN(n22743) );
  NAND4_X1 U26576 ( .A1(n22746), .A2(n22745), .A3(n22744), .A4(n22743), .ZN(
        n22767) );
  AOI22_X1 U26577 ( .A1(n27918), .A2(\xmem_data[8][0] ), .B1(n23802), .B2(
        \xmem_data[9][0] ), .ZN(n22750) );
  AOI22_X1 U26578 ( .A1(n29238), .A2(\xmem_data[10][0] ), .B1(n28428), .B2(
        \xmem_data[11][0] ), .ZN(n22749) );
  AOI22_X1 U26579 ( .A1(n20506), .A2(\xmem_data[12][0] ), .B1(n20984), .B2(
        \xmem_data[13][0] ), .ZN(n22748) );
  AOI22_X1 U26580 ( .A1(n28098), .A2(\xmem_data[14][0] ), .B1(n20782), .B2(
        \xmem_data[15][0] ), .ZN(n22747) );
  NAND4_X1 U26581 ( .A1(n22750), .A2(n22749), .A3(n22748), .A4(n22747), .ZN(
        n22766) );
  AOI22_X1 U26582 ( .A1(n22751), .A2(\xmem_data[16][0] ), .B1(n14982), .B2(
        \xmem_data[17][0] ), .ZN(n22757) );
  AOI22_X1 U26583 ( .A1(n30900), .A2(\xmem_data[18][0] ), .B1(n20986), .B2(
        \xmem_data[19][0] ), .ZN(n22756) );
  AOI22_X1 U26584 ( .A1(n22752), .A2(\xmem_data[20][0] ), .B1(n3335), .B2(
        \xmem_data[21][0] ), .ZN(n22755) );
  AOI22_X1 U26585 ( .A1(n22753), .A2(\xmem_data[22][0] ), .B1(n29064), .B2(
        \xmem_data[23][0] ), .ZN(n22754) );
  NAND4_X1 U26586 ( .A1(n22757), .A2(n22756), .A3(n22755), .A4(n22754), .ZN(
        n22765) );
  AOI22_X1 U26587 ( .A1(n3222), .A2(\xmem_data[24][0] ), .B1(n25693), .B2(
        \xmem_data[25][0] ), .ZN(n22763) );
  AOI22_X1 U26588 ( .A1(n30534), .A2(\xmem_data[26][0] ), .B1(n22758), .B2(
        \xmem_data[27][0] ), .ZN(n22762) );
  AOI22_X1 U26589 ( .A1(n22759), .A2(\xmem_data[28][0] ), .B1(n28952), .B2(
        \xmem_data[29][0] ), .ZN(n22761) );
  AOI22_X1 U26590 ( .A1(n13474), .A2(\xmem_data[30][0] ), .B1(n25422), .B2(
        \xmem_data[31][0] ), .ZN(n22760) );
  NAND4_X1 U26591 ( .A1(n22763), .A2(n22762), .A3(n22761), .A4(n22760), .ZN(
        n22764) );
  OR4_X1 U26592 ( .A1(n22767), .A2(n22766), .A3(n22765), .A4(n22764), .ZN(
        n22769) );
  XNOR2_X1 U26593 ( .A(n34623), .B(\fmem_data[5][7] ), .ZN(n22774) );
  XNOR2_X1 U26594 ( .A(n3354), .B(\fmem_data[2][7] ), .ZN(n22776) );
  XNOR2_X1 U26595 ( .A(n32419), .B(\fmem_data[5][5] ), .ZN(n31884) );
  XNOR2_X1 U26596 ( .A(n22779), .B(n24841), .ZN(n27317) );
  FA_X1 U26597 ( .A(n22782), .B(n22781), .CI(n22780), .CO(n23580), .S(n33888)
         );
  AOI22_X1 U26598 ( .A1(n23740), .A2(\xmem_data[120][1] ), .B1(n23739), .B2(
        \xmem_data[121][1] ), .ZN(n22786) );
  AOI22_X1 U26599 ( .A1(n23741), .A2(\xmem_data[122][1] ), .B1(n17061), .B2(
        \xmem_data[123][1] ), .ZN(n22785) );
  AOI22_X1 U26600 ( .A1(n23742), .A2(\xmem_data[124][1] ), .B1(n29103), .B2(
        \xmem_data[125][1] ), .ZN(n22784) );
  AOI22_X1 U26601 ( .A1(n27447), .A2(\xmem_data[126][1] ), .B1(n20546), .B2(
        \xmem_data[127][1] ), .ZN(n22783) );
  NAND4_X1 U26602 ( .A1(n22786), .A2(n22785), .A3(n22784), .A4(n22783), .ZN(
        n22803) );
  AOI22_X1 U26603 ( .A1(n23730), .A2(\xmem_data[112][1] ), .B1(n20707), .B2(
        \xmem_data[113][1] ), .ZN(n22790) );
  AOI22_X1 U26604 ( .A1(n29124), .A2(\xmem_data[114][1] ), .B1(n31309), .B2(
        \xmem_data[115][1] ), .ZN(n22789) );
  AOI22_X1 U26605 ( .A1(n23732), .A2(\xmem_data[116][1] ), .B1(n23731), .B2(
        \xmem_data[117][1] ), .ZN(n22788) );
  AOI22_X1 U26606 ( .A1(n23734), .A2(\xmem_data[118][1] ), .B1(n3221), .B2(
        \xmem_data[119][1] ), .ZN(n22787) );
  NAND4_X1 U26607 ( .A1(n22790), .A2(n22789), .A3(n22788), .A4(n22787), .ZN(
        n22801) );
  AOI22_X1 U26608 ( .A1(n23722), .A2(\xmem_data[104][1] ), .B1(n29049), .B2(
        \xmem_data[105][1] ), .ZN(n22794) );
  AOI22_X1 U26609 ( .A1(n24615), .A2(\xmem_data[106][1] ), .B1(n25364), .B2(
        \xmem_data[107][1] ), .ZN(n22793) );
  AOI22_X1 U26610 ( .A1(n23724), .A2(\xmem_data[108][1] ), .B1(n23723), .B2(
        \xmem_data[109][1] ), .ZN(n22792) );
  AOI22_X1 U26611 ( .A1(n25582), .A2(\xmem_data[110][1] ), .B1(n23725), .B2(
        \xmem_data[111][1] ), .ZN(n22791) );
  NAND4_X1 U26612 ( .A1(n22794), .A2(n22793), .A3(n22792), .A4(n22791), .ZN(
        n22800) );
  AOI22_X1 U26613 ( .A1(n17013), .A2(\xmem_data[96][1] ), .B1(n22675), .B2(
        \xmem_data[97][1] ), .ZN(n22798) );
  AOI22_X1 U26614 ( .A1(n25710), .A2(\xmem_data[98][1] ), .B1(n23715), .B2(
        \xmem_data[99][1] ), .ZN(n22797) );
  AOI22_X1 U26615 ( .A1(n16988), .A2(\xmem_data[100][1] ), .B1(n23716), .B2(
        \xmem_data[101][1] ), .ZN(n22796) );
  AOI22_X1 U26616 ( .A1(n23717), .A2(\xmem_data[102][1] ), .B1(n21006), .B2(
        \xmem_data[103][1] ), .ZN(n22795) );
  NAND4_X1 U26617 ( .A1(n22798), .A2(n22797), .A3(n22796), .A4(n22795), .ZN(
        n22799) );
  OR3_X1 U26618 ( .A1(n22801), .A2(n22800), .A3(n22799), .ZN(n22802) );
  OAI21_X1 U26619 ( .B1(n22803), .B2(n22802), .A(n23751), .ZN(n22886) );
  AOI22_X1 U26620 ( .A1(n23740), .A2(\xmem_data[88][1] ), .B1(n23739), .B2(
        \xmem_data[89][1] ), .ZN(n22807) );
  AOI22_X1 U26621 ( .A1(n23741), .A2(\xmem_data[90][1] ), .B1(n20806), .B2(
        \xmem_data[91][1] ), .ZN(n22806) );
  AOI22_X1 U26622 ( .A1(n23742), .A2(\xmem_data[92][1] ), .B1(n27446), .B2(
        \xmem_data[93][1] ), .ZN(n22805) );
  AOI22_X1 U26623 ( .A1(n27447), .A2(\xmem_data[94][1] ), .B1(n30884), .B2(
        \xmem_data[95][1] ), .ZN(n22804) );
  NAND4_X1 U26624 ( .A1(n22807), .A2(n22806), .A3(n22805), .A4(n22804), .ZN(
        n22824) );
  AOI22_X1 U26625 ( .A1(n23730), .A2(\xmem_data[80][1] ), .B1(n20951), .B2(
        \xmem_data[81][1] ), .ZN(n22811) );
  AOI22_X1 U26626 ( .A1(n20953), .A2(\xmem_data[82][1] ), .B1(n28075), .B2(
        \xmem_data[83][1] ), .ZN(n22810) );
  AOI22_X1 U26627 ( .A1(n23732), .A2(\xmem_data[84][1] ), .B1(n23731), .B2(
        \xmem_data[85][1] ), .ZN(n22809) );
  AOI22_X1 U26628 ( .A1(n23734), .A2(\xmem_data[86][1] ), .B1(n3221), .B2(
        \xmem_data[87][1] ), .ZN(n22808) );
  NAND4_X1 U26629 ( .A1(n22811), .A2(n22810), .A3(n22809), .A4(n22808), .ZN(
        n22822) );
  AOI22_X1 U26630 ( .A1(n23722), .A2(\xmem_data[72][1] ), .B1(n30871), .B2(
        \xmem_data[73][1] ), .ZN(n22815) );
  AOI22_X1 U26631 ( .A1(n3178), .A2(\xmem_data[74][1] ), .B1(n20816), .B2(
        \xmem_data[75][1] ), .ZN(n22814) );
  AOI22_X1 U26632 ( .A1(n23724), .A2(\xmem_data[76][1] ), .B1(n23723), .B2(
        \xmem_data[77][1] ), .ZN(n22813) );
  AOI22_X1 U26633 ( .A1(n24685), .A2(\xmem_data[78][1] ), .B1(n23725), .B2(
        \xmem_data[79][1] ), .ZN(n22812) );
  NAND4_X1 U26634 ( .A1(n22815), .A2(n22814), .A3(n22813), .A4(n22812), .ZN(
        n22821) );
  AOI22_X1 U26635 ( .A1(n30608), .A2(\xmem_data[64][1] ), .B1(n30552), .B2(
        \xmem_data[65][1] ), .ZN(n22819) );
  AOI22_X1 U26636 ( .A1(n30614), .A2(\xmem_data[66][1] ), .B1(n23715), .B2(
        \xmem_data[67][1] ), .ZN(n22818) );
  AOI22_X1 U26637 ( .A1(n30666), .A2(\xmem_data[68][1] ), .B1(n23716), .B2(
        \xmem_data[69][1] ), .ZN(n22817) );
  AOI22_X1 U26638 ( .A1(n23717), .A2(\xmem_data[70][1] ), .B1(n29048), .B2(
        \xmem_data[71][1] ), .ZN(n22816) );
  NAND4_X1 U26639 ( .A1(n22819), .A2(n22818), .A3(n22817), .A4(n22816), .ZN(
        n22820) );
  OR3_X1 U26640 ( .A1(n22822), .A2(n22821), .A3(n22820), .ZN(n22823) );
  OAI21_X1 U26641 ( .B1(n22824), .B2(n22823), .A(n23713), .ZN(n22885) );
  NAND2_X1 U26642 ( .A1(n25450), .A2(\xmem_data[61][1] ), .ZN(n22850) );
  AOI22_X1 U26643 ( .A1(n23753), .A2(\xmem_data[48][1] ), .B1(n30524), .B2(
        \xmem_data[49][1] ), .ZN(n22828) );
  AOI22_X1 U26644 ( .A1(n17056), .A2(\xmem_data[50][1] ), .B1(n20709), .B2(
        \xmem_data[51][1] ), .ZN(n22827) );
  AOI22_X1 U26645 ( .A1(n23754), .A2(\xmem_data[52][1] ), .B1(n29286), .B2(
        \xmem_data[53][1] ), .ZN(n22826) );
  AOI22_X1 U26646 ( .A1(n23756), .A2(\xmem_data[54][1] ), .B1(n3221), .B2(
        \xmem_data[55][1] ), .ZN(n22825) );
  NAND4_X1 U26647 ( .A1(n22828), .A2(n22827), .A3(n22826), .A4(n22825), .ZN(
        n22847) );
  AOI22_X1 U26648 ( .A1(n23762), .A2(\xmem_data[32][1] ), .B1(n23761), .B2(
        \xmem_data[33][1] ), .ZN(n22832) );
  AOI22_X1 U26649 ( .A1(n23763), .A2(\xmem_data[34][1] ), .B1(n20798), .B2(
        \xmem_data[35][1] ), .ZN(n22831) );
  AOI22_X1 U26650 ( .A1(n30746), .A2(\xmem_data[36][1] ), .B1(n3212), .B2(
        \xmem_data[37][1] ), .ZN(n22830) );
  AOI22_X1 U26651 ( .A1(n23764), .A2(\xmem_data[38][1] ), .B1(n27918), .B2(
        \xmem_data[39][1] ), .ZN(n22829) );
  NAND4_X1 U26652 ( .A1(n22832), .A2(n22831), .A3(n22830), .A4(n22829), .ZN(
        n22846) );
  AOI22_X1 U26653 ( .A1(n23777), .A2(\xmem_data[40][1] ), .B1(n23776), .B2(
        \xmem_data[41][1] ), .ZN(n22836) );
  AOI22_X1 U26654 ( .A1(n25575), .A2(\xmem_data[42][1] ), .B1(n23778), .B2(
        \xmem_data[43][1] ), .ZN(n22835) );
  AOI22_X1 U26655 ( .A1(n23780), .A2(\xmem_data[44][1] ), .B1(n23779), .B2(
        \xmem_data[45][1] ), .ZN(n22834) );
  AOI22_X1 U26656 ( .A1(n21058), .A2(\xmem_data[46][1] ), .B1(n23781), .B2(
        \xmem_data[47][1] ), .ZN(n22833) );
  NAND4_X1 U26657 ( .A1(n22836), .A2(n22835), .A3(n22834), .A4(n22833), .ZN(
        n22845) );
  AOI22_X1 U26658 ( .A1(n23770), .A2(\xmem_data[56][1] ), .B1(n23769), .B2(
        \xmem_data[57][1] ), .ZN(n22837) );
  INV_X1 U26659 ( .A(n22837), .ZN(n22841) );
  AOI22_X1 U26660 ( .A1(n27447), .A2(\xmem_data[62][1] ), .B1(n24130), .B2(
        \xmem_data[63][1] ), .ZN(n22838) );
  INV_X1 U26661 ( .A(n22838), .ZN(n22840) );
  AND2_X1 U26662 ( .A1(n3140), .A2(\xmem_data[60][1] ), .ZN(n22839) );
  NOR3_X1 U26663 ( .A1(n22841), .A2(n22840), .A3(n22839), .ZN(n22843) );
  AOI22_X1 U26664 ( .A1(n27938), .A2(\xmem_data[58][1] ), .B1(n24633), .B2(
        \xmem_data[59][1] ), .ZN(n22842) );
  NAND2_X1 U26665 ( .A1(n22843), .A2(n22842), .ZN(n22844) );
  NOR4_X1 U26666 ( .A1(n22847), .A2(n22846), .A3(n22845), .A4(n22844), .ZN(
        n22849) );
  INV_X1 U26667 ( .A(n23790), .ZN(n22848) );
  AOI21_X1 U26668 ( .B1(n22850), .B2(n22849), .A(n22848), .ZN(n22851) );
  INV_X1 U26669 ( .A(n22851), .ZN(n22884) );
  AOI22_X1 U26670 ( .A1(n23812), .A2(\xmem_data[26][1] ), .B1(n23811), .B2(
        \xmem_data[27][1] ), .ZN(n22853) );
  AND2_X1 U26671 ( .A1(n22853), .A2(n22852), .ZN(n22858) );
  AOI22_X1 U26672 ( .A1(n29026), .A2(\xmem_data[24][1] ), .B1(n25491), .B2(
        \xmem_data[25][1] ), .ZN(n22854) );
  AOI22_X1 U26673 ( .A1(n29820), .A2(\xmem_data[16][1] ), .B1(n30601), .B2(
        \xmem_data[17][1] ), .ZN(n22862) );
  AOI22_X1 U26674 ( .A1(n28076), .A2(\xmem_data[18][1] ), .B1(n28317), .B2(
        \xmem_data[19][1] ), .ZN(n22861) );
  AOI22_X1 U26675 ( .A1(n23754), .A2(\xmem_data[20][1] ), .B1(n29253), .B2(
        \xmem_data[21][1] ), .ZN(n22860) );
  AOI22_X1 U26676 ( .A1(n27902), .A2(\xmem_data[22][1] ), .B1(n3220), .B2(
        \xmem_data[23][1] ), .ZN(n22859) );
  NAND4_X1 U26677 ( .A1(n22862), .A2(n22861), .A3(n22860), .A4(n22859), .ZN(
        n22863) );
  AOI22_X1 U26678 ( .A1(n23802), .A2(\xmem_data[8][1] ), .B1(n23801), .B2(
        \xmem_data[9][1] ), .ZN(n22868) );
  AOI22_X1 U26679 ( .A1(n28493), .A2(\xmem_data[10][1] ), .B1(n28494), .B2(
        \xmem_data[11][1] ), .ZN(n22867) );
  AOI22_X1 U26680 ( .A1(n25718), .A2(\xmem_data[12][1] ), .B1(n28983), .B2(
        \xmem_data[13][1] ), .ZN(n22866) );
  AOI22_X1 U26681 ( .A1(n20734), .A2(\xmem_data[14][1] ), .B1(n27981), .B2(
        \xmem_data[15][1] ), .ZN(n22865) );
  NAND4_X1 U26682 ( .A1(n22868), .A2(n22867), .A3(n22866), .A4(n22865), .ZN(
        n22874) );
  AOI22_X1 U26683 ( .A1(n23792), .A2(\xmem_data[0][1] ), .B1(n20775), .B2(
        \xmem_data[1][1] ), .ZN(n22872) );
  AOI22_X1 U26684 ( .A1(n28298), .A2(\xmem_data[2][1] ), .B1(n23793), .B2(
        \xmem_data[3][1] ), .ZN(n22871) );
  AOI22_X1 U26685 ( .A1(n30303), .A2(\xmem_data[4][1] ), .B1(n3208), .B2(
        \xmem_data[5][1] ), .ZN(n22870) );
  AOI22_X1 U26686 ( .A1(n30949), .A2(\xmem_data[6][1] ), .B1(n23796), .B2(
        \xmem_data[7][1] ), .ZN(n22869) );
  NAND4_X1 U26687 ( .A1(n22872), .A2(n22871), .A3(n22870), .A4(n22869), .ZN(
        n22873) );
  NOR2_X1 U26688 ( .A1(n22874), .A2(n22873), .ZN(n22875) );
  NAND2_X1 U26689 ( .A1(n22876), .A2(n22875), .ZN(n22882) );
  INV_X1 U26690 ( .A(n23822), .ZN(n22877) );
  NOR2_X1 U26691 ( .A1(n22877), .A2(n39028), .ZN(n22878) );
  AND2_X1 U26692 ( .A1(n3126), .A2(\xmem_data[28][1] ), .ZN(n22879) );
  XNOR2_X1 U26693 ( .A(n32979), .B(\fmem_data[4][5] ), .ZN(n31445) );
  AOI22_X1 U26694 ( .A1(n23762), .A2(\xmem_data[32][2] ), .B1(n23761), .B2(
        \xmem_data[33][2] ), .ZN(n22890) );
  AOI22_X1 U26695 ( .A1(n23763), .A2(\xmem_data[34][2] ), .B1(n28090), .B2(
        \xmem_data[35][2] ), .ZN(n22889) );
  AOI22_X1 U26696 ( .A1(n28516), .A2(\xmem_data[36][2] ), .B1(n3213), .B2(
        \xmem_data[37][2] ), .ZN(n22888) );
  AOI22_X1 U26697 ( .A1(n23764), .A2(\xmem_data[38][2] ), .B1(n24707), .B2(
        \xmem_data[39][2] ), .ZN(n22887) );
  NAND4_X1 U26698 ( .A1(n22890), .A2(n22889), .A3(n22888), .A4(n22887), .ZN(
        n22906) );
  AOI22_X1 U26699 ( .A1(n23777), .A2(\xmem_data[40][2] ), .B1(n23776), .B2(
        \xmem_data[41][2] ), .ZN(n22894) );
  AOI22_X1 U26700 ( .A1(n28385), .A2(\xmem_data[42][2] ), .B1(n23778), .B2(
        \xmem_data[43][2] ), .ZN(n22893) );
  AOI22_X1 U26701 ( .A1(n23780), .A2(\xmem_data[44][2] ), .B1(n23779), .B2(
        \xmem_data[45][2] ), .ZN(n22892) );
  AOI22_X1 U26702 ( .A1(n25582), .A2(\xmem_data[46][2] ), .B1(n23781), .B2(
        \xmem_data[47][2] ), .ZN(n22891) );
  NAND4_X1 U26703 ( .A1(n22894), .A2(n22893), .A3(n22892), .A4(n22891), .ZN(
        n22905) );
  AOI22_X1 U26704 ( .A1(n23753), .A2(\xmem_data[48][2] ), .B1(n28329), .B2(
        \xmem_data[49][2] ), .ZN(n22898) );
  AOI22_X1 U26705 ( .A1(n29057), .A2(\xmem_data[50][2] ), .B1(n20578), .B2(
        \xmem_data[51][2] ), .ZN(n22897) );
  AOI22_X1 U26706 ( .A1(n23754), .A2(\xmem_data[52][2] ), .B1(n25485), .B2(
        \xmem_data[53][2] ), .ZN(n22896) );
  AOI22_X1 U26707 ( .A1(n23756), .A2(\xmem_data[54][2] ), .B1(n3221), .B2(
        \xmem_data[55][2] ), .ZN(n22895) );
  NAND4_X1 U26708 ( .A1(n22898), .A2(n22897), .A3(n22896), .A4(n22895), .ZN(
        n22904) );
  AOI22_X1 U26709 ( .A1(n23770), .A2(\xmem_data[56][2] ), .B1(n23769), .B2(
        \xmem_data[57][2] ), .ZN(n22902) );
  AOI22_X1 U26710 ( .A1(n25617), .A2(\xmem_data[58][2] ), .B1(n30882), .B2(
        \xmem_data[59][2] ), .ZN(n22901) );
  AOI22_X1 U26711 ( .A1(n25732), .A2(\xmem_data[60][2] ), .B1(n25450), .B2(
        \xmem_data[61][2] ), .ZN(n22900) );
  AOI22_X1 U26712 ( .A1(n27447), .A2(\xmem_data[62][2] ), .B1(n30884), .B2(
        \xmem_data[63][2] ), .ZN(n22899) );
  NAND4_X1 U26713 ( .A1(n22902), .A2(n22901), .A3(n22900), .A4(n22899), .ZN(
        n22903) );
  OR4_X1 U26714 ( .A1(n22906), .A2(n22905), .A3(n22904), .A4(n22903), .ZN(
        n22933) );
  NAND2_X1 U26715 ( .A1(n25450), .A2(\xmem_data[29][2] ), .ZN(n22931) );
  AOI22_X1 U26716 ( .A1(n29657), .A2(\xmem_data[16][2] ), .B1(n20769), .B2(
        \xmem_data[17][2] ), .ZN(n22910) );
  AOI22_X1 U26717 ( .A1(n28038), .A2(\xmem_data[18][2] ), .B1(n28317), .B2(
        \xmem_data[19][2] ), .ZN(n22909) );
  AOI22_X1 U26718 ( .A1(n3317), .A2(\xmem_data[20][2] ), .B1(n3247), .B2(
        \xmem_data[21][2] ), .ZN(n22908) );
  AOI22_X1 U26719 ( .A1(n28355), .A2(\xmem_data[22][2] ), .B1(n3217), .B2(
        \xmem_data[23][2] ), .ZN(n22907) );
  NAND4_X1 U26720 ( .A1(n22910), .A2(n22909), .A3(n22908), .A4(n22907), .ZN(
        n22929) );
  AOI22_X1 U26721 ( .A1(n23792), .A2(\xmem_data[0][2] ), .B1(n27452), .B2(
        \xmem_data[1][2] ), .ZN(n22914) );
  AOI22_X1 U26722 ( .A1(n20541), .A2(\xmem_data[2][2] ), .B1(n23793), .B2(
        \xmem_data[3][2] ), .ZN(n22913) );
  AOI22_X1 U26723 ( .A1(n30948), .A2(\xmem_data[4][2] ), .B1(n3208), .B2(
        \xmem_data[5][2] ), .ZN(n22912) );
  AOI22_X1 U26724 ( .A1(n25434), .A2(\xmem_data[6][2] ), .B1(n23796), .B2(
        \xmem_data[7][2] ), .ZN(n22911) );
  NAND4_X1 U26725 ( .A1(n22914), .A2(n22913), .A3(n22912), .A4(n22911), .ZN(
        n22928) );
  AOI22_X1 U26726 ( .A1(n23802), .A2(\xmem_data[8][2] ), .B1(n23801), .B2(
        \xmem_data[9][2] ), .ZN(n22918) );
  AOI22_X1 U26727 ( .A1(n30557), .A2(\xmem_data[10][2] ), .B1(n28291), .B2(
        \xmem_data[11][2] ), .ZN(n22917) );
  AOI22_X1 U26728 ( .A1(n20950), .A2(\xmem_data[12][2] ), .B1(n20553), .B2(
        \xmem_data[13][2] ), .ZN(n22916) );
  AOI22_X1 U26729 ( .A1(n27847), .A2(\xmem_data[14][2] ), .B1(n30496), .B2(
        \xmem_data[15][2] ), .ZN(n22915) );
  NAND4_X1 U26730 ( .A1(n22918), .A2(n22917), .A3(n22916), .A4(n22915), .ZN(
        n22927) );
  AOI22_X1 U26731 ( .A1(n23812), .A2(\xmem_data[26][2] ), .B1(n23811), .B2(
        \xmem_data[27][2] ), .ZN(n22925) );
  AOI22_X1 U26732 ( .A1(n28367), .A2(\xmem_data[24][2] ), .B1(n20500), .B2(
        \xmem_data[25][2] ), .ZN(n22919) );
  INV_X1 U26733 ( .A(n22919), .ZN(n22923) );
  AND2_X1 U26734 ( .A1(n3134), .A2(\xmem_data[28][2] ), .ZN(n22922) );
  AOI22_X1 U26735 ( .A1(n23813), .A2(\xmem_data[30][2] ), .B1(n13475), .B2(
        \xmem_data[31][2] ), .ZN(n22920) );
  INV_X1 U26736 ( .A(n22920), .ZN(n22921) );
  NOR3_X1 U26737 ( .A1(n22923), .A2(n22922), .A3(n22921), .ZN(n22924) );
  NAND2_X1 U26738 ( .A1(n22925), .A2(n22924), .ZN(n22926) );
  NOR4_X1 U26739 ( .A1(n22929), .A2(n22928), .A3(n22927), .A4(n22926), .ZN(
        n22930) );
  AOI21_X1 U26740 ( .B1(n22931), .B2(n22930), .A(n22877), .ZN(n22932) );
  AOI21_X1 U26741 ( .B1(n22933), .B2(n23790), .A(n22932), .ZN(n22977) );
  AOI22_X1 U26742 ( .A1(n28671), .A2(\xmem_data[96][2] ), .B1(n21015), .B2(
        \xmem_data[97][2] ), .ZN(n22937) );
  AOI22_X1 U26743 ( .A1(n3175), .A2(\xmem_data[98][2] ), .B1(n23715), .B2(
        \xmem_data[99][2] ), .ZN(n22936) );
  AOI22_X1 U26744 ( .A1(n28516), .A2(\xmem_data[100][2] ), .B1(n23716), .B2(
        \xmem_data[101][2] ), .ZN(n22935) );
  AOI22_X1 U26745 ( .A1(n23717), .A2(\xmem_data[102][2] ), .B1(n24707), .B2(
        \xmem_data[103][2] ), .ZN(n22934) );
  NAND4_X1 U26746 ( .A1(n22937), .A2(n22936), .A3(n22935), .A4(n22934), .ZN(
        n22953) );
  AOI22_X1 U26747 ( .A1(n23722), .A2(\xmem_data[104][2] ), .B1(n29318), .B2(
        \xmem_data[105][2] ), .ZN(n22941) );
  AOI22_X1 U26748 ( .A1(n24220), .A2(\xmem_data[106][2] ), .B1(n25581), .B2(
        \xmem_data[107][2] ), .ZN(n22940) );
  AOI22_X1 U26749 ( .A1(n23724), .A2(\xmem_data[108][2] ), .B1(n23723), .B2(
        \xmem_data[109][2] ), .ZN(n22939) );
  AOI22_X1 U26750 ( .A1(n27847), .A2(\xmem_data[110][2] ), .B1(n23725), .B2(
        \xmem_data[111][2] ), .ZN(n22938) );
  NAND4_X1 U26751 ( .A1(n22941), .A2(n22940), .A3(n22939), .A4(n22938), .ZN(
        n22952) );
  AOI22_X1 U26752 ( .A1(n23730), .A2(\xmem_data[112][2] ), .B1(n20579), .B2(
        \xmem_data[113][2] ), .ZN(n22945) );
  AOI22_X1 U26753 ( .A1(n20986), .A2(\xmem_data[114][2] ), .B1(n27563), .B2(
        \xmem_data[115][2] ), .ZN(n22944) );
  AOI22_X1 U26754 ( .A1(n23732), .A2(\xmem_data[116][2] ), .B1(n23731), .B2(
        \xmem_data[117][2] ), .ZN(n22943) );
  AOI22_X1 U26755 ( .A1(n23734), .A2(\xmem_data[118][2] ), .B1(n3217), .B2(
        \xmem_data[119][2] ), .ZN(n22942) );
  NAND4_X1 U26756 ( .A1(n22945), .A2(n22944), .A3(n22943), .A4(n22942), .ZN(
        n22951) );
  AOI22_X1 U26757 ( .A1(n23740), .A2(\xmem_data[120][2] ), .B1(n23739), .B2(
        \xmem_data[121][2] ), .ZN(n22949) );
  AOI22_X1 U26758 ( .A1(n23741), .A2(\xmem_data[122][2] ), .B1(n27994), .B2(
        \xmem_data[123][2] ), .ZN(n22948) );
  AOI22_X1 U26759 ( .A1(n23742), .A2(\xmem_data[124][2] ), .B1(n28510), .B2(
        \xmem_data[125][2] ), .ZN(n22947) );
  AOI22_X1 U26760 ( .A1(n27447), .A2(\xmem_data[126][2] ), .B1(n27863), .B2(
        \xmem_data[127][2] ), .ZN(n22946) );
  NAND4_X1 U26761 ( .A1(n22949), .A2(n22948), .A3(n22947), .A4(n22946), .ZN(
        n22950) );
  OR4_X1 U26762 ( .A1(n22953), .A2(n22952), .A3(n22951), .A4(n22950), .ZN(
        n22975) );
  AOI22_X1 U26763 ( .A1(n31353), .A2(\xmem_data[64][2] ), .B1(n29232), .B2(
        \xmem_data[65][2] ), .ZN(n22957) );
  AOI22_X1 U26764 ( .A1(n3176), .A2(\xmem_data[66][2] ), .B1(n23715), .B2(
        \xmem_data[67][2] ), .ZN(n22956) );
  AOI22_X1 U26765 ( .A1(n29008), .A2(\xmem_data[68][2] ), .B1(n23716), .B2(
        \xmem_data[69][2] ), .ZN(n22955) );
  AOI22_X1 U26766 ( .A1(n23717), .A2(\xmem_data[70][2] ), .B1(n29048), .B2(
        \xmem_data[71][2] ), .ZN(n22954) );
  NAND4_X1 U26767 ( .A1(n22957), .A2(n22956), .A3(n22955), .A4(n22954), .ZN(
        n22973) );
  AOI22_X1 U26768 ( .A1(n23722), .A2(\xmem_data[72][2] ), .B1(n31360), .B2(
        \xmem_data[73][2] ), .ZN(n22961) );
  AOI22_X1 U26769 ( .A1(n27974), .A2(\xmem_data[74][2] ), .B1(n30898), .B2(
        \xmem_data[75][2] ), .ZN(n22960) );
  AOI22_X1 U26770 ( .A1(n23724), .A2(\xmem_data[76][2] ), .B1(n23723), .B2(
        \xmem_data[77][2] ), .ZN(n22959) );
  AOI22_X1 U26771 ( .A1(n20782), .A2(\xmem_data[78][2] ), .B1(n23725), .B2(
        \xmem_data[79][2] ), .ZN(n22958) );
  NAND4_X1 U26772 ( .A1(n22961), .A2(n22960), .A3(n22959), .A4(n22958), .ZN(
        n22972) );
  AOI22_X1 U26773 ( .A1(n23730), .A2(\xmem_data[80][2] ), .B1(n20769), .B2(
        \xmem_data[81][2] ), .ZN(n22965) );
  AOI22_X1 U26774 ( .A1(n25686), .A2(\xmem_data[82][2] ), .B1(n12471), .B2(
        \xmem_data[83][2] ), .ZN(n22964) );
  AOI22_X1 U26775 ( .A1(n23732), .A2(\xmem_data[84][2] ), .B1(n23731), .B2(
        \xmem_data[85][2] ), .ZN(n22963) );
  AOI22_X1 U26776 ( .A1(n23734), .A2(\xmem_data[86][2] ), .B1(n3218), .B2(
        \xmem_data[87][2] ), .ZN(n22962) );
  NAND4_X1 U26777 ( .A1(n22965), .A2(n22964), .A3(n22963), .A4(n22962), .ZN(
        n22971) );
  AOI22_X1 U26778 ( .A1(n23740), .A2(\xmem_data[88][2] ), .B1(n23739), .B2(
        \xmem_data[89][2] ), .ZN(n22969) );
  AOI22_X1 U26779 ( .A1(n23741), .A2(\xmem_data[90][2] ), .B1(n29181), .B2(
        \xmem_data[91][2] ), .ZN(n22968) );
  AOI22_X1 U26780 ( .A1(n23742), .A2(\xmem_data[92][2] ), .B1(n28045), .B2(
        \xmem_data[93][2] ), .ZN(n22967) );
  AOI22_X1 U26781 ( .A1(n27447), .A2(\xmem_data[94][2] ), .B1(n28481), .B2(
        \xmem_data[95][2] ), .ZN(n22966) );
  NAND4_X1 U26782 ( .A1(n22969), .A2(n22968), .A3(n22967), .A4(n22966), .ZN(
        n22970) );
  OR4_X1 U26783 ( .A1(n22973), .A2(n22972), .A3(n22971), .A4(n22970), .ZN(
        n22974) );
  AOI22_X1 U26784 ( .A1(n23751), .A2(n22975), .B1(n23713), .B2(n22974), .ZN(
        n22976) );
  AOI22_X1 U26785 ( .A1(n29419), .A2(\xmem_data[80][1] ), .B1(n29418), .B2(
        \xmem_data[81][1] ), .ZN(n22982) );
  AOI22_X1 U26786 ( .A1(n29420), .A2(\xmem_data[82][1] ), .B1(n23754), .B2(
        \xmem_data[83][1] ), .ZN(n22981) );
  AOI22_X1 U26787 ( .A1(n28136), .A2(\xmem_data[84][1] ), .B1(n27832), .B2(
        \xmem_data[85][1] ), .ZN(n22980) );
  AND2_X1 U26788 ( .A1(n29422), .A2(\xmem_data[87][1] ), .ZN(n22978) );
  AOI21_X1 U26789 ( .B1(n29628), .B2(\xmem_data[86][1] ), .A(n22978), .ZN(
        n22979) );
  NAND4_X1 U26790 ( .A1(n22982), .A2(n22981), .A3(n22980), .A4(n22979), .ZN(
        n22998) );
  AOI22_X1 U26791 ( .A1(n27703), .A2(\xmem_data[92][1] ), .B1(n28665), .B2(
        \xmem_data[93][1] ), .ZN(n22986) );
  AOI22_X1 U26792 ( .A1(n29402), .A2(\xmem_data[90][1] ), .B1(n29350), .B2(
        \xmem_data[91][1] ), .ZN(n22985) );
  AOI22_X1 U26793 ( .A1(n29400), .A2(\xmem_data[88][1] ), .B1(n27833), .B2(
        \xmem_data[89][1] ), .ZN(n22984) );
  AOI22_X1 U26794 ( .A1(n29404), .A2(\xmem_data[94][1] ), .B1(n29403), .B2(
        \xmem_data[95][1] ), .ZN(n22983) );
  NAND4_X1 U26795 ( .A1(n22986), .A2(n22985), .A3(n22984), .A4(n22983), .ZN(
        n22997) );
  AOI22_X1 U26796 ( .A1(n29604), .A2(\xmem_data[64][1] ), .B1(n30084), .B2(
        \xmem_data[65][1] ), .ZN(n22990) );
  AOI22_X1 U26797 ( .A1(n29397), .A2(\xmem_data[66][1] ), .B1(n27818), .B2(
        \xmem_data[67][1] ), .ZN(n22989) );
  AOI22_X1 U26798 ( .A1(n3168), .A2(\xmem_data[68][1] ), .B1(n3187), .B2(
        \xmem_data[69][1] ), .ZN(n22988) );
  AOI22_X1 U26799 ( .A1(n30684), .A2(\xmem_data[70][1] ), .B1(n29410), .B2(
        \xmem_data[71][1] ), .ZN(n22987) );
  NAND4_X1 U26800 ( .A1(n22990), .A2(n22989), .A3(n22988), .A4(n22987), .ZN(
        n22996) );
  AOI22_X1 U26801 ( .A1(n30766), .A2(\xmem_data[72][1] ), .B1(n30685), .B2(
        \xmem_data[73][1] ), .ZN(n22994) );
  AOI22_X1 U26802 ( .A1(n29380), .A2(\xmem_data[74][1] ), .B1(n29379), .B2(
        \xmem_data[75][1] ), .ZN(n22993) );
  AOI22_X1 U26803 ( .A1(n29382), .A2(\xmem_data[76][1] ), .B1(n29381), .B2(
        \xmem_data[77][1] ), .ZN(n22992) );
  AOI22_X1 U26804 ( .A1(n29384), .A2(\xmem_data[78][1] ), .B1(n29383), .B2(
        \xmem_data[79][1] ), .ZN(n22991) );
  NAND4_X1 U26805 ( .A1(n22994), .A2(n22993), .A3(n22992), .A4(n22991), .ZN(
        n22995) );
  AOI22_X1 U26806 ( .A1(n29447), .A2(\xmem_data[48][1] ), .B1(n3124), .B2(
        \xmem_data[49][1] ), .ZN(n23003) );
  AOI22_X1 U26807 ( .A1(n29449), .A2(\xmem_data[50][1] ), .B1(n20828), .B2(
        \xmem_data[51][1] ), .ZN(n23002) );
  AOI22_X1 U26808 ( .A1(n30291), .A2(\xmem_data[52][1] ), .B1(n30707), .B2(
        \xmem_data[53][1] ), .ZN(n23001) );
  AOI22_X1 U26809 ( .A1(n29790), .A2(\xmem_data[54][1] ), .B1(n29431), .B2(
        \xmem_data[55][1] ), .ZN(n23000) );
  NAND4_X1 U26810 ( .A1(n23003), .A2(n23002), .A3(n23001), .A4(n23000), .ZN(
        n23020) );
  AOI22_X1 U26811 ( .A1(n30697), .A2(\xmem_data[56][1] ), .B1(n30293), .B2(
        \xmem_data[57][1] ), .ZN(n23007) );
  AOI22_X1 U26812 ( .A1(n29450), .A2(\xmem_data[58][1] ), .B1(n29350), .B2(
        \xmem_data[59][1] ), .ZN(n23006) );
  AOI22_X1 U26813 ( .A1(n27703), .A2(\xmem_data[60][1] ), .B1(n28738), .B2(
        \xmem_data[61][1] ), .ZN(n23005) );
  AOI22_X1 U26814 ( .A1(n29802), .A2(\xmem_data[62][1] ), .B1(n29451), .B2(
        \xmem_data[63][1] ), .ZN(n23004) );
  NAND4_X1 U26815 ( .A1(n23007), .A2(n23006), .A3(n23005), .A4(n23004), .ZN(
        n23019) );
  AOI22_X1 U26816 ( .A1(n3162), .A2(\xmem_data[36][1] ), .B1(n3188), .B2(
        \xmem_data[37][1] ), .ZN(n23012) );
  AOI22_X1 U26817 ( .A1(n29436), .A2(\xmem_data[32][1] ), .B1(n30301), .B2(
        \xmem_data[33][1] ), .ZN(n23011) );
  AOI22_X1 U26818 ( .A1(n29438), .A2(\xmem_data[34][1] ), .B1(n3157), .B2(
        \xmem_data[35][1] ), .ZN(n23010) );
  AND2_X1 U26819 ( .A1(n29439), .A2(\xmem_data[39][1] ), .ZN(n23008) );
  AOI21_X1 U26820 ( .B1(n26812), .B2(\xmem_data[38][1] ), .A(n23008), .ZN(
        n23009) );
  NAND4_X1 U26821 ( .A1(n23012), .A2(n23011), .A3(n23010), .A4(n23009), .ZN(
        n23018) );
  AOI22_X1 U26822 ( .A1(n29547), .A2(\xmem_data[40][1] ), .B1(n30765), .B2(
        \xmem_data[41][1] ), .ZN(n23016) );
  AOI22_X1 U26823 ( .A1(n29461), .A2(\xmem_data[42][1] ), .B1(n3151), .B2(
        \xmem_data[43][1] ), .ZN(n23015) );
  AOI22_X1 U26824 ( .A1(n29463), .A2(\xmem_data[44][1] ), .B1(n29462), .B2(
        \xmem_data[45][1] ), .ZN(n23014) );
  AOI22_X1 U26825 ( .A1(n29464), .A2(\xmem_data[46][1] ), .B1(n20826), .B2(
        \xmem_data[47][1] ), .ZN(n23013) );
  NAND4_X1 U26826 ( .A1(n23016), .A2(n23015), .A3(n23014), .A4(n23013), .ZN(
        n23017) );
  NAND2_X1 U26827 ( .A1(n23021), .A2(n29471), .ZN(n23073) );
  AOI22_X1 U26828 ( .A1(n29419), .A2(\xmem_data[112][1] ), .B1(n29418), .B2(
        \xmem_data[113][1] ), .ZN(n23026) );
  AOI22_X1 U26829 ( .A1(n29420), .A2(\xmem_data[114][1] ), .B1(n3318), .B2(
        \xmem_data[115][1] ), .ZN(n23025) );
  AOI22_X1 U26830 ( .A1(n29788), .A2(\xmem_data[116][1] ), .B1(n30222), .B2(
        \xmem_data[117][1] ), .ZN(n23024) );
  AND2_X1 U26831 ( .A1(n29422), .A2(\xmem_data[119][1] ), .ZN(n23022) );
  AOI21_X1 U26832 ( .B1(n28138), .B2(\xmem_data[118][1] ), .A(n23022), .ZN(
        n23023) );
  NAND4_X1 U26833 ( .A1(n23026), .A2(n23025), .A3(n23024), .A4(n23023), .ZN(
        n23043) );
  AOI22_X1 U26834 ( .A1(n29400), .A2(\xmem_data[120][1] ), .B1(n3197), .B2(
        \xmem_data[121][1] ), .ZN(n23030) );
  AOI22_X1 U26835 ( .A1(n29402), .A2(\xmem_data[122][1] ), .B1(n23742), .B2(
        \xmem_data[123][1] ), .ZN(n23029) );
  AOI22_X1 U26836 ( .A1(n29602), .A2(\xmem_data[124][1] ), .B1(n29347), .B2(
        \xmem_data[125][1] ), .ZN(n23028) );
  AOI22_X1 U26837 ( .A1(n29404), .A2(\xmem_data[126][1] ), .B1(n29403), .B2(
        \xmem_data[127][1] ), .ZN(n23027) );
  NAND4_X1 U26838 ( .A1(n23030), .A2(n23029), .A3(n23028), .A4(n23027), .ZN(
        n23042) );
  AOI22_X1 U26839 ( .A1(n3162), .A2(\xmem_data[100][1] ), .B1(n3188), .B2(
        \xmem_data[101][1] ), .ZN(n23035) );
  AOI22_X1 U26840 ( .A1(n29397), .A2(\xmem_data[98][1] ), .B1(n27945), .B2(
        \xmem_data[99][1] ), .ZN(n23034) );
  AOI22_X1 U26841 ( .A1(n29714), .A2(\xmem_data[96][1] ), .B1(n30301), .B2(
        \xmem_data[97][1] ), .ZN(n23033) );
  AND2_X1 U26842 ( .A1(n29410), .A2(\xmem_data[103][1] ), .ZN(n23031) );
  NAND4_X1 U26843 ( .A1(n23035), .A2(n23034), .A3(n23033), .A4(n23032), .ZN(
        n23041) );
  AOI22_X1 U26844 ( .A1(n30063), .A2(\xmem_data[104][1] ), .B1(n30266), .B2(
        \xmem_data[105][1] ), .ZN(n23039) );
  AOI22_X1 U26845 ( .A1(n29380), .A2(\xmem_data[106][1] ), .B1(n29379), .B2(
        \xmem_data[107][1] ), .ZN(n23038) );
  AOI22_X1 U26846 ( .A1(n29382), .A2(\xmem_data[108][1] ), .B1(n29381), .B2(
        \xmem_data[109][1] ), .ZN(n23037) );
  AOI22_X1 U26847 ( .A1(n29384), .A2(\xmem_data[110][1] ), .B1(n29383), .B2(
        \xmem_data[111][1] ), .ZN(n23036) );
  NAND4_X1 U26848 ( .A1(n23039), .A2(n23038), .A3(n23037), .A4(n23036), .ZN(
        n23040) );
  NAND2_X1 U26849 ( .A1(n23044), .A2(n29428), .ZN(n23072) );
  AOI22_X1 U26850 ( .A1(n3164), .A2(\xmem_data[4][1] ), .B1(n3187), .B2(
        \xmem_data[5][1] ), .ZN(n23051) );
  AOI22_X1 U26851 ( .A1(n29501), .A2(\xmem_data[26][1] ), .B1(n3375), .B2(
        \xmem_data[27][1] ), .ZN(n23047) );
  AOI22_X1 U26852 ( .A1(n29500), .A2(\xmem_data[30][1] ), .B1(n28233), .B2(
        \xmem_data[31][1] ), .ZN(n23046) );
  AOI22_X1 U26853 ( .A1(n7275), .A2(\xmem_data[16][1] ), .B1(n29497), .B2(
        \xmem_data[17][1] ), .ZN(n23045) );
  NAND3_X1 U26854 ( .A1(n23047), .A2(n23046), .A3(n23045), .ZN(n23048) );
  AOI21_X1 U26855 ( .B1(n29810), .B2(\xmem_data[6][1] ), .A(n23048), .ZN(
        n23050) );
  AOI22_X1 U26856 ( .A1(n28136), .A2(\xmem_data[20][1] ), .B1(n30293), .B2(
        \xmem_data[25][1] ), .ZN(n23049) );
  AOI22_X1 U26857 ( .A1(n29547), .A2(\xmem_data[8][1] ), .B1(n30266), .B2(
        \xmem_data[9][1] ), .ZN(n23055) );
  AOI22_X1 U26858 ( .A1(n7270), .A2(\xmem_data[10][1] ), .B1(n3307), .B2(
        \xmem_data[11][1] ), .ZN(n23054) );
  AOI22_X1 U26859 ( .A1(n29724), .A2(\xmem_data[12][1] ), .B1(n29462), .B2(
        \xmem_data[13][1] ), .ZN(n23053) );
  AOI22_X1 U26860 ( .A1(n29489), .A2(\xmem_data[14][1] ), .B1(n27568), .B2(
        \xmem_data[15][1] ), .ZN(n23052) );
  NAND2_X1 U26861 ( .A1(n3392), .A2(\xmem_data[22][1] ), .ZN(n23057) );
  AOI22_X1 U26862 ( .A1(n27754), .A2(\xmem_data[0][1] ), .B1(n26884), .B2(
        \xmem_data[1][1] ), .ZN(n23056) );
  NAND2_X1 U26863 ( .A1(n23057), .A2(n23056), .ZN(n23066) );
  NAND2_X1 U26864 ( .A1(n28209), .A2(\xmem_data[24][1] ), .ZN(n23064) );
  AOI22_X1 U26865 ( .A1(n29499), .A2(\xmem_data[18][1] ), .B1(n3149), .B2(
        \xmem_data[19][1] ), .ZN(n23063) );
  AOI22_X1 U26866 ( .A1(n29475), .A2(\xmem_data[2][1] ), .B1(n29315), .B2(
        \xmem_data[3][1] ), .ZN(n23058) );
  NAND2_X1 U26867 ( .A1(n29494), .A2(\xmem_data[23][1] ), .ZN(n23060) );
  NAND2_X1 U26868 ( .A1(n28754), .A2(\xmem_data[7][1] ), .ZN(n23059) );
  NAND2_X1 U26869 ( .A1(n23060), .A2(n23059), .ZN(n23061) );
  AOI21_X1 U26870 ( .B1(n30222), .B2(\xmem_data[21][1] ), .A(n23061), .ZN(
        n23062) );
  NAND4_X1 U26871 ( .A1(n23064), .A2(n23063), .A3(n23058), .A4(n23062), .ZN(
        n23065) );
  NOR2_X1 U26872 ( .A1(n23066), .A2(n23065), .ZN(n23068) );
  AOI22_X1 U26873 ( .A1(n30248), .A2(\xmem_data[28][1] ), .B1(n30190), .B2(
        \xmem_data[29][1] ), .ZN(n23067) );
  NAND4_X1 U26874 ( .A1(n23069), .A2(n3820), .A3(n23068), .A4(n23067), .ZN(
        n23070) );
  NAND2_X1 U26875 ( .A1(n23070), .A2(n29511), .ZN(n23071) );
  NAND4_X2 U26876 ( .A1(n23074), .A2(n23073), .A3(n23072), .A4(n23071), .ZN(
        n34783) );
  XNOR2_X1 U26877 ( .A(n34783), .B(\fmem_data[3][5] ), .ZN(n31174) );
  XNOR2_X1 U26878 ( .A(n33720), .B(\fmem_data[3][5] ), .ZN(n32153) );
  OAI22_X1 U26879 ( .A1(n34918), .A2(n31174), .B1(n32153), .B2(n34919), .ZN(
        n28537) );
  NAND2_X1 U26880 ( .A1(n28535), .A2(n28537), .ZN(n23165) );
  XNOR2_X1 U26881 ( .A(n31492), .B(\fmem_data[25][3] ), .ZN(n31443) );
  AOI22_X1 U26882 ( .A1(n29089), .A2(\xmem_data[64][4] ), .B1(n3301), .B2(
        \xmem_data[65][4] ), .ZN(n23078) );
  AOI22_X1 U26883 ( .A1(n28098), .A2(\xmem_data[66][4] ), .B1(n29151), .B2(
        \xmem_data[67][4] ), .ZN(n23077) );
  AOI22_X1 U26884 ( .A1(n29086), .A2(\xmem_data[68][4] ), .B1(n28772), .B2(
        \xmem_data[69][4] ), .ZN(n23076) );
  AOI22_X1 U26885 ( .A1(n22727), .A2(\xmem_data[70][4] ), .B1(n28076), .B2(
        \xmem_data[71][4] ), .ZN(n23075) );
  NAND4_X1 U26886 ( .A1(n23078), .A2(n23077), .A3(n23076), .A4(n23075), .ZN(
        n23095) );
  AND2_X1 U26887 ( .A1(n30863), .A2(\xmem_data[74][4] ), .ZN(n23079) );
  AOI21_X1 U26888 ( .B1(n27502), .B2(\xmem_data[75][4] ), .A(n23079), .ZN(
        n23083) );
  AOI22_X1 U26889 ( .A1(n21309), .A2(\xmem_data[72][4] ), .B1(n28039), .B2(
        \xmem_data[73][4] ), .ZN(n23082) );
  AOI22_X1 U26890 ( .A1(n3219), .A2(\xmem_data[76][4] ), .B1(n30964), .B2(
        \xmem_data[77][4] ), .ZN(n23081) );
  AOI22_X1 U26891 ( .A1(n29095), .A2(\xmem_data[78][4] ), .B1(n29027), .B2(
        \xmem_data[79][4] ), .ZN(n23080) );
  NAND4_X1 U26892 ( .A1(n23083), .A2(n23082), .A3(n23081), .A4(n23080), .ZN(
        n23094) );
  AOI22_X1 U26893 ( .A1(n29104), .A2(\xmem_data[80][4] ), .B1(n29157), .B2(
        \xmem_data[81][4] ), .ZN(n23087) );
  AOI22_X1 U26894 ( .A1(n29103), .A2(\xmem_data[82][4] ), .B1(n25422), .B2(
        \xmem_data[83][4] ), .ZN(n23086) );
  AOI22_X1 U26895 ( .A1(n25456), .A2(\xmem_data[84][4] ), .B1(n24640), .B2(
        \xmem_data[85][4] ), .ZN(n23085) );
  AOI22_X1 U26896 ( .A1(n24516), .A2(\xmem_data[86][4] ), .B1(n29109), .B2(
        \xmem_data[87][4] ), .ZN(n23084) );
  NAND4_X1 U26897 ( .A1(n23087), .A2(n23086), .A3(n23085), .A4(n23084), .ZN(
        n23093) );
  AOI22_X1 U26898 ( .A1(n30513), .A2(\xmem_data[88][4] ), .B1(n29187), .B2(
        \xmem_data[89][4] ), .ZN(n23091) );
  AOI22_X1 U26899 ( .A1(n25574), .A2(\xmem_data[90][4] ), .B1(n20585), .B2(
        \xmem_data[91][4] ), .ZN(n23090) );
  AOI22_X1 U26900 ( .A1(n25398), .A2(\xmem_data[92][4] ), .B1(n20815), .B2(
        \xmem_data[93][4] ), .ZN(n23089) );
  AOI22_X1 U26901 ( .A1(n29101), .A2(\xmem_data[94][4] ), .B1(n30899), .B2(
        \xmem_data[95][4] ), .ZN(n23088) );
  NAND4_X1 U26902 ( .A1(n23091), .A2(n23090), .A3(n23089), .A4(n23088), .ZN(
        n23092) );
  OR4_X1 U26903 ( .A1(n23095), .A2(n23094), .A3(n23093), .A4(n23092), .ZN(
        n23117) );
  AOI22_X1 U26904 ( .A1(n24470), .A2(\xmem_data[104][4] ), .B1(n23732), .B2(
        \xmem_data[105][4] ), .ZN(n23099) );
  AOI22_X1 U26905 ( .A1(n29173), .A2(\xmem_data[106][4] ), .B1(n24694), .B2(
        \xmem_data[107][4] ), .ZN(n23098) );
  AOI22_X1 U26906 ( .A1(n3217), .A2(\xmem_data[108][4] ), .B1(n29431), .B2(
        \xmem_data[109][4] ), .ZN(n23097) );
  AOI22_X1 U26907 ( .A1(n22710), .A2(\xmem_data[110][4] ), .B1(n29174), .B2(
        \xmem_data[111][4] ), .ZN(n23096) );
  NAND4_X1 U26908 ( .A1(n23099), .A2(n23098), .A3(n23097), .A4(n23096), .ZN(
        n23115) );
  AOI22_X1 U26909 ( .A1(n28327), .A2(\xmem_data[96][4] ), .B1(n3307), .B2(
        \xmem_data[97][4] ), .ZN(n23103) );
  AOI22_X1 U26910 ( .A1(n29126), .A2(\xmem_data[98][4] ), .B1(n29151), .B2(
        \xmem_data[99][4] ), .ZN(n23102) );
  AOI22_X1 U26911 ( .A1(n28500), .A2(\xmem_data[100][4] ), .B1(n27852), .B2(
        \xmem_data[101][4] ), .ZN(n23101) );
  AOI22_X1 U26912 ( .A1(n20951), .A2(\xmem_data[102][4] ), .B1(n24688), .B2(
        \xmem_data[103][4] ), .ZN(n23100) );
  NAND4_X1 U26913 ( .A1(n23103), .A2(n23102), .A3(n23101), .A4(n23100), .ZN(
        n23114) );
  AOI22_X1 U26914 ( .A1(n29181), .A2(\xmem_data[112][4] ), .B1(n27396), .B2(
        \xmem_data[113][4] ), .ZN(n23107) );
  AOI22_X1 U26915 ( .A1(n28045), .A2(\xmem_data[114][4] ), .B1(n30885), .B2(
        \xmem_data[115][4] ), .ZN(n23106) );
  AOI22_X1 U26916 ( .A1(n29180), .A2(\xmem_data[116][4] ), .B1(n29179), .B2(
        \xmem_data[117][4] ), .ZN(n23105) );
  AOI22_X1 U26917 ( .A1(n22702), .A2(\xmem_data[118][4] ), .B1(n28298), .B2(
        \xmem_data[119][4] ), .ZN(n23104) );
  NAND4_X1 U26918 ( .A1(n23107), .A2(n23106), .A3(n23105), .A4(n23104), .ZN(
        n23113) );
  AOI22_X1 U26919 ( .A1(n22741), .A2(\xmem_data[120][4] ), .B1(n29187), .B2(
        \xmem_data[121][4] ), .ZN(n23111) );
  AOI22_X1 U26920 ( .A1(n20543), .A2(\xmem_data[122][4] ), .B1(n20585), .B2(
        \xmem_data[123][4] ), .ZN(n23110) );
  AOI22_X1 U26921 ( .A1(n16989), .A2(\xmem_data[124][4] ), .B1(n24710), .B2(
        \xmem_data[125][4] ), .ZN(n23109) );
  AOI22_X1 U26922 ( .A1(n29190), .A2(\xmem_data[126][4] ), .B1(n3205), .B2(
        \xmem_data[127][4] ), .ZN(n23108) );
  NAND4_X1 U26923 ( .A1(n23111), .A2(n23110), .A3(n23109), .A4(n23108), .ZN(
        n23112) );
  OR4_X1 U26924 ( .A1(n23115), .A2(n23114), .A3(n23113), .A4(n23112), .ZN(
        n23116) );
  AOI22_X1 U26925 ( .A1(n23117), .A2(n29201), .B1(n23116), .B2(n29171), .ZN(
        n23163) );
  AOI22_X1 U26926 ( .A1(n28517), .A2(\xmem_data[24][4] ), .B1(n29187), .B2(
        \xmem_data[25][4] ), .ZN(n23121) );
  AOI22_X1 U26927 ( .A1(n29188), .A2(\xmem_data[26][4] ), .B1(n24708), .B2(
        \xmem_data[27][4] ), .ZN(n23120) );
  AOI22_X1 U26928 ( .A1(n25398), .A2(\xmem_data[28][4] ), .B1(n28687), .B2(
        \xmem_data[29][4] ), .ZN(n23119) );
  AOI22_X1 U26929 ( .A1(n27523), .A2(\xmem_data[30][4] ), .B1(n20593), .B2(
        \xmem_data[31][4] ), .ZN(n23118) );
  AOI22_X1 U26930 ( .A1(n13444), .A2(\xmem_data[16][4] ), .B1(n27396), .B2(
        \xmem_data[17][4] ), .ZN(n23125) );
  AOI22_X1 U26931 ( .A1(n28007), .A2(\xmem_data[18][4] ), .B1(n23813), .B2(
        \xmem_data[19][4] ), .ZN(n23124) );
  AOI22_X1 U26932 ( .A1(n24158), .A2(\xmem_data[20][4] ), .B1(n20545), .B2(
        \xmem_data[21][4] ), .ZN(n23123) );
  AOI22_X1 U26933 ( .A1(n13168), .A2(\xmem_data[22][4] ), .B1(n16986), .B2(
        \xmem_data[23][4] ), .ZN(n23122) );
  AOI22_X1 U26934 ( .A1(n20711), .A2(\xmem_data[10][4] ), .B1(n28044), .B2(
        \xmem_data[11][4] ), .ZN(n23138) );
  AOI22_X1 U26935 ( .A1(n29125), .A2(\xmem_data[6][4] ), .B1(n29124), .B2(
        \xmem_data[7][4] ), .ZN(n23129) );
  AOI22_X1 U26936 ( .A1(n27365), .A2(\xmem_data[2][4] ), .B1(n21058), .B2(
        \xmem_data[3][4] ), .ZN(n23128) );
  AOI22_X1 U26937 ( .A1(n25562), .A2(\xmem_data[14][4] ), .B1(n22709), .B2(
        \xmem_data[15][4] ), .ZN(n23127) );
  AOI22_X1 U26938 ( .A1(n3219), .A2(\xmem_data[12][4] ), .B1(n30593), .B2(
        \xmem_data[13][4] ), .ZN(n23126) );
  NAND4_X1 U26939 ( .A1(n23129), .A2(n23128), .A3(n23127), .A4(n23126), .ZN(
        n23136) );
  AOI22_X1 U26940 ( .A1(n21009), .A2(\xmem_data[0][4] ), .B1(n3330), .B2(
        \xmem_data[1][4] ), .ZN(n23131) );
  NAND2_X1 U26941 ( .A1(n29136), .A2(\xmem_data[4][4] ), .ZN(n23130) );
  NAND2_X1 U26942 ( .A1(n23131), .A2(n23130), .ZN(n23135) );
  AOI21_X1 U26943 ( .B1(n29118), .B2(\xmem_data[8][4] ), .A(n3737), .ZN(n23133) );
  NAND2_X1 U26944 ( .A1(n28772), .A2(\xmem_data[5][4] ), .ZN(n23132) );
  NAND2_X1 U26945 ( .A1(n23133), .A2(n23132), .ZN(n23134) );
  NOR3_X1 U26946 ( .A1(n23136), .A2(n23135), .A3(n23134), .ZN(n23137) );
  NAND4_X1 U26947 ( .A1(n3831), .A2(n3533), .A3(n23138), .A4(n23137), .ZN(
        n23161) );
  AND2_X1 U26948 ( .A1(n28501), .A2(\xmem_data[42][4] ), .ZN(n23139) );
  AOI21_X1 U26949 ( .B1(n24631), .B2(\xmem_data[43][4] ), .A(n23139), .ZN(
        n23143) );
  AOI22_X1 U26950 ( .A1(n28037), .A2(\xmem_data[40][4] ), .B1(n27813), .B2(
        \xmem_data[41][4] ), .ZN(n23142) );
  AOI22_X1 U26951 ( .A1(n3222), .A2(\xmem_data[44][4] ), .B1(n24533), .B2(
        \xmem_data[45][4] ), .ZN(n23141) );
  AOI22_X1 U26952 ( .A1(n29095), .A2(\xmem_data[46][4] ), .B1(n22758), .B2(
        \xmem_data[47][4] ), .ZN(n23140) );
  NAND4_X1 U26953 ( .A1(n23143), .A2(n23142), .A3(n23141), .A4(n23140), .ZN(
        n23159) );
  AOI22_X1 U26954 ( .A1(n29089), .A2(\xmem_data[32][4] ), .B1(n24522), .B2(
        \xmem_data[33][4] ), .ZN(n23147) );
  AOI22_X1 U26955 ( .A1(n27975), .A2(\xmem_data[34][4] ), .B1(n30497), .B2(
        \xmem_data[35][4] ), .ZN(n23146) );
  AOI22_X1 U26956 ( .A1(n29086), .A2(\xmem_data[36][4] ), .B1(n29327), .B2(
        \xmem_data[37][4] ), .ZN(n23145) );
  AOI22_X1 U26957 ( .A1(n25528), .A2(\xmem_data[38][4] ), .B1(n27959), .B2(
        \xmem_data[39][4] ), .ZN(n23144) );
  NAND4_X1 U26958 ( .A1(n23147), .A2(n23146), .A3(n23145), .A4(n23144), .ZN(
        n23158) );
  AOI22_X1 U26959 ( .A1(n29104), .A2(\xmem_data[48][4] ), .B1(n27396), .B2(
        \xmem_data[49][4] ), .ZN(n23151) );
  AOI22_X1 U26960 ( .A1(n29103), .A2(\xmem_data[50][4] ), .B1(n27447), .B2(
        \xmem_data[51][4] ), .ZN(n23150) );
  AOI22_X1 U26961 ( .A1(n3357), .A2(\xmem_data[52][4] ), .B1(n30508), .B2(
        \xmem_data[53][4] ), .ZN(n23149) );
  AOI22_X1 U26962 ( .A1(n28375), .A2(\xmem_data[54][4] ), .B1(n29109), .B2(
        \xmem_data[55][4] ), .ZN(n23148) );
  NAND4_X1 U26963 ( .A1(n23151), .A2(n23150), .A3(n23149), .A4(n23148), .ZN(
        n23157) );
  AOI22_X1 U26964 ( .A1(n25671), .A2(\xmem_data[56][4] ), .B1(n3464), .B2(
        \xmem_data[57][4] ), .ZN(n23155) );
  AOI22_X1 U26965 ( .A1(n29188), .A2(\xmem_data[58][4] ), .B1(n24509), .B2(
        \xmem_data[59][4] ), .ZN(n23154) );
  AOI22_X1 U26966 ( .A1(n31270), .A2(\xmem_data[60][4] ), .B1(n27855), .B2(
        \xmem_data[61][4] ), .ZN(n23153) );
  AOI22_X1 U26967 ( .A1(n29101), .A2(\xmem_data[62][4] ), .B1(n24615), .B2(
        \xmem_data[63][4] ), .ZN(n23152) );
  NAND4_X1 U26968 ( .A1(n23155), .A2(n23154), .A3(n23153), .A4(n23152), .ZN(
        n23156) );
  OR4_X1 U26969 ( .A1(n23159), .A2(n23158), .A3(n23157), .A4(n23156), .ZN(
        n23160) );
  AOI22_X1 U26970 ( .A1(n23161), .A2(n29143), .B1(n23160), .B2(n29145), .ZN(
        n23162) );
  XNOR2_X1 U26971 ( .A(n33246), .B(\fmem_data[25][3] ), .ZN(n29209) );
  OAI21_X1 U26972 ( .B1(n28537), .B2(n28535), .A(n28536), .ZN(n23164) );
  NAND2_X1 U26973 ( .A1(n23165), .A2(n23164), .ZN(n33887) );
  FA_X1 U26974 ( .A(n23168), .B(n23167), .CI(n23166), .CO(n23175), .S(n33886)
         );
  XNOR2_X1 U26975 ( .A(n23170), .B(n23169), .ZN(n23172) );
  XNOR2_X1 U26976 ( .A(n23172), .B(n23171), .ZN(n34147) );
  XNOR2_X1 U26977 ( .A(n23176), .B(n23175), .ZN(n34148) );
  OAI21_X1 U26978 ( .B1(n34149), .B2(n34147), .A(n34148), .ZN(n23178) );
  NAND2_X1 U26979 ( .A1(n34149), .A2(n34147), .ZN(n23177) );
  NAND2_X1 U26980 ( .A1(n23178), .A2(n23177), .ZN(n27318) );
  OAI21_X1 U26981 ( .B1(n27316), .B2(n27317), .A(n27318), .ZN(n23180) );
  NAND2_X1 U26982 ( .A1(n27316), .A2(n27317), .ZN(n23179) );
  NAND2_X1 U26983 ( .A1(n23180), .A2(n23179), .ZN(n27315) );
  FA_X1 U26984 ( .A(n23183), .B(n23182), .CI(n23181), .CO(n26260), .S(n34165)
         );
  FA_X1 U26985 ( .A(n23186), .B(n23185), .CI(n23184), .CO(n26261), .S(n34164)
         );
  FA_X1 U26986 ( .A(n23189), .B(n23188), .CI(n23187), .CO(n23174), .S(n28920)
         );
  AOI22_X1 U26987 ( .A1(n24623), .A2(\xmem_data[32][1] ), .B1(n24622), .B2(
        \xmem_data[33][1] ), .ZN(n23195) );
  AOI22_X1 U26988 ( .A1(n20552), .A2(\xmem_data[34][1] ), .B1(n28292), .B2(
        \xmem_data[35][1] ), .ZN(n23194) );
  AND2_X1 U26989 ( .A1(n24624), .A2(\xmem_data[37][1] ), .ZN(n23190) );
  AOI21_X1 U26990 ( .B1(n29298), .B2(\xmem_data[36][1] ), .A(n23190), .ZN(
        n23193) );
  AND2_X1 U26991 ( .A1(n25358), .A2(\xmem_data[38][1] ), .ZN(n23191) );
  AOI21_X1 U26992 ( .B1(n3203), .B2(\xmem_data[39][1] ), .A(n23191), .ZN(
        n23192) );
  AND4_X1 U26993 ( .A1(n23195), .A2(n23194), .A3(n23193), .A4(n23192), .ZN(
        n23204) );
  AOI22_X1 U26994 ( .A1(n28053), .A2(\xmem_data[56][1] ), .B1(n23716), .B2(
        \xmem_data[57][1] ), .ZN(n23199) );
  AOI22_X1 U26995 ( .A1(n24647), .A2(\xmem_data[62][1] ), .B1(n20816), .B2(
        \xmem_data[63][1] ), .ZN(n23198) );
  AOI22_X1 U26996 ( .A1(n29319), .A2(\xmem_data[60][1] ), .B1(n24646), .B2(
        \xmem_data[61][1] ), .ZN(n23197) );
  AOI22_X1 U26997 ( .A1(n24214), .A2(\xmem_data[58][1] ), .B1(n24645), .B2(
        \xmem_data[59][1] ), .ZN(n23196) );
  NAND4_X1 U26998 ( .A1(n23199), .A2(n23198), .A3(n23197), .A4(n23196), .ZN(
        n23202) );
  AOI22_X1 U26999 ( .A1(n3282), .A2(\xmem_data[48][1] ), .B1(n25492), .B2(
        \xmem_data[49][1] ), .ZN(n23200) );
  INV_X1 U27000 ( .A(n23200), .ZN(n23201) );
  NOR2_X1 U27001 ( .A1(n23202), .A2(n23201), .ZN(n23203) );
  NAND2_X1 U27002 ( .A1(n23204), .A2(n23203), .ZN(n23216) );
  AOI22_X1 U27003 ( .A1(n24630), .A2(\xmem_data[40][1] ), .B1(n3247), .B2(
        \xmem_data[41][1] ), .ZN(n23209) );
  AND2_X1 U27004 ( .A1(n3219), .A2(\xmem_data[43][1] ), .ZN(n23205) );
  AOI21_X1 U27005 ( .B1(n24631), .B2(\xmem_data[42][1] ), .A(n23205), .ZN(
        n23208) );
  AOI22_X1 U27006 ( .A1(n24632), .A2(\xmem_data[44][1] ), .B1(n25491), .B2(
        \xmem_data[45][1] ), .ZN(n23207) );
  AOI22_X1 U27007 ( .A1(n3341), .A2(\xmem_data[46][1] ), .B1(n24633), .B2(
        \xmem_data[47][1] ), .ZN(n23206) );
  NAND4_X1 U27008 ( .A1(n23209), .A2(n23208), .A3(n23207), .A4(n23206), .ZN(
        n23214) );
  AOI22_X1 U27009 ( .A1(n24640), .A2(\xmem_data[52][1] ), .B1(n24639), .B2(
        \xmem_data[53][1] ), .ZN(n23212) );
  AOI22_X1 U27010 ( .A1(n20541), .A2(\xmem_data[54][1] ), .B1(n29271), .B2(
        \xmem_data[55][1] ), .ZN(n23211) );
  AOI22_X1 U27011 ( .A1(n24638), .A2(\xmem_data[50][1] ), .B1(n28373), .B2(
        \xmem_data[51][1] ), .ZN(n23210) );
  NAND3_X1 U27012 ( .A1(n23212), .A2(n23211), .A3(n23210), .ZN(n23213) );
  OR2_X1 U27013 ( .A1(n23214), .A2(n23213), .ZN(n23215) );
  OAI21_X1 U27014 ( .B1(n23216), .B2(n23215), .A(n24659), .ZN(n23241) );
  AOI22_X1 U27015 ( .A1(n30295), .A2(\xmem_data[16][1] ), .B1(n28045), .B2(
        \xmem_data[17][1] ), .ZN(n23218) );
  AOI22_X1 U27016 ( .A1(n25717), .A2(\xmem_data[30][1] ), .B1(n28462), .B2(
        \xmem_data[31][1] ), .ZN(n23217) );
  NAND3_X1 U27017 ( .A1(n23241), .A2(n23218), .A3(n23217), .ZN(n23244) );
  NAND2_X1 U27018 ( .A1(n27910), .A2(\xmem_data[18][1] ), .ZN(n23240) );
  AOI22_X1 U27019 ( .A1(n29439), .A2(\xmem_data[28][1] ), .B1(n24592), .B2(
        \xmem_data[29][1] ), .ZN(n23224) );
  AOI22_X1 U27020 ( .A1(n30943), .A2(\xmem_data[20][1] ), .B1(n13168), .B2(
        \xmem_data[21][1] ), .ZN(n23223) );
  NAND2_X1 U27021 ( .A1(n24590), .A2(\xmem_data[19][1] ), .ZN(n23220) );
  NAND2_X1 U27022 ( .A1(n28516), .A2(\xmem_data[24][1] ), .ZN(n23219) );
  NAND2_X1 U27023 ( .A1(n23220), .A2(n23219), .ZN(n23221) );
  AOI21_X1 U27024 ( .B1(\xmem_data[23][1] ), .B2(n24597), .A(n23221), .ZN(
        n23222) );
  NAND3_X1 U27025 ( .A1(n23224), .A2(n23223), .A3(n23222), .ZN(n23235) );
  AOI22_X1 U27026 ( .A1(n27813), .A2(\xmem_data[8][1] ), .B1(n3247), .B2(
        \xmem_data[9][1] ), .ZN(n23228) );
  AOI22_X1 U27027 ( .A1(n24694), .A2(\xmem_data[10][1] ), .B1(n3217), .B2(
        \xmem_data[11][1] ), .ZN(n23227) );
  AOI22_X1 U27028 ( .A1(n30593), .A2(\xmem_data[12][1] ), .B1(n28476), .B2(
        \xmem_data[13][1] ), .ZN(n23226) );
  AOI22_X1 U27029 ( .A1(n3340), .A2(\xmem_data[14][1] ), .B1(n30882), .B2(
        \xmem_data[15][1] ), .ZN(n23225) );
  NAND4_X1 U27030 ( .A1(n23228), .A2(n23227), .A3(n23226), .A4(n23225), .ZN(
        n23234) );
  AOI22_X1 U27031 ( .A1(n30269), .A2(\xmem_data[0][1] ), .B1(n24622), .B2(
        \xmem_data[1][1] ), .ZN(n23232) );
  AOI22_X1 U27032 ( .A1(n24606), .A2(\xmem_data[2][1] ), .B1(n30496), .B2(
        \xmem_data[3][1] ), .ZN(n23231) );
  AOI22_X1 U27033 ( .A1(n20567), .A2(\xmem_data[4][1] ), .B1(n20707), .B2(
        \xmem_data[5][1] ), .ZN(n23230) );
  AOI22_X1 U27034 ( .A1(n24607), .A2(\xmem_data[6][1] ), .B1(n30571), .B2(
        \xmem_data[7][1] ), .ZN(n23229) );
  NAND4_X1 U27035 ( .A1(n23232), .A2(n23231), .A3(n23230), .A4(n23229), .ZN(
        n23233) );
  OR3_X1 U27036 ( .A1(n23235), .A2(n23234), .A3(n23233), .ZN(n23236) );
  AOI21_X1 U27037 ( .B1(n25383), .B2(\xmem_data[25][1] ), .A(n23236), .ZN(
        n23239) );
  AOI22_X1 U27038 ( .A1(n24593), .A2(\xmem_data[26][1] ), .B1(n14912), .B2(
        \xmem_data[27][1] ), .ZN(n23238) );
  NAND2_X1 U27039 ( .A1(n30614), .A2(\xmem_data[22][1] ), .ZN(n23237) );
  NAND4_X1 U27040 ( .A1(n23240), .A2(n23239), .A3(n23238), .A4(n23237), .ZN(
        n23243) );
  NAND2_X1 U27041 ( .A1(n23241), .A2(n24662), .ZN(n23242) );
  OAI21_X1 U27042 ( .B1(n23244), .B2(n23243), .A(n23242), .ZN(n23288) );
  AOI22_X1 U27043 ( .A1(n29246), .A2(\xmem_data[96][1] ), .B1(n23779), .B2(
        \xmem_data[97][1] ), .ZN(n23248) );
  AOI22_X1 U27044 ( .A1(n24685), .A2(\xmem_data[98][1] ), .B1(n28468), .B2(
        \xmem_data[99][1] ), .ZN(n23247) );
  AOI22_X1 U27045 ( .A1(n24687), .A2(\xmem_data[100][1] ), .B1(n24686), .B2(
        \xmem_data[101][1] ), .ZN(n23246) );
  AOI22_X1 U27046 ( .A1(n24688), .A2(\xmem_data[102][1] ), .B1(n31346), .B2(
        \xmem_data[103][1] ), .ZN(n23245) );
  NAND4_X1 U27047 ( .A1(n23248), .A2(n23247), .A3(n23246), .A4(n23245), .ZN(
        n23264) );
  AOI22_X1 U27048 ( .A1(n24693), .A2(\xmem_data[104][1] ), .B1(n30863), .B2(
        \xmem_data[105][1] ), .ZN(n23252) );
  AOI22_X1 U27049 ( .A1(n24694), .A2(\xmem_data[106][1] ), .B1(n3219), .B2(
        \xmem_data[107][1] ), .ZN(n23251) );
  AOI22_X1 U27050 ( .A1(n24696), .A2(\xmem_data[108][1] ), .B1(n24695), .B2(
        \xmem_data[109][1] ), .ZN(n23250) );
  AOI22_X1 U27051 ( .A1(n24697), .A2(\xmem_data[110][1] ), .B1(n17061), .B2(
        \xmem_data[111][1] ), .ZN(n23249) );
  NAND4_X1 U27052 ( .A1(n23252), .A2(n23251), .A3(n23250), .A4(n23249), .ZN(
        n23263) );
  AOI22_X1 U27053 ( .A1(n24702), .A2(\xmem_data[112][1] ), .B1(n25450), .B2(
        \xmem_data[113][1] ), .ZN(n23256) );
  AOI22_X1 U27054 ( .A1(n27447), .A2(\xmem_data[114][1] ), .B1(n28481), .B2(
        \xmem_data[115][1] ), .ZN(n23255) );
  AOI22_X1 U27055 ( .A1(n29308), .A2(\xmem_data[116][1] ), .B1(n13168), .B2(
        \xmem_data[117][1] ), .ZN(n23254) );
  AOI22_X1 U27056 ( .A1(n16986), .A2(\xmem_data[118][1] ), .B1(n27912), .B2(
        \xmem_data[119][1] ), .ZN(n23253) );
  NAND4_X1 U27057 ( .A1(n23256), .A2(n23255), .A3(n23254), .A4(n23253), .ZN(
        n23262) );
  AOI22_X1 U27058 ( .A1(n28752), .A2(\xmem_data[120][1] ), .B1(n27864), .B2(
        \xmem_data[121][1] ), .ZN(n23260) );
  AOI22_X1 U27059 ( .A1(n24708), .A2(\xmem_data[122][1] ), .B1(n24707), .B2(
        \xmem_data[123][1] ), .ZN(n23259) );
  AOI22_X1 U27060 ( .A1(n24710), .A2(\xmem_data[124][1] ), .B1(n24709), .B2(
        \xmem_data[125][1] ), .ZN(n23258) );
  AOI22_X1 U27061 ( .A1(n28385), .A2(\xmem_data[126][1] ), .B1(n17001), .B2(
        \xmem_data[127][1] ), .ZN(n23257) );
  NAND4_X1 U27062 ( .A1(n23260), .A2(n23259), .A3(n23258), .A4(n23257), .ZN(
        n23261) );
  OR4_X1 U27063 ( .A1(n23264), .A2(n23263), .A3(n23262), .A4(n23261), .ZN(
        n23286) );
  AOI22_X1 U27064 ( .A1(n29573), .A2(\xmem_data[64][1] ), .B1(n20553), .B2(
        \xmem_data[65][1] ), .ZN(n23268) );
  AOI22_X1 U27065 ( .A1(n24685), .A2(\xmem_data[66][1] ), .B1(n22751), .B2(
        \xmem_data[67][1] ), .ZN(n23267) );
  AOI22_X1 U27066 ( .A1(n24687), .A2(\xmem_data[68][1] ), .B1(n24686), .B2(
        \xmem_data[69][1] ), .ZN(n23266) );
  AOI22_X1 U27067 ( .A1(n24688), .A2(\xmem_data[70][1] ), .B1(n20489), .B2(
        \xmem_data[71][1] ), .ZN(n23265) );
  NAND4_X1 U27068 ( .A1(n23268), .A2(n23267), .A3(n23266), .A4(n23265), .ZN(
        n23284) );
  AOI22_X1 U27069 ( .A1(n24693), .A2(\xmem_data[72][1] ), .B1(n23731), .B2(
        \xmem_data[73][1] ), .ZN(n23272) );
  AOI22_X1 U27070 ( .A1(n24694), .A2(\xmem_data[74][1] ), .B1(n3222), .B2(
        \xmem_data[75][1] ), .ZN(n23271) );
  AOI22_X1 U27071 ( .A1(n24696), .A2(\xmem_data[76][1] ), .B1(n24695), .B2(
        \xmem_data[77][1] ), .ZN(n23270) );
  AOI22_X1 U27072 ( .A1(n24697), .A2(\xmem_data[78][1] ), .B1(n3255), .B2(
        \xmem_data[79][1] ), .ZN(n23269) );
  NAND4_X1 U27073 ( .A1(n23272), .A2(n23271), .A3(n23270), .A4(n23269), .ZN(
        n23283) );
  AOI22_X1 U27074 ( .A1(n24702), .A2(\xmem_data[80][1] ), .B1(n25450), .B2(
        \xmem_data[81][1] ), .ZN(n23276) );
  AOI22_X1 U27075 ( .A1(n25422), .A2(\xmem_data[82][1] ), .B1(n29307), .B2(
        \xmem_data[83][1] ), .ZN(n23275) );
  AOI22_X1 U27076 ( .A1(n29179), .A2(\xmem_data[84][1] ), .B1(n28416), .B2(
        \xmem_data[85][1] ), .ZN(n23274) );
  AOI22_X1 U27077 ( .A1(n17041), .A2(\xmem_data[86][1] ), .B1(n22674), .B2(
        \xmem_data[87][1] ), .ZN(n23273) );
  NAND4_X1 U27078 ( .A1(n23276), .A2(n23275), .A3(n23274), .A4(n23273), .ZN(
        n23282) );
  AOI22_X1 U27079 ( .A1(n31354), .A2(\xmem_data[88][1] ), .B1(n3207), .B2(
        \xmem_data[89][1] ), .ZN(n23280) );
  AOI22_X1 U27080 ( .A1(n24708), .A2(\xmem_data[90][1] ), .B1(n24707), .B2(
        \xmem_data[91][1] ), .ZN(n23279) );
  AOI22_X1 U27081 ( .A1(n24710), .A2(\xmem_data[92][1] ), .B1(n24709), .B2(
        \xmem_data[93][1] ), .ZN(n23278) );
  AOI22_X1 U27082 ( .A1(n29100), .A2(\xmem_data[94][1] ), .B1(n23778), .B2(
        \xmem_data[95][1] ), .ZN(n23277) );
  NAND4_X1 U27083 ( .A1(n23280), .A2(n23279), .A3(n23278), .A4(n23277), .ZN(
        n23281) );
  OR4_X1 U27084 ( .A1(n23284), .A2(n23283), .A3(n23282), .A4(n23281), .ZN(
        n23285) );
  AOI22_X1 U27085 ( .A1(n24722), .A2(n23286), .B1(n24720), .B2(n23285), .ZN(
        n23287) );
  XNOR2_X1 U27086 ( .A(n33683), .B(\fmem_data[24][5] ), .ZN(n31167) );
  AOI22_X1 U27087 ( .A1(n24623), .A2(\xmem_data[32][2] ), .B1(n24622), .B2(
        \xmem_data[33][2] ), .ZN(n23292) );
  AOI22_X1 U27088 ( .A1(n3172), .A2(\xmem_data[34][2] ), .B1(n28468), .B2(
        \xmem_data[35][2] ), .ZN(n23291) );
  AOI22_X1 U27089 ( .A1(n25684), .A2(\xmem_data[36][2] ), .B1(n24624), .B2(
        \xmem_data[37][2] ), .ZN(n23290) );
  AOI22_X1 U27090 ( .A1(n30909), .A2(\xmem_data[38][2] ), .B1(n3203), .B2(
        \xmem_data[39][2] ), .ZN(n23289) );
  NAND4_X1 U27091 ( .A1(n23292), .A2(n23291), .A3(n23290), .A4(n23289), .ZN(
        n23308) );
  AOI22_X1 U27092 ( .A1(n24630), .A2(\xmem_data[40][2] ), .B1(n3247), .B2(
        \xmem_data[41][2] ), .ZN(n23296) );
  AOI22_X1 U27093 ( .A1(n24631), .A2(\xmem_data[42][2] ), .B1(n3217), .B2(
        \xmem_data[43][2] ), .ZN(n23295) );
  AOI22_X1 U27094 ( .A1(n24632), .A2(\xmem_data[44][2] ), .B1(n24207), .B2(
        \xmem_data[45][2] ), .ZN(n23294) );
  AOI22_X1 U27095 ( .A1(n3341), .A2(\xmem_data[46][2] ), .B1(n24633), .B2(
        \xmem_data[47][2] ), .ZN(n23293) );
  NAND4_X1 U27096 ( .A1(n23296), .A2(n23295), .A3(n23294), .A4(n23293), .ZN(
        n23307) );
  AOI22_X1 U27097 ( .A1(n3281), .A2(\xmem_data[48][2] ), .B1(n25492), .B2(
        \xmem_data[49][2] ), .ZN(n23300) );
  AOI22_X1 U27098 ( .A1(n24638), .A2(\xmem_data[50][2] ), .B1(n28373), .B2(
        \xmem_data[51][2] ), .ZN(n23299) );
  AOI22_X1 U27099 ( .A1(n24640), .A2(\xmem_data[52][2] ), .B1(n24639), .B2(
        \xmem_data[53][2] ), .ZN(n23298) );
  AOI22_X1 U27100 ( .A1(n16986), .A2(\xmem_data[54][2] ), .B1(n29009), .B2(
        \xmem_data[55][2] ), .ZN(n23297) );
  NAND4_X1 U27101 ( .A1(n23300), .A2(n23299), .A3(n23298), .A4(n23297), .ZN(
        n23306) );
  AOI22_X1 U27102 ( .A1(n28516), .A2(\xmem_data[56][2] ), .B1(n27454), .B2(
        \xmem_data[57][2] ), .ZN(n23304) );
  AOI22_X1 U27103 ( .A1(n29317), .A2(\xmem_data[58][2] ), .B1(n24645), .B2(
        \xmem_data[59][2] ), .ZN(n23303) );
  AOI22_X1 U27104 ( .A1(n29012), .A2(\xmem_data[60][2] ), .B1(n24646), .B2(
        \xmem_data[61][2] ), .ZN(n23302) );
  AOI22_X1 U27105 ( .A1(n24647), .A2(\xmem_data[62][2] ), .B1(n25581), .B2(
        \xmem_data[63][2] ), .ZN(n23301) );
  NAND4_X1 U27106 ( .A1(n23304), .A2(n23303), .A3(n23302), .A4(n23301), .ZN(
        n23305) );
  OR4_X1 U27107 ( .A1(n23308), .A2(n23307), .A3(n23306), .A4(n23305), .ZN(
        n23337) );
  AOI22_X1 U27108 ( .A1(n28152), .A2(\xmem_data[20][2] ), .B1(n13168), .B2(
        \xmem_data[21][2] ), .ZN(n23315) );
  AOI22_X1 U27109 ( .A1(n27515), .A2(\xmem_data[22][2] ), .B1(n24597), .B2(
        \xmem_data[23][2] ), .ZN(n23309) );
  INV_X1 U27110 ( .A(n23309), .ZN(n23313) );
  AOI22_X1 U27111 ( .A1(n27551), .A2(\xmem_data[18][2] ), .B1(n24590), .B2(
        \xmem_data[19][2] ), .ZN(n23311) );
  NAND2_X1 U27112 ( .A1(n25377), .A2(\xmem_data[16][2] ), .ZN(n23310) );
  NAND2_X1 U27113 ( .A1(n23311), .A2(n23310), .ZN(n23312) );
  NOR2_X1 U27114 ( .A1(n23313), .A2(n23312), .ZN(n23314) );
  NAND2_X1 U27115 ( .A1(n23315), .A2(n23314), .ZN(n23326) );
  AOI22_X1 U27116 ( .A1(n30746), .A2(\xmem_data[24][2] ), .B1(n27989), .B2(
        \xmem_data[25][2] ), .ZN(n23319) );
  AOI22_X1 U27117 ( .A1(n24593), .A2(\xmem_data[26][2] ), .B1(n28492), .B2(
        \xmem_data[27][2] ), .ZN(n23318) );
  AOI22_X1 U27118 ( .A1(n27825), .A2(\xmem_data[28][2] ), .B1(n24592), .B2(
        \xmem_data[29][2] ), .ZN(n23317) );
  AOI22_X1 U27119 ( .A1(n29100), .A2(\xmem_data[30][2] ), .B1(n28429), .B2(
        \xmem_data[31][2] ), .ZN(n23316) );
  NAND4_X1 U27120 ( .A1(n23319), .A2(n23318), .A3(n23317), .A4(n23316), .ZN(
        n23325) );
  AOI22_X1 U27121 ( .A1(n3317), .A2(\xmem_data[8][2] ), .B1(n3247), .B2(
        \xmem_data[9][2] ), .ZN(n23323) );
  AOI22_X1 U27122 ( .A1(n20576), .A2(\xmem_data[10][2] ), .B1(n3219), .B2(
        \xmem_data[11][2] ), .ZN(n23322) );
  AOI22_X1 U27123 ( .A1(n20724), .A2(\xmem_data[12][2] ), .B1(n25491), .B2(
        \xmem_data[13][2] ), .ZN(n23321) );
  AOI22_X1 U27124 ( .A1(n28475), .A2(\xmem_data[14][2] ), .B1(n20993), .B2(
        \xmem_data[15][2] ), .ZN(n23320) );
  NAND4_X1 U27125 ( .A1(n23323), .A2(n23322), .A3(n23321), .A4(n23320), .ZN(
        n23324) );
  OR3_X1 U27126 ( .A1(n23326), .A2(n23325), .A3(n23324), .ZN(n23332) );
  AOI22_X1 U27127 ( .A1(n3151), .A2(\xmem_data[0][2] ), .B1(n27975), .B2(
        \xmem_data[1][2] ), .ZN(n23330) );
  AOI22_X1 U27128 ( .A1(n24606), .A2(\xmem_data[2][2] ), .B1(n20488), .B2(
        \xmem_data[3][2] ), .ZN(n23329) );
  AOI22_X1 U27129 ( .A1(n27852), .A2(\xmem_data[4][2] ), .B1(n20707), .B2(
        \xmem_data[5][2] ), .ZN(n23328) );
  AOI22_X1 U27130 ( .A1(n24607), .A2(\xmem_data[6][2] ), .B1(n28317), .B2(
        \xmem_data[7][2] ), .ZN(n23327) );
  NAND4_X1 U27131 ( .A1(n23330), .A2(n23329), .A3(n23328), .A4(n23327), .ZN(
        n23331) );
  NOR2_X1 U27132 ( .A1(n23332), .A2(n23331), .ZN(n23333) );
  NOR2_X1 U27133 ( .A1(n23333), .A2(n24662), .ZN(n23336) );
  NOR2_X1 U27134 ( .A1(n24662), .A2(n39007), .ZN(n23334) );
  AND2_X1 U27135 ( .A1(n31252), .A2(n23334), .ZN(n23335) );
  AOI211_X1 U27136 ( .C1(n23337), .C2(n24659), .A(n23336), .B(n23335), .ZN(
        n23381) );
  AOI22_X1 U27137 ( .A1(n24522), .A2(\xmem_data[96][2] ), .B1(n20553), .B2(
        \xmem_data[97][2] ), .ZN(n23341) );
  AOI22_X1 U27138 ( .A1(n24685), .A2(\xmem_data[98][2] ), .B1(n23781), .B2(
        \xmem_data[99][2] ), .ZN(n23340) );
  AOI22_X1 U27139 ( .A1(n24687), .A2(\xmem_data[100][2] ), .B1(n24686), .B2(
        \xmem_data[101][2] ), .ZN(n23339) );
  AOI22_X1 U27140 ( .A1(n24688), .A2(\xmem_data[102][2] ), .B1(n28366), .B2(
        \xmem_data[103][2] ), .ZN(n23338) );
  NAND4_X1 U27141 ( .A1(n23341), .A2(n23340), .A3(n23339), .A4(n23338), .ZN(
        n23357) );
  AOI22_X1 U27142 ( .A1(n24693), .A2(\xmem_data[104][2] ), .B1(n25360), .B2(
        \xmem_data[105][2] ), .ZN(n23345) );
  AOI22_X1 U27143 ( .A1(n24694), .A2(\xmem_data[106][2] ), .B1(n3218), .B2(
        \xmem_data[107][2] ), .ZN(n23344) );
  AOI22_X1 U27144 ( .A1(n24696), .A2(\xmem_data[108][2] ), .B1(n24695), .B2(
        \xmem_data[109][2] ), .ZN(n23343) );
  AOI22_X1 U27145 ( .A1(n24697), .A2(\xmem_data[110][2] ), .B1(n27550), .B2(
        \xmem_data[111][2] ), .ZN(n23342) );
  NAND4_X1 U27146 ( .A1(n23345), .A2(n23344), .A3(n23343), .A4(n23342), .ZN(
        n23356) );
  AOI22_X1 U27147 ( .A1(n24702), .A2(\xmem_data[112][2] ), .B1(n28510), .B2(
        \xmem_data[113][2] ), .ZN(n23349) );
  AOI22_X1 U27148 ( .A1(n23813), .A2(\xmem_data[114][2] ), .B1(n27988), .B2(
        \xmem_data[115][2] ), .ZN(n23348) );
  AOI22_X1 U27149 ( .A1(n28346), .A2(\xmem_data[116][2] ), .B1(n13168), .B2(
        \xmem_data[117][2] ), .ZN(n23347) );
  AOI22_X1 U27150 ( .A1(n10977), .A2(\xmem_data[118][2] ), .B1(n20584), .B2(
        \xmem_data[119][2] ), .ZN(n23346) );
  NAND4_X1 U27151 ( .A1(n23349), .A2(n23348), .A3(n23347), .A4(n23346), .ZN(
        n23355) );
  AOI22_X1 U27152 ( .A1(n29605), .A2(\xmem_data[120][2] ), .B1(n3207), .B2(
        \xmem_data[121][2] ), .ZN(n23353) );
  AOI22_X1 U27153 ( .A1(n24708), .A2(\xmem_data[122][2] ), .B1(n24707), .B2(
        \xmem_data[123][2] ), .ZN(n23352) );
  AOI22_X1 U27154 ( .A1(n24710), .A2(\xmem_data[124][2] ), .B1(n24709), .B2(
        \xmem_data[125][2] ), .ZN(n23351) );
  AOI22_X1 U27155 ( .A1(n27952), .A2(\xmem_data[126][2] ), .B1(n21009), .B2(
        \xmem_data[127][2] ), .ZN(n23350) );
  NAND4_X1 U27156 ( .A1(n23353), .A2(n23352), .A3(n23351), .A4(n23350), .ZN(
        n23354) );
  OR4_X1 U27157 ( .A1(n23357), .A2(n23356), .A3(n23355), .A4(n23354), .ZN(
        n23379) );
  AOI22_X1 U27158 ( .A1(n29324), .A2(\xmem_data[64][2] ), .B1(n14975), .B2(
        \xmem_data[65][2] ), .ZN(n23361) );
  AOI22_X1 U27159 ( .A1(n24685), .A2(\xmem_data[66][2] ), .B1(n30496), .B2(
        \xmem_data[67][2] ), .ZN(n23360) );
  AOI22_X1 U27160 ( .A1(n24687), .A2(\xmem_data[68][2] ), .B1(n24686), .B2(
        \xmem_data[69][2] ), .ZN(n23359) );
  AOI22_X1 U27161 ( .A1(n24688), .A2(\xmem_data[70][2] ), .B1(n28317), .B2(
        \xmem_data[71][2] ), .ZN(n23358) );
  NAND4_X1 U27162 ( .A1(n23361), .A2(n23360), .A3(n23359), .A4(n23358), .ZN(
        n23377) );
  AOI22_X1 U27163 ( .A1(n24693), .A2(\xmem_data[72][2] ), .B1(n25360), .B2(
        \xmem_data[73][2] ), .ZN(n23365) );
  AOI22_X1 U27164 ( .A1(n24694), .A2(\xmem_data[74][2] ), .B1(n3222), .B2(
        \xmem_data[75][2] ), .ZN(n23364) );
  AOI22_X1 U27165 ( .A1(n24696), .A2(\xmem_data[76][2] ), .B1(n24695), .B2(
        \xmem_data[77][2] ), .ZN(n23363) );
  AOI22_X1 U27166 ( .A1(n24697), .A2(\xmem_data[78][2] ), .B1(n31275), .B2(
        \xmem_data[79][2] ), .ZN(n23362) );
  NAND4_X1 U27167 ( .A1(n23365), .A2(n23364), .A3(n23363), .A4(n23362), .ZN(
        n23376) );
  AOI22_X1 U27168 ( .A1(n24702), .A2(\xmem_data[80][2] ), .B1(n28343), .B2(
        \xmem_data[81][2] ), .ZN(n23369) );
  AOI22_X1 U27169 ( .A1(n27447), .A2(\xmem_data[82][2] ), .B1(n20588), .B2(
        \xmem_data[83][2] ), .ZN(n23368) );
  AOI22_X1 U27170 ( .A1(n31327), .A2(\xmem_data[84][2] ), .B1(n13168), .B2(
        \xmem_data[85][2] ), .ZN(n23367) );
  AOI22_X1 U27171 ( .A1(n29109), .A2(\xmem_data[86][2] ), .B1(n29309), .B2(
        \xmem_data[87][2] ), .ZN(n23366) );
  NAND4_X1 U27172 ( .A1(n23369), .A2(n23368), .A3(n23367), .A4(n23366), .ZN(
        n23375) );
  AOI22_X1 U27173 ( .A1(n30948), .A2(\xmem_data[88][2] ), .B1(n27864), .B2(
        \xmem_data[89][2] ), .ZN(n23373) );
  AOI22_X1 U27174 ( .A1(n24708), .A2(\xmem_data[90][2] ), .B1(n24707), .B2(
        \xmem_data[91][2] ), .ZN(n23372) );
  AOI22_X1 U27175 ( .A1(n24710), .A2(\xmem_data[92][2] ), .B1(n24709), .B2(
        \xmem_data[93][2] ), .ZN(n23371) );
  AOI22_X1 U27176 ( .A1(n29100), .A2(\xmem_data[94][2] ), .B1(n29055), .B2(
        \xmem_data[95][2] ), .ZN(n23370) );
  NAND4_X1 U27177 ( .A1(n23373), .A2(n23372), .A3(n23371), .A4(n23370), .ZN(
        n23374) );
  OR4_X1 U27178 ( .A1(n23377), .A2(n23376), .A3(n23375), .A4(n23374), .ZN(
        n23378) );
  AOI22_X1 U27179 ( .A1(n24722), .A2(n23379), .B1(n24720), .B2(n23378), .ZN(
        n23380) );
  NAND2_X1 U27180 ( .A1(n23381), .A2(n23380), .ZN(n33803) );
  XNOR2_X1 U27181 ( .A(n33803), .B(\fmem_data[24][5] ), .ZN(n27582) );
  OAI22_X1 U27182 ( .A1(n31167), .A2(n34041), .B1(n27582), .B2(n34039), .ZN(
        n28903) );
  AOI22_X1 U27183 ( .A1(n21007), .A2(\xmem_data[96][1] ), .B1(n25398), .B2(
        \xmem_data[97][1] ), .ZN(n23385) );
  AOI22_X1 U27184 ( .A1(n25400), .A2(\xmem_data[98][1] ), .B1(n25399), .B2(
        \xmem_data[99][1] ), .ZN(n23384) );
  AOI22_X1 U27185 ( .A1(n3178), .A2(\xmem_data[100][1] ), .B1(n28462), .B2(
        \xmem_data[101][1] ), .ZN(n23383) );
  AOI22_X1 U27186 ( .A1(n25401), .A2(\xmem_data[102][1] ), .B1(n14975), .B2(
        \xmem_data[103][1] ), .ZN(n23382) );
  NAND4_X1 U27187 ( .A1(n23385), .A2(n23384), .A3(n23383), .A4(n23382), .ZN(
        n23401) );
  AOI22_X1 U27188 ( .A1(n20782), .A2(\xmem_data[104][1] ), .B1(n25406), .B2(
        \xmem_data[105][1] ), .ZN(n23389) );
  AOI22_X1 U27189 ( .A1(n25407), .A2(\xmem_data[106][1] ), .B1(n31261), .B2(
        \xmem_data[107][1] ), .ZN(n23388) );
  AOI22_X1 U27190 ( .A1(n25408), .A2(\xmem_data[108][1] ), .B1(n12471), .B2(
        \xmem_data[109][1] ), .ZN(n23387) );
  AOI22_X1 U27191 ( .A1(n3318), .A2(\xmem_data[110][1] ), .B1(n30863), .B2(
        \xmem_data[111][1] ), .ZN(n23386) );
  NAND4_X1 U27192 ( .A1(n23389), .A2(n23388), .A3(n23387), .A4(n23386), .ZN(
        n23400) );
  AOI22_X1 U27193 ( .A1(n25413), .A2(\xmem_data[112][1] ), .B1(n3219), .B2(
        \xmem_data[113][1] ), .ZN(n23393) );
  AOI22_X1 U27194 ( .A1(n25414), .A2(\xmem_data[114][1] ), .B1(n25491), .B2(
        \xmem_data[115][1] ), .ZN(n23392) );
  AOI22_X1 U27195 ( .A1(n25416), .A2(\xmem_data[116][1] ), .B1(n25415), .B2(
        \xmem_data[117][1] ), .ZN(n23391) );
  AOI22_X1 U27196 ( .A1(n25417), .A2(\xmem_data[118][1] ), .B1(n25450), .B2(
        \xmem_data[119][1] ), .ZN(n23390) );
  NAND4_X1 U27197 ( .A1(n23393), .A2(n23392), .A3(n23391), .A4(n23390), .ZN(
        n23399) );
  AOI22_X1 U27198 ( .A1(n25422), .A2(\xmem_data[120][1] ), .B1(n24158), .B2(
        \xmem_data[121][1] ), .ZN(n23397) );
  AOI22_X1 U27199 ( .A1(n25424), .A2(\xmem_data[122][1] ), .B1(n25423), .B2(
        \xmem_data[123][1] ), .ZN(n23396) );
  AOI22_X1 U27200 ( .A1(n25425), .A2(\xmem_data[124][1] ), .B1(n22674), .B2(
        \xmem_data[125][1] ), .ZN(n23395) );
  AOI22_X1 U27201 ( .A1(n30892), .A2(\xmem_data[126][1] ), .B1(n30615), .B2(
        \xmem_data[127][1] ), .ZN(n23394) );
  NAND4_X1 U27202 ( .A1(n23397), .A2(n23396), .A3(n23395), .A4(n23394), .ZN(
        n23398) );
  OR4_X1 U27203 ( .A1(n23401), .A2(n23400), .A3(n23399), .A4(n23398), .ZN(
        n23423) );
  AOI22_X1 U27204 ( .A1(n23717), .A2(\xmem_data[64][1] ), .B1(n25398), .B2(
        \xmem_data[65][1] ), .ZN(n23405) );
  AOI22_X1 U27205 ( .A1(n25400), .A2(\xmem_data[66][1] ), .B1(n25399), .B2(
        \xmem_data[67][1] ), .ZN(n23404) );
  AOI22_X1 U27206 ( .A1(n27974), .A2(\xmem_data[68][1] ), .B1(n28060), .B2(
        \xmem_data[69][1] ), .ZN(n23403) );
  AOI22_X1 U27207 ( .A1(n25401), .A2(\xmem_data[70][1] ), .B1(n14975), .B2(
        \xmem_data[71][1] ), .ZN(n23402) );
  NAND4_X1 U27208 ( .A1(n23405), .A2(n23404), .A3(n23403), .A4(n23402), .ZN(
        n23421) );
  AOI22_X1 U27209 ( .A1(n29325), .A2(\xmem_data[72][1] ), .B1(n25406), .B2(
        \xmem_data[73][1] ), .ZN(n23409) );
  AOI22_X1 U27210 ( .A1(n25407), .A2(\xmem_data[74][1] ), .B1(n24524), .B2(
        \xmem_data[75][1] ), .ZN(n23408) );
  AOI22_X1 U27211 ( .A1(n25408), .A2(\xmem_data[76][1] ), .B1(n20709), .B2(
        \xmem_data[77][1] ), .ZN(n23407) );
  AOI22_X1 U27212 ( .A1(n3318), .A2(\xmem_data[78][1] ), .B1(n27501), .B2(
        \xmem_data[79][1] ), .ZN(n23406) );
  NAND4_X1 U27213 ( .A1(n23409), .A2(n23408), .A3(n23407), .A4(n23406), .ZN(
        n23420) );
  AOI22_X1 U27214 ( .A1(n25413), .A2(\xmem_data[80][1] ), .B1(n3220), .B2(
        \xmem_data[81][1] ), .ZN(n23413) );
  AOI22_X1 U27215 ( .A1(n25414), .A2(\xmem_data[82][1] ), .B1(n20787), .B2(
        \xmem_data[83][1] ), .ZN(n23412) );
  AOI22_X1 U27216 ( .A1(n25416), .A2(\xmem_data[84][1] ), .B1(n25415), .B2(
        \xmem_data[85][1] ), .ZN(n23411) );
  AOI22_X1 U27217 ( .A1(n25417), .A2(\xmem_data[86][1] ), .B1(n25492), .B2(
        \xmem_data[87][1] ), .ZN(n23410) );
  NAND4_X1 U27218 ( .A1(n23413), .A2(n23412), .A3(n23411), .A4(n23410), .ZN(
        n23419) );
  AOI22_X1 U27219 ( .A1(n25422), .A2(\xmem_data[88][1] ), .B1(n20588), .B2(
        \xmem_data[89][1] ), .ZN(n23417) );
  AOI22_X1 U27220 ( .A1(n25424), .A2(\xmem_data[90][1] ), .B1(n25423), .B2(
        \xmem_data[91][1] ), .ZN(n23416) );
  AOI22_X1 U27221 ( .A1(n25425), .A2(\xmem_data[92][1] ), .B1(n24160), .B2(
        \xmem_data[93][1] ), .ZN(n23415) );
  AOI22_X1 U27222 ( .A1(n29437), .A2(\xmem_data[94][1] ), .B1(n22742), .B2(
        \xmem_data[95][1] ), .ZN(n23414) );
  NAND4_X1 U27223 ( .A1(n23417), .A2(n23416), .A3(n23415), .A4(n23414), .ZN(
        n23418) );
  OR4_X1 U27224 ( .A1(n23421), .A2(n23420), .A3(n23419), .A4(n23418), .ZN(
        n23422) );
  AOI22_X1 U27225 ( .A1(n25473), .A2(n23423), .B1(n25471), .B2(n23422), .ZN(
        n23477) );
  AOI22_X1 U27226 ( .A1(n27919), .A2(\xmem_data[0][1] ), .B1(n25520), .B2(
        \xmem_data[1][1] ), .ZN(n23427) );
  AOI22_X1 U27227 ( .A1(n30872), .A2(\xmem_data[2][1] ), .B1(n25367), .B2(
        \xmem_data[3][1] ), .ZN(n23426) );
  AOI22_X1 U27228 ( .A1(n20593), .A2(\xmem_data[4][1] ), .B1(n25364), .B2(
        \xmem_data[5][1] ), .ZN(n23425) );
  AOI22_X1 U27229 ( .A1(n20984), .A2(\xmem_data[6][1] ), .B1(n22685), .B2(
        \xmem_data[7][1] ), .ZN(n23424) );
  NAND4_X1 U27230 ( .A1(n23427), .A2(n23426), .A3(n23425), .A4(n23424), .ZN(
        n23433) );
  AOI22_X1 U27231 ( .A1(n28293), .A2(\xmem_data[8][1] ), .B1(n25359), .B2(
        \xmem_data[9][1] ), .ZN(n23431) );
  AOI22_X1 U27232 ( .A1(n30257), .A2(\xmem_data[10][1] ), .B1(n25388), .B2(
        \xmem_data[11][1] ), .ZN(n23430) );
  AOI22_X1 U27233 ( .A1(n25358), .A2(\xmem_data[12][1] ), .B1(n25357), .B2(
        \xmem_data[13][1] ), .ZN(n23429) );
  AOI22_X1 U27234 ( .A1(n21308), .A2(\xmem_data[14][1] ), .B1(n25360), .B2(
        \xmem_data[15][1] ), .ZN(n23428) );
  NAND4_X1 U27235 ( .A1(n23431), .A2(n23430), .A3(n23429), .A4(n23428), .ZN(
        n23432) );
  OR2_X1 U27236 ( .A1(n23433), .A2(n23432), .ZN(n23450) );
  NAND2_X1 U27237 ( .A1(n25354), .A2(\xmem_data[16][1] ), .ZN(n23435) );
  NAND2_X1 U27238 ( .A1(n3221), .A2(\xmem_data[17][1] ), .ZN(n23434) );
  NAND2_X1 U27239 ( .A1(n23435), .A2(n23434), .ZN(n23439) );
  AOI22_X1 U27240 ( .A1(n3342), .A2(\xmem_data[20][1] ), .B1(n28372), .B2(
        \xmem_data[21][1] ), .ZN(n23437) );
  NAND2_X1 U27241 ( .A1(n25377), .A2(\xmem_data[22][1] ), .ZN(n23436) );
  NAND2_X1 U27242 ( .A1(n23437), .A2(n23436), .ZN(n23438) );
  NOR2_X1 U27243 ( .A1(n23439), .A2(n23438), .ZN(n23448) );
  AOI22_X1 U27244 ( .A1(n28374), .A2(\xmem_data[24][1] ), .B1(n20982), .B2(
        \xmem_data[25][1] ), .ZN(n23443) );
  AOI22_X1 U27245 ( .A1(n17013), .A2(\xmem_data[26][1] ), .B1(n24159), .B2(
        \xmem_data[27][1] ), .ZN(n23442) );
  AOI22_X1 U27246 ( .A1(n31268), .A2(\xmem_data[28][1] ), .B1(n25382), .B2(
        \xmem_data[29][1] ), .ZN(n23441) );
  AOI22_X1 U27247 ( .A1(n17018), .A2(\xmem_data[30][1] ), .B1(n25383), .B2(
        \xmem_data[31][1] ), .ZN(n23440) );
  NAND4_X1 U27248 ( .A1(n23443), .A2(n23442), .A3(n23441), .A4(n23440), .ZN(
        n23446) );
  AOI22_X1 U27249 ( .A1(n29422), .A2(\xmem_data[18][1] ), .B1(n23769), .B2(
        \xmem_data[19][1] ), .ZN(n23444) );
  NAND2_X1 U27250 ( .A1(n23448), .A2(n23447), .ZN(n23449) );
  NOR2_X1 U27251 ( .A1(n23450), .A2(n23449), .ZN(n23452) );
  NAND2_X1 U27252 ( .A1(n30877), .A2(\xmem_data[23][1] ), .ZN(n23451) );
  AOI21_X1 U27253 ( .B1(n23452), .B2(n23451), .A(n25392), .ZN(n23475) );
  AOI22_X1 U27254 ( .A1(n25434), .A2(\xmem_data[32][1] ), .B1(n28427), .B2(
        \xmem_data[33][1] ), .ZN(n23456) );
  AOI22_X1 U27255 ( .A1(n29047), .A2(\xmem_data[34][1] ), .B1(n25435), .B2(
        \xmem_data[35][1] ), .ZN(n23455) );
  AOI22_X1 U27256 ( .A1(n3178), .A2(\xmem_data[36][1] ), .B1(n30495), .B2(
        \xmem_data[37][1] ), .ZN(n23454) );
  AOI22_X1 U27257 ( .A1(n3308), .A2(\xmem_data[38][1] ), .B1(n28098), .B2(
        \xmem_data[39][1] ), .ZN(n23453) );
  NAND4_X1 U27258 ( .A1(n23456), .A2(n23455), .A3(n23454), .A4(n23453), .ZN(
        n23472) );
  AOI22_X1 U27259 ( .A1(n13486), .A2(\xmem_data[40][1] ), .B1(n20488), .B2(
        \xmem_data[41][1] ), .ZN(n23460) );
  AOI22_X1 U27260 ( .A1(n30754), .A2(\xmem_data[42][1] ), .B1(n25440), .B2(
        \xmem_data[43][1] ), .ZN(n23459) );
  AOI22_X1 U27261 ( .A1(n25441), .A2(\xmem_data[44][1] ), .B1(n31309), .B2(
        \xmem_data[45][1] ), .ZN(n23458) );
  AOI22_X1 U27262 ( .A1(n25443), .A2(\xmem_data[46][1] ), .B1(n25442), .B2(
        \xmem_data[47][1] ), .ZN(n23457) );
  NAND4_X1 U27263 ( .A1(n23460), .A2(n23459), .A3(n23458), .A4(n23457), .ZN(
        n23471) );
  AOI22_X1 U27264 ( .A1(n30503), .A2(\xmem_data[48][1] ), .B1(n3218), .B2(
        \xmem_data[49][1] ), .ZN(n23464) );
  AOI22_X1 U27265 ( .A1(n25448), .A2(\xmem_data[50][1] ), .B1(n29095), .B2(
        \xmem_data[51][1] ), .ZN(n23463) );
  AOI22_X1 U27266 ( .A1(n25449), .A2(\xmem_data[52][1] ), .B1(n21068), .B2(
        \xmem_data[53][1] ), .ZN(n23462) );
  AOI22_X1 U27267 ( .A1(n25451), .A2(\xmem_data[54][1] ), .B1(n25450), .B2(
        \xmem_data[55][1] ), .ZN(n23461) );
  NAND4_X1 U27268 ( .A1(n23464), .A2(n23463), .A3(n23462), .A4(n23461), .ZN(
        n23470) );
  AOI22_X1 U27269 ( .A1(n27447), .A2(\xmem_data[56][1] ), .B1(n30854), .B2(
        \xmem_data[57][1] ), .ZN(n23468) );
  AOI22_X1 U27270 ( .A1(n25457), .A2(\xmem_data[58][1] ), .B1(n27535), .B2(
        \xmem_data[59][1] ), .ZN(n23467) );
  AOI22_X1 U27271 ( .A1(n25459), .A2(\xmem_data[60][1] ), .B1(n25458), .B2(
        \xmem_data[61][1] ), .ZN(n23466) );
  AOI22_X1 U27272 ( .A1(n25461), .A2(\xmem_data[62][1] ), .B1(n25460), .B2(
        \xmem_data[63][1] ), .ZN(n23465) );
  NAND4_X1 U27273 ( .A1(n23468), .A2(n23467), .A3(n23466), .A4(n23465), .ZN(
        n23469) );
  OR4_X1 U27274 ( .A1(n23472), .A2(n23471), .A3(n23470), .A4(n23469), .ZN(
        n23473) );
  AND2_X1 U27275 ( .A1(n23473), .A2(n25396), .ZN(n23474) );
  NOR2_X1 U27276 ( .A1(n23475), .A2(n23474), .ZN(n23476) );
  XNOR2_X1 U27277 ( .A(n33677), .B(\fmem_data[30][5] ), .ZN(n31169) );
  AOI22_X1 U27278 ( .A1(n25434), .A2(\xmem_data[32][2] ), .B1(n28492), .B2(
        \xmem_data[33][2] ), .ZN(n23481) );
  AOI22_X1 U27279 ( .A1(n14971), .A2(\xmem_data[34][2] ), .B1(n25435), .B2(
        \xmem_data[35][2] ), .ZN(n23480) );
  AOI22_X1 U27280 ( .A1(n27462), .A2(\xmem_data[36][2] ), .B1(n20943), .B2(
        \xmem_data[37][2] ), .ZN(n23479) );
  AOI22_X1 U27281 ( .A1(n3308), .A2(\xmem_data[38][2] ), .B1(n28062), .B2(
        \xmem_data[39][2] ), .ZN(n23478) );
  NAND4_X1 U27282 ( .A1(n23481), .A2(n23480), .A3(n23479), .A4(n23478), .ZN(
        n23497) );
  AOI22_X1 U27283 ( .A1(n24572), .A2(\xmem_data[40][2] ), .B1(n20488), .B2(
        \xmem_data[41][2] ), .ZN(n23485) );
  AOI22_X1 U27284 ( .A1(n20577), .A2(\xmem_data[42][2] ), .B1(n25440), .B2(
        \xmem_data[43][2] ), .ZN(n23484) );
  AOI22_X1 U27285 ( .A1(n25441), .A2(\xmem_data[44][2] ), .B1(n25629), .B2(
        \xmem_data[45][2] ), .ZN(n23483) );
  AOI22_X1 U27286 ( .A1(n25443), .A2(\xmem_data[46][2] ), .B1(n25442), .B2(
        \xmem_data[47][2] ), .ZN(n23482) );
  NAND4_X1 U27287 ( .A1(n23485), .A2(n23484), .A3(n23483), .A4(n23482), .ZN(
        n23496) );
  AOI22_X1 U27288 ( .A1(n25692), .A2(\xmem_data[48][2] ), .B1(n3217), .B2(
        \xmem_data[49][2] ), .ZN(n23489) );
  AOI22_X1 U27289 ( .A1(n25448), .A2(\xmem_data[50][2] ), .B1(n27444), .B2(
        \xmem_data[51][2] ), .ZN(n23488) );
  AOI22_X1 U27290 ( .A1(n25449), .A2(\xmem_data[52][2] ), .B1(n25616), .B2(
        \xmem_data[53][2] ), .ZN(n23487) );
  AOI22_X1 U27291 ( .A1(n25451), .A2(\xmem_data[54][2] ), .B1(n28307), .B2(
        \xmem_data[55][2] ), .ZN(n23486) );
  NAND4_X1 U27292 ( .A1(n23489), .A2(n23488), .A3(n23487), .A4(n23486), .ZN(
        n23495) );
  AOI22_X1 U27293 ( .A1(n22712), .A2(\xmem_data[56][2] ), .B1(n3357), .B2(
        \xmem_data[57][2] ), .ZN(n23493) );
  AOI22_X1 U27294 ( .A1(n25457), .A2(\xmem_data[58][2] ), .B1(n21075), .B2(
        \xmem_data[59][2] ), .ZN(n23492) );
  AOI22_X1 U27295 ( .A1(n25459), .A2(\xmem_data[60][2] ), .B1(n25458), .B2(
        \xmem_data[61][2] ), .ZN(n23491) );
  AOI22_X1 U27296 ( .A1(n29396), .A2(\xmem_data[62][2] ), .B1(n25460), .B2(
        \xmem_data[63][2] ), .ZN(n23490) );
  NAND4_X1 U27297 ( .A1(n23493), .A2(n23492), .A3(n23491), .A4(n23490), .ZN(
        n23494) );
  OR4_X1 U27298 ( .A1(n23497), .A2(n23496), .A3(n23495), .A4(n23494), .ZN(
        n23528) );
  AOI22_X1 U27299 ( .A1(n28096), .A2(\xmem_data[0][2] ), .B1(n28058), .B2(
        \xmem_data[1][2] ), .ZN(n23501) );
  AOI22_X1 U27300 ( .A1(n27825), .A2(\xmem_data[2][2] ), .B1(n25367), .B2(
        \xmem_data[3][2] ), .ZN(n23500) );
  AOI22_X1 U27301 ( .A1(n3325), .A2(\xmem_data[4][2] ), .B1(n25364), .B2(
        \xmem_data[5][2] ), .ZN(n23499) );
  AOI22_X1 U27302 ( .A1(n17004), .A2(\xmem_data[6][2] ), .B1(n28098), .B2(
        \xmem_data[7][2] ), .ZN(n23498) );
  NAND4_X1 U27303 ( .A1(n23501), .A2(n23500), .A3(n23499), .A4(n23498), .ZN(
        n23507) );
  AOI22_X1 U27304 ( .A1(n31316), .A2(\xmem_data[8][2] ), .B1(n25359), .B2(
        \xmem_data[9][2] ), .ZN(n23505) );
  AOI22_X1 U27305 ( .A1(n27852), .A2(\xmem_data[10][2] ), .B1(n25388), .B2(
        \xmem_data[11][2] ), .ZN(n23504) );
  AOI22_X1 U27306 ( .A1(n25358), .A2(\xmem_data[12][2] ), .B1(n25357), .B2(
        \xmem_data[13][2] ), .ZN(n23503) );
  AOI22_X1 U27307 ( .A1(n3306), .A2(\xmem_data[14][2] ), .B1(n25360), .B2(
        \xmem_data[15][2] ), .ZN(n23502) );
  NAND4_X1 U27308 ( .A1(n23505), .A2(n23504), .A3(n23503), .A4(n23502), .ZN(
        n23506) );
  OR2_X1 U27309 ( .A1(n23507), .A2(n23506), .ZN(n23524) );
  NAND2_X1 U27310 ( .A1(n25354), .A2(\xmem_data[16][2] ), .ZN(n23509) );
  NAND2_X1 U27311 ( .A1(n3221), .A2(\xmem_data[17][2] ), .ZN(n23508) );
  NAND2_X1 U27312 ( .A1(n23509), .A2(n23508), .ZN(n23513) );
  AOI22_X1 U27313 ( .A1(n30883), .A2(\xmem_data[20][2] ), .B1(n24140), .B2(
        \xmem_data[21][2] ), .ZN(n23511) );
  NAND2_X1 U27314 ( .A1(n25377), .A2(\xmem_data[22][2] ), .ZN(n23510) );
  NAND2_X1 U27315 ( .A1(n23511), .A2(n23510), .ZN(n23512) );
  NOR2_X1 U27316 ( .A1(n23513), .A2(n23512), .ZN(n23522) );
  AOI22_X1 U27317 ( .A1(n28374), .A2(\xmem_data[24][2] ), .B1(n13475), .B2(
        \xmem_data[25][2] ), .ZN(n23517) );
  AOI22_X1 U27318 ( .A1(n31353), .A2(\xmem_data[26][2] ), .B1(n23761), .B2(
        \xmem_data[27][2] ), .ZN(n23516) );
  AOI22_X1 U27319 ( .A1(n17041), .A2(\xmem_data[28][2] ), .B1(n25382), .B2(
        \xmem_data[29][2] ), .ZN(n23515) );
  AOI22_X1 U27320 ( .A1(n27455), .A2(\xmem_data[30][2] ), .B1(n25383), .B2(
        \xmem_data[31][2] ), .ZN(n23514) );
  NAND4_X1 U27321 ( .A1(n23517), .A2(n23516), .A3(n23515), .A4(n23514), .ZN(
        n23520) );
  AOI22_X1 U27322 ( .A1(n27831), .A2(\xmem_data[18][2] ), .B1(n20500), .B2(
        \xmem_data[19][2] ), .ZN(n23518) );
  NOR2_X1 U27323 ( .A1(n23524), .A2(n23523), .ZN(n23526) );
  NAND2_X1 U27324 ( .A1(n27547), .A2(\xmem_data[23][2] ), .ZN(n23525) );
  AOI21_X1 U27325 ( .B1(n23526), .B2(n23525), .A(n25392), .ZN(n23527) );
  AOI21_X1 U27326 ( .B1(n23528), .B2(n25396), .A(n23527), .ZN(n23572) );
  AOI22_X1 U27327 ( .A1(n25573), .A2(\xmem_data[96][2] ), .B1(n25398), .B2(
        \xmem_data[97][2] ), .ZN(n23532) );
  AOI22_X1 U27328 ( .A1(n25400), .A2(\xmem_data[98][2] ), .B1(n25399), .B2(
        \xmem_data[99][2] ), .ZN(n23531) );
  AOI22_X1 U27329 ( .A1(n29240), .A2(\xmem_data[100][2] ), .B1(n27461), .B2(
        \xmem_data[101][2] ), .ZN(n23530) );
  AOI22_X1 U27330 ( .A1(n25401), .A2(\xmem_data[102][2] ), .B1(n14975), .B2(
        \xmem_data[103][2] ), .ZN(n23529) );
  NAND4_X1 U27331 ( .A1(n23532), .A2(n23531), .A3(n23530), .A4(n23529), .ZN(
        n23548) );
  AOI22_X1 U27332 ( .A1(n14976), .A2(\xmem_data[104][2] ), .B1(n25406), .B2(
        \xmem_data[105][2] ), .ZN(n23536) );
  AOI22_X1 U27333 ( .A1(n25407), .A2(\xmem_data[106][2] ), .B1(n25440), .B2(
        \xmem_data[107][2] ), .ZN(n23535) );
  AOI22_X1 U27334 ( .A1(n25408), .A2(\xmem_data[108][2] ), .B1(n25357), .B2(
        \xmem_data[109][2] ), .ZN(n23534) );
  AOI22_X1 U27335 ( .A1(n3318), .A2(\xmem_data[110][2] ), .B1(n25360), .B2(
        \xmem_data[111][2] ), .ZN(n23533) );
  NAND4_X1 U27336 ( .A1(n23536), .A2(n23535), .A3(n23534), .A4(n23533), .ZN(
        n23547) );
  AOI22_X1 U27337 ( .A1(n25413), .A2(\xmem_data[112][2] ), .B1(n3218), .B2(
        \xmem_data[113][2] ), .ZN(n23540) );
  AOI22_X1 U27338 ( .A1(n25414), .A2(\xmem_data[114][2] ), .B1(n20723), .B2(
        \xmem_data[115][2] ), .ZN(n23539) );
  AOI22_X1 U27339 ( .A1(n25416), .A2(\xmem_data[116][2] ), .B1(n25415), .B2(
        \xmem_data[117][2] ), .ZN(n23538) );
  AOI22_X1 U27340 ( .A1(n25417), .A2(\xmem_data[118][2] ), .B1(n25450), .B2(
        \xmem_data[119][2] ), .ZN(n23537) );
  NAND4_X1 U27341 ( .A1(n23540), .A2(n23539), .A3(n23538), .A4(n23537), .ZN(
        n23546) );
  AOI22_X1 U27342 ( .A1(n25422), .A2(\xmem_data[120][2] ), .B1(n22739), .B2(
        \xmem_data[121][2] ), .ZN(n23544) );
  AOI22_X1 U27343 ( .A1(n25424), .A2(\xmem_data[122][2] ), .B1(n25423), .B2(
        \xmem_data[123][2] ), .ZN(n23543) );
  AOI22_X1 U27344 ( .A1(n25425), .A2(\xmem_data[124][2] ), .B1(n20584), .B2(
        \xmem_data[125][2] ), .ZN(n23542) );
  AOI22_X1 U27345 ( .A1(n20939), .A2(\xmem_data[126][2] ), .B1(n27516), .B2(
        \xmem_data[127][2] ), .ZN(n23541) );
  NAND4_X1 U27346 ( .A1(n23544), .A2(n23543), .A3(n23542), .A4(n23541), .ZN(
        n23545) );
  OR4_X1 U27347 ( .A1(n23548), .A2(n23547), .A3(n23546), .A4(n23545), .ZN(
        n23570) );
  AOI22_X1 U27348 ( .A1(n23717), .A2(\xmem_data[64][2] ), .B1(n25398), .B2(
        \xmem_data[65][2] ), .ZN(n23552) );
  AOI22_X1 U27349 ( .A1(n25400), .A2(\xmem_data[66][2] ), .B1(n25399), .B2(
        \xmem_data[67][2] ), .ZN(n23551) );
  AOI22_X1 U27350 ( .A1(n25521), .A2(\xmem_data[68][2] ), .B1(n30598), .B2(
        \xmem_data[69][2] ), .ZN(n23550) );
  AOI22_X1 U27351 ( .A1(n25401), .A2(\xmem_data[70][2] ), .B1(n14975), .B2(
        \xmem_data[71][2] ), .ZN(n23549) );
  NAND4_X1 U27352 ( .A1(n23552), .A2(n23551), .A3(n23550), .A4(n23549), .ZN(
        n23568) );
  AOI22_X1 U27353 ( .A1(n3179), .A2(\xmem_data[72][2] ), .B1(n25406), .B2(
        \xmem_data[73][2] ), .ZN(n23556) );
  AOI22_X1 U27354 ( .A1(n25407), .A2(\xmem_data[74][2] ), .B1(n31261), .B2(
        \xmem_data[75][2] ), .ZN(n23555) );
  AOI22_X1 U27355 ( .A1(n25408), .A2(\xmem_data[76][2] ), .B1(n3203), .B2(
        \xmem_data[77][2] ), .ZN(n23554) );
  AOI22_X1 U27356 ( .A1(n3318), .A2(\xmem_data[78][2] ), .B1(n23731), .B2(
        \xmem_data[79][2] ), .ZN(n23553) );
  NAND4_X1 U27357 ( .A1(n23556), .A2(n23555), .A3(n23554), .A4(n23553), .ZN(
        n23567) );
  AOI22_X1 U27358 ( .A1(n25413), .A2(\xmem_data[80][2] ), .B1(n3219), .B2(
        \xmem_data[81][2] ), .ZN(n23560) );
  AOI22_X1 U27359 ( .A1(n25414), .A2(\xmem_data[82][2] ), .B1(n20723), .B2(
        \xmem_data[83][2] ), .ZN(n23559) );
  AOI22_X1 U27360 ( .A1(n25416), .A2(\xmem_data[84][2] ), .B1(n25415), .B2(
        \xmem_data[85][2] ), .ZN(n23558) );
  AOI22_X1 U27361 ( .A1(n25417), .A2(\xmem_data[86][2] ), .B1(n29103), .B2(
        \xmem_data[87][2] ), .ZN(n23557) );
  NAND4_X1 U27362 ( .A1(n23560), .A2(n23559), .A3(n23558), .A4(n23557), .ZN(
        n23566) );
  AOI22_X1 U27363 ( .A1(n25422), .A2(\xmem_data[88][2] ), .B1(n24130), .B2(
        \xmem_data[89][2] ), .ZN(n23564) );
  AOI22_X1 U27364 ( .A1(n25424), .A2(\xmem_data[90][2] ), .B1(n25423), .B2(
        \xmem_data[91][2] ), .ZN(n23563) );
  AOI22_X1 U27365 ( .A1(n25425), .A2(\xmem_data[92][2] ), .B1(n30613), .B2(
        \xmem_data[93][2] ), .ZN(n23562) );
  AOI22_X1 U27366 ( .A1(n20718), .A2(\xmem_data[94][2] ), .B1(n25460), .B2(
        \xmem_data[95][2] ), .ZN(n23561) );
  NAND4_X1 U27367 ( .A1(n23564), .A2(n23563), .A3(n23562), .A4(n23561), .ZN(
        n23565) );
  OR4_X1 U27368 ( .A1(n23568), .A2(n23567), .A3(n23566), .A4(n23565), .ZN(
        n23569) );
  AOI22_X1 U27369 ( .A1(n25473), .A2(n23570), .B1(n25471), .B2(n23569), .ZN(
        n23571) );
  OAI22_X1 U27370 ( .A1(n31169), .A2(n33103), .B1(n30997), .B2(n33105), .ZN(
        n28902) );
  XNOR2_X1 U27371 ( .A(n23577), .B(n23576), .ZN(n28921) );
  OAI21_X1 U27372 ( .B1(n28920), .B2(n28922), .A(n28921), .ZN(n23579) );
  NAND2_X1 U27373 ( .A1(n23579), .A2(n23578), .ZN(n34171) );
  FA_X1 U27374 ( .A(n23582), .B(n23581), .CI(n23580), .CO(n22154), .S(n34170)
         );
  FA_X1 U27375 ( .A(n23585), .B(n23584), .CI(n23583), .CO(n26804), .S(n28915)
         );
  FA_X1 U27376 ( .A(n23588), .B(n23587), .CI(n23586), .CO(n23173), .S(n28914)
         );
  FA_X1 U27377 ( .A(n23591), .B(n23590), .CI(n23589), .CO(n23171), .S(n28913)
         );
  FA_X1 U27378 ( .A(n23594), .B(n23593), .CI(n23592), .CO(n35209), .S(n27313)
         );
  FA_X1 U27379 ( .A(n23597), .B(n23596), .CI(n23595), .CO(n35174), .S(n24848)
         );
  FA_X1 U27380 ( .A(n3493), .B(n23599), .CI(n23598), .CO(n31833), .S(n24847)
         );
  FA_X1 U27381 ( .A(n23602), .B(n23601), .CI(n23600), .CO(n24850), .S(n22153)
         );
  OAI21_X1 U27382 ( .B1(n24848), .B2(n24847), .A(n24850), .ZN(n23604) );
  NAND2_X1 U27383 ( .A1(n24847), .A2(n24848), .ZN(n23603) );
  NAND2_X1 U27384 ( .A1(n23604), .A2(n23603), .ZN(n31807) );
  XNOR2_X1 U27385 ( .A(n32211), .B(\fmem_data[15][5] ), .ZN(n30384) );
  XOR2_X1 U27386 ( .A(\fmem_data[15][4] ), .B(\fmem_data[15][5] ), .Z(n23605)
         );
  AOI22_X1 U27387 ( .A1(n30223), .A2(\xmem_data[64][6] ), .B1(n29697), .B2(
        \xmem_data[65][6] ), .ZN(n23609) );
  AOI22_X1 U27388 ( .A1(n29790), .A2(\xmem_data[66][6] ), .B1(n28218), .B2(
        \xmem_data[67][6] ), .ZN(n23608) );
  AOI22_X1 U27389 ( .A1(n30294), .A2(\xmem_data[68][6] ), .B1(n30776), .B2(
        \xmem_data[69][6] ), .ZN(n23607) );
  AOI22_X1 U27390 ( .A1(n30219), .A2(\xmem_data[70][6] ), .B1(n30295), .B2(
        \xmem_data[71][6] ), .ZN(n23606) );
  NAND4_X1 U27391 ( .A1(n23609), .A2(n23608), .A3(n23607), .A4(n23606), .ZN(
        n23625) );
  AOI22_X1 U27392 ( .A1(n30248), .A2(\xmem_data[72][6] ), .B1(n29589), .B2(
        \xmem_data[73][6] ), .ZN(n23613) );
  AOI22_X1 U27393 ( .A1(n30171), .A2(\xmem_data[74][6] ), .B1(n30083), .B2(
        \xmem_data[75][6] ), .ZN(n23612) );
  AOI22_X1 U27394 ( .A1(n27754), .A2(\xmem_data[76][6] ), .B1(n30084), .B2(
        \xmem_data[77][6] ), .ZN(n23611) );
  AOI22_X1 U27395 ( .A1(n30304), .A2(\xmem_data[78][6] ), .B1(n27945), .B2(
        \xmem_data[79][6] ), .ZN(n23610) );
  NAND4_X1 U27396 ( .A1(n23613), .A2(n23612), .A3(n23611), .A4(n23610), .ZN(
        n23624) );
  AOI22_X1 U27397 ( .A1(n3161), .A2(\xmem_data[80][6] ), .B1(n3183), .B2(
        \xmem_data[81][6] ), .ZN(n23617) );
  AOI22_X1 U27398 ( .A1(n30715), .A2(\xmem_data[82][6] ), .B1(n30309), .B2(
        \xmem_data[83][6] ), .ZN(n23616) );
  AOI22_X1 U27399 ( .A1(n30063), .A2(\xmem_data[84][6] ), .B1(n30170), .B2(
        \xmem_data[85][6] ), .ZN(n23615) );
  AOI22_X1 U27400 ( .A1(n30270), .A2(\xmem_data[86][6] ), .B1(n30311), .B2(
        \xmem_data[87][6] ), .ZN(n23614) );
  NAND4_X1 U27401 ( .A1(n23617), .A2(n23616), .A3(n23615), .A4(n23614), .ZN(
        n23623) );
  AOI22_X1 U27402 ( .A1(n3211), .A2(\xmem_data[88][6] ), .B1(n3193), .B2(
        \xmem_data[89][6] ), .ZN(n23621) );
  AOI22_X1 U27403 ( .A1(n30258), .A2(\xmem_data[90][6] ), .B1(n27852), .B2(
        \xmem_data[91][6] ), .ZN(n23620) );
  AOI22_X1 U27404 ( .A1(n30318), .A2(\xmem_data[92][6] ), .B1(n3420), .B2(
        \xmem_data[93][6] ), .ZN(n23619) );
  AOI22_X1 U27405 ( .A1(n30200), .A2(\xmem_data[94][6] ), .B1(n3153), .B2(
        \xmem_data[95][6] ), .ZN(n23618) );
  NAND4_X1 U27406 ( .A1(n23621), .A2(n23620), .A3(n23619), .A4(n23618), .ZN(
        n23622) );
  OR4_X1 U27407 ( .A1(n23625), .A2(n23624), .A3(n23623), .A4(n23622), .ZN(
        n23647) );
  AOI22_X1 U27408 ( .A1(n29788), .A2(\xmem_data[96][6] ), .B1(n30775), .B2(
        \xmem_data[97][6] ), .ZN(n23629) );
  AOI22_X1 U27409 ( .A1(n30279), .A2(\xmem_data[98][6] ), .B1(n30278), .B2(
        \xmem_data[99][6] ), .ZN(n23628) );
  AOI22_X1 U27410 ( .A1(n30280), .A2(\xmem_data[100][6] ), .B1(n27833), .B2(
        \xmem_data[101][6] ), .ZN(n23627) );
  AOI22_X1 U27411 ( .A1(n30282), .A2(\xmem_data[102][6] ), .B1(n3138), .B2(
        \xmem_data[103][6] ), .ZN(n23626) );
  NAND4_X1 U27412 ( .A1(n23629), .A2(n23628), .A3(n23627), .A4(n23626), .ZN(
        n23645) );
  AOI22_X1 U27413 ( .A1(n28146), .A2(\xmem_data[104][6] ), .B1(n30190), .B2(
        \xmem_data[105][6] ), .ZN(n23633) );
  AOI22_X1 U27414 ( .A1(n30300), .A2(\xmem_data[106][6] ), .B1(n29451), .B2(
        \xmem_data[107][6] ), .ZN(n23632) );
  AOI22_X1 U27415 ( .A1(n28779), .A2(\xmem_data[108][6] ), .B1(n27728), .B2(
        \xmem_data[109][6] ), .ZN(n23631) );
  AOI22_X1 U27416 ( .A1(n30251), .A2(\xmem_data[110][6] ), .B1(n3120), .B2(
        \xmem_data[111][6] ), .ZN(n23630) );
  NAND4_X1 U27417 ( .A1(n23633), .A2(n23632), .A3(n23631), .A4(n23630), .ZN(
        n23644) );
  AOI22_X1 U27418 ( .A1(n3161), .A2(\xmem_data[112][6] ), .B1(n3187), .B2(
        \xmem_data[113][6] ), .ZN(n23637) );
  AOI22_X1 U27419 ( .A1(n29810), .A2(\xmem_data[114][6] ), .B1(n29439), .B2(
        \xmem_data[115][6] ), .ZN(n23636) );
  AOI22_X1 U27420 ( .A1(n29363), .A2(\xmem_data[116][6] ), .B1(n29721), .B2(
        \xmem_data[117][6] ), .ZN(n23635) );
  AOI22_X1 U27421 ( .A1(n30270), .A2(\xmem_data[118][6] ), .B1(n30269), .B2(
        \xmem_data[119][6] ), .ZN(n23634) );
  NAND4_X1 U27422 ( .A1(n23637), .A2(n23636), .A3(n23635), .A4(n23634), .ZN(
        n23643) );
  AOI22_X1 U27423 ( .A1(n3211), .A2(\xmem_data[120][6] ), .B1(n30256), .B2(
        \xmem_data[121][6] ), .ZN(n23641) );
  AOI22_X1 U27424 ( .A1(n30048), .A2(\xmem_data[122][6] ), .B1(n30257), .B2(
        \xmem_data[123][6] ), .ZN(n23640) );
  AOI22_X1 U27425 ( .A1(n30260), .A2(\xmem_data[124][6] ), .B1(n3420), .B2(
        \xmem_data[125][6] ), .ZN(n23639) );
  AOI22_X1 U27426 ( .A1(n30200), .A2(\xmem_data[126][6] ), .B1(n3350), .B2(
        \xmem_data[127][6] ), .ZN(n23638) );
  NAND4_X1 U27427 ( .A1(n23641), .A2(n23640), .A3(n23639), .A4(n23638), .ZN(
        n23642) );
  AOI22_X1 U27428 ( .A1(n27710), .A2(\xmem_data[32][6] ), .B1(n30695), .B2(
        \xmem_data[33][6] ), .ZN(n23651) );
  AOI22_X1 U27429 ( .A1(n28207), .A2(\xmem_data[34][6] ), .B1(n29832), .B2(
        \xmem_data[35][6] ), .ZN(n23650) );
  AOI22_X1 U27430 ( .A1(n30294), .A2(\xmem_data[36][6] ), .B1(n29798), .B2(
        \xmem_data[37][6] ), .ZN(n23649) );
  AOI22_X1 U27431 ( .A1(n30219), .A2(\xmem_data[38][6] ), .B1(n30295), .B2(
        \xmem_data[39][6] ), .ZN(n23648) );
  NAND4_X1 U27432 ( .A1(n23651), .A2(n23650), .A3(n23649), .A4(n23648), .ZN(
        n23667) );
  AOI22_X1 U27433 ( .A1(n29590), .A2(\xmem_data[40][6] ), .B1(n29589), .B2(
        \xmem_data[41][6] ), .ZN(n23655) );
  AOI22_X1 U27434 ( .A1(n30300), .A2(\xmem_data[42][6] ), .B1(n30083), .B2(
        \xmem_data[43][6] ), .ZN(n23654) );
  AOI22_X1 U27435 ( .A1(n29436), .A2(\xmem_data[44][6] ), .B1(n26884), .B2(
        \xmem_data[45][6] ), .ZN(n23653) );
  AOI22_X1 U27436 ( .A1(n30304), .A2(\xmem_data[46][6] ), .B1(n30746), .B2(
        \xmem_data[47][6] ), .ZN(n23652) );
  NAND4_X1 U27437 ( .A1(n23655), .A2(n23654), .A3(n23653), .A4(n23652), .ZN(
        n23666) );
  AOI22_X1 U27438 ( .A1(n3167), .A2(\xmem_data[48][6] ), .B1(n3191), .B2(
        \xmem_data[49][6] ), .ZN(n23659) );
  AOI22_X1 U27439 ( .A1(n30764), .A2(\xmem_data[50][6] ), .B1(n30309), .B2(
        \xmem_data[51][6] ), .ZN(n23658) );
  AOI22_X1 U27440 ( .A1(n28680), .A2(\xmem_data[52][6] ), .B1(n29721), .B2(
        \xmem_data[53][6] ), .ZN(n23657) );
  AOI22_X1 U27441 ( .A1(n30270), .A2(\xmem_data[54][6] ), .B1(n30311), .B2(
        \xmem_data[55][6] ), .ZN(n23656) );
  NAND4_X1 U27442 ( .A1(n23659), .A2(n23658), .A3(n23657), .A4(n23656), .ZN(
        n23665) );
  AOI22_X1 U27443 ( .A1(n3211), .A2(\xmem_data[56][6] ), .B1(n3193), .B2(
        \xmem_data[57][6] ), .ZN(n23663) );
  AOI22_X1 U27444 ( .A1(n30258), .A2(\xmem_data[58][6] ), .B1(n27568), .B2(
        \xmem_data[59][6] ), .ZN(n23662) );
  AOI22_X1 U27445 ( .A1(n30318), .A2(\xmem_data[60][6] ), .B1(n30317), .B2(
        \xmem_data[61][6] ), .ZN(n23661) );
  AOI22_X1 U27446 ( .A1(n30320), .A2(\xmem_data[62][6] ), .B1(n3153), .B2(
        \xmem_data[63][6] ), .ZN(n23660) );
  NAND4_X1 U27447 ( .A1(n23663), .A2(n23662), .A3(n23661), .A4(n23660), .ZN(
        n23664) );
  OR4_X1 U27448 ( .A1(n23667), .A2(n23666), .A3(n23665), .A4(n23664), .ZN(
        n23689) );
  AOI22_X1 U27449 ( .A1(n29421), .A2(\xmem_data[0][6] ), .B1(n27013), .B2(
        \xmem_data[1][6] ), .ZN(n23671) );
  AOI22_X1 U27450 ( .A1(n30279), .A2(\xmem_data[2][6] ), .B1(n30278), .B2(
        \xmem_data[3][6] ), .ZN(n23670) );
  AOI22_X1 U27451 ( .A1(n28219), .A2(\xmem_data[4][6] ), .B1(n30696), .B2(
        \xmem_data[5][6] ), .ZN(n23669) );
  AOI22_X1 U27452 ( .A1(n30219), .A2(\xmem_data[6][6] ), .B1(n3132), .B2(
        \xmem_data[7][6] ), .ZN(n23668) );
  NAND4_X1 U27453 ( .A1(n23671), .A2(n23670), .A3(n23669), .A4(n23668), .ZN(
        n23687) );
  AOI22_X1 U27454 ( .A1(n30191), .A2(\xmem_data[8][6] ), .B1(n29482), .B2(
        \xmem_data[9][6] ), .ZN(n23675) );
  AOI22_X1 U27455 ( .A1(n3214), .A2(\xmem_data[10][6] ), .B1(n28743), .B2(
        \xmem_data[11][6] ), .ZN(n23674) );
  AOI22_X1 U27456 ( .A1(n29395), .A2(\xmem_data[12][6] ), .B1(n26884), .B2(
        \xmem_data[13][6] ), .ZN(n23673) );
  AOI22_X1 U27457 ( .A1(n30304), .A2(\xmem_data[14][6] ), .B1(n31354), .B2(
        \xmem_data[15][6] ), .ZN(n23672) );
  NAND4_X1 U27458 ( .A1(n23675), .A2(n23674), .A3(n23673), .A4(n23672), .ZN(
        n23686) );
  AOI22_X1 U27459 ( .A1(n3167), .A2(\xmem_data[16][6] ), .B1(n3191), .B2(
        \xmem_data[17][6] ), .ZN(n23679) );
  AOI22_X1 U27460 ( .A1(n28689), .A2(\xmem_data[18][6] ), .B1(n21050), .B2(
        \xmem_data[19][6] ), .ZN(n23678) );
  AOI22_X1 U27461 ( .A1(n30198), .A2(\xmem_data[20][6] ), .B1(n30170), .B2(
        \xmem_data[21][6] ), .ZN(n23677) );
  AOI22_X1 U27462 ( .A1(n30205), .A2(\xmem_data[22][6] ), .B1(n31315), .B2(
        \xmem_data[23][6] ), .ZN(n23676) );
  NAND4_X1 U27463 ( .A1(n23679), .A2(n23678), .A3(n23677), .A4(n23676), .ZN(
        n23685) );
  AOI22_X1 U27464 ( .A1(n3210), .A2(\xmem_data[24][6] ), .B1(n3193), .B2(
        \xmem_data[25][6] ), .ZN(n23683) );
  AOI22_X1 U27465 ( .A1(n30258), .A2(\xmem_data[26][6] ), .B1(n20985), .B2(
        \xmem_data[27][6] ), .ZN(n23682) );
  AOI22_X1 U27466 ( .A1(n30199), .A2(\xmem_data[28][6] ), .B1(n3420), .B2(
        \xmem_data[29][6] ), .ZN(n23681) );
  AOI22_X1 U27467 ( .A1(n30200), .A2(\xmem_data[30][6] ), .B1(n3434), .B2(
        \xmem_data[31][6] ), .ZN(n23680) );
  NAND4_X1 U27468 ( .A1(n23683), .A2(n23682), .A3(n23681), .A4(n23680), .ZN(
        n23684) );
  OR4_X1 U27469 ( .A1(n23687), .A2(n23686), .A3(n23685), .A4(n23684), .ZN(
        n23688) );
  AOI22_X1 U27470 ( .A1(n30329), .A2(n23689), .B1(n30228), .B2(n23688), .ZN(
        n23690) );
  AOI22_X1 U27471 ( .A1(n23762), .A2(\xmem_data[64][7] ), .B1(n23761), .B2(
        \xmem_data[65][7] ), .ZN(n23695) );
  AOI22_X1 U27472 ( .A1(n23763), .A2(\xmem_data[66][7] ), .B1(n22703), .B2(
        \xmem_data[67][7] ), .ZN(n23694) );
  AOI22_X1 U27473 ( .A1(n30948), .A2(\xmem_data[68][7] ), .B1(n3213), .B2(
        \xmem_data[69][7] ), .ZN(n23693) );
  AOI22_X1 U27474 ( .A1(n23764), .A2(\xmem_data[70][7] ), .B1(n14970), .B2(
        \xmem_data[71][7] ), .ZN(n23692) );
  NAND4_X1 U27475 ( .A1(n23695), .A2(n23694), .A3(n23693), .A4(n23692), .ZN(
        n23712) );
  AOI22_X1 U27476 ( .A1(n23777), .A2(\xmem_data[72][7] ), .B1(n23776), .B2(
        \xmem_data[73][7] ), .ZN(n23699) );
  AOI22_X1 U27477 ( .A1(n3325), .A2(\xmem_data[74][7] ), .B1(n23778), .B2(
        \xmem_data[75][7] ), .ZN(n23698) );
  AOI22_X1 U27478 ( .A1(n23780), .A2(\xmem_data[76][7] ), .B1(n23779), .B2(
        \xmem_data[77][7] ), .ZN(n23697) );
  AOI22_X1 U27479 ( .A1(n21058), .A2(\xmem_data[78][7] ), .B1(n23781), .B2(
        \xmem_data[79][7] ), .ZN(n23696) );
  NAND4_X1 U27480 ( .A1(n23699), .A2(n23698), .A3(n23697), .A4(n23696), .ZN(
        n23711) );
  AOI22_X1 U27481 ( .A1(n23753), .A2(\xmem_data[80][7] ), .B1(n30524), .B2(
        \xmem_data[81][7] ), .ZN(n23704) );
  AOI22_X1 U27482 ( .A1(n17030), .A2(\xmem_data[82][7] ), .B1(n24625), .B2(
        \xmem_data[83][7] ), .ZN(n23703) );
  AOI22_X1 U27483 ( .A1(n23754), .A2(\xmem_data[84][7] ), .B1(n20568), .B2(
        \xmem_data[85][7] ), .ZN(n23702) );
  AND2_X1 U27484 ( .A1(n3219), .A2(\xmem_data[87][7] ), .ZN(n23700) );
  AOI21_X1 U27485 ( .B1(n23756), .B2(\xmem_data[86][7] ), .A(n23700), .ZN(
        n23701) );
  NAND4_X1 U27486 ( .A1(n23704), .A2(n23703), .A3(n23702), .A4(n23701), .ZN(
        n23710) );
  AOI22_X1 U27487 ( .A1(n23770), .A2(\xmem_data[88][7] ), .B1(n23769), .B2(
        \xmem_data[89][7] ), .ZN(n23708) );
  AOI22_X1 U27488 ( .A1(n29289), .A2(\xmem_data[90][7] ), .B1(n13444), .B2(
        \xmem_data[91][7] ), .ZN(n23707) );
  AOI22_X1 U27489 ( .A1(n29157), .A2(\xmem_data[92][7] ), .B1(n25450), .B2(
        \xmem_data[93][7] ), .ZN(n23706) );
  AOI22_X1 U27490 ( .A1(n27447), .A2(\xmem_data[94][7] ), .B1(n14933), .B2(
        \xmem_data[95][7] ), .ZN(n23705) );
  NAND4_X1 U27491 ( .A1(n23708), .A2(n23707), .A3(n23706), .A4(n23705), .ZN(
        n23709) );
  OR4_X1 U27492 ( .A1(n23712), .A2(n23711), .A3(n23710), .A4(n23709), .ZN(
        n23714) );
  NAND2_X1 U27493 ( .A1(n23714), .A2(n23713), .ZN(n23827) );
  AOI22_X1 U27494 ( .A1(n31327), .A2(\xmem_data[96][7] ), .B1(n13168), .B2(
        \xmem_data[97][7] ), .ZN(n23721) );
  AOI22_X1 U27495 ( .A1(n24131), .A2(\xmem_data[98][7] ), .B1(n23715), .B2(
        \xmem_data[99][7] ), .ZN(n23720) );
  AOI22_X1 U27496 ( .A1(n29807), .A2(\xmem_data[100][7] ), .B1(n23716), .B2(
        \xmem_data[101][7] ), .ZN(n23719) );
  AOI22_X1 U27497 ( .A1(n23717), .A2(\xmem_data[102][7] ), .B1(n31355), .B2(
        \xmem_data[103][7] ), .ZN(n23718) );
  NAND4_X1 U27498 ( .A1(n23721), .A2(n23720), .A3(n23719), .A4(n23718), .ZN(
        n23750) );
  AOI22_X1 U27499 ( .A1(n23722), .A2(\xmem_data[104][7] ), .B1(n23776), .B2(
        \xmem_data[105][7] ), .ZN(n23729) );
  AOI22_X1 U27500 ( .A1(n28428), .A2(\xmem_data[106][7] ), .B1(n25716), .B2(
        \xmem_data[107][7] ), .ZN(n23728) );
  AOI22_X1 U27501 ( .A1(n23724), .A2(\xmem_data[108][7] ), .B1(n23723), .B2(
        \xmem_data[109][7] ), .ZN(n23727) );
  AOI22_X1 U27502 ( .A1(n20782), .A2(\xmem_data[110][7] ), .B1(n23725), .B2(
        \xmem_data[111][7] ), .ZN(n23726) );
  NAND4_X1 U27503 ( .A1(n23729), .A2(n23728), .A3(n23727), .A4(n23726), .ZN(
        n23749) );
  AOI22_X1 U27504 ( .A1(n23730), .A2(\xmem_data[112][7] ), .B1(n31261), .B2(
        \xmem_data[113][7] ), .ZN(n23738) );
  AOI22_X1 U27505 ( .A1(n17056), .A2(\xmem_data[114][7] ), .B1(n24625), .B2(
        \xmem_data[115][7] ), .ZN(n23737) );
  AOI22_X1 U27506 ( .A1(n23732), .A2(\xmem_data[116][7] ), .B1(n23731), .B2(
        \xmem_data[117][7] ), .ZN(n23736) );
  AND2_X1 U27507 ( .A1(n3219), .A2(\xmem_data[119][7] ), .ZN(n23733) );
  AOI21_X1 U27508 ( .B1(n23734), .B2(\xmem_data[118][7] ), .A(n23733), .ZN(
        n23735) );
  NAND4_X1 U27509 ( .A1(n23738), .A2(n23737), .A3(n23736), .A4(n23735), .ZN(
        n23748) );
  AOI22_X1 U27510 ( .A1(n23740), .A2(\xmem_data[120][7] ), .B1(n23739), .B2(
        \xmem_data[121][7] ), .ZN(n23746) );
  AOI22_X1 U27511 ( .A1(n23741), .A2(\xmem_data[122][7] ), .B1(n20993), .B2(
        \xmem_data[123][7] ), .ZN(n23745) );
  AOI22_X1 U27512 ( .A1(n23742), .A2(\xmem_data[124][7] ), .B1(n28510), .B2(
        \xmem_data[125][7] ), .ZN(n23744) );
  AOI22_X1 U27513 ( .A1(n27447), .A2(\xmem_data[126][7] ), .B1(n29180), .B2(
        \xmem_data[127][7] ), .ZN(n23743) );
  NAND4_X1 U27514 ( .A1(n23746), .A2(n23745), .A3(n23744), .A4(n23743), .ZN(
        n23747) );
  OR4_X1 U27515 ( .A1(n23750), .A2(n23749), .A3(n23748), .A4(n23747), .ZN(
        n23752) );
  NAND2_X1 U27516 ( .A1(n23752), .A2(n23751), .ZN(n23826) );
  AOI22_X1 U27517 ( .A1(n23753), .A2(\xmem_data[48][7] ), .B1(n20769), .B2(
        \xmem_data[49][7] ), .ZN(n23760) );
  AOI22_X1 U27518 ( .A1(n25408), .A2(\xmem_data[50][7] ), .B1(n20489), .B2(
        \xmem_data[51][7] ), .ZN(n23759) );
  AOI22_X1 U27519 ( .A1(n23754), .A2(\xmem_data[52][7] ), .B1(n29286), .B2(
        \xmem_data[53][7] ), .ZN(n23758) );
  AND2_X1 U27520 ( .A1(n3221), .A2(\xmem_data[55][7] ), .ZN(n23755) );
  AOI21_X1 U27521 ( .B1(n23756), .B2(\xmem_data[54][7] ), .A(n23755), .ZN(
        n23757) );
  NAND4_X1 U27522 ( .A1(n23760), .A2(n23759), .A3(n23758), .A4(n23757), .ZN(
        n23789) );
  AOI22_X1 U27523 ( .A1(n23762), .A2(\xmem_data[32][7] ), .B1(n23761), .B2(
        \xmem_data[33][7] ), .ZN(n23768) );
  AOI22_X1 U27524 ( .A1(n23763), .A2(\xmem_data[34][7] ), .B1(n28052), .B2(
        \xmem_data[35][7] ), .ZN(n23767) );
  AOI22_X1 U27525 ( .A1(n16988), .A2(\xmem_data[36][7] ), .B1(n25460), .B2(
        \xmem_data[37][7] ), .ZN(n23766) );
  AOI22_X1 U27526 ( .A1(n23764), .A2(\xmem_data[38][7] ), .B1(n22718), .B2(
        \xmem_data[39][7] ), .ZN(n23765) );
  NAND4_X1 U27527 ( .A1(n23768), .A2(n23767), .A3(n23766), .A4(n23765), .ZN(
        n23788) );
  AOI22_X1 U27528 ( .A1(n23770), .A2(\xmem_data[56][7] ), .B1(n23769), .B2(
        \xmem_data[57][7] ), .ZN(n23775) );
  AOI22_X1 U27529 ( .A1(n24534), .A2(\xmem_data[58][7] ), .B1(n3255), .B2(
        \xmem_data[59][7] ), .ZN(n23774) );
  AOI22_X1 U27530 ( .A1(n30698), .A2(\xmem_data[60][7] ), .B1(n25450), .B2(
        \xmem_data[61][7] ), .ZN(n23773) );
  AOI22_X1 U27531 ( .A1(n27447), .A2(\xmem_data[62][7] ), .B1(n20588), .B2(
        \xmem_data[63][7] ), .ZN(n23772) );
  NAND4_X1 U27532 ( .A1(n23775), .A2(n23774), .A3(n23773), .A4(n23772), .ZN(
        n23787) );
  AOI22_X1 U27533 ( .A1(n23777), .A2(\xmem_data[40][7] ), .B1(n23776), .B2(
        \xmem_data[41][7] ), .ZN(n23785) );
  AOI22_X1 U27534 ( .A1(n25575), .A2(\xmem_data[42][7] ), .B1(n23778), .B2(
        \xmem_data[43][7] ), .ZN(n23784) );
  AOI22_X1 U27535 ( .A1(n23780), .A2(\xmem_data[44][7] ), .B1(n23779), .B2(
        \xmem_data[45][7] ), .ZN(n23783) );
  AOI22_X1 U27536 ( .A1(n20818), .A2(\xmem_data[46][7] ), .B1(n23781), .B2(
        \xmem_data[47][7] ), .ZN(n23782) );
  NAND4_X1 U27537 ( .A1(n23785), .A2(n23784), .A3(n23783), .A4(n23782), .ZN(
        n23786) );
  OR4_X1 U27538 ( .A1(n23789), .A2(n23788), .A3(n23787), .A4(n23786), .ZN(
        n23791) );
  NAND2_X1 U27539 ( .A1(n23791), .A2(n23790), .ZN(n23825) );
  AOI22_X1 U27540 ( .A1(n23792), .A2(\xmem_data[0][7] ), .B1(n24212), .B2(
        \xmem_data[1][7] ), .ZN(n23800) );
  AOI22_X1 U27541 ( .A1(n17041), .A2(\xmem_data[2][7] ), .B1(n23793), .B2(
        \xmem_data[3][7] ), .ZN(n23799) );
  AOI22_X1 U27542 ( .A1(n30746), .A2(\xmem_data[4][7] ), .B1(n3208), .B2(
        \xmem_data[5][7] ), .ZN(n23798) );
  AOI22_X1 U27543 ( .A1(n24509), .A2(\xmem_data[6][7] ), .B1(n23796), .B2(
        \xmem_data[7][7] ), .ZN(n23797) );
  NAND4_X1 U27544 ( .A1(n23800), .A2(n23799), .A3(n23798), .A4(n23797), .ZN(
        n23821) );
  AOI22_X1 U27545 ( .A1(n23802), .A2(\xmem_data[8][7] ), .B1(n23801), .B2(
        \xmem_data[9][7] ), .ZN(n23806) );
  AOI22_X1 U27546 ( .A1(n30557), .A2(\xmem_data[10][7] ), .B1(n20506), .B2(
        \xmem_data[11][7] ), .ZN(n23805) );
  AOI22_X1 U27547 ( .A1(n3307), .A2(\xmem_data[12][7] ), .B1(n27365), .B2(
        \xmem_data[13][7] ), .ZN(n23804) );
  AOI22_X1 U27548 ( .A1(n20782), .A2(\xmem_data[14][7] ), .B1(n21057), .B2(
        \xmem_data[15][7] ), .ZN(n23803) );
  NAND4_X1 U27549 ( .A1(n23806), .A2(n23805), .A3(n23804), .A4(n23803), .ZN(
        n23820) );
  AOI22_X1 U27550 ( .A1(n30674), .A2(\xmem_data[16][7] ), .B1(n31261), .B2(
        \xmem_data[17][7] ), .ZN(n23810) );
  AOI22_X1 U27551 ( .A1(n27564), .A2(\xmem_data[18][7] ), .B1(n24625), .B2(
        \xmem_data[19][7] ), .ZN(n23809) );
  AOI22_X1 U27552 ( .A1(n3228), .A2(\xmem_data[20][7] ), .B1(n28501), .B2(
        \xmem_data[21][7] ), .ZN(n23808) );
  AOI22_X1 U27553 ( .A1(n28364), .A2(\xmem_data[22][7] ), .B1(n3218), .B2(
        \xmem_data[23][7] ), .ZN(n23807) );
  NAND4_X1 U27554 ( .A1(n23810), .A2(n23809), .A3(n23808), .A4(n23807), .ZN(
        n23819) );
  AOI22_X1 U27555 ( .A1(n20805), .A2(\xmem_data[24][7] ), .B1(n31367), .B2(
        \xmem_data[25][7] ), .ZN(n23817) );
  AOI22_X1 U27556 ( .A1(n23812), .A2(\xmem_data[26][7] ), .B1(n23811), .B2(
        \xmem_data[27][7] ), .ZN(n23816) );
  AOI22_X1 U27557 ( .A1(n29706), .A2(\xmem_data[28][7] ), .B1(n13474), .B2(
        \xmem_data[29][7] ), .ZN(n23815) );
  AOI22_X1 U27558 ( .A1(n23813), .A2(\xmem_data[30][7] ), .B1(n13475), .B2(
        \xmem_data[31][7] ), .ZN(n23814) );
  NAND4_X1 U27559 ( .A1(n23817), .A2(n23816), .A3(n23815), .A4(n23814), .ZN(
        n23818) );
  OR4_X1 U27560 ( .A1(n23821), .A2(n23820), .A3(n23819), .A4(n23818), .ZN(
        n23823) );
  NAND2_X1 U27561 ( .A1(n23823), .A2(n23822), .ZN(n23824) );
  XNOR2_X1 U27562 ( .A(n35324), .B(\fmem_data[4][3] ), .ZN(n33056) );
  XNOR2_X1 U27563 ( .A(n31882), .B(\fmem_data[21][5] ), .ZN(n30436) );
  XNOR2_X1 U27564 ( .A(n31660), .B(\fmem_data[21][5] ), .ZN(n33303) );
  OAI22_X1 U27565 ( .A1(n30436), .A2(n34194), .B1(n33303), .B2(n34195), .ZN(
        n26030) );
  XNOR2_X1 U27566 ( .A(n28539), .B(\fmem_data[13][7] ), .ZN(n33132) );
  FA_X1 U27567 ( .A(n23830), .B(n23829), .CI(n23828), .CO(n24838), .S(n26795)
         );
  XNOR2_X1 U27568 ( .A(n31807), .B(n31806), .ZN(n23924) );
  AOI22_X1 U27569 ( .A1(n29421), .A2(\xmem_data[32][7] ), .B1(n29753), .B2(
        \xmem_data[33][7] ), .ZN(n23834) );
  AOI22_X1 U27570 ( .A1(n29628), .A2(\xmem_data[34][7] ), .B1(n30292), .B2(
        \xmem_data[35][7] ), .ZN(n23833) );
  AOI22_X1 U27571 ( .A1(n30294), .A2(\xmem_data[36][7] ), .B1(n3170), .B2(
        \xmem_data[37][7] ), .ZN(n23832) );
  AOI22_X1 U27572 ( .A1(n30219), .A2(\xmem_data[38][7] ), .B1(n30295), .B2(
        \xmem_data[39][7] ), .ZN(n23831) );
  NAND4_X1 U27573 ( .A1(n23834), .A2(n23833), .A3(n23832), .A4(n23831), .ZN(
        n23850) );
  AOI22_X1 U27574 ( .A1(n3249), .A2(\xmem_data[40][7] ), .B1(n30190), .B2(
        \xmem_data[41][7] ), .ZN(n23838) );
  AOI22_X1 U27575 ( .A1(n3214), .A2(\xmem_data[42][7] ), .B1(n27763), .B2(
        \xmem_data[43][7] ), .ZN(n23837) );
  AOI22_X1 U27576 ( .A1(n3174), .A2(\xmem_data[44][7] ), .B1(n28110), .B2(
        \xmem_data[45][7] ), .ZN(n23836) );
  AOI22_X1 U27577 ( .A1(n30304), .A2(\xmem_data[46][7] ), .B1(n29396), .B2(
        \xmem_data[47][7] ), .ZN(n23835) );
  NAND4_X1 U27578 ( .A1(n23838), .A2(n23837), .A3(n23836), .A4(n23835), .ZN(
        n23849) );
  AOI22_X1 U27579 ( .A1(n3165), .A2(\xmem_data[48][7] ), .B1(n3191), .B2(
        \xmem_data[49][7] ), .ZN(n23842) );
  AOI22_X1 U27580 ( .A1(n26812), .A2(\xmem_data[50][7] ), .B1(n30309), .B2(
        \xmem_data[51][7] ), .ZN(n23841) );
  AOI22_X1 U27581 ( .A1(n29815), .A2(\xmem_data[52][7] ), .B1(n29487), .B2(
        \xmem_data[53][7] ), .ZN(n23840) );
  AOI22_X1 U27582 ( .A1(n30270), .A2(\xmem_data[54][7] ), .B1(n30311), .B2(
        \xmem_data[55][7] ), .ZN(n23839) );
  NAND4_X1 U27583 ( .A1(n23842), .A2(n23841), .A3(n23840), .A4(n23839), .ZN(
        n23848) );
  AOI22_X1 U27584 ( .A1(n3211), .A2(\xmem_data[56][7] ), .B1(n3193), .B2(
        \xmem_data[57][7] ), .ZN(n23846) );
  AOI22_X1 U27585 ( .A1(n30258), .A2(\xmem_data[58][7] ), .B1(n29298), .B2(
        \xmem_data[59][7] ), .ZN(n23845) );
  AOI22_X1 U27586 ( .A1(n30318), .A2(\xmem_data[60][7] ), .B1(n30317), .B2(
        \xmem_data[61][7] ), .ZN(n23844) );
  AOI22_X1 U27587 ( .A1(n30320), .A2(\xmem_data[62][7] ), .B1(n3153), .B2(
        \xmem_data[63][7] ), .ZN(n23843) );
  NAND4_X1 U27588 ( .A1(n23846), .A2(n23845), .A3(n23844), .A4(n23843), .ZN(
        n23847) );
  OR4_X1 U27589 ( .A1(n23850), .A2(n23849), .A3(n23848), .A4(n23847), .ZN(
        n23872) );
  AOI22_X1 U27590 ( .A1(n28136), .A2(\xmem_data[0][7] ), .B1(n30182), .B2(
        \xmem_data[1][7] ), .ZN(n23854) );
  AOI22_X1 U27591 ( .A1(n3392), .A2(\xmem_data[2][7] ), .B1(n30292), .B2(
        \xmem_data[3][7] ), .ZN(n23853) );
  AOI22_X1 U27592 ( .A1(n30294), .A2(\xmem_data[4][7] ), .B1(n28786), .B2(
        \xmem_data[5][7] ), .ZN(n23852) );
  AOI22_X1 U27593 ( .A1(n30219), .A2(\xmem_data[6][7] ), .B1(n3131), .B2(
        \xmem_data[7][7] ), .ZN(n23851) );
  NAND4_X1 U27594 ( .A1(n23854), .A2(n23853), .A3(n23852), .A4(n23851), .ZN(
        n23870) );
  AOI22_X1 U27595 ( .A1(n3249), .A2(\xmem_data[8][7] ), .B1(n28665), .B2(
        \xmem_data[9][7] ), .ZN(n23858) );
  AOI22_X1 U27596 ( .A1(n30192), .A2(\xmem_data[10][7] ), .B1(n28152), .B2(
        \xmem_data[11][7] ), .ZN(n23857) );
  AOI22_X1 U27597 ( .A1(n28685), .A2(\xmem_data[12][7] ), .B1(n30301), .B2(
        \xmem_data[13][7] ), .ZN(n23856) );
  AOI22_X1 U27598 ( .A1(n30304), .A2(\xmem_data[14][7] ), .B1(n28752), .B2(
        \xmem_data[15][7] ), .ZN(n23855) );
  NAND4_X1 U27599 ( .A1(n23858), .A2(n23857), .A3(n23856), .A4(n23855), .ZN(
        n23869) );
  AOI22_X1 U27600 ( .A1(n23901), .A2(\xmem_data[18][7] ), .B1(n30309), .B2(
        \xmem_data[19][7] ), .ZN(n23862) );
  AOI22_X1 U27601 ( .A1(n3164), .A2(\xmem_data[16][7] ), .B1(n3183), .B2(
        \xmem_data[17][7] ), .ZN(n23861) );
  AOI22_X1 U27602 ( .A1(n30198), .A2(\xmem_data[20][7] ), .B1(n29487), .B2(
        \xmem_data[21][7] ), .ZN(n23860) );
  AOI22_X1 U27603 ( .A1(n30205), .A2(\xmem_data[22][7] ), .B1(n28701), .B2(
        \xmem_data[23][7] ), .ZN(n23859) );
  NAND4_X1 U27604 ( .A1(n23862), .A2(n23861), .A3(n23860), .A4(n23859), .ZN(
        n23868) );
  AOI22_X1 U27605 ( .A1(n3210), .A2(\xmem_data[24][7] ), .B1(n3193), .B2(
        \xmem_data[25][7] ), .ZN(n23866) );
  AOI22_X1 U27606 ( .A1(n30258), .A2(\xmem_data[26][7] ), .B1(n28036), .B2(
        \xmem_data[27][7] ), .ZN(n23865) );
  AOI22_X1 U27607 ( .A1(n30199), .A2(\xmem_data[28][7] ), .B1(n3420), .B2(
        \xmem_data[29][7] ), .ZN(n23864) );
  AOI22_X1 U27608 ( .A1(n30200), .A2(\xmem_data[30][7] ), .B1(n3153), .B2(
        \xmem_data[31][7] ), .ZN(n23863) );
  NAND4_X1 U27609 ( .A1(n23866), .A2(n23865), .A3(n23864), .A4(n23863), .ZN(
        n23867) );
  AOI22_X1 U27610 ( .A1(n30329), .A2(n23872), .B1(n30228), .B2(n23871), .ZN(
        n23917) );
  AOI22_X1 U27611 ( .A1(n28734), .A2(\xmem_data[64][7] ), .B1(n30290), .B2(
        \xmem_data[65][7] ), .ZN(n23876) );
  AOI22_X1 U27612 ( .A1(n30279), .A2(\xmem_data[66][7] ), .B1(n30278), .B2(
        \xmem_data[67][7] ), .ZN(n23875) );
  AOI22_X1 U27613 ( .A1(n30294), .A2(\xmem_data[68][7] ), .B1(n30696), .B2(
        \xmem_data[69][7] ), .ZN(n23874) );
  AOI22_X1 U27614 ( .A1(n30219), .A2(\xmem_data[70][7] ), .B1(n30295), .B2(
        \xmem_data[71][7] ), .ZN(n23873) );
  NAND4_X1 U27615 ( .A1(n23876), .A2(n23875), .A3(n23874), .A4(n23873), .ZN(
        n23892) );
  AOI22_X1 U27616 ( .A1(n29705), .A2(\xmem_data[72][7] ), .B1(n30730), .B2(
        \xmem_data[73][7] ), .ZN(n23880) );
  AOI22_X1 U27617 ( .A1(n30171), .A2(\xmem_data[74][7] ), .B1(n31353), .B2(
        \xmem_data[75][7] ), .ZN(n23879) );
  AOI22_X1 U27618 ( .A1(n30665), .A2(\xmem_data[76][7] ), .B1(n29768), .B2(
        \xmem_data[77][7] ), .ZN(n23878) );
  AOI22_X1 U27619 ( .A1(n30304), .A2(\xmem_data[78][7] ), .B1(n29315), .B2(
        \xmem_data[79][7] ), .ZN(n23877) );
  NAND4_X1 U27620 ( .A1(n23880), .A2(n23879), .A3(n23878), .A4(n23877), .ZN(
        n23891) );
  AOI22_X1 U27621 ( .A1(n3166), .A2(\xmem_data[80][7] ), .B1(n3184), .B2(
        \xmem_data[81][7] ), .ZN(n23884) );
  AOI22_X1 U27622 ( .A1(n29716), .A2(\xmem_data[82][7] ), .B1(n30309), .B2(
        \xmem_data[83][7] ), .ZN(n23883) );
  AOI22_X1 U27623 ( .A1(n28173), .A2(\xmem_data[84][7] ), .B1(n30170), .B2(
        \xmem_data[85][7] ), .ZN(n23882) );
  AOI22_X1 U27624 ( .A1(n30270), .A2(\xmem_data[86][7] ), .B1(n30311), .B2(
        \xmem_data[87][7] ), .ZN(n23881) );
  NAND4_X1 U27625 ( .A1(n23884), .A2(n23883), .A3(n23882), .A4(n23881), .ZN(
        n23890) );
  AOI22_X1 U27626 ( .A1(n3210), .A2(\xmem_data[88][7] ), .B1(n3193), .B2(
        \xmem_data[89][7] ), .ZN(n23888) );
  AOI22_X1 U27627 ( .A1(n30048), .A2(\xmem_data[90][7] ), .B1(n21060), .B2(
        \xmem_data[91][7] ), .ZN(n23887) );
  AOI22_X1 U27628 ( .A1(n30318), .A2(\xmem_data[92][7] ), .B1(n3420), .B2(
        \xmem_data[93][7] ), .ZN(n23886) );
  AOI22_X1 U27629 ( .A1(n30200), .A2(\xmem_data[94][7] ), .B1(n3153), .B2(
        \xmem_data[95][7] ), .ZN(n23885) );
  NAND4_X1 U27630 ( .A1(n23888), .A2(n23887), .A3(n23886), .A4(n23885), .ZN(
        n23889) );
  OR4_X1 U27631 ( .A1(n23892), .A2(n23891), .A3(n23890), .A4(n23889), .ZN(
        n23915) );
  AOI22_X1 U27632 ( .A1(n29433), .A2(\xmem_data[96][7] ), .B1(n30290), .B2(
        \xmem_data[97][7] ), .ZN(n23896) );
  AOI22_X1 U27633 ( .A1(n28700), .A2(\xmem_data[98][7] ), .B1(n30278), .B2(
        \xmem_data[99][7] ), .ZN(n23895) );
  AOI22_X1 U27634 ( .A1(n30280), .A2(\xmem_data[100][7] ), .B1(n29629), .B2(
        \xmem_data[101][7] ), .ZN(n23894) );
  AOI22_X1 U27635 ( .A1(n30282), .A2(\xmem_data[102][7] ), .B1(n3137), .B2(
        \xmem_data[103][7] ), .ZN(n23893) );
  NAND4_X1 U27636 ( .A1(n23896), .A2(n23895), .A3(n23894), .A4(n23893), .ZN(
        n23913) );
  AOI22_X1 U27637 ( .A1(n30248), .A2(\xmem_data[104][7] ), .B1(n29347), .B2(
        \xmem_data[105][7] ), .ZN(n23900) );
  AOI22_X1 U27638 ( .A1(n30300), .A2(\xmem_data[106][7] ), .B1(n30083), .B2(
        \xmem_data[107][7] ), .ZN(n23899) );
  AOI22_X1 U27639 ( .A1(n27754), .A2(\xmem_data[108][7] ), .B1(n30249), .B2(
        \xmem_data[109][7] ), .ZN(n23898) );
  AOI22_X1 U27640 ( .A1(n30251), .A2(\xmem_data[110][7] ), .B1(n29437), .B2(
        \xmem_data[111][7] ), .ZN(n23897) );
  NAND4_X1 U27641 ( .A1(n23900), .A2(n23899), .A3(n23898), .A4(n23897), .ZN(
        n23912) );
  AOI22_X1 U27642 ( .A1(n23901), .A2(\xmem_data[114][7] ), .B1(n27825), .B2(
        \xmem_data[115][7] ), .ZN(n23905) );
  AOI22_X1 U27643 ( .A1(n3161), .A2(\xmem_data[112][7] ), .B1(n3191), .B2(
        \xmem_data[113][7] ), .ZN(n23904) );
  AOI22_X1 U27644 ( .A1(n27713), .A2(\xmem_data[116][7] ), .B1(n30685), .B2(
        \xmem_data[117][7] ), .ZN(n23903) );
  AOI22_X1 U27645 ( .A1(n30270), .A2(\xmem_data[118][7] ), .B1(n30269), .B2(
        \xmem_data[119][7] ), .ZN(n23902) );
  NAND4_X1 U27646 ( .A1(n23905), .A2(n23904), .A3(n23903), .A4(n23902), .ZN(
        n23911) );
  AOI22_X1 U27647 ( .A1(n3210), .A2(\xmem_data[120][7] ), .B1(n30256), .B2(
        \xmem_data[121][7] ), .ZN(n23909) );
  AOI22_X1 U27648 ( .A1(n30258), .A2(\xmem_data[122][7] ), .B1(n30257), .B2(
        \xmem_data[123][7] ), .ZN(n23908) );
  AOI22_X1 U27649 ( .A1(n30260), .A2(\xmem_data[124][7] ), .B1(n3420), .B2(
        \xmem_data[125][7] ), .ZN(n23907) );
  AOI22_X1 U27650 ( .A1(n30200), .A2(\xmem_data[126][7] ), .B1(n3305), .B2(
        \xmem_data[127][7] ), .ZN(n23906) );
  NAND4_X1 U27651 ( .A1(n23909), .A2(n23908), .A3(n23907), .A4(n23906), .ZN(
        n23910) );
  XOR2_X1 U27652 ( .A(\fmem_data[9][4] ), .B(\fmem_data[9][5] ), .Z(n23919) );
  XNOR2_X1 U27653 ( .A(n35021), .B(\fmem_data[9][5] ), .ZN(n34861) );
  XNOR2_X1 U27654 ( .A(n32228), .B(\fmem_data[5][7] ), .ZN(n30357) );
  OAI22_X1 U27655 ( .A1(n30357), .A2(n35497), .B1(n23920), .B2(n35498), .ZN(
        n25600) );
  XNOR2_X1 U27656 ( .A(n31897), .B(\fmem_data[28][7] ), .ZN(n30354) );
  FA_X1 U27657 ( .A(n23923), .B(n23922), .CI(n23921), .CO(n31783), .S(n16355)
         );
  XNOR2_X1 U27658 ( .A(n23924), .B(n31805), .ZN(n31848) );
  XNOR2_X1 U27659 ( .A(n35270), .B(\fmem_data[19][5] ), .ZN(n34921) );
  XNOR2_X1 U27660 ( .A(n31246), .B(\fmem_data[11][7] ), .ZN(n35113) );
  OAI22_X1 U27661 ( .A1(n35113), .A2(n35634), .B1(n23925), .B2(n35633), .ZN(
        n31781) );
  XNOR2_X1 U27662 ( .A(n3321), .B(\fmem_data[27][7] ), .ZN(n35146) );
  AOI22_X1 U27663 ( .A1(n27834), .A2(\xmem_data[112][4] ), .B1(n28208), .B2(
        \xmem_data[113][4] ), .ZN(n23929) );
  AOI22_X1 U27664 ( .A1(n3223), .A2(\xmem_data[114][4] ), .B1(n3140), .B2(
        \xmem_data[115][4] ), .ZN(n23928) );
  AOI22_X1 U27665 ( .A1(n27703), .A2(\xmem_data[116][4] ), .B1(n29389), .B2(
        \xmem_data[117][4] ), .ZN(n23927) );
  AOI22_X1 U27666 ( .A1(n29709), .A2(\xmem_data[118][4] ), .B1(n25457), .B2(
        \xmem_data[119][4] ), .ZN(n23926) );
  NAND4_X1 U27667 ( .A1(n23929), .A2(n23928), .A3(n23927), .A4(n23926), .ZN(
        n23945) );
  AOI22_X1 U27668 ( .A1(n7451), .A2(\xmem_data[104][4] ), .B1(n27812), .B2(
        \xmem_data[105][4] ), .ZN(n23933) );
  AOI22_X1 U27669 ( .A1(n27814), .A2(\xmem_data[106][4] ), .B1(n27813), .B2(
        \xmem_data[107][4] ), .ZN(n23932) );
  AOI22_X1 U27670 ( .A1(n27741), .A2(\xmem_data[108][4] ), .B1(n30654), .B2(
        \xmem_data[109][4] ), .ZN(n23931) );
  AOI22_X1 U27671 ( .A1(n28207), .A2(\xmem_data[110][4] ), .B1(n27831), .B2(
        \xmem_data[111][4] ), .ZN(n23930) );
  NAND4_X1 U27672 ( .A1(n23933), .A2(n23932), .A3(n23931), .A4(n23930), .ZN(
        n23944) );
  AOI22_X1 U27673 ( .A1(n3174), .A2(\xmem_data[120][4] ), .B1(n30237), .B2(
        \xmem_data[121][4] ), .ZN(n23937) );
  AOI22_X1 U27674 ( .A1(n27819), .A2(\xmem_data[122][4] ), .B1(n28752), .B2(
        \xmem_data[123][4] ), .ZN(n23936) );
  AOI22_X1 U27675 ( .A1(n3167), .A2(\xmem_data[124][4] ), .B1(n3191), .B2(
        \xmem_data[125][4] ), .ZN(n23935) );
  AOI22_X1 U27676 ( .A1(n23901), .A2(\xmem_data[126][4] ), .B1(n28147), .B2(
        \xmem_data[127][4] ), .ZN(n23934) );
  NAND4_X1 U27677 ( .A1(n23937), .A2(n23936), .A3(n23935), .A4(n23934), .ZN(
        n23943) );
  AOI22_X1 U27678 ( .A1(n30076), .A2(\xmem_data[96][4] ), .B1(n29487), .B2(
        \xmem_data[97][4] ), .ZN(n23941) );
  AOI22_X1 U27679 ( .A1(n27804), .A2(\xmem_data[98][4] ), .B1(n23724), .B2(
        \xmem_data[99][4] ), .ZN(n23940) );
  AOI22_X1 U27680 ( .A1(n29724), .A2(\xmem_data[100][4] ), .B1(n27805), .B2(
        \xmem_data[101][4] ), .ZN(n23939) );
  AOI22_X1 U27681 ( .A1(n27806), .A2(\xmem_data[102][4] ), .B1(n29383), .B2(
        \xmem_data[103][4] ), .ZN(n23938) );
  NAND4_X1 U27682 ( .A1(n23941), .A2(n23940), .A3(n23939), .A4(n23938), .ZN(
        n23942) );
  OR4_X1 U27683 ( .A1(n23945), .A2(n23944), .A3(n23943), .A4(n23942), .ZN(
        n23946) );
  NAND2_X1 U27684 ( .A1(n23946), .A2(n27801), .ZN(n24014) );
  AOI22_X1 U27685 ( .A1(n27701), .A2(\xmem_data[48][4] ), .B1(n28667), .B2(
        \xmem_data[49][4] ), .ZN(n23950) );
  AOI22_X1 U27686 ( .A1(n27702), .A2(\xmem_data[50][4] ), .B1(n3140), .B2(
        \xmem_data[51][4] ), .ZN(n23949) );
  AOI22_X1 U27687 ( .A1(n30633), .A2(\xmem_data[52][4] ), .B1(n29347), .B2(
        \xmem_data[53][4] ), .ZN(n23948) );
  AOI22_X1 U27688 ( .A1(n29802), .A2(\xmem_data[54][4] ), .B1(n28051), .B2(
        \xmem_data[55][4] ), .ZN(n23947) );
  NAND4_X1 U27689 ( .A1(n23948), .A2(n23949), .A3(n23950), .A4(n23947), .ZN(
        n23966) );
  AOI22_X1 U27690 ( .A1(n28765), .A2(\xmem_data[40][4] ), .B1(n27723), .B2(
        \xmem_data[41][4] ), .ZN(n23954) );
  AOI22_X1 U27691 ( .A1(n27742), .A2(\xmem_data[42][4] ), .B1(n3149), .B2(
        \xmem_data[43][4] ), .ZN(n23953) );
  AOI22_X1 U27692 ( .A1(n29626), .A2(\xmem_data[44][4] ), .B1(n28206), .B2(
        \xmem_data[45][4] ), .ZN(n23952) );
  AOI22_X1 U27693 ( .A1(n3392), .A2(\xmem_data[46][4] ), .B1(n27708), .B2(
        \xmem_data[47][4] ), .ZN(n23951) );
  NAND4_X1 U27694 ( .A1(n23954), .A2(n23953), .A3(n23952), .A4(n23951), .ZN(
        n23965) );
  AOI22_X1 U27695 ( .A1(n3174), .A2(\xmem_data[56][4] ), .B1(n30090), .B2(
        \xmem_data[57][4] ), .ZN(n23958) );
  AOI22_X1 U27696 ( .A1(n27729), .A2(\xmem_data[58][4] ), .B1(n24213), .B2(
        \xmem_data[59][4] ), .ZN(n23957) );
  AOI22_X1 U27697 ( .A1(n3161), .A2(\xmem_data[60][4] ), .B1(n3187), .B2(
        \xmem_data[61][4] ), .ZN(n23956) );
  AOI22_X1 U27698 ( .A1(n23901), .A2(\xmem_data[62][4] ), .B1(n25400), .B2(
        \xmem_data[63][4] ), .ZN(n23955) );
  NAND4_X1 U27699 ( .A1(n23958), .A2(n23957), .A3(n23956), .A4(n23955), .ZN(
        n23964) );
  AOI22_X1 U27700 ( .A1(n28680), .A2(\xmem_data[32][4] ), .B1(n30266), .B2(
        \xmem_data[33][4] ), .ZN(n23962) );
  AOI22_X1 U27701 ( .A1(n27714), .A2(\xmem_data[34][4] ), .B1(n3328), .B2(
        \xmem_data[35][4] ), .ZN(n23961) );
  AOI22_X1 U27702 ( .A1(n27716), .A2(\xmem_data[36][4] ), .B1(n27715), .B2(
        \xmem_data[37][4] ), .ZN(n23960) );
  AOI22_X1 U27703 ( .A1(n27718), .A2(\xmem_data[38][4] ), .B1(n27717), .B2(
        \xmem_data[39][4] ), .ZN(n23959) );
  NAND4_X1 U27704 ( .A1(n23962), .A2(n23961), .A3(n23960), .A4(n23959), .ZN(
        n23963) );
  OR4_X1 U27705 ( .A1(n23964), .A2(n23965), .A3(n23966), .A4(n23963), .ZN(
        n23967) );
  NAND2_X1 U27706 ( .A1(n23967), .A2(n27737), .ZN(n24013) );
  AOI22_X1 U27707 ( .A1(n28765), .A2(\xmem_data[72][4] ), .B1(n27723), .B2(
        \xmem_data[73][4] ), .ZN(n23971) );
  AOI22_X1 U27708 ( .A1(n11850), .A2(\xmem_data[74][4] ), .B1(n3149), .B2(
        \xmem_data[75][4] ), .ZN(n23970) );
  AOI22_X1 U27709 ( .A1(n28734), .A2(\xmem_data[76][4] ), .B1(n30182), .B2(
        \xmem_data[77][4] ), .ZN(n23969) );
  AOI22_X1 U27710 ( .A1(n3392), .A2(\xmem_data[78][4] ), .B1(n27708), .B2(
        \xmem_data[79][4] ), .ZN(n23968) );
  NAND4_X1 U27711 ( .A1(n23971), .A2(n23970), .A3(n23969), .A4(n23968), .ZN(
        n23989) );
  AOI22_X1 U27712 ( .A1(n30302), .A2(\xmem_data[88][4] ), .B1(n30193), .B2(
        \xmem_data[89][4] ), .ZN(n23976) );
  AOI22_X1 U27713 ( .A1(n27729), .A2(\xmem_data[90][4] ), .B1(n3121), .B2(
        \xmem_data[91][4] ), .ZN(n23975) );
  AOI22_X1 U27714 ( .A1(n3167), .A2(\xmem_data[92][4] ), .B1(n3188), .B2(
        \xmem_data[93][4] ), .ZN(n23974) );
  AND2_X1 U27715 ( .A1(n28232), .A2(\xmem_data[95][4] ), .ZN(n23972) );
  AOI21_X1 U27716 ( .B1(n30684), .B2(\xmem_data[94][4] ), .A(n23972), .ZN(
        n23973) );
  NAND4_X1 U27717 ( .A1(n23976), .A2(n23975), .A3(n23974), .A4(n23973), .ZN(
        n23987) );
  AOI22_X1 U27718 ( .A1(n27701), .A2(\xmem_data[80][4] ), .B1(n29798), .B2(
        \xmem_data[81][4] ), .ZN(n23980) );
  AOI22_X1 U27719 ( .A1(n27702), .A2(\xmem_data[82][4] ), .B1(n3147), .B2(
        \xmem_data[83][4] ), .ZN(n23979) );
  AOI22_X1 U27720 ( .A1(n30248), .A2(\xmem_data[84][4] ), .B1(n29589), .B2(
        \xmem_data[85][4] ), .ZN(n23978) );
  AOI22_X1 U27721 ( .A1(n26879), .A2(\xmem_data[86][4] ), .B1(n30508), .B2(
        \xmem_data[87][4] ), .ZN(n23977) );
  NAND4_X1 U27722 ( .A1(n23980), .A2(n23979), .A3(n23978), .A4(n23977), .ZN(
        n23986) );
  AOI22_X1 U27723 ( .A1(n29488), .A2(\xmem_data[64][4] ), .B1(n30716), .B2(
        \xmem_data[65][4] ), .ZN(n23984) );
  AOI22_X1 U27724 ( .A1(n27714), .A2(\xmem_data[66][4] ), .B1(n29246), .B2(
        \xmem_data[67][4] ), .ZN(n23983) );
  AOI22_X1 U27725 ( .A1(n27716), .A2(\xmem_data[68][4] ), .B1(n27715), .B2(
        \xmem_data[69][4] ), .ZN(n23982) );
  AOI22_X1 U27726 ( .A1(n27718), .A2(\xmem_data[70][4] ), .B1(n27717), .B2(
        \xmem_data[71][4] ), .ZN(n23981) );
  NAND4_X1 U27727 ( .A1(n23984), .A2(n23983), .A3(n23982), .A4(n23981), .ZN(
        n23985) );
  OR3_X1 U27728 ( .A1(n23987), .A2(n23986), .A3(n23985), .ZN(n23988) );
  OAI21_X1 U27729 ( .B1(n23989), .B2(n23988), .A(n27839), .ZN(n24012) );
  AOI22_X1 U27730 ( .A1(n28717), .A2(\xmem_data[8][4] ), .B1(n27743), .B2(
        \xmem_data[9][4] ), .ZN(n23993) );
  AOI22_X1 U27731 ( .A1(n27742), .A2(\xmem_data[10][4] ), .B1(n28245), .B2(
        \xmem_data[11][4] ), .ZN(n23992) );
  AOI22_X1 U27732 ( .A1(n27710), .A2(\xmem_data[12][4] ), .B1(n26616), .B2(
        \xmem_data[13][4] ), .ZN(n23991) );
  AOI22_X1 U27733 ( .A1(n30279), .A2(\xmem_data[14][4] ), .B1(n30278), .B2(
        \xmem_data[15][4] ), .ZN(n23990) );
  NAND4_X1 U27734 ( .A1(n23993), .A2(n23992), .A3(n23991), .A4(n23990), .ZN(
        n24009) );
  AOI22_X1 U27735 ( .A1(n27771), .A2(\xmem_data[16][4] ), .B1(n29708), .B2(
        \xmem_data[17][4] ), .ZN(n23997) );
  AOI22_X1 U27736 ( .A1(n3223), .A2(\xmem_data[18][4] ), .B1(n3146), .B2(
        \xmem_data[19][4] ), .ZN(n23996) );
  AOI22_X1 U27737 ( .A1(n28739), .A2(\xmem_data[20][4] ), .B1(n29704), .B2(
        \xmem_data[21][4] ), .ZN(n23995) );
  AOI22_X1 U27738 ( .A1(n29500), .A2(\xmem_data[22][4] ), .B1(n23762), .B2(
        \xmem_data[23][4] ), .ZN(n23994) );
  NAND4_X1 U27739 ( .A1(n23997), .A2(n23996), .A3(n23995), .A4(n23994), .ZN(
        n24008) );
  AOI22_X1 U27740 ( .A1(n3165), .A2(\xmem_data[28][4] ), .B1(n3184), .B2(
        \xmem_data[29][4] ), .ZN(n24001) );
  AOI22_X1 U27741 ( .A1(n27756), .A2(\xmem_data[26][4] ), .B1(n25672), .B2(
        \xmem_data[27][4] ), .ZN(n24000) );
  AOI22_X1 U27742 ( .A1(n28779), .A2(\xmem_data[24][4] ), .B1(n29648), .B2(
        \xmem_data[25][4] ), .ZN(n23999) );
  AOI22_X1 U27743 ( .A1(n28689), .A2(\xmem_data[30][4] ), .B1(n27825), .B2(
        \xmem_data[31][4] ), .ZN(n23998) );
  NAND4_X1 U27744 ( .A1(n24001), .A2(n24000), .A3(n23999), .A4(n23998), .ZN(
        n24007) );
  AOI22_X1 U27745 ( .A1(n29488), .A2(\xmem_data[0][4] ), .B1(n30170), .B2(
        \xmem_data[1][4] ), .ZN(n24005) );
  AOI22_X1 U27746 ( .A1(n27804), .A2(\xmem_data[2][4] ), .B1(n3151), .B2(
        \xmem_data[3][4] ), .ZN(n24004) );
  AOI22_X1 U27747 ( .A1(n29724), .A2(\xmem_data[4][4] ), .B1(n29462), .B2(
        \xmem_data[5][4] ), .ZN(n24003) );
  AOI22_X1 U27748 ( .A1(n27806), .A2(\xmem_data[6][4] ), .B1(n25407), .B2(
        \xmem_data[7][4] ), .ZN(n24002) );
  NAND4_X1 U27749 ( .A1(n24005), .A2(n24004), .A3(n24003), .A4(n24002), .ZN(
        n24006) );
  XNOR2_X1 U27750 ( .A(n31893), .B(\fmem_data[27][7] ), .ZN(n31936) );
  OAI22_X1 U27751 ( .A1(n35146), .A2(n35642), .B1(n31936), .B2(n35641), .ZN(
        n31780) );
  NAND2_X1 U27752 ( .A1(n25450), .A2(\xmem_data[15][2] ), .ZN(n24045) );
  AOI22_X1 U27753 ( .A1(n28337), .A2(\xmem_data[24][2] ), .B1(n29316), .B2(
        \xmem_data[25][2] ), .ZN(n24020) );
  AOI22_X1 U27754 ( .A1(n28754), .A2(\xmem_data[26][2] ), .B1(n24116), .B2(
        \xmem_data[27][2] ), .ZN(n24019) );
  AOI22_X1 U27755 ( .A1(n27974), .A2(\xmem_data[28][2] ), .B1(n21009), .B2(
        \xmem_data[29][2] ), .ZN(n24018) );
  AOI22_X1 U27756 ( .A1(n3329), .A2(\xmem_data[30][2] ), .B1(n27975), .B2(
        \xmem_data[31][2] ), .ZN(n24017) );
  NAND4_X1 U27757 ( .A1(n24020), .A2(n24019), .A3(n24018), .A4(n24017), .ZN(
        n24026) );
  AOI22_X1 U27758 ( .A1(n20734), .A2(\xmem_data[0][2] ), .B1(n27981), .B2(
        \xmem_data[1][2] ), .ZN(n24024) );
  AOI22_X1 U27759 ( .A1(n20985), .A2(\xmem_data[2][2] ), .B1(n17050), .B2(
        \xmem_data[3][2] ), .ZN(n24023) );
  AOI22_X1 U27760 ( .A1(n25630), .A2(\xmem_data[4][2] ), .B1(n21309), .B2(
        \xmem_data[5][2] ), .ZN(n24022) );
  AOI22_X1 U27761 ( .A1(n3449), .A2(\xmem_data[6][2] ), .B1(n25360), .B2(
        \xmem_data[7][2] ), .ZN(n24021) );
  NAND4_X1 U27762 ( .A1(n24024), .A2(n24023), .A3(n24022), .A4(n24021), .ZN(
        n24025) );
  OR2_X1 U27763 ( .A1(n24026), .A2(n24025), .ZN(n24042) );
  AOI22_X1 U27764 ( .A1(n20991), .A2(\xmem_data[8][2] ), .B1(n3217), .B2(
        \xmem_data[9][2] ), .ZN(n24027) );
  INV_X1 U27765 ( .A(n24027), .ZN(n24031) );
  AOI22_X1 U27766 ( .A1(n3340), .A2(\xmem_data[12][2] ), .B1(n27994), .B2(
        \xmem_data[13][2] ), .ZN(n24029) );
  NAND2_X1 U27767 ( .A1(n3128), .A2(\xmem_data[14][2] ), .ZN(n24028) );
  NAND2_X1 U27768 ( .A1(n24029), .A2(n24028), .ZN(n24030) );
  NOR2_X1 U27769 ( .A1(n24031), .A2(n24030), .ZN(n24040) );
  AOI22_X1 U27770 ( .A1(n20961), .A2(\xmem_data[16][2] ), .B1(n27988), .B2(
        \xmem_data[17][2] ), .ZN(n24035) );
  AOI22_X1 U27771 ( .A1(n24556), .A2(\xmem_data[18][2] ), .B1(n28416), .B2(
        \xmem_data[19][2] ), .ZN(n24034) );
  AOI22_X1 U27772 ( .A1(n27515), .A2(\xmem_data[20][2] ), .B1(n24160), .B2(
        \xmem_data[21][2] ), .ZN(n24033) );
  AOI22_X1 U27773 ( .A1(n17018), .A2(\xmem_data[22][2] ), .B1(n27989), .B2(
        \xmem_data[23][2] ), .ZN(n24032) );
  NAND4_X1 U27774 ( .A1(n24035), .A2(n24034), .A3(n24033), .A4(n24032), .ZN(
        n24038) );
  AOI22_X1 U27775 ( .A1(n27831), .A2(\xmem_data[10][2] ), .B1(n30534), .B2(
        \xmem_data[11][2] ), .ZN(n24036) );
  NAND2_X1 U27776 ( .A1(n24040), .A2(n24039), .ZN(n24041) );
  NOR2_X1 U27777 ( .A1(n24042), .A2(n24041), .ZN(n24044) );
  AOI21_X1 U27778 ( .B1(n24045), .B2(n24044), .A(n24043), .ZN(n24068) );
  AOI22_X1 U27779 ( .A1(n29325), .A2(\xmem_data[32][2] ), .B1(n20488), .B2(
        \xmem_data[33][2] ), .ZN(n24049) );
  AOI22_X1 U27780 ( .A1(n30901), .A2(\xmem_data[34][2] ), .B1(n25440), .B2(
        \xmem_data[35][2] ), .ZN(n24048) );
  AOI22_X1 U27781 ( .A1(n28076), .A2(\xmem_data[36][2] ), .B1(n28075), .B2(
        \xmem_data[37][2] ), .ZN(n24047) );
  AOI22_X1 U27782 ( .A1(n3434), .A2(\xmem_data[38][2] ), .B1(n3247), .B2(
        \xmem_data[39][2] ), .ZN(n24046) );
  NAND4_X1 U27783 ( .A1(n24049), .A2(n24048), .A3(n24047), .A4(n24046), .ZN(
        n24065) );
  AOI22_X1 U27784 ( .A1(n28082), .A2(\xmem_data[40][2] ), .B1(n3221), .B2(
        \xmem_data[41][2] ), .ZN(n24053) );
  AOI22_X1 U27785 ( .A1(n22708), .A2(\xmem_data[42][2] ), .B1(n30534), .B2(
        \xmem_data[43][2] ), .ZN(n24052) );
  AOI22_X1 U27786 ( .A1(n28083), .A2(\xmem_data[44][2] ), .B1(n22669), .B2(
        \xmem_data[45][2] ), .ZN(n24051) );
  AOI22_X1 U27787 ( .A1(n28084), .A2(\xmem_data[46][2] ), .B1(n25514), .B2(
        \xmem_data[47][2] ), .ZN(n24050) );
  NAND4_X1 U27788 ( .A1(n24053), .A2(n24052), .A3(n24051), .A4(n24050), .ZN(
        n24064) );
  AOI22_X1 U27789 ( .A1(n27551), .A2(\xmem_data[48][2] ), .B1(n13475), .B2(
        \xmem_data[49][2] ), .ZN(n24057) );
  AOI22_X1 U27790 ( .A1(n28089), .A2(\xmem_data[50][2] ), .B1(n29232), .B2(
        \xmem_data[51][2] ), .ZN(n24056) );
  AOI22_X1 U27791 ( .A1(n17041), .A2(\xmem_data[52][2] ), .B1(n28090), .B2(
        \xmem_data[53][2] ), .ZN(n24055) );
  AOI22_X1 U27792 ( .A1(n20776), .A2(\xmem_data[54][2] ), .B1(n27989), .B2(
        \xmem_data[55][2] ), .ZN(n24054) );
  NAND4_X1 U27793 ( .A1(n24057), .A2(n24056), .A3(n24055), .A4(n24054), .ZN(
        n24063) );
  AOI22_X1 U27794 ( .A1(n28096), .A2(\xmem_data[56][2] ), .B1(n22718), .B2(
        \xmem_data[57][2] ), .ZN(n24061) );
  AOI22_X1 U27795 ( .A1(n28302), .A2(\xmem_data[58][2] ), .B1(n28097), .B2(
        \xmem_data[59][2] ), .ZN(n24060) );
  AOI22_X1 U27796 ( .A1(n30956), .A2(\xmem_data[60][2] ), .B1(n28291), .B2(
        \xmem_data[61][2] ), .ZN(n24059) );
  AOI22_X1 U27797 ( .A1(n30686), .A2(\xmem_data[62][2] ), .B1(n28098), .B2(
        \xmem_data[63][2] ), .ZN(n24058) );
  NAND4_X1 U27798 ( .A1(n24061), .A2(n24060), .A3(n24059), .A4(n24058), .ZN(
        n24062) );
  OR4_X1 U27799 ( .A1(n24065), .A2(n24064), .A3(n24063), .A4(n24062), .ZN(
        n24066) );
  AND2_X1 U27800 ( .A1(n24066), .A2(n28107), .ZN(n24067) );
  NOR2_X1 U27801 ( .A1(n24068), .A2(n24067), .ZN(n31588) );
  AOI22_X1 U27802 ( .A1(n3171), .A2(\xmem_data[96][2] ), .B1(n23781), .B2(
        \xmem_data[97][2] ), .ZN(n24072) );
  AOI22_X1 U27803 ( .A1(n28036), .A2(\xmem_data[98][2] ), .B1(n28035), .B2(
        \xmem_data[99][2] ), .ZN(n24071) );
  AOI22_X1 U27804 ( .A1(n28038), .A2(\xmem_data[100][2] ), .B1(n28037), .B2(
        \xmem_data[101][2] ), .ZN(n24070) );
  AOI22_X1 U27805 ( .A1(n28039), .A2(\xmem_data[102][2] ), .B1(n28501), .B2(
        \xmem_data[103][2] ), .ZN(n24069) );
  NAND4_X1 U27806 ( .A1(n24072), .A2(n24071), .A3(n24070), .A4(n24069), .ZN(
        n24088) );
  AOI22_X1 U27807 ( .A1(n28044), .A2(\xmem_data[104][2] ), .B1(n3222), .B2(
        \xmem_data[105][2] ), .ZN(n24076) );
  AOI22_X1 U27808 ( .A1(n25414), .A2(\xmem_data[106][2] ), .B1(n24695), .B2(
        \xmem_data[107][2] ), .ZN(n24075) );
  AOI22_X1 U27809 ( .A1(n25617), .A2(\xmem_data[108][2] ), .B1(n28342), .B2(
        \xmem_data[109][2] ), .ZN(n24074) );
  AOI22_X1 U27810 ( .A1(n30710), .A2(\xmem_data[110][2] ), .B1(n28007), .B2(
        \xmem_data[111][2] ), .ZN(n24073) );
  NAND4_X1 U27811 ( .A1(n24076), .A2(n24075), .A3(n24074), .A4(n24073), .ZN(
        n24087) );
  AOI22_X1 U27812 ( .A1(n28050), .A2(\xmem_data[112][2] ), .B1(n27943), .B2(
        \xmem_data[113][2] ), .ZN(n24080) );
  AOI22_X1 U27813 ( .A1(n28051), .A2(\xmem_data[114][2] ), .B1(n24212), .B2(
        \xmem_data[115][2] ), .ZN(n24079) );
  AOI22_X1 U27814 ( .A1(n25425), .A2(\xmem_data[116][2] ), .B1(n28052), .B2(
        \xmem_data[117][2] ), .ZN(n24078) );
  AOI22_X1 U27815 ( .A1(n3158), .A2(\xmem_data[118][2] ), .B1(n3213), .B2(
        \xmem_data[119][2] ), .ZN(n24077) );
  NAND4_X1 U27816 ( .A1(n24080), .A2(n24079), .A3(n24078), .A4(n24077), .ZN(
        n24086) );
  AOI22_X1 U27817 ( .A1(n28059), .A2(\xmem_data[120][2] ), .B1(n28058), .B2(
        \xmem_data[121][2] ), .ZN(n24084) );
  AOI22_X1 U27818 ( .A1(n28781), .A2(\xmem_data[122][2] ), .B1(n21049), .B2(
        \xmem_data[123][2] ), .ZN(n24083) );
  AOI22_X1 U27819 ( .A1(n28061), .A2(\xmem_data[124][2] ), .B1(n28060), .B2(
        \xmem_data[125][2] ), .ZN(n24082) );
  AOI22_X1 U27820 ( .A1(n28226), .A2(\xmem_data[126][2] ), .B1(n28062), .B2(
        \xmem_data[127][2] ), .ZN(n24081) );
  NAND4_X1 U27821 ( .A1(n24084), .A2(n24083), .A3(n24082), .A4(n24081), .ZN(
        n24085) );
  OR4_X1 U27822 ( .A1(n24088), .A2(n24087), .A3(n24086), .A4(n24085), .ZN(
        n24110) );
  AOI22_X1 U27823 ( .A1(n3209), .A2(\xmem_data[64][2] ), .B1(n28328), .B2(
        \xmem_data[65][2] ), .ZN(n24092) );
  AOI22_X1 U27824 ( .A1(n28036), .A2(\xmem_data[66][2] ), .B1(n28035), .B2(
        \xmem_data[67][2] ), .ZN(n24091) );
  AOI22_X1 U27825 ( .A1(n28038), .A2(\xmem_data[68][2] ), .B1(n28037), .B2(
        \xmem_data[69][2] ), .ZN(n24090) );
  AOI22_X1 U27826 ( .A1(n28039), .A2(\xmem_data[70][2] ), .B1(n30863), .B2(
        \xmem_data[71][2] ), .ZN(n24089) );
  NAND4_X1 U27827 ( .A1(n24092), .A2(n24091), .A3(n24090), .A4(n24089), .ZN(
        n24108) );
  AOI22_X1 U27828 ( .A1(n28044), .A2(\xmem_data[72][2] ), .B1(n3221), .B2(
        \xmem_data[73][2] ), .ZN(n24096) );
  AOI22_X1 U27829 ( .A1(n28137), .A2(\xmem_data[74][2] ), .B1(n24207), .B2(
        \xmem_data[75][2] ), .ZN(n24095) );
  AOI22_X1 U27830 ( .A1(n17010), .A2(\xmem_data[76][2] ), .B1(n25616), .B2(
        \xmem_data[77][2] ), .ZN(n24094) );
  AOI22_X1 U27831 ( .A1(n24702), .A2(\xmem_data[78][2] ), .B1(n28343), .B2(
        \xmem_data[79][2] ), .ZN(n24093) );
  NAND4_X1 U27832 ( .A1(n24096), .A2(n24095), .A3(n24094), .A4(n24093), .ZN(
        n24107) );
  AOI22_X1 U27833 ( .A1(n28050), .A2(\xmem_data[80][2] ), .B1(n28415), .B2(
        \xmem_data[81][2] ), .ZN(n24100) );
  AOI22_X1 U27834 ( .A1(n28051), .A2(\xmem_data[82][2] ), .B1(n22740), .B2(
        \xmem_data[83][2] ), .ZN(n24099) );
  AOI22_X1 U27835 ( .A1(n20959), .A2(\xmem_data[84][2] ), .B1(n28052), .B2(
        \xmem_data[85][2] ), .ZN(n24098) );
  AOI22_X1 U27836 ( .A1(n3121), .A2(\xmem_data[86][2] ), .B1(n29279), .B2(
        \xmem_data[87][2] ), .ZN(n24097) );
  NAND4_X1 U27837 ( .A1(n24100), .A2(n24099), .A3(n24098), .A4(n24097), .ZN(
        n24106) );
  AOI22_X1 U27838 ( .A1(n28059), .A2(\xmem_data[88][2] ), .B1(n28058), .B2(
        \xmem_data[89][2] ), .ZN(n24104) );
  AOI22_X1 U27839 ( .A1(n29012), .A2(\xmem_data[90][2] ), .B1(n24510), .B2(
        \xmem_data[91][2] ), .ZN(n24103) );
  AOI22_X1 U27840 ( .A1(n28061), .A2(\xmem_data[92][2] ), .B1(n28060), .B2(
        \xmem_data[93][2] ), .ZN(n24102) );
  AOI22_X1 U27841 ( .A1(n29324), .A2(\xmem_data[94][2] ), .B1(n28062), .B2(
        \xmem_data[95][2] ), .ZN(n24101) );
  NAND4_X1 U27842 ( .A1(n24104), .A2(n24103), .A3(n24102), .A4(n24101), .ZN(
        n24105) );
  OR4_X1 U27843 ( .A1(n24108), .A2(n24107), .A3(n24106), .A4(n24105), .ZN(
        n24109) );
  AOI22_X1 U27844 ( .A1(n28071), .A2(n24110), .B1(n28033), .B2(n24109), .ZN(
        n31585) );
  NAND2_X1 U27845 ( .A1(n31588), .A2(n31585), .ZN(n32124) );
  XNOR2_X1 U27846 ( .A(n32124), .B(\fmem_data[22][7] ), .ZN(n31947) );
  XNOR2_X1 U27847 ( .A(n35316), .B(\fmem_data[15][3] ), .ZN(n33170) );
  XOR2_X1 U27848 ( .A(\fmem_data[15][2] ), .B(\fmem_data[15][3] ), .Z(n24113)
         );
  NOR2_X1 U27849 ( .A1(n30138), .A2(n3618), .ZN(n24434) );
  AOI22_X1 U27850 ( .A1(n29048), .A2(\xmem_data[16][7] ), .B1(n24115), .B2(
        \xmem_data[17][7] ), .ZN(n24121) );
  AOI22_X1 U27851 ( .A1(n24116), .A2(\xmem_data[18][7] ), .B1(n24190), .B2(
        \xmem_data[19][7] ), .ZN(n24120) );
  AOI22_X1 U27852 ( .A1(n24117), .A2(\xmem_data[20][7] ), .B1(n30269), .B2(
        \xmem_data[21][7] ), .ZN(n24119) );
  AOI22_X1 U27853 ( .A1(n20983), .A2(\xmem_data[22][7] ), .B1(n20782), .B2(
        \xmem_data[23][7] ), .ZN(n24118) );
  NAND4_X1 U27854 ( .A1(n24121), .A2(n24120), .A3(n24119), .A4(n24118), .ZN(
        n24129) );
  AOI22_X1 U27855 ( .A1(n28979), .A2(\xmem_data[24][7] ), .B1(n28241), .B2(
        \xmem_data[25][7] ), .ZN(n24127) );
  AOI22_X1 U27856 ( .A1(n24122), .A2(\xmem_data[26][7] ), .B1(n28354), .B2(
        \xmem_data[27][7] ), .ZN(n24126) );
  AOI22_X1 U27857 ( .A1(n20709), .A2(\xmem_data[28][7] ), .B1(n24693), .B2(
        \xmem_data[29][7] ), .ZN(n24125) );
  AND2_X1 U27858 ( .A1(n30589), .A2(\xmem_data[30][7] ), .ZN(n24123) );
  AOI21_X1 U27859 ( .B1(n27439), .B2(\xmem_data[31][7] ), .A(n24123), .ZN(
        n24124) );
  NAND4_X1 U27860 ( .A1(n24127), .A2(n24126), .A3(n24125), .A4(n24124), .ZN(
        n24128) );
  OR2_X1 U27861 ( .A1(n24129), .A2(n24128), .ZN(n24150) );
  AOI22_X1 U27862 ( .A1(n24130), .A2(\xmem_data[8][7] ), .B1(n27763), .B2(
        \xmem_data[9][7] ), .ZN(n24138) );
  AOI22_X1 U27863 ( .A1(n24132), .A2(\xmem_data[10][7] ), .B1(n28980), .B2(
        \xmem_data[11][7] ), .ZN(n24137) );
  AOI22_X1 U27864 ( .A1(n22703), .A2(\xmem_data[12][7] ), .B1(n30543), .B2(
        \xmem_data[13][7] ), .ZN(n24136) );
  AOI22_X1 U27865 ( .A1(n24134), .A2(\xmem_data[14][7] ), .B1(n24133), .B2(
        \xmem_data[15][7] ), .ZN(n24135) );
  NAND4_X1 U27866 ( .A1(n24138), .A2(n24137), .A3(n24136), .A4(n24135), .ZN(
        n24148) );
  AOI22_X1 U27867 ( .A1(n3217), .A2(\xmem_data[0][7] ), .B1(n24139), .B2(
        \xmem_data[1][7] ), .ZN(n24144) );
  AOI22_X1 U27868 ( .A1(n24140), .A2(\xmem_data[4][7] ), .B1(n3126), .B2(
        \xmem_data[5][7] ), .ZN(n24143) );
  AOI22_X1 U27869 ( .A1(n28508), .A2(\xmem_data[2][7] ), .B1(n24141), .B2(
        \xmem_data[3][7] ), .ZN(n24142) );
  NAND3_X1 U27870 ( .A1(n24144), .A2(n24143), .A3(n24142), .ZN(n24147) );
  AND2_X1 U27871 ( .A1(n23813), .A2(\xmem_data[7][7] ), .ZN(n24145) );
  NOR2_X1 U27872 ( .A1(n24150), .A2(n24149), .ZN(n24152) );
  OR2_X1 U27873 ( .A1(n24152), .A2(n24151), .ZN(n24240) );
  AOI22_X1 U27874 ( .A1(n3218), .A2(\xmem_data[96][7] ), .B1(n20724), .B2(
        \xmem_data[97][7] ), .ZN(n24156) );
  AOI22_X1 U27875 ( .A1(n20598), .A2(\xmem_data[98][7] ), .B1(n24697), .B2(
        \xmem_data[99][7] ), .ZN(n24155) );
  AOI22_X1 U27876 ( .A1(n13444), .A2(\xmem_data[100][7] ), .B1(n3135), .B2(
        \xmem_data[101][7] ), .ZN(n24154) );
  AOI22_X1 U27877 ( .A1(n25514), .A2(\xmem_data[102][7] ), .B1(n28374), .B2(
        \xmem_data[103][7] ), .ZN(n24153) );
  NAND4_X1 U27878 ( .A1(n24156), .A2(n24155), .A3(n24154), .A4(n24153), .ZN(
        n24180) );
  AOI22_X1 U27879 ( .A1(n24158), .A2(\xmem_data[104][7] ), .B1(n24157), .B2(
        \xmem_data[105][7] ), .ZN(n24164) );
  AOI22_X1 U27880 ( .A1(n24159), .A2(\xmem_data[106][7] ), .B1(n30514), .B2(
        \xmem_data[107][7] ), .ZN(n24163) );
  AOI22_X1 U27881 ( .A1(n24160), .A2(\xmem_data[108][7] ), .B1(n30543), .B2(
        \xmem_data[109][7] ), .ZN(n24162) );
  AOI22_X1 U27882 ( .A1(n3212), .A2(\xmem_data[110][7] ), .B1(n29010), .B2(
        \xmem_data[111][7] ), .ZN(n24161) );
  NAND4_X1 U27883 ( .A1(n24164), .A2(n24163), .A3(n24162), .A4(n24161), .ZN(
        n24179) );
  AOI22_X1 U27884 ( .A1(n30544), .A2(\xmem_data[112][7] ), .B1(n17044), .B2(
        \xmem_data[113][7] ), .ZN(n24171) );
  AOI22_X1 U27885 ( .A1(n24165), .A2(\xmem_data[114][7] ), .B1(n20593), .B2(
        \xmem_data[115][7] ), .ZN(n24170) );
  AOI22_X1 U27886 ( .A1(n28429), .A2(\xmem_data[116][7] ), .B1(n3300), .B2(
        \xmem_data[117][7] ), .ZN(n24169) );
  AOI22_X1 U27887 ( .A1(n24167), .A2(\xmem_data[118][7] ), .B1(n24166), .B2(
        \xmem_data[119][7] ), .ZN(n24168) );
  NAND4_X1 U27888 ( .A1(n24171), .A2(n24170), .A3(n24169), .A4(n24168), .ZN(
        n24178) );
  AOI22_X1 U27889 ( .A1(n23781), .A2(\xmem_data[120][7] ), .B1(n27568), .B2(
        \xmem_data[121][7] ), .ZN(n24176) );
  AOI22_X1 U27890 ( .A1(n20707), .A2(\xmem_data[122][7] ), .B1(n27959), .B2(
        \xmem_data[123][7] ), .ZN(n24175) );
  AOI22_X1 U27891 ( .A1(n25685), .A2(\xmem_data[124][7] ), .B1(n25725), .B2(
        \xmem_data[125][7] ), .ZN(n24174) );
  AOI22_X1 U27892 ( .A1(n24172), .A2(\xmem_data[126][7] ), .B1(n31348), .B2(
        \xmem_data[127][7] ), .ZN(n24173) );
  NAND4_X1 U27893 ( .A1(n24176), .A2(n24175), .A3(n24174), .A4(n24173), .ZN(
        n24177) );
  OR4_X1 U27894 ( .A1(n24180), .A2(n24179), .A3(n24178), .A4(n24177), .ZN(
        n24206) );
  AOI22_X1 U27895 ( .A1(n29017), .A2(\xmem_data[88][7] ), .B1(n29298), .B2(
        \xmem_data[89][7] ), .ZN(n24185) );
  AOI22_X1 U27896 ( .A1(n31344), .A2(\xmem_data[90][7] ), .B1(n25408), .B2(
        \xmem_data[91][7] ), .ZN(n24184) );
  AOI22_X1 U27897 ( .A1(n24573), .A2(\xmem_data[92][7] ), .B1(n3317), .B2(
        \xmem_data[93][7] ), .ZN(n24183) );
  AND2_X1 U27898 ( .A1(n24439), .A2(\xmem_data[94][7] ), .ZN(n24181) );
  AOI21_X1 U27899 ( .B1(n25730), .B2(\xmem_data[95][7] ), .A(n24181), .ZN(
        n24182) );
  NAND4_X1 U27900 ( .A1(n24185), .A2(n24184), .A3(n24183), .A4(n24182), .ZN(
        n24202) );
  AOI22_X1 U27901 ( .A1(n3358), .A2(\xmem_data[72][7] ), .B1(n17064), .B2(
        \xmem_data[73][7] ), .ZN(n24189) );
  AOI22_X1 U27902 ( .A1(n24212), .A2(\xmem_data[74][7] ), .B1(n20541), .B2(
        \xmem_data[75][7] ), .ZN(n24188) );
  AOI22_X1 U27903 ( .A1(n25382), .A2(\xmem_data[76][7] ), .B1(n30746), .B2(
        \xmem_data[77][7] ), .ZN(n24187) );
  AOI22_X1 U27904 ( .A1(n31269), .A2(\xmem_data[78][7] ), .B1(n24214), .B2(
        \xmem_data[79][7] ), .ZN(n24186) );
  NAND4_X1 U27905 ( .A1(n24189), .A2(n24188), .A3(n24187), .A4(n24186), .ZN(
        n24201) );
  AOI22_X1 U27906 ( .A1(n24219), .A2(\xmem_data[80][7] ), .B1(n23777), .B2(
        \xmem_data[81][7] ), .ZN(n24194) );
  AOI22_X1 U27907 ( .A1(n24221), .A2(\xmem_data[82][7] ), .B1(n24190), .B2(
        \xmem_data[83][7] ), .ZN(n24193) );
  AOI22_X1 U27908 ( .A1(n24222), .A2(\xmem_data[84][7] ), .B1(n3337), .B2(
        \xmem_data[85][7] ), .ZN(n24192) );
  AOI22_X1 U27909 ( .A1(n24223), .A2(\xmem_data[86][7] ), .B1(n29325), .B2(
        \xmem_data[87][7] ), .ZN(n24191) );
  NAND4_X1 U27910 ( .A1(n24194), .A2(n24193), .A3(n24192), .A4(n24191), .ZN(
        n24200) );
  AOI22_X1 U27911 ( .A1(n3218), .A2(\xmem_data[64][7] ), .B1(n21067), .B2(
        \xmem_data[65][7] ), .ZN(n24198) );
  AOI22_X1 U27912 ( .A1(n24207), .A2(\xmem_data[66][7] ), .B1(n20969), .B2(
        \xmem_data[67][7] ), .ZN(n24197) );
  AOI22_X1 U27913 ( .A1(n23811), .A2(\xmem_data[68][7] ), .B1(n21074), .B2(
        \xmem_data[69][7] ), .ZN(n24196) );
  AOI22_X1 U27914 ( .A1(n28045), .A2(\xmem_data[70][7] ), .B1(n25604), .B2(
        \xmem_data[71][7] ), .ZN(n24195) );
  NAND4_X1 U27915 ( .A1(n24198), .A2(n24197), .A3(n24196), .A4(n24195), .ZN(
        n24199) );
  OR4_X1 U27916 ( .A1(n24202), .A2(n24201), .A3(n24200), .A4(n24199), .ZN(
        n24203) );
  AOI22_X1 U27917 ( .A1(n24206), .A2(n24205), .B1(n24204), .B2(n24203), .ZN(
        n24239) );
  AOI22_X1 U27918 ( .A1(n3219), .A2(\xmem_data[32][7] ), .B1(n27708), .B2(
        \xmem_data[33][7] ), .ZN(n24211) );
  AOI22_X1 U27919 ( .A1(n24207), .A2(\xmem_data[34][7] ), .B1(n3322), .B2(
        \xmem_data[35][7] ), .ZN(n24210) );
  AOI22_X1 U27920 ( .A1(n3256), .A2(\xmem_data[36][7] ), .B1(n3126), .B2(
        \xmem_data[37][7] ), .ZN(n24209) );
  AOI22_X1 U27921 ( .A1(n28007), .A2(\xmem_data[38][7] ), .B1(n25604), .B2(
        \xmem_data[39][7] ), .ZN(n24208) );
  NAND4_X1 U27922 ( .A1(n24211), .A2(n24210), .A3(n24209), .A4(n24208), .ZN(
        n24235) );
  AOI22_X1 U27923 ( .A1(n27863), .A2(\xmem_data[40][7] ), .B1(n31353), .B2(
        \xmem_data[41][7] ), .ZN(n24218) );
  AOI22_X1 U27924 ( .A1(n24212), .A2(\xmem_data[42][7] ), .B1(n30514), .B2(
        \xmem_data[43][7] ), .ZN(n24217) );
  AOI22_X1 U27925 ( .A1(n25709), .A2(\xmem_data[44][7] ), .B1(n27945), .B2(
        \xmem_data[45][7] ), .ZN(n24216) );
  AOI22_X1 U27926 ( .A1(n3213), .A2(\xmem_data[46][7] ), .B1(n24214), .B2(
        \xmem_data[47][7] ), .ZN(n24215) );
  NAND4_X1 U27927 ( .A1(n24218), .A2(n24217), .A3(n24216), .A4(n24215), .ZN(
        n24234) );
  AOI22_X1 U27928 ( .A1(n24219), .A2(\xmem_data[48][7] ), .B1(n27825), .B2(
        \xmem_data[49][7] ), .ZN(n24227) );
  AOI22_X1 U27929 ( .A1(n24221), .A2(\xmem_data[50][7] ), .B1(n25717), .B2(
        \xmem_data[51][7] ), .ZN(n24226) );
  AOI22_X1 U27930 ( .A1(n24222), .A2(\xmem_data[52][7] ), .B1(n17004), .B2(
        \xmem_data[53][7] ), .ZN(n24225) );
  AOI22_X1 U27931 ( .A1(n24223), .A2(\xmem_data[54][7] ), .B1(n3179), .B2(
        \xmem_data[55][7] ), .ZN(n24224) );
  NAND4_X1 U27932 ( .A1(n24227), .A2(n24226), .A3(n24225), .A4(n24224), .ZN(
        n24233) );
  AOI22_X1 U27933 ( .A1(n17049), .A2(\xmem_data[56][7] ), .B1(n27568), .B2(
        \xmem_data[57][7] ), .ZN(n24231) );
  AOI22_X1 U27934 ( .A1(n24686), .A2(\xmem_data[58][7] ), .B1(n27500), .B2(
        \xmem_data[59][7] ), .ZN(n24230) );
  AOI22_X1 U27935 ( .A1(n28075), .A2(\xmem_data[60][7] ), .B1(n3305), .B2(
        \xmem_data[61][7] ), .ZN(n24229) );
  AOI22_X1 U27936 ( .A1(n25360), .A2(\xmem_data[62][7] ), .B1(n20991), .B2(
        \xmem_data[63][7] ), .ZN(n24228) );
  NAND4_X1 U27937 ( .A1(n24231), .A2(n24230), .A3(n24229), .A4(n24228), .ZN(
        n24232) );
  OR4_X1 U27938 ( .A1(n24235), .A2(n24234), .A3(n24233), .A4(n24232), .ZN(
        n24237) );
  NAND2_X1 U27939 ( .A1(n24237), .A2(n24236), .ZN(n24238) );
  AOI22_X1 U27940 ( .A1(n30964), .A2(\xmem_data[32][2] ), .B1(n23739), .B2(
        \xmem_data[33][2] ), .ZN(n24244) );
  AOI22_X1 U27941 ( .A1(n24534), .A2(\xmem_data[34][2] ), .B1(n28372), .B2(
        \xmem_data[35][2] ), .ZN(n24243) );
  AOI22_X1 U27942 ( .A1(n25451), .A2(\xmem_data[36][2] ), .B1(n24657), .B2(
        \xmem_data[37][2] ), .ZN(n24242) );
  AOI22_X1 U27943 ( .A1(n31321), .A2(\xmem_data[38][2] ), .B1(n3358), .B2(
        \xmem_data[39][2] ), .ZN(n24241) );
  NAND4_X1 U27944 ( .A1(n24244), .A2(n24243), .A3(n24242), .A4(n24241), .ZN(
        n24260) );
  AOI22_X1 U27945 ( .A1(n31327), .A2(\xmem_data[40][2] ), .B1(n31326), .B2(
        \xmem_data[41][2] ), .ZN(n24248) );
  AOI22_X1 U27946 ( .A1(n20959), .A2(\xmem_data[42][2] ), .B1(n25671), .B2(
        \xmem_data[43][2] ), .ZN(n24247) );
  AOI22_X1 U27947 ( .A1(n31328), .A2(\xmem_data[44][2] ), .B1(n31269), .B2(
        \xmem_data[45][2] ), .ZN(n24246) );
  AOI22_X1 U27948 ( .A1(n31330), .A2(\xmem_data[46][2] ), .B1(n31329), .B2(
        \xmem_data[47][2] ), .ZN(n24245) );
  NAND4_X1 U27949 ( .A1(n24248), .A2(n24247), .A3(n24246), .A4(n24245), .ZN(
        n24259) );
  AOI22_X1 U27950 ( .A1(n24710), .A2(\xmem_data[48][2] ), .B1(n29190), .B2(
        \xmem_data[49][2] ), .ZN(n24252) );
  AOI22_X1 U27951 ( .A1(n24220), .A2(\xmem_data[50][2] ), .B1(n25581), .B2(
        \xmem_data[51][2] ), .ZN(n24251) );
  AOI22_X1 U27952 ( .A1(n31315), .A2(\xmem_data[52][2] ), .B1(n31314), .B2(
        \xmem_data[53][2] ), .ZN(n24250) );
  AOI22_X1 U27953 ( .A1(n31316), .A2(\xmem_data[54][2] ), .B1(n11008), .B2(
        \xmem_data[55][2] ), .ZN(n24249) );
  NAND4_X1 U27954 ( .A1(n24252), .A2(n24251), .A3(n24250), .A4(n24249), .ZN(
        n24258) );
  AOI22_X1 U27955 ( .A1(n31308), .A2(\xmem_data[56][2] ), .B1(n20769), .B2(
        \xmem_data[57][2] ), .ZN(n24256) );
  AOI22_X1 U27956 ( .A1(n27959), .A2(\xmem_data[58][2] ), .B1(n31309), .B2(
        \xmem_data[59][2] ), .ZN(n24255) );
  AOI22_X1 U27957 ( .A1(n3332), .A2(\xmem_data[60][2] ), .B1(n25485), .B2(
        \xmem_data[61][2] ), .ZN(n24254) );
  AOI22_X1 U27958 ( .A1(n28364), .A2(\xmem_data[62][2] ), .B1(n3218), .B2(
        \xmem_data[63][2] ), .ZN(n24253) );
  NAND4_X1 U27959 ( .A1(n24256), .A2(n24255), .A3(n24254), .A4(n24253), .ZN(
        n24257) );
  OR4_X1 U27960 ( .A1(n24260), .A2(n24259), .A3(n24258), .A4(n24257), .ZN(
        n24261) );
  AND2_X1 U27961 ( .A1(n24261), .A2(n31340), .ZN(n24290) );
  AOI22_X1 U27962 ( .A1(n30608), .A2(\xmem_data[8][2] ), .B1(n29232), .B2(
        \xmem_data[9][2] ), .ZN(n24265) );
  AOI22_X1 U27963 ( .A1(n31268), .A2(\xmem_data[10][2] ), .B1(n23715), .B2(
        \xmem_data[11][2] ), .ZN(n24264) );
  AOI22_X1 U27964 ( .A1(n28752), .A2(\xmem_data[12][2] ), .B1(n31269), .B2(
        \xmem_data[13][2] ), .ZN(n24263) );
  AOI22_X1 U27965 ( .A1(n28096), .A2(\xmem_data[14][2] ), .B1(n31270), .B2(
        \xmem_data[15][2] ), .ZN(n24262) );
  AOI22_X1 U27966 ( .A1(n31255), .A2(\xmem_data[16][2] ), .B1(n31254), .B2(
        \xmem_data[17][2] ), .ZN(n24269) );
  AOI22_X1 U27967 ( .A1(n3205), .A2(\xmem_data[18][2] ), .B1(n25364), .B2(
        \xmem_data[19][2] ), .ZN(n24268) );
  AOI22_X1 U27968 ( .A1(n23780), .A2(\xmem_data[20][2] ), .B1(n24622), .B2(
        \xmem_data[21][2] ), .ZN(n24267) );
  AOI22_X1 U27969 ( .A1(n29325), .A2(\xmem_data[22][2] ), .B1(n31256), .B2(
        \xmem_data[23][2] ), .ZN(n24266) );
  NAND2_X1 U27970 ( .A1(n25450), .A2(\xmem_data[5][2] ), .ZN(n24270) );
  AOI22_X1 U27971 ( .A1(n29494), .A2(\xmem_data[0][2] ), .B1(n20500), .B2(
        \xmem_data[1][2] ), .ZN(n24274) );
  AOI22_X1 U27972 ( .A1(n31276), .A2(\xmem_data[6][2] ), .B1(n27943), .B2(
        \xmem_data[7][2] ), .ZN(n24273) );
  AOI22_X1 U27973 ( .A1(n25416), .A2(\xmem_data[2][2] ), .B1(n31275), .B2(
        \xmem_data[3][2] ), .ZN(n24272) );
  NAND3_X1 U27974 ( .A1(n24274), .A2(n24273), .A3(n24272), .ZN(n24276) );
  AND2_X1 U27975 ( .A1(n29350), .A2(\xmem_data[4][2] ), .ZN(n24275) );
  NOR2_X1 U27976 ( .A1(n24277), .A2(n4004), .ZN(n24288) );
  AOI22_X1 U27977 ( .A1(n29657), .A2(\xmem_data[24][2] ), .B1(n31261), .B2(
        \xmem_data[25][2] ), .ZN(n24279) );
  AOI22_X1 U27978 ( .A1(n28164), .A2(\xmem_data[28][2] ), .B1(n30589), .B2(
        \xmem_data[29][2] ), .ZN(n24278) );
  NAND2_X1 U27979 ( .A1(n24279), .A2(n24278), .ZN(n24286) );
  AND2_X1 U27980 ( .A1(n27502), .A2(\xmem_data[30][2] ), .ZN(n24285) );
  NAND2_X1 U27981 ( .A1(n3219), .A2(\xmem_data[31][2] ), .ZN(n24281) );
  NAND2_X1 U27982 ( .A1(n3380), .A2(\xmem_data[26][2] ), .ZN(n24280) );
  NAND2_X1 U27983 ( .A1(n24281), .A2(n24280), .ZN(n24282) );
  AOI21_X1 U27984 ( .B1(n31262), .B2(\xmem_data[27][2] ), .A(n24282), .ZN(
        n24283) );
  INV_X1 U27985 ( .A(n24283), .ZN(n24284) );
  NOR3_X1 U27986 ( .A1(n24286), .A2(n24285), .A3(n24284), .ZN(n24287) );
  AOI21_X1 U27987 ( .B1(n24288), .B2(n24287), .A(n31041), .ZN(n24289) );
  NOR2_X1 U27988 ( .A1(n24290), .A2(n24289), .ZN(n24334) );
  AOI22_X1 U27989 ( .A1(n31368), .A2(\xmem_data[64][2] ), .B1(n31367), .B2(
        \xmem_data[65][2] ), .ZN(n24294) );
  AOI22_X1 U27990 ( .A1(n24697), .A2(\xmem_data[66][2] ), .B1(n14890), .B2(
        \xmem_data[67][2] ), .ZN(n24293) );
  AOI22_X1 U27991 ( .A1(n28344), .A2(\xmem_data[68][2] ), .B1(n29045), .B2(
        \xmem_data[69][2] ), .ZN(n24292) );
  AOI22_X1 U27992 ( .A1(n23813), .A2(\xmem_data[70][2] ), .B1(n3358), .B2(
        \xmem_data[71][2] ), .ZN(n24291) );
  NAND4_X1 U27993 ( .A1(n24294), .A2(n24293), .A3(n24292), .A4(n24291), .ZN(
        n24310) );
  AOI22_X1 U27994 ( .A1(n31353), .A2(\xmem_data[72][2] ), .B1(n29232), .B2(
        \xmem_data[73][2] ), .ZN(n24298) );
  AOI22_X1 U27995 ( .A1(n28298), .A2(\xmem_data[74][2] ), .B1(n20544), .B2(
        \xmem_data[75][2] ), .ZN(n24297) );
  AOI22_X1 U27996 ( .A1(n3120), .A2(\xmem_data[76][2] ), .B1(n29188), .B2(
        \xmem_data[77][2] ), .ZN(n24296) );
  AOI22_X1 U27997 ( .A1(n28337), .A2(\xmem_data[78][2] ), .B1(n31355), .B2(
        \xmem_data[79][2] ), .ZN(n24295) );
  NAND4_X1 U27998 ( .A1(n24298), .A2(n24297), .A3(n24296), .A4(n24295), .ZN(
        n24309) );
  AOI22_X1 U27999 ( .A1(n17021), .A2(\xmem_data[80][2] ), .B1(n31360), .B2(
        \xmem_data[81][2] ), .ZN(n24302) );
  AOI22_X1 U28000 ( .A1(n24647), .A2(\xmem_data[82][2] ), .B1(n31361), .B2(
        \xmem_data[83][2] ), .ZN(n24301) );
  AOI22_X1 U28001 ( .A1(n29573), .A2(\xmem_data[84][2] ), .B1(n31362), .B2(
        \xmem_data[85][2] ), .ZN(n24300) );
  AOI22_X1 U28002 ( .A1(n24685), .A2(\xmem_data[86][2] ), .B1(n28468), .B2(
        \xmem_data[87][2] ), .ZN(n24299) );
  NAND4_X1 U28003 ( .A1(n24302), .A2(n24301), .A3(n24300), .A4(n24299), .ZN(
        n24308) );
  AOI22_X1 U28004 ( .A1(n31345), .A2(\xmem_data[88][2] ), .B1(n31344), .B2(
        \xmem_data[89][2] ), .ZN(n24306) );
  AOI22_X1 U28005 ( .A1(n25358), .A2(\xmem_data[90][2] ), .B1(n31346), .B2(
        \xmem_data[91][2] ), .ZN(n24305) );
  AOI22_X1 U28006 ( .A1(n3414), .A2(\xmem_data[92][2] ), .B1(n31347), .B2(
        \xmem_data[93][2] ), .ZN(n24304) );
  AOI22_X1 U28007 ( .A1(n31348), .A2(\xmem_data[94][2] ), .B1(n3218), .B2(
        \xmem_data[95][2] ), .ZN(n24303) );
  NAND4_X1 U28008 ( .A1(n24306), .A2(n24305), .A3(n24304), .A4(n24303), .ZN(
        n24307) );
  OR4_X1 U28009 ( .A1(n24310), .A2(n24309), .A3(n24308), .A4(n24307), .ZN(
        n24332) );
  AOI22_X1 U28010 ( .A1(n31368), .A2(\xmem_data[96][2] ), .B1(n31367), .B2(
        \xmem_data[97][2] ), .ZN(n24314) );
  AOI22_X1 U28011 ( .A1(n25694), .A2(\xmem_data[98][2] ), .B1(n20806), .B2(
        \xmem_data[99][2] ), .ZN(n24313) );
  AOI22_X1 U28012 ( .A1(n3135), .A2(\xmem_data[100][2] ), .B1(n24657), .B2(
        \xmem_data[101][2] ), .ZN(n24312) );
  AOI22_X1 U28013 ( .A1(n28050), .A2(\xmem_data[102][2] ), .B1(n29180), .B2(
        \xmem_data[103][2] ), .ZN(n24311) );
  NAND4_X1 U28014 ( .A1(n24314), .A2(n24313), .A3(n24312), .A4(n24311), .ZN(
        n24330) );
  AOI22_X1 U28015 ( .A1(n31353), .A2(\xmem_data[104][2] ), .B1(n24516), .B2(
        \xmem_data[105][2] ), .ZN(n24318) );
  AOI22_X1 U28016 ( .A1(n25425), .A2(\xmem_data[106][2] ), .B1(n25606), .B2(
        \xmem_data[107][2] ), .ZN(n24317) );
  AOI22_X1 U28017 ( .A1(n3466), .A2(\xmem_data[108][2] ), .B1(n27989), .B2(
        \xmem_data[109][2] ), .ZN(n24316) );
  AOI22_X1 U28018 ( .A1(n21007), .A2(\xmem_data[110][2] ), .B1(n31355), .B2(
        \xmem_data[111][2] ), .ZN(n24315) );
  NAND4_X1 U28019 ( .A1(n24318), .A2(n24317), .A3(n24316), .A4(n24315), .ZN(
        n24329) );
  AOI22_X1 U28020 ( .A1(n30872), .A2(\xmem_data[112][2] ), .B1(n31360), .B2(
        \xmem_data[113][2] ), .ZN(n24322) );
  AOI22_X1 U28021 ( .A1(n24511), .A2(\xmem_data[114][2] ), .B1(n31361), .B2(
        \xmem_data[115][2] ), .ZN(n24321) );
  AOI22_X1 U28022 ( .A1(n30645), .A2(\xmem_data[116][2] ), .B1(n31362), .B2(
        \xmem_data[117][2] ), .ZN(n24320) );
  AOI22_X1 U28023 ( .A1(n3179), .A2(\xmem_data[118][2] ), .B1(n28328), .B2(
        \xmem_data[119][2] ), .ZN(n24319) );
  NAND4_X1 U28024 ( .A1(n24322), .A2(n24321), .A3(n24320), .A4(n24319), .ZN(
        n24328) );
  AOI22_X1 U28025 ( .A1(n31345), .A2(\xmem_data[120][2] ), .B1(n31344), .B2(
        \xmem_data[121][2] ), .ZN(n24326) );
  AOI22_X1 U28026 ( .A1(n17030), .A2(\xmem_data[122][2] ), .B1(n31346), .B2(
        \xmem_data[123][2] ), .ZN(n24325) );
  AOI22_X1 U28027 ( .A1(n20828), .A2(\xmem_data[124][2] ), .B1(n31347), .B2(
        \xmem_data[125][2] ), .ZN(n24324) );
  AOI22_X1 U28028 ( .A1(n31348), .A2(\xmem_data[126][2] ), .B1(n3219), .B2(
        \xmem_data[127][2] ), .ZN(n24323) );
  NAND4_X1 U28029 ( .A1(n24326), .A2(n24325), .A3(n24324), .A4(n24323), .ZN(
        n24327) );
  OR4_X1 U28030 ( .A1(n24330), .A2(n24329), .A3(n24328), .A4(n24327), .ZN(
        n24331) );
  XNOR2_X1 U28031 ( .A(n32235), .B(\fmem_data[12][7] ), .ZN(n33182) );
  AOI22_X1 U28032 ( .A1(n25561), .A2(\xmem_data[32][2] ), .B1(n3306), .B2(
        \xmem_data[33][2] ), .ZN(n24339) );
  AOI22_X1 U28033 ( .A1(n31347), .A2(\xmem_data[34][2] ), .B1(n25508), .B2(
        \xmem_data[35][2] ), .ZN(n24338) );
  AOI22_X1 U28034 ( .A1(n3221), .A2(\xmem_data[36][2] ), .B1(n25414), .B2(
        \xmem_data[37][2] ), .ZN(n24337) );
  AOI22_X1 U28035 ( .A1(n25562), .A2(\xmem_data[38][2] ), .B1(n3342), .B2(
        \xmem_data[39][2] ), .ZN(n24336) );
  NAND4_X1 U28036 ( .A1(n24339), .A2(n24338), .A3(n24337), .A4(n24336), .ZN(
        n24355) );
  AOI22_X1 U28037 ( .A1(n20806), .A2(\xmem_data[40][2] ), .B1(n3147), .B2(
        \xmem_data[41][2] ), .ZN(n24343) );
  AOI22_X1 U28038 ( .A1(n28007), .A2(\xmem_data[42][2] ), .B1(n30885), .B2(
        \xmem_data[43][2] ), .ZN(n24342) );
  AOI22_X1 U28039 ( .A1(n3357), .A2(\xmem_data[44][2] ), .B1(n28743), .B2(
        \xmem_data[45][2] ), .ZN(n24341) );
  AOI22_X1 U28040 ( .A1(n14998), .A2(\xmem_data[46][2] ), .B1(n25567), .B2(
        \xmem_data[47][2] ), .ZN(n24340) );
  NAND4_X1 U28041 ( .A1(n24343), .A2(n24342), .A3(n24341), .A4(n24340), .ZN(
        n24354) );
  AOI22_X1 U28042 ( .A1(n29271), .A2(\xmem_data[48][2] ), .B1(n3120), .B2(
        \xmem_data[49][2] ), .ZN(n24347) );
  AOI22_X1 U28043 ( .A1(n25574), .A2(\xmem_data[50][2] ), .B1(n25573), .B2(
        \xmem_data[51][2] ), .ZN(n24346) );
  AOI22_X1 U28044 ( .A1(n14970), .A2(\xmem_data[52][2] ), .B1(n20815), .B2(
        \xmem_data[53][2] ), .ZN(n24345) );
  AOI22_X1 U28045 ( .A1(n25576), .A2(\xmem_data[54][2] ), .B1(n25575), .B2(
        \xmem_data[55][2] ), .ZN(n24344) );
  NAND4_X1 U28046 ( .A1(n24347), .A2(n24346), .A3(n24345), .A4(n24344), .ZN(
        n24353) );
  AOI22_X1 U28047 ( .A1(n14882), .A2(\xmem_data[56][2] ), .B1(n28461), .B2(
        \xmem_data[57][2] ), .ZN(n24351) );
  AOI22_X1 U28048 ( .A1(n25583), .A2(\xmem_data[58][2] ), .B1(n25582), .B2(
        \xmem_data[59][2] ), .ZN(n24350) );
  AOI22_X1 U28049 ( .A1(n27526), .A2(\xmem_data[60][2] ), .B1(n25584), .B2(
        \xmem_data[61][2] ), .ZN(n24349) );
  AOI22_X1 U28050 ( .A1(n29326), .A2(\xmem_data[62][2] ), .B1(n27500), .B2(
        \xmem_data[63][2] ), .ZN(n24348) );
  NAND4_X1 U28051 ( .A1(n24351), .A2(n24350), .A3(n24349), .A4(n24348), .ZN(
        n24352) );
  OR4_X1 U28052 ( .A1(n24355), .A2(n24354), .A3(n24353), .A4(n24352), .ZN(
        n24385) );
  AOI22_X1 U28053 ( .A1(n25481), .A2(\xmem_data[12][2] ), .B1(n27763), .B2(
        \xmem_data[13][2] ), .ZN(n24362) );
  AOI22_X1 U28054 ( .A1(n25486), .A2(\xmem_data[8][2] ), .B1(n21074), .B2(
        \xmem_data[9][2] ), .ZN(n24356) );
  INV_X1 U28055 ( .A(n24356), .ZN(n24360) );
  AOI22_X1 U28056 ( .A1(n28375), .A2(\xmem_data[14][2] ), .B1(n28334), .B2(
        \xmem_data[15][2] ), .ZN(n24358) );
  NAND2_X1 U28057 ( .A1(n27447), .A2(\xmem_data[11][2] ), .ZN(n24357) );
  NAND2_X1 U28058 ( .A1(n24358), .A2(n24357), .ZN(n24359) );
  NOR2_X1 U28059 ( .A1(n24360), .A2(n24359), .ZN(n24361) );
  NAND2_X1 U28060 ( .A1(n24362), .A2(n24361), .ZN(n24374) );
  AOI22_X1 U28061 ( .A1(n14935), .A2(\xmem_data[16][2] ), .B1(n28053), .B2(
        \xmem_data[17][2] ), .ZN(n24366) );
  AOI22_X1 U28062 ( .A1(n27516), .A2(\xmem_data[18][2] ), .B1(n25434), .B2(
        \xmem_data[19][2] ), .ZN(n24365) );
  AOI22_X1 U28063 ( .A1(n24219), .A2(\xmem_data[20][2] ), .B1(n28687), .B2(
        \xmem_data[21][2] ), .ZN(n24364) );
  AOI22_X1 U28064 ( .A1(n27523), .A2(\xmem_data[22][2] ), .B1(n3325), .B2(
        \xmem_data[23][2] ), .ZN(n24363) );
  NAND4_X1 U28065 ( .A1(n24366), .A2(n24365), .A3(n24364), .A4(n24363), .ZN(
        n24373) );
  AOI22_X1 U28066 ( .A1(n25581), .A2(\xmem_data[24][2] ), .B1(n30269), .B2(
        \xmem_data[25][2] ), .ZN(n24371) );
  AOI22_X1 U28067 ( .A1(n24570), .A2(\xmem_data[26][2] ), .B1(n14976), .B2(
        \xmem_data[27][2] ), .ZN(n24370) );
  AND2_X1 U28068 ( .A1(n31256), .A2(\xmem_data[28][2] ), .ZN(n24367) );
  AOI21_X1 U28069 ( .B1(n28772), .B2(\xmem_data[29][2] ), .A(n24367), .ZN(
        n24369) );
  AOI22_X1 U28070 ( .A1(n27957), .A2(\xmem_data[30][2] ), .B1(n24607), .B2(
        \xmem_data[31][2] ), .ZN(n24368) );
  NAND4_X1 U28071 ( .A1(n24371), .A2(n24370), .A3(n24369), .A4(n24368), .ZN(
        n24372) );
  AOI22_X1 U28072 ( .A1(n29328), .A2(\xmem_data[0][2] ), .B1(n3433), .B2(
        \xmem_data[1][2] ), .ZN(n24380) );
  AND2_X1 U28073 ( .A1(n25485), .A2(\xmem_data[2][2] ), .ZN(n24378) );
  AOI22_X1 U28074 ( .A1(n25491), .A2(\xmem_data[6][2] ), .B1(n25490), .B2(
        \xmem_data[7][2] ), .ZN(n24376) );
  AOI22_X1 U28075 ( .A1(n3219), .A2(\xmem_data[4][2] ), .B1(n21067), .B2(
        \xmem_data[5][2] ), .ZN(n24375) );
  NAND2_X1 U28076 ( .A1(n24376), .A2(n24375), .ZN(n24377) );
  AOI211_X1 U28077 ( .C1(n24694), .C2(\xmem_data[3][2] ), .A(n24378), .B(
        n24377), .ZN(n24379) );
  NAND2_X1 U28078 ( .A1(n24380), .A2(n24379), .ZN(n24381) );
  NOR2_X1 U28079 ( .A1(n24381), .A2(n3805), .ZN(n24382) );
  AOI21_X1 U28080 ( .B1(n24383), .B2(n24382), .A(n25505), .ZN(n24384) );
  AOI21_X1 U28081 ( .B1(n24385), .B2(n25593), .A(n24384), .ZN(n24430) );
  AOI22_X1 U28082 ( .A1(n27501), .A2(\xmem_data[98][2] ), .B1(n25508), .B2(
        \xmem_data[99][2] ), .ZN(n24389) );
  AOI22_X1 U28083 ( .A1(n28317), .A2(\xmem_data[96][2] ), .B1(n24630), .B2(
        \xmem_data[97][2] ), .ZN(n24388) );
  AOI22_X1 U28084 ( .A1(n3219), .A2(\xmem_data[100][2] ), .B1(n29256), .B2(
        \xmem_data[101][2] ), .ZN(n24387) );
  AOI22_X1 U28085 ( .A1(n25509), .A2(\xmem_data[102][2] ), .B1(n25416), .B2(
        \xmem_data[103][2] ), .ZN(n24386) );
  NAND4_X1 U28086 ( .A1(n24389), .A2(n24388), .A3(n24387), .A4(n24386), .ZN(
        n24405) );
  AOI22_X1 U28087 ( .A1(n30550), .A2(\xmem_data[104][2] ), .B1(n28084), .B2(
        \xmem_data[105][2] ), .ZN(n24393) );
  AOI22_X1 U28088 ( .A1(n25514), .A2(\xmem_data[106][2] ), .B1(n27447), .B2(
        \xmem_data[107][2] ), .ZN(n24392) );
  AOI22_X1 U28089 ( .A1(n27988), .A2(\xmem_data[108][2] ), .B1(n28743), .B2(
        \xmem_data[109][2] ), .ZN(n24391) );
  AOI22_X1 U28090 ( .A1(n21075), .A2(\xmem_data[110][2] ), .B1(n28298), .B2(
        \xmem_data[111][2] ), .ZN(n24390) );
  NAND4_X1 U28091 ( .A1(n24393), .A2(n24392), .A3(n24391), .A4(n24390), .ZN(
        n24404) );
  AOI22_X1 U28092 ( .A1(n25709), .A2(\xmem_data[112][2] ), .B1(n25519), .B2(
        \xmem_data[113][2] ), .ZN(n24397) );
  AOI22_X1 U28093 ( .A1(n3208), .A2(\xmem_data[114][2] ), .B1(n20585), .B2(
        \xmem_data[115][2] ), .ZN(n24396) );
  AOI22_X1 U28094 ( .A1(n25520), .A2(\xmem_data[116][2] ), .B1(n30950), .B2(
        \xmem_data[117][2] ), .ZN(n24395) );
  AOI22_X1 U28095 ( .A1(n24221), .A2(\xmem_data[118][2] ), .B1(n25521), .B2(
        \xmem_data[119][2] ), .ZN(n24394) );
  NAND4_X1 U28096 ( .A1(n24397), .A2(n24396), .A3(n24395), .A4(n24394), .ZN(
        n24403) );
  AOI22_X1 U28097 ( .A1(n28462), .A2(\xmem_data[120][2] ), .B1(n24623), .B2(
        \xmem_data[121][2] ), .ZN(n24401) );
  AOI22_X1 U28098 ( .A1(n28983), .A2(\xmem_data[122][2] ), .B1(n25526), .B2(
        \xmem_data[123][2] ), .ZN(n24400) );
  AOI22_X1 U28099 ( .A1(n25527), .A2(\xmem_data[124][2] ), .B1(n30674), .B2(
        \xmem_data[125][2] ), .ZN(n24399) );
  AOI22_X1 U28100 ( .A1(n25528), .A2(\xmem_data[126][2] ), .B1(n25724), .B2(
        \xmem_data[127][2] ), .ZN(n24398) );
  NAND4_X1 U28101 ( .A1(n24401), .A2(n24400), .A3(n24399), .A4(n24398), .ZN(
        n24402) );
  OR4_X1 U28102 ( .A1(n24405), .A2(n24404), .A3(n24403), .A4(n24402), .ZN(
        n24428) );
  AND2_X1 U28103 ( .A1(n20711), .A2(\xmem_data[66][2] ), .ZN(n24406) );
  AOI21_X1 U28104 ( .B1(n25508), .B2(\xmem_data[67][2] ), .A(n24406), .ZN(
        n24410) );
  AOI22_X1 U28105 ( .A1(n28075), .A2(\xmem_data[64][2] ), .B1(n3229), .B2(
        \xmem_data[65][2] ), .ZN(n24409) );
  AOI22_X1 U28106 ( .A1(n3221), .A2(\xmem_data[68][2] ), .B1(n23740), .B2(
        \xmem_data[69][2] ), .ZN(n24408) );
  AOI22_X1 U28107 ( .A1(n25509), .A2(\xmem_data[70][2] ), .B1(n29174), .B2(
        \xmem_data[71][2] ), .ZN(n24407) );
  NAND4_X1 U28108 ( .A1(n24410), .A2(n24409), .A3(n24408), .A4(n24407), .ZN(
        n24426) );
  AOI22_X1 U28109 ( .A1(n24633), .A2(\xmem_data[72][2] ), .B1(n3375), .B2(
        \xmem_data[73][2] ), .ZN(n24414) );
  AOI22_X1 U28110 ( .A1(n25514), .A2(\xmem_data[74][2] ), .B1(n27447), .B2(
        \xmem_data[75][2] ), .ZN(n24413) );
  AOI22_X1 U28111 ( .A1(n24130), .A2(\xmem_data[76][2] ), .B1(n28671), .B2(
        \xmem_data[77][2] ), .ZN(n24412) );
  AOI22_X1 U28112 ( .A1(n24212), .A2(\xmem_data[78][2] ), .B1(n31268), .B2(
        \xmem_data[79][2] ), .ZN(n24411) );
  NAND4_X1 U28113 ( .A1(n24414), .A2(n24413), .A3(n24412), .A4(n24411), .ZN(
        n24425) );
  AOI22_X1 U28114 ( .A1(n25606), .A2(\xmem_data[80][2] ), .B1(n25519), .B2(
        \xmem_data[81][2] ), .ZN(n24418) );
  AOI22_X1 U28115 ( .A1(n29188), .A2(\xmem_data[82][2] ), .B1(n21007), .B2(
        \xmem_data[83][2] ), .ZN(n24417) );
  AOI22_X1 U28116 ( .A1(n25520), .A2(\xmem_data[84][2] ), .B1(n30893), .B2(
        \xmem_data[85][2] ), .ZN(n24416) );
  AOI22_X1 U28117 ( .A1(n13481), .A2(\xmem_data[86][2] ), .B1(n25521), .B2(
        \xmem_data[87][2] ), .ZN(n24415) );
  NAND4_X1 U28118 ( .A1(n24418), .A2(n24417), .A3(n24416), .A4(n24415), .ZN(
        n24424) );
  AOI22_X1 U28119 ( .A1(n25581), .A2(\xmem_data[88][2] ), .B1(n3302), .B2(
        \xmem_data[89][2] ), .ZN(n24422) );
  AOI22_X1 U28120 ( .A1(n24223), .A2(\xmem_data[90][2] ), .B1(n25526), .B2(
        \xmem_data[91][2] ), .ZN(n24421) );
  AOI22_X1 U28121 ( .A1(n25527), .A2(\xmem_data[92][2] ), .B1(n20770), .B2(
        \xmem_data[93][2] ), .ZN(n24420) );
  AOI22_X1 U28122 ( .A1(n25528), .A2(\xmem_data[94][2] ), .B1(n25630), .B2(
        \xmem_data[95][2] ), .ZN(n24419) );
  NAND4_X1 U28123 ( .A1(n24422), .A2(n24421), .A3(n24420), .A4(n24419), .ZN(
        n24423) );
  OR4_X1 U28124 ( .A1(n24426), .A2(n24425), .A3(n24424), .A4(n24423), .ZN(
        n24427) );
  AOI22_X1 U28125 ( .A1(n25560), .A2(n24428), .B1(n25558), .B2(n24427), .ZN(
        n24429) );
  NAND2_X1 U28126 ( .A1(n24430), .A2(n24429), .ZN(n31512) );
  XNOR2_X1 U28127 ( .A(n31512), .B(\fmem_data[17][7] ), .ZN(n31989) );
  INV_X1 U28128 ( .A(n30139), .ZN(n24433) );
  NAND2_X1 U28129 ( .A1(n30138), .A2(n3618), .ZN(n24432) );
  OAI21_X1 U28130 ( .B1(n24434), .B2(n24433), .A(n24432), .ZN(n31793) );
  XNOR2_X1 U28131 ( .A(n32283), .B(\fmem_data[18][7] ), .ZN(n33038) );
  XOR2_X1 U28132 ( .A(\fmem_data[18][6] ), .B(\fmem_data[18][7] ), .Z(n24435)
         );
  XNOR2_X1 U28133 ( .A(n3442), .B(\fmem_data[18][7] ), .ZN(n31820) );
  XNOR2_X1 U28134 ( .A(n32163), .B(\fmem_data[26][5] ), .ZN(n33046) );
  OAI22_X1 U28135 ( .A1(n33046), .A2(n35033), .B1(n24436), .B2(n35034), .ZN(
        n26025) );
  XOR2_X1 U28136 ( .A(\fmem_data[16][5] ), .B(\fmem_data[16][4] ), .Z(n24437)
         );
  AOI22_X1 U28137 ( .A1(n28218), .A2(\xmem_data[4][6] ), .B1(n27444), .B2(
        \xmem_data[5][6] ), .ZN(n24447) );
  AOI22_X1 U28138 ( .A1(n24438), .A2(\xmem_data[6][6] ), .B1(n22669), .B2(
        \xmem_data[7][6] ), .ZN(n24446) );
  AOI22_X1 U28139 ( .A1(n20828), .A2(\xmem_data[0][6] ), .B1(n24439), .B2(
        \xmem_data[1][6] ), .ZN(n24440) );
  INV_X1 U28140 ( .A(n24440), .ZN(n24442) );
  AND2_X1 U28141 ( .A1(n3222), .A2(\xmem_data[3][6] ), .ZN(n24441) );
  NOR2_X1 U28142 ( .A1(n24442), .A2(n24441), .ZN(n24445) );
  NAND2_X1 U28143 ( .A1(n24443), .A2(\xmem_data[2][6] ), .ZN(n24444) );
  NAND4_X1 U28144 ( .A1(n24447), .A2(n24446), .A3(n24445), .A4(n24444), .ZN(
        n24478) );
  AOI22_X1 U28145 ( .A1(n28743), .A2(\xmem_data[12][6] ), .B1(n24448), .B2(
        \xmem_data[13][6] ), .ZN(n24456) );
  AOI22_X1 U28146 ( .A1(n16986), .A2(\xmem_data[14][6] ), .B1(n24160), .B2(
        \xmem_data[15][6] ), .ZN(n24449) );
  INV_X1 U28147 ( .A(n24449), .ZN(n24454) );
  AOI22_X1 U28148 ( .A1(n24450), .A2(\xmem_data[10][6] ), .B1(n22701), .B2(
        \xmem_data[11][6] ), .ZN(n24452) );
  NAND2_X1 U28149 ( .A1(n30710), .A2(\xmem_data[8][6] ), .ZN(n24451) );
  NAND2_X1 U28150 ( .A1(n24452), .A2(n24451), .ZN(n24453) );
  NOR2_X1 U28151 ( .A1(n24454), .A2(n24453), .ZN(n24455) );
  NAND2_X1 U28152 ( .A1(n24456), .A2(n24455), .ZN(n24477) );
  AOI22_X1 U28153 ( .A1(n24458), .A2(\xmem_data[16][6] ), .B1(n24457), .B2(
        \xmem_data[17][6] ), .ZN(n24465) );
  AOI22_X1 U28154 ( .A1(n24133), .A2(\xmem_data[18][6] ), .B1(n24459), .B2(
        \xmem_data[19][6] ), .ZN(n24464) );
  AOI22_X1 U28155 ( .A1(n30309), .A2(\xmem_data[20][6] ), .B1(n24460), .B2(
        \xmem_data[21][6] ), .ZN(n24463) );
  AOI22_X1 U28156 ( .A1(n3178), .A2(\xmem_data[22][6] ), .B1(n28462), .B2(
        \xmem_data[23][6] ), .ZN(n24462) );
  NAND4_X1 U28157 ( .A1(n24465), .A2(n24464), .A3(n24463), .A4(n24462), .ZN(
        n24476) );
  AOI22_X1 U28158 ( .A1(n3338), .A2(\xmem_data[24][6] ), .B1(n23779), .B2(
        \xmem_data[25][6] ), .ZN(n24474) );
  AOI22_X1 U28159 ( .A1(n24467), .A2(\xmem_data[26][6] ), .B1(n28468), .B2(
        \xmem_data[27][6] ), .ZN(n24473) );
  AOI22_X1 U28160 ( .A1(n28467), .A2(\xmem_data[28][6] ), .B1(n24468), .B2(
        \xmem_data[29][6] ), .ZN(n24472) );
  AND2_X1 U28161 ( .A1(n20986), .A2(\xmem_data[30][6] ), .ZN(n24469) );
  AOI21_X1 U28162 ( .B1(n24470), .B2(\xmem_data[31][6] ), .A(n24469), .ZN(
        n24471) );
  NAND4_X1 U28163 ( .A1(n24474), .A2(n24473), .A3(n24472), .A4(n24471), .ZN(
        n24475) );
  NAND2_X1 U28164 ( .A1(n25450), .A2(\xmem_data[9][6] ), .ZN(n24479) );
  AOI21_X1 U28165 ( .B1(n24480), .B2(n24479), .A(n22298), .ZN(n24589) );
  AND2_X1 U28166 ( .A1(n25441), .A2(\xmem_data[62][6] ), .ZN(n24481) );
  AOI21_X1 U28167 ( .B1(n24573), .B2(\xmem_data[63][6] ), .A(n24481), .ZN(
        n24482) );
  AOI22_X1 U28168 ( .A1(n24545), .A2(\xmem_data[48][6] ), .B1(n23716), .B2(
        \xmem_data[49][6] ), .ZN(n24483) );
  INV_X1 U28169 ( .A(n24483), .ZN(n24484) );
  AOI22_X1 U28170 ( .A1(n24571), .A2(\xmem_data[56][6] ), .B1(n24570), .B2(
        \xmem_data[57][6] ), .ZN(n24486) );
  INV_X1 U28171 ( .A(n24486), .ZN(n24497) );
  AOI22_X1 U28172 ( .A1(n29298), .A2(\xmem_data[60][6] ), .B1(n13487), .B2(
        \xmem_data[61][6] ), .ZN(n24487) );
  INV_X1 U28173 ( .A(n24487), .ZN(n24493) );
  AOI22_X1 U28174 ( .A1(n14971), .A2(\xmem_data[52][6] ), .B1(n14913), .B2(
        \xmem_data[53][6] ), .ZN(n24488) );
  INV_X1 U28175 ( .A(n24488), .ZN(n24492) );
  AOI22_X1 U28176 ( .A1(n24547), .A2(\xmem_data[50][6] ), .B1(n24546), .B2(
        \xmem_data[51][6] ), .ZN(n24490) );
  AOI22_X1 U28177 ( .A1(n30525), .A2(\xmem_data[58][6] ), .B1(n29086), .B2(
        \xmem_data[59][6] ), .ZN(n24489) );
  NAND2_X1 U28178 ( .A1(n24490), .A2(n24489), .ZN(n24491) );
  NOR3_X1 U28179 ( .A1(n24493), .A2(n24492), .A3(n24491), .ZN(n24495) );
  AOI22_X1 U28180 ( .A1(n24220), .A2(\xmem_data[54][6] ), .B1(n3372), .B2(
        \xmem_data[55][6] ), .ZN(n24494) );
  NAND2_X1 U28181 ( .A1(n24495), .A2(n24494), .ZN(n24496) );
  AOI22_X1 U28182 ( .A1(n27396), .A2(\xmem_data[40][6] ), .B1(n24553), .B2(
        \xmem_data[41][6] ), .ZN(n24501) );
  AOI22_X1 U28183 ( .A1(n24554), .A2(\xmem_data[42][6] ), .B1(n25456), .B2(
        \xmem_data[43][6] ), .ZN(n24500) );
  AOI22_X1 U28184 ( .A1(n24556), .A2(\xmem_data[44][6] ), .B1(n24555), .B2(
        \xmem_data[45][6] ), .ZN(n24499) );
  AOI22_X1 U28185 ( .A1(n25425), .A2(\xmem_data[46][6] ), .B1(n30541), .B2(
        \xmem_data[47][6] ), .ZN(n24498) );
  AOI22_X1 U28186 ( .A1(n25624), .A2(\xmem_data[32][6] ), .B1(n31347), .B2(
        \xmem_data[33][6] ), .ZN(n24505) );
  AOI22_X1 U28187 ( .A1(n24562), .A2(\xmem_data[34][6] ), .B1(n3219), .B2(
        \xmem_data[35][6] ), .ZN(n24504) );
  AOI22_X1 U28188 ( .A1(n24563), .A2(\xmem_data[36][6] ), .B1(n20500), .B2(
        \xmem_data[37][6] ), .ZN(n24503) );
  AOI22_X1 U28189 ( .A1(n24565), .A2(\xmem_data[38][6] ), .B1(n24564), .B2(
        \xmem_data[39][6] ), .ZN(n24502) );
  NAND2_X1 U28190 ( .A1(n3818), .A2(n3514), .ZN(n24506) );
  NOR3_X1 U28191 ( .A1(n3965), .A2(n24507), .A3(n24506), .ZN(n24587) );
  INV_X1 U28192 ( .A(n24508), .ZN(n24586) );
  AOI22_X1 U28193 ( .A1(n29237), .A2(\xmem_data[112][6] ), .B1(n28335), .B2(
        \xmem_data[113][6] ), .ZN(n24515) );
  AOI22_X1 U28194 ( .A1(n24509), .A2(\xmem_data[114][6] ), .B1(n14912), .B2(
        \xmem_data[115][6] ), .ZN(n24514) );
  AOI22_X1 U28195 ( .A1(n14971), .A2(\xmem_data[116][6] ), .B1(n24510), .B2(
        \xmem_data[117][6] ), .ZN(n24513) );
  AOI22_X1 U28196 ( .A1(n24511), .A2(\xmem_data[118][6] ), .B1(n30898), .B2(
        \xmem_data[119][6] ), .ZN(n24512) );
  NAND4_X1 U28197 ( .A1(n24515), .A2(n24514), .A3(n24513), .A4(n24512), .ZN(
        n24544) );
  AOI22_X1 U28198 ( .A1(n28308), .A2(\xmem_data[104][6] ), .B1(n25514), .B2(
        \xmem_data[105][6] ), .ZN(n24520) );
  AOI22_X1 U28199 ( .A1(n20809), .A2(\xmem_data[106][6] ), .B1(n29307), .B2(
        \xmem_data[107][6] ), .ZN(n24519) );
  AOI22_X1 U28200 ( .A1(n31353), .A2(\xmem_data[108][6] ), .B1(n24516), .B2(
        \xmem_data[109][6] ), .ZN(n24518) );
  AOI22_X1 U28201 ( .A1(n3175), .A2(\xmem_data[110][6] ), .B1(n25671), .B2(
        \xmem_data[111][6] ), .ZN(n24517) );
  NAND4_X1 U28202 ( .A1(n24520), .A2(n24519), .A3(n24518), .A4(n24517), .ZN(
        n24541) );
  AOI22_X1 U28203 ( .A1(n24522), .A2(\xmem_data[120][6] ), .B1(n24521), .B2(
        \xmem_data[121][6] ), .ZN(n24530) );
  AOI22_X1 U28204 ( .A1(n3209), .A2(\xmem_data[122][6] ), .B1(n23725), .B2(
        \xmem_data[123][6] ), .ZN(n24529) );
  AOI22_X1 U28205 ( .A1(n31308), .A2(\xmem_data[124][6] ), .B1(n24524), .B2(
        \xmem_data[125][6] ), .ZN(n24528) );
  AOI22_X1 U28206 ( .A1(n24526), .A2(\xmem_data[126][6] ), .B1(n24525), .B2(
        \xmem_data[127][6] ), .ZN(n24527) );
  NAND4_X1 U28207 ( .A1(n24530), .A2(n24529), .A3(n24528), .A4(n24527), .ZN(
        n24540) );
  AOI22_X1 U28208 ( .A1(n25624), .A2(\xmem_data[96][6] ), .B1(n25687), .B2(
        \xmem_data[97][6] ), .ZN(n24538) );
  AND2_X1 U28209 ( .A1(n3217), .A2(\xmem_data[99][6] ), .ZN(n24531) );
  AOI21_X1 U28210 ( .B1(n24532), .B2(\xmem_data[98][6] ), .A(n24531), .ZN(
        n24537) );
  AOI22_X1 U28211 ( .A1(n24533), .A2(\xmem_data[100][6] ), .B1(n20500), .B2(
        \xmem_data[101][6] ), .ZN(n24536) );
  AOI22_X1 U28212 ( .A1(n24534), .A2(\xmem_data[102][6] ), .B1(n25486), .B2(
        \xmem_data[103][6] ), .ZN(n24535) );
  NAND4_X1 U28213 ( .A1(n24538), .A2(n24537), .A3(n24536), .A4(n24535), .ZN(
        n24539) );
  OR3_X1 U28214 ( .A1(n24541), .A2(n24540), .A3(n24539), .ZN(n24543) );
  OAI21_X1 U28215 ( .B1(n24544), .B2(n24543), .A(n24542), .ZN(n24585) );
  AOI22_X1 U28216 ( .A1(n24545), .A2(\xmem_data[80][6] ), .B1(n25460), .B2(
        \xmem_data[81][6] ), .ZN(n24552) );
  AOI22_X1 U28217 ( .A1(n24547), .A2(\xmem_data[82][6] ), .B1(n24546), .B2(
        \xmem_data[83][6] ), .ZN(n24551) );
  AOI22_X1 U28218 ( .A1(n30617), .A2(\xmem_data[84][6] ), .B1(n25576), .B2(
        \xmem_data[85][6] ), .ZN(n24550) );
  AOI22_X1 U28219 ( .A1(n29100), .A2(\xmem_data[86][6] ), .B1(n28327), .B2(
        \xmem_data[87][6] ), .ZN(n24549) );
  NAND4_X1 U28220 ( .A1(n24552), .A2(n24551), .A3(n24550), .A4(n24549), .ZN(
        n24583) );
  AOI22_X1 U28221 ( .A1(n3281), .A2(\xmem_data[72][6] ), .B1(n24553), .B2(
        \xmem_data[73][6] ), .ZN(n24560) );
  AOI22_X1 U28222 ( .A1(n24554), .A2(\xmem_data[74][6] ), .B1(n27943), .B2(
        \xmem_data[75][6] ), .ZN(n24559) );
  AOI22_X1 U28223 ( .A1(n24556), .A2(\xmem_data[76][6] ), .B1(n24555), .B2(
        \xmem_data[77][6] ), .ZN(n24558) );
  AOI22_X1 U28224 ( .A1(n16986), .A2(\xmem_data[78][6] ), .B1(n29309), .B2(
        \xmem_data[79][6] ), .ZN(n24557) );
  NAND4_X1 U28225 ( .A1(n24560), .A2(n24559), .A3(n24558), .A4(n24557), .ZN(
        n24580) );
  AOI22_X1 U28226 ( .A1(n25443), .A2(\xmem_data[64][6] ), .B1(n31347), .B2(
        \xmem_data[65][6] ), .ZN(n24569) );
  AND2_X1 U28227 ( .A1(n3220), .A2(\xmem_data[67][6] ), .ZN(n24561) );
  AOI21_X1 U28228 ( .B1(n24562), .B2(\xmem_data[66][6] ), .A(n24561), .ZN(
        n24568) );
  AOI22_X1 U28229 ( .A1(n24563), .A2(\xmem_data[68][6] ), .B1(n24695), .B2(
        \xmem_data[69][6] ), .ZN(n24567) );
  AOI22_X1 U28230 ( .A1(n24565), .A2(\xmem_data[70][6] ), .B1(n24564), .B2(
        \xmem_data[71][6] ), .ZN(n24566) );
  NAND4_X1 U28231 ( .A1(n24569), .A2(n24568), .A3(n24567), .A4(n24566), .ZN(
        n24579) );
  AOI22_X1 U28232 ( .A1(n24571), .A2(\xmem_data[88][6] ), .B1(n24570), .B2(
        \xmem_data[89][6] ), .ZN(n24577) );
  AOI22_X1 U28233 ( .A1(n24572), .A2(\xmem_data[90][6] ), .B1(n21057), .B2(
        \xmem_data[91][6] ), .ZN(n24576) );
  AOI22_X1 U28234 ( .A1(n31308), .A2(\xmem_data[92][6] ), .B1(n24122), .B2(
        \xmem_data[93][6] ), .ZN(n24575) );
  AOI22_X1 U28235 ( .A1(n17056), .A2(\xmem_data[94][6] ), .B1(n24573), .B2(
        \xmem_data[95][6] ), .ZN(n24574) );
  NAND4_X1 U28236 ( .A1(n24577), .A2(n24576), .A3(n24575), .A4(n24574), .ZN(
        n24578) );
  OAI21_X1 U28237 ( .B1(n24583), .B2(n24582), .A(n24581), .ZN(n24584) );
  OAI211_X1 U28238 ( .C1(n24587), .C2(n24586), .A(n24585), .B(n24584), .ZN(
        n24588) );
  XNOR2_X1 U28239 ( .A(n34980), .B(\fmem_data[16][5] ), .ZN(n33327) );
  OAI22_X1 U28240 ( .A1(n32017), .A2(n33326), .B1(n33327), .B2(n33328), .ZN(
        n26024) );
  AOI22_X1 U28241 ( .A1(n25422), .A2(\xmem_data[18][3] ), .B1(n24590), .B2(
        \xmem_data[19][3] ), .ZN(n24591) );
  AOI22_X1 U28242 ( .A1(n25400), .A2(\xmem_data[28][3] ), .B1(n24592), .B2(
        \xmem_data[29][3] ), .ZN(n24596) );
  AOI22_X1 U28243 ( .A1(n27944), .A2(\xmem_data[20][3] ), .B1(n13168), .B2(
        \xmem_data[21][3] ), .ZN(n24595) );
  AOI22_X1 U28244 ( .A1(n24593), .A2(\xmem_data[26][3] ), .B1(n25677), .B2(
        \xmem_data[27][3] ), .ZN(n24594) );
  NAND4_X1 U28245 ( .A1(n24591), .A2(n24596), .A3(n24595), .A4(n24594), .ZN(
        n24601) );
  AOI22_X1 U28246 ( .A1(n25461), .A2(\xmem_data[24][3] ), .B1(n29188), .B2(
        \xmem_data[25][3] ), .ZN(n24599) );
  AOI22_X1 U28247 ( .A1(n24597), .A2(\xmem_data[23][3] ), .B1(n20506), .B2(
        \xmem_data[31][3] ), .ZN(n24598) );
  NAND2_X1 U28248 ( .A1(n24599), .A2(n24598), .ZN(n24600) );
  OR2_X1 U28249 ( .A1(n24601), .A2(n24600), .ZN(n24614) );
  AOI22_X1 U28250 ( .A1(n3142), .A2(\xmem_data[8][3] ), .B1(n3247), .B2(
        \xmem_data[9][3] ), .ZN(n24605) );
  AOI22_X1 U28251 ( .A1(n28318), .A2(\xmem_data[10][3] ), .B1(n3219), .B2(
        \xmem_data[11][3] ), .ZN(n24604) );
  AOI22_X1 U28252 ( .A1(n29832), .A2(\xmem_data[12][3] ), .B1(n23769), .B2(
        \xmem_data[13][3] ), .ZN(n24603) );
  AOI22_X1 U28253 ( .A1(n24697), .A2(\xmem_data[14][3] ), .B1(n27994), .B2(
        \xmem_data[15][3] ), .ZN(n24602) );
  NAND4_X1 U28254 ( .A1(n24605), .A2(n24604), .A3(n24603), .A4(n24602), .ZN(
        n24613) );
  AOI22_X1 U28255 ( .A1(n3329), .A2(\xmem_data[0][3] ), .B1(n27365), .B2(
        \xmem_data[1][3] ), .ZN(n24611) );
  AOI22_X1 U28256 ( .A1(n24606), .A2(\xmem_data[2][3] ), .B1(n28500), .B2(
        \xmem_data[3][3] ), .ZN(n24610) );
  AOI22_X1 U28257 ( .A1(n30674), .A2(\xmem_data[4][3] ), .B1(n30524), .B2(
        \xmem_data[5][3] ), .ZN(n24609) );
  AOI22_X1 U28258 ( .A1(n24607), .A2(\xmem_data[6][3] ), .B1(n27958), .B2(
        \xmem_data[7][3] ), .ZN(n24608) );
  NAND4_X1 U28259 ( .A1(n24611), .A2(n24610), .A3(n24609), .A4(n24608), .ZN(
        n24612) );
  OR3_X1 U28260 ( .A1(n24614), .A2(n24613), .A3(n24612), .ZN(n24619) );
  NAND2_X1 U28261 ( .A1(n25567), .A2(\xmem_data[22][3] ), .ZN(n24617) );
  AND2_X1 U28262 ( .A1(n3131), .A2(\xmem_data[16][3] ), .ZN(n24620) );
  NOR2_X1 U28263 ( .A1(n24621), .A2(n24620), .ZN(n24663) );
  AOI22_X1 U28264 ( .A1(n24623), .A2(\xmem_data[32][3] ), .B1(n24622), .B2(
        \xmem_data[33][3] ), .ZN(n24629) );
  AOI22_X1 U28265 ( .A1(n3179), .A2(\xmem_data[34][3] ), .B1(n27463), .B2(
        \xmem_data[35][3] ), .ZN(n24628) );
  AOI22_X1 U28266 ( .A1(n20770), .A2(\xmem_data[36][3] ), .B1(n24624), .B2(
        \xmem_data[37][3] ), .ZN(n24627) );
  AOI22_X1 U28267 ( .A1(n24526), .A2(\xmem_data[38][3] ), .B1(n3203), .B2(
        \xmem_data[39][3] ), .ZN(n24626) );
  NAND4_X1 U28268 ( .A1(n24629), .A2(n24628), .A3(n24627), .A4(n24626), .ZN(
        n24655) );
  AOI22_X1 U28269 ( .A1(n24630), .A2(\xmem_data[40][3] ), .B1(n3247), .B2(
        \xmem_data[41][3] ), .ZN(n24637) );
  AOI22_X1 U28270 ( .A1(n24631), .A2(\xmem_data[42][3] ), .B1(n3222), .B2(
        \xmem_data[43][3] ), .ZN(n24636) );
  AOI22_X1 U28271 ( .A1(n24632), .A2(\xmem_data[44][3] ), .B1(n22667), .B2(
        \xmem_data[45][3] ), .ZN(n24635) );
  AOI22_X1 U28272 ( .A1(n3340), .A2(\xmem_data[46][3] ), .B1(n24633), .B2(
        \xmem_data[47][3] ), .ZN(n24634) );
  NAND4_X1 U28273 ( .A1(n24637), .A2(n24636), .A3(n24635), .A4(n24634), .ZN(
        n24654) );
  AOI22_X1 U28274 ( .A1(n3282), .A2(\xmem_data[48][3] ), .B1(n29103), .B2(
        \xmem_data[49][3] ), .ZN(n24644) );
  AOI22_X1 U28275 ( .A1(n24638), .A2(\xmem_data[50][3] ), .B1(n28415), .B2(
        \xmem_data[51][3] ), .ZN(n24643) );
  AOI22_X1 U28276 ( .A1(n24640), .A2(\xmem_data[52][3] ), .B1(n24639), .B2(
        \xmem_data[53][3] ), .ZN(n24642) );
  AOI22_X1 U28277 ( .A1(n28334), .A2(\xmem_data[54][3] ), .B1(n29009), .B2(
        \xmem_data[55][3] ), .ZN(n24641) );
  NAND4_X1 U28278 ( .A1(n24644), .A2(n24643), .A3(n24642), .A4(n24641), .ZN(
        n24653) );
  AOI22_X1 U28279 ( .A1(n24213), .A2(\xmem_data[56][3] ), .B1(n24134), .B2(
        \xmem_data[57][3] ), .ZN(n24651) );
  AOI22_X1 U28280 ( .A1(n23717), .A2(\xmem_data[58][3] ), .B1(n24645), .B2(
        \xmem_data[59][3] ), .ZN(n24650) );
  AOI22_X1 U28281 ( .A1(n20730), .A2(\xmem_data[60][3] ), .B1(n24646), .B2(
        \xmem_data[61][3] ), .ZN(n24649) );
  AOI22_X1 U28282 ( .A1(n24647), .A2(\xmem_data[62][3] ), .B1(n27951), .B2(
        \xmem_data[63][3] ), .ZN(n24648) );
  NAND4_X1 U28283 ( .A1(n24651), .A2(n24650), .A3(n24649), .A4(n24648), .ZN(
        n24652) );
  OR4_X1 U28284 ( .A1(n24655), .A2(n24654), .A3(n24653), .A4(n24652), .ZN(
        n24660) );
  NOR2_X1 U28285 ( .A1(n24662), .A2(n39009), .ZN(n24656) );
  AND2_X1 U28286 ( .A1(n28007), .A2(n24656), .ZN(n24658) );
  AOI22_X1 U28287 ( .A1(n17004), .A2(\xmem_data[96][3] ), .B1(n20781), .B2(
        \xmem_data[97][3] ), .ZN(n24668) );
  AOI22_X1 U28288 ( .A1(n24685), .A2(\xmem_data[98][3] ), .B1(n25359), .B2(
        \xmem_data[99][3] ), .ZN(n24667) );
  AOI22_X1 U28289 ( .A1(n24687), .A2(\xmem_data[100][3] ), .B1(n24686), .B2(
        \xmem_data[101][3] ), .ZN(n24666) );
  AOI22_X1 U28290 ( .A1(n24688), .A2(\xmem_data[102][3] ), .B1(n31262), .B2(
        \xmem_data[103][3] ), .ZN(n24665) );
  NAND4_X1 U28291 ( .A1(n24668), .A2(n24667), .A3(n24666), .A4(n24665), .ZN(
        n24684) );
  AOI22_X1 U28292 ( .A1(n24693), .A2(\xmem_data[104][3] ), .B1(n30863), .B2(
        \xmem_data[105][3] ), .ZN(n24672) );
  AOI22_X1 U28293 ( .A1(n24694), .A2(\xmem_data[106][3] ), .B1(n3221), .B2(
        \xmem_data[107][3] ), .ZN(n24671) );
  AOI22_X1 U28294 ( .A1(n24696), .A2(\xmem_data[108][3] ), .B1(n24695), .B2(
        \xmem_data[109][3] ), .ZN(n24670) );
  AOI22_X1 U28295 ( .A1(n24697), .A2(\xmem_data[110][3] ), .B1(n24140), .B2(
        \xmem_data[111][3] ), .ZN(n24669) );
  NAND4_X1 U28296 ( .A1(n24672), .A2(n24671), .A3(n24670), .A4(n24669), .ZN(
        n24683) );
  AOI22_X1 U28297 ( .A1(n24702), .A2(\xmem_data[112][3] ), .B1(n27446), .B2(
        \xmem_data[113][3] ), .ZN(n24676) );
  AOI22_X1 U28298 ( .A1(n30885), .A2(\xmem_data[114][3] ), .B1(n27863), .B2(
        \xmem_data[115][3] ), .ZN(n24675) );
  AOI22_X1 U28299 ( .A1(n30508), .A2(\xmem_data[116][3] ), .B1(n27452), .B2(
        \xmem_data[117][3] ), .ZN(n24674) );
  AOI22_X1 U28300 ( .A1(n30514), .A2(\xmem_data[118][3] ), .B1(n29046), .B2(
        \xmem_data[119][3] ), .ZN(n24673) );
  NAND4_X1 U28301 ( .A1(n24676), .A2(n24675), .A3(n24674), .A4(n24673), .ZN(
        n24682) );
  AOI22_X1 U28302 ( .A1(n3158), .A2(\xmem_data[120][3] ), .B1(n25383), .B2(
        \xmem_data[121][3] ), .ZN(n24680) );
  AOI22_X1 U28303 ( .A1(n24708), .A2(\xmem_data[122][3] ), .B1(n24707), .B2(
        \xmem_data[123][3] ), .ZN(n24679) );
  AOI22_X1 U28304 ( .A1(n24710), .A2(\xmem_data[124][3] ), .B1(n24709), .B2(
        \xmem_data[125][3] ), .ZN(n24678) );
  AOI22_X1 U28305 ( .A1(n20593), .A2(\xmem_data[126][3] ), .B1(n3372), .B2(
        \xmem_data[127][3] ), .ZN(n24677) );
  NAND4_X1 U28306 ( .A1(n24680), .A2(n24679), .A3(n24678), .A4(n24677), .ZN(
        n24681) );
  OR4_X1 U28307 ( .A1(n24684), .A2(n24683), .A3(n24682), .A4(n24681), .ZN(
        n24721) );
  AOI22_X1 U28308 ( .A1(n14974), .A2(\xmem_data[64][3] ), .B1(n24570), .B2(
        \xmem_data[65][3] ), .ZN(n24692) );
  AOI22_X1 U28309 ( .A1(n24685), .A2(\xmem_data[66][3] ), .B1(n28500), .B2(
        \xmem_data[67][3] ), .ZN(n24691) );
  AOI22_X1 U28310 ( .A1(n24687), .A2(\xmem_data[68][3] ), .B1(n24686), .B2(
        \xmem_data[69][3] ), .ZN(n24690) );
  AOI22_X1 U28311 ( .A1(n24688), .A2(\xmem_data[70][3] ), .B1(n27958), .B2(
        \xmem_data[71][3] ), .ZN(n24689) );
  NAND4_X1 U28312 ( .A1(n24692), .A2(n24691), .A3(n24690), .A4(n24689), .ZN(
        n24718) );
  AOI22_X1 U28313 ( .A1(n24693), .A2(\xmem_data[72][3] ), .B1(n25360), .B2(
        \xmem_data[73][3] ), .ZN(n24701) );
  AOI22_X1 U28314 ( .A1(n24694), .A2(\xmem_data[74][3] ), .B1(n3218), .B2(
        \xmem_data[75][3] ), .ZN(n24700) );
  AOI22_X1 U28315 ( .A1(n24696), .A2(\xmem_data[76][3] ), .B1(n24695), .B2(
        \xmem_data[77][3] ), .ZN(n24699) );
  AOI22_X1 U28316 ( .A1(n24697), .A2(\xmem_data[78][3] ), .B1(n30882), .B2(
        \xmem_data[79][3] ), .ZN(n24698) );
  NAND4_X1 U28317 ( .A1(n24701), .A2(n24700), .A3(n24699), .A4(n24698), .ZN(
        n24717) );
  AOI22_X1 U28318 ( .A1(n24702), .A2(\xmem_data[80][3] ), .B1(n25450), .B2(
        \xmem_data[81][3] ), .ZN(n24706) );
  AOI22_X1 U28319 ( .A1(n30607), .A2(\xmem_data[82][3] ), .B1(n20546), .B2(
        \xmem_data[83][3] ), .ZN(n24705) );
  AOI22_X1 U28320 ( .A1(n20545), .A2(\xmem_data[84][3] ), .B1(n28416), .B2(
        \xmem_data[85][3] ), .ZN(n24704) );
  AOI22_X1 U28321 ( .A1(n3176), .A2(\xmem_data[86][3] ), .B1(n20584), .B2(
        \xmem_data[87][3] ), .ZN(n24703) );
  NAND4_X1 U28322 ( .A1(n24706), .A2(n24705), .A3(n24704), .A4(n24703), .ZN(
        n24716) );
  AOI22_X1 U28323 ( .A1(n27755), .A2(\xmem_data[88][3] ), .B1(n3208), .B2(
        \xmem_data[89][3] ), .ZN(n24714) );
  AOI22_X1 U28324 ( .A1(n24708), .A2(\xmem_data[90][3] ), .B1(n24707), .B2(
        \xmem_data[91][3] ), .ZN(n24713) );
  AOI22_X1 U28325 ( .A1(n24710), .A2(\xmem_data[92][3] ), .B1(n24709), .B2(
        \xmem_data[93][3] ), .ZN(n24712) );
  AOI22_X1 U28326 ( .A1(n28428), .A2(\xmem_data[94][3] ), .B1(n24222), .B2(
        \xmem_data[95][3] ), .ZN(n24711) );
  NAND4_X1 U28327 ( .A1(n24714), .A2(n24713), .A3(n24712), .A4(n24711), .ZN(
        n24715) );
  OR4_X1 U28328 ( .A1(n24718), .A2(n24717), .A3(n24716), .A4(n24715), .ZN(
        n24719) );
  AOI22_X1 U28329 ( .A1(n24722), .A2(n24721), .B1(n24720), .B2(n24719), .ZN(
        n24723) );
  NAND2_X1 U28330 ( .A1(n24724), .A2(n24723), .ZN(n32614) );
  XOR2_X1 U28331 ( .A(\fmem_data[24][6] ), .B(\fmem_data[24][7] ), .Z(n24725)
         );
  AOI22_X1 U28332 ( .A1(n28740), .A2(\xmem_data[64][2] ), .B1(n29798), .B2(
        \xmem_data[65][2] ), .ZN(n24728) );
  INV_X1 U28333 ( .A(n24728), .ZN(n24734) );
  AOI22_X1 U28334 ( .A1(n29705), .A2(\xmem_data[68][2] ), .B1(n28665), .B2(
        \xmem_data[69][2] ), .ZN(n24729) );
  INV_X1 U28335 ( .A(n24729), .ZN(n24733) );
  AOI22_X1 U28336 ( .A1(n3244), .A2(\xmem_data[66][2] ), .B1(n3126), .B2(
        \xmem_data[67][2] ), .ZN(n24731) );
  AOI22_X1 U28337 ( .A1(n28744), .A2(\xmem_data[70][2] ), .B1(n28743), .B2(
        \xmem_data[71][2] ), .ZN(n24730) );
  NAND2_X1 U28338 ( .A1(n24731), .A2(n24730), .ZN(n24732) );
  NOR3_X1 U28339 ( .A1(n24734), .A2(n24733), .A3(n24732), .ZN(n24754) );
  AOI22_X1 U28340 ( .A1(n30250), .A2(\xmem_data[72][2] ), .B1(n28110), .B2(
        \xmem_data[73][2] ), .ZN(n24738) );
  AOI22_X1 U28341 ( .A1(n28753), .A2(\xmem_data[74][2] ), .B1(n29396), .B2(
        \xmem_data[75][2] ), .ZN(n24737) );
  AOI22_X1 U28342 ( .A1(n3164), .A2(\xmem_data[76][2] ), .B1(n3190), .B2(
        \xmem_data[77][2] ), .ZN(n24736) );
  AOI22_X1 U28343 ( .A1(n29476), .A2(\xmem_data[78][2] ), .B1(n28781), .B2(
        \xmem_data[79][2] ), .ZN(n24735) );
  NAND4_X1 U28344 ( .A1(n24738), .A2(n24737), .A3(n24736), .A4(n24735), .ZN(
        n24747) );
  AND2_X1 U28345 ( .A1(n30775), .A2(\xmem_data[93][2] ), .ZN(n24739) );
  AOI21_X1 U28346 ( .B1(n29626), .B2(\xmem_data[92][2] ), .A(n24739), .ZN(
        n24745) );
  AOI22_X1 U28347 ( .A1(n29786), .A2(\xmem_data[88][2] ), .B1(n3124), .B2(
        \xmem_data[89][2] ), .ZN(n24740) );
  AOI22_X1 U28348 ( .A1(n28719), .A2(\xmem_data[90][2] ), .B1(n28718), .B2(
        \xmem_data[91][2] ), .ZN(n24741) );
  NAND2_X1 U28349 ( .A1(n24745), .A2(n24744), .ZN(n24746) );
  NOR2_X1 U28350 ( .A1(n24747), .A2(n24746), .ZN(n24753) );
  AOI22_X1 U28351 ( .A1(n27740), .A2(\xmem_data[94][2] ), .B1(n28733), .B2(
        \xmem_data[95][2] ), .ZN(n24752) );
  AOI22_X1 U28352 ( .A1(n30198), .A2(\xmem_data[80][2] ), .B1(n30170), .B2(
        \xmem_data[81][2] ), .ZN(n24751) );
  AOI22_X1 U28353 ( .A1(n28720), .A2(\xmem_data[82][2] ), .B1(n24623), .B2(
        \xmem_data[83][2] ), .ZN(n24750) );
  AOI22_X1 U28354 ( .A1(n28725), .A2(\xmem_data[84][2] ), .B1(n28724), .B2(
        \xmem_data[85][2] ), .ZN(n24749) );
  AOI22_X1 U28355 ( .A1(n28727), .A2(\xmem_data[86][2] ), .B1(n20708), .B2(
        \xmem_data[87][2] ), .ZN(n24748) );
  NAND4_X1 U28356 ( .A1(n24754), .A2(n24753), .A3(n24752), .A4(n3764), .ZN(
        n24755) );
  NAND2_X1 U28357 ( .A1(n24755), .A2(n28662), .ZN(n24834) );
  AOI22_X1 U28358 ( .A1(n28146), .A2(\xmem_data[100][2] ), .B1(n29389), .B2(
        \xmem_data[101][2] ), .ZN(n24756) );
  INV_X1 U28359 ( .A(n24756), .ZN(n24762) );
  AOI22_X1 U28360 ( .A1(n28740), .A2(\xmem_data[96][2] ), .B1(n30217), .B2(
        \xmem_data[97][2] ), .ZN(n24757) );
  INV_X1 U28361 ( .A(n24757), .ZN(n24761) );
  AOI22_X1 U28362 ( .A1(n3244), .A2(\xmem_data[98][2] ), .B1(n3126), .B2(
        \xmem_data[99][2] ), .ZN(n24759) );
  AOI22_X1 U28363 ( .A1(n28744), .A2(\xmem_data[102][2] ), .B1(n28743), .B2(
        \xmem_data[103][2] ), .ZN(n24758) );
  NAND2_X1 U28364 ( .A1(n24759), .A2(n24758), .ZN(n24760) );
  NOR3_X1 U28365 ( .A1(n24762), .A2(n24761), .A3(n24760), .ZN(n24779) );
  AND2_X1 U28366 ( .A1(n28733), .A2(\xmem_data[127][2] ), .ZN(n24763) );
  AOI21_X1 U28367 ( .B1(n28138), .B2(\xmem_data[126][2] ), .A(n24763), .ZN(
        n24764) );
  INV_X1 U28368 ( .A(n24764), .ZN(n24769) );
  AOI22_X1 U28369 ( .A1(n29433), .A2(\xmem_data[124][2] ), .B1(n28766), .B2(
        \xmem_data[125][2] ), .ZN(n24767) );
  AOI22_X1 U28370 ( .A1(n28719), .A2(\xmem_data[122][2] ), .B1(n28718), .B2(
        \xmem_data[123][2] ), .ZN(n24766) );
  AOI22_X1 U28371 ( .A1(n29829), .A2(\xmem_data[120][2] ), .B1(n3124), .B2(
        \xmem_data[121][2] ), .ZN(n24765) );
  NOR2_X1 U28372 ( .A1(n24769), .A2(n24768), .ZN(n24778) );
  AOI22_X1 U28373 ( .A1(n28680), .A2(\xmem_data[112][2] ), .B1(n29721), .B2(
        \xmem_data[113][2] ), .ZN(n24773) );
  AOI22_X1 U28374 ( .A1(n28720), .A2(\xmem_data[114][2] ), .B1(n24571), .B2(
        \xmem_data[115][2] ), .ZN(n24772) );
  AOI22_X1 U28375 ( .A1(n28725), .A2(\xmem_data[116][2] ), .B1(n28724), .B2(
        \xmem_data[117][2] ), .ZN(n24771) );
  AOI22_X1 U28376 ( .A1(n28727), .A2(\xmem_data[118][2] ), .B1(n21060), .B2(
        \xmem_data[119][2] ), .ZN(n24770) );
  AOI22_X1 U28377 ( .A1(n29395), .A2(\xmem_data[104][2] ), .B1(n26884), .B2(
        \xmem_data[105][2] ), .ZN(n24777) );
  AOI22_X1 U28378 ( .A1(n28753), .A2(\xmem_data[106][2] ), .B1(n29315), .B2(
        \xmem_data[107][2] ), .ZN(n24776) );
  AOI22_X1 U28379 ( .A1(n3166), .A2(\xmem_data[108][2] ), .B1(n3189), .B2(
        \xmem_data[109][2] ), .ZN(n24775) );
  AOI22_X1 U28380 ( .A1(n27031), .A2(\xmem_data[110][2] ), .B1(n28687), .B2(
        \xmem_data[111][2] ), .ZN(n24774) );
  NAND4_X1 U28381 ( .A1(n24779), .A2(n24778), .A3(n3789), .A4(n3508), .ZN(
        n24780) );
  NAND2_X1 U28382 ( .A1(n24780), .A2(n28762), .ZN(n24833) );
  AOI22_X1 U28383 ( .A1(n30635), .A2(\xmem_data[40][2] ), .B1(n28110), .B2(
        \xmem_data[41][2] ), .ZN(n24784) );
  AOI22_X1 U28384 ( .A1(n28686), .A2(\xmem_data[42][2] ), .B1(n23795), .B2(
        \xmem_data[43][2] ), .ZN(n24783) );
  AOI22_X1 U28385 ( .A1(n3164), .A2(\xmem_data[44][2] ), .B1(n3182), .B2(
        \xmem_data[45][2] ), .ZN(n24782) );
  AOI22_X1 U28386 ( .A1(n30062), .A2(\xmem_data[46][2] ), .B1(n28781), .B2(
        \xmem_data[47][2] ), .ZN(n24781) );
  NAND4_X1 U28387 ( .A1(n24784), .A2(n24783), .A3(n24782), .A4(n24781), .ZN(
        n24793) );
  AND2_X1 U28388 ( .A1(n30106), .A2(\xmem_data[61][2] ), .ZN(n24785) );
  AOI21_X1 U28389 ( .B1(n27710), .B2(\xmem_data[60][2] ), .A(n24785), .ZN(
        n24791) );
  AOI22_X1 U28390 ( .A1(n29829), .A2(\xmem_data[56][2] ), .B1(n29497), .B2(
        \xmem_data[57][2] ), .ZN(n24786) );
  AOI22_X1 U28391 ( .A1(n3227), .A2(\xmem_data[58][2] ), .B1(n28677), .B2(
        \xmem_data[59][2] ), .ZN(n24787) );
  NAND2_X1 U28392 ( .A1(n24791), .A2(n24790), .ZN(n24792) );
  NOR2_X1 U28393 ( .A1(n24793), .A2(n24792), .ZN(n24807) );
  AOI22_X1 U28394 ( .A1(n28219), .A2(\xmem_data[32][2] ), .B1(n29798), .B2(
        \xmem_data[33][2] ), .ZN(n24800) );
  AOI22_X1 U28395 ( .A1(n28739), .A2(\xmem_data[36][2] ), .B1(n29389), .B2(
        \xmem_data[37][2] ), .ZN(n24799) );
  AOI22_X1 U28396 ( .A1(n28670), .A2(\xmem_data[34][2] ), .B1(n28308), .B2(
        \xmem_data[35][2] ), .ZN(n24794) );
  AOI22_X1 U28397 ( .A1(n28744), .A2(\xmem_data[38][2] ), .B1(n28671), .B2(
        \xmem_data[39][2] ), .ZN(n24795) );
  AND3_X1 U28398 ( .A1(n24800), .A2(n24799), .A3(n24798), .ZN(n24806) );
  AOI22_X1 U28399 ( .A1(n29628), .A2(\xmem_data[62][2] ), .B1(n29565), .B2(
        \xmem_data[63][2] ), .ZN(n24805) );
  AOI22_X1 U28400 ( .A1(n30198), .A2(\xmem_data[48][2] ), .B1(n29640), .B2(
        \xmem_data[49][2] ), .ZN(n24804) );
  AOI22_X1 U28401 ( .A1(n28702), .A2(\xmem_data[50][2] ), .B1(n28701), .B2(
        \xmem_data[51][2] ), .ZN(n24803) );
  AOI22_X1 U28402 ( .A1(n28725), .A2(\xmem_data[52][2] ), .B1(n28696), .B2(
        \xmem_data[53][2] ), .ZN(n24802) );
  AOI22_X1 U28403 ( .A1(n28681), .A2(\xmem_data[54][2] ), .B1(n29327), .B2(
        \xmem_data[55][2] ), .ZN(n24801) );
  NAND4_X1 U28404 ( .A1(n24807), .A2(n24806), .A3(n24805), .A4(n3762), .ZN(
        n24831) );
  AOI22_X1 U28405 ( .A1(n30302), .A2(\xmem_data[8][2] ), .B1(n28778), .B2(
        \xmem_data[9][2] ), .ZN(n24811) );
  AOI22_X1 U28406 ( .A1(n28753), .A2(\xmem_data[10][2] ), .B1(n30303), .B2(
        \xmem_data[11][2] ), .ZN(n24810) );
  AOI22_X1 U28407 ( .A1(n3166), .A2(\xmem_data[12][2] ), .B1(n3187), .B2(
        \xmem_data[13][2] ), .ZN(n24809) );
  AOI22_X1 U28408 ( .A1(n30070), .A2(\xmem_data[14][2] ), .B1(n28754), .B2(
        \xmem_data[15][2] ), .ZN(n24808) );
  NAND4_X1 U28409 ( .A1(n24808), .A2(n24810), .A3(n24809), .A4(n24811), .ZN(
        n24814) );
  AOI22_X1 U28410 ( .A1(n28700), .A2(\xmem_data[30][2] ), .B1(n30292), .B2(
        \xmem_data[31][2] ), .ZN(n24812) );
  INV_X1 U28411 ( .A(n24812), .ZN(n24813) );
  NOR2_X1 U28412 ( .A1(n24814), .A2(n24813), .ZN(n24829) );
  AOI22_X1 U28413 ( .A1(n28173), .A2(\xmem_data[16][2] ), .B1(n30644), .B2(
        \xmem_data[17][2] ), .ZN(n24818) );
  AOI22_X1 U28414 ( .A1(n28702), .A2(\xmem_data[18][2] ), .B1(n3151), .B2(
        \xmem_data[19][2] ), .ZN(n24817) );
  AOI22_X1 U28415 ( .A1(n28725), .A2(\xmem_data[20][2] ), .B1(n28724), .B2(
        \xmem_data[21][2] ), .ZN(n24816) );
  AOI22_X1 U28416 ( .A1(n29489), .A2(\xmem_data[22][2] ), .B1(n28772), .B2(
        \xmem_data[23][2] ), .ZN(n24815) );
  AOI22_X1 U28417 ( .A1(n28787), .A2(\xmem_data[0][2] ), .B1(n29556), .B2(
        \xmem_data[1][2] ), .ZN(n24822) );
  AOI22_X1 U28418 ( .A1(n3244), .A2(\xmem_data[2][2] ), .B1(n29762), .B2(
        \xmem_data[3][2] ), .ZN(n24821) );
  AOI22_X1 U28419 ( .A1(n30633), .A2(\xmem_data[4][2] ), .B1(n28665), .B2(
        \xmem_data[5][2] ), .ZN(n24820) );
  AOI22_X1 U28420 ( .A1(n28788), .A2(\xmem_data[6][2] ), .B1(n30663), .B2(
        \xmem_data[7][2] ), .ZN(n24819) );
  AOI22_X1 U28421 ( .A1(n27741), .A2(\xmem_data[28][2] ), .B1(n30100), .B2(
        \xmem_data[29][2] ), .ZN(n24823) );
  INV_X1 U28422 ( .A(n24823), .ZN(n24827) );
  AOI22_X1 U28423 ( .A1(n29786), .A2(\xmem_data[24][2] ), .B1(n27723), .B2(
        \xmem_data[25][2] ), .ZN(n24825) );
  AOI22_X1 U28424 ( .A1(n3227), .A2(\xmem_data[26][2] ), .B1(n3149), .B2(
        \xmem_data[27][2] ), .ZN(n24824) );
  NAND2_X1 U28425 ( .A1(n24825), .A2(n24824), .ZN(n24826) );
  NOR2_X1 U28426 ( .A1(n24827), .A2(n24826), .ZN(n24828) );
  NAND4_X1 U28427 ( .A1(n24829), .A2(n3821), .A3(n3521), .A4(n24828), .ZN(
        n24830) );
  AOI22_X1 U28428 ( .A1(n24831), .A2(n28713), .B1(n28794), .B2(n24830), .ZN(
        n24832) );
  NAND3_X1 U28429 ( .A1(n24834), .A2(n24833), .A3(n24832), .ZN(n32233) );
  XNOR2_X1 U28430 ( .A(n32233), .B(\fmem_data[11][7] ), .ZN(n30385) );
  OAI22_X1 U28431 ( .A1(n30385), .A2(n35633), .B1(n24835), .B2(n35634), .ZN(
        n27330) );
  NAND2_X1 U28432 ( .A1(n26038), .A2(n26037), .ZN(n24836) );
  NAND2_X1 U28433 ( .A1(n24837), .A2(n24836), .ZN(n31792) );
  XNOR2_X1 U28434 ( .A(n31848), .B(n31847), .ZN(n24851) );
  FA_X1 U28435 ( .A(n24840), .B(n24839), .CI(n24838), .CO(n31806), .S(n28928)
         );
  INV_X1 U28436 ( .A(n24841), .ZN(n24846) );
  NOR2_X1 U28437 ( .A1(n24842), .A2(n24843), .ZN(n24845) );
  NAND2_X1 U28438 ( .A1(n24843), .A2(n24842), .ZN(n24844) );
  OAI21_X1 U28439 ( .B1(n24846), .B2(n24845), .A(n24844), .ZN(n28927) );
  XNOR2_X1 U28440 ( .A(n24848), .B(n24847), .ZN(n24849) );
  XNOR2_X1 U28441 ( .A(n24850), .B(n24849), .ZN(n28926) );
  XNOR2_X1 U28442 ( .A(n24851), .B(n31846), .ZN(n31774) );
  XNOR2_X1 U28443 ( .A(n32176), .B(\fmem_data[1][7] ), .ZN(n33217) );
  AOI22_X1 U28444 ( .A1(n29790), .A2(\xmem_data[122][5] ), .B1(n29565), .B2(
        \xmem_data[123][5] ), .ZN(n24855) );
  AOI22_X1 U28445 ( .A1(n28734), .A2(\xmem_data[120][5] ), .B1(n29831), .B2(
        \xmem_data[121][5] ), .ZN(n24854) );
  AOI22_X1 U28446 ( .A1(n29630), .A2(\xmem_data[124][5] ), .B1(n28667), .B2(
        \xmem_data[125][5] ), .ZN(n24853) );
  AOI22_X1 U28447 ( .A1(n29568), .A2(\xmem_data[126][5] ), .B1(n3345), .B2(
        \xmem_data[127][5] ), .ZN(n24852) );
  NAND4_X1 U28448 ( .A1(n24855), .A2(n24854), .A3(n24853), .A4(n24852), .ZN(
        n24871) );
  AOI22_X1 U28449 ( .A1(n29616), .A2(\xmem_data[112][5] ), .B1(n29579), .B2(
        \xmem_data[113][5] ), .ZN(n24859) );
  AOI22_X1 U28450 ( .A1(n29617), .A2(\xmem_data[114][5] ), .B1(n27852), .B2(
        \xmem_data[115][5] ), .ZN(n24858) );
  AOI22_X1 U28451 ( .A1(n29583), .A2(\xmem_data[116][5] ), .B1(n29582), .B2(
        \xmem_data[117][5] ), .ZN(n24857) );
  AOI22_X1 U28452 ( .A1(n29584), .A2(\xmem_data[118][5] ), .B1(n28718), .B2(
        \xmem_data[119][5] ), .ZN(n24856) );
  NAND4_X1 U28453 ( .A1(n24859), .A2(n24858), .A3(n24857), .A4(n24856), .ZN(
        n24870) );
  AOI22_X1 U28454 ( .A1(n3163), .A2(\xmem_data[104][5] ), .B1(n3183), .B2(
        \xmem_data[105][5] ), .ZN(n24863) );
  AOI22_X1 U28455 ( .A1(n29476), .A2(\xmem_data[106][5] ), .B1(n29410), .B2(
        \xmem_data[107][5] ), .ZN(n24862) );
  AOI22_X1 U28456 ( .A1(n30717), .A2(\xmem_data[108][5] ), .B1(n29487), .B2(
        \xmem_data[109][5] ), .ZN(n24861) );
  AOI22_X1 U28457 ( .A1(n29574), .A2(\xmem_data[110][5] ), .B1(n29573), .B2(
        \xmem_data[111][5] ), .ZN(n24860) );
  NAND4_X1 U28458 ( .A1(n24863), .A2(n24862), .A3(n24861), .A4(n24860), .ZN(
        n24869) );
  AOI22_X1 U28459 ( .A1(n30633), .A2(\xmem_data[96][5] ), .B1(n28145), .B2(
        \xmem_data[97][5] ), .ZN(n24867) );
  AOI22_X1 U28460 ( .A1(n3239), .A2(\xmem_data[98][5] ), .B1(n29591), .B2(
        \xmem_data[99][5] ), .ZN(n24866) );
  AOI22_X1 U28461 ( .A1(n30250), .A2(\xmem_data[100][5] ), .B1(n29768), .B2(
        \xmem_data[101][5] ), .ZN(n24865) );
  AOI22_X1 U28462 ( .A1(n29593), .A2(\xmem_data[102][5] ), .B1(n27517), .B2(
        \xmem_data[103][5] ), .ZN(n24864) );
  NAND4_X1 U28463 ( .A1(n24867), .A2(n24866), .A3(n24865), .A4(n24864), .ZN(
        n24868) );
  OR4_X2 U28464 ( .A1(n24871), .A2(n24868), .A3(n24869), .A4(n24870), .ZN(
        n24872) );
  NAND2_X1 U28465 ( .A1(n24872), .A2(n29598), .ZN(n24947) );
  AOI22_X1 U28466 ( .A1(n28138), .A2(\xmem_data[90][5] ), .B1(n29627), .B2(
        \xmem_data[91][5] ), .ZN(n24875) );
  AOI22_X1 U28467 ( .A1(n29667), .A2(\xmem_data[94][5] ), .B1(n30698), .B2(
        \xmem_data[95][5] ), .ZN(n24874) );
  AOI22_X1 U28468 ( .A1(n28751), .A2(\xmem_data[68][5] ), .B1(n28778), .B2(
        \xmem_data[69][5] ), .ZN(n24873) );
  NAND2_X1 U28469 ( .A1(n30293), .A2(\xmem_data[93][5] ), .ZN(n24877) );
  NAND2_X1 U28470 ( .A1(n29566), .A2(\xmem_data[92][5] ), .ZN(n24876) );
  AOI22_X1 U28471 ( .A1(n29641), .A2(\xmem_data[78][5] ), .B1(n30645), .B2(
        \xmem_data[79][5] ), .ZN(n24880) );
  AOI22_X1 U28472 ( .A1(n29603), .A2(\xmem_data[66][5] ), .B1(n27911), .B2(
        \xmem_data[67][5] ), .ZN(n24879) );
  AOI22_X1 U28473 ( .A1(n29649), .A2(\xmem_data[70][5] ), .B1(n24545), .B2(
        \xmem_data[71][5] ), .ZN(n24878) );
  AOI22_X1 U28474 ( .A1(n3168), .A2(\xmem_data[72][5] ), .B1(n3186), .B2(
        \xmem_data[73][5] ), .ZN(n24882) );
  AOI22_X1 U28475 ( .A1(n29810), .A2(\xmem_data[74][5] ), .B1(n29639), .B2(
        \xmem_data[75][5] ), .ZN(n24881) );
  NAND4_X1 U28476 ( .A1(n3481), .A2(n3954), .A3(n3554), .A4(n24883), .ZN(
        n24895) );
  AOI22_X1 U28477 ( .A1(n29590), .A2(\xmem_data[64][5] ), .B1(n29646), .B2(
        \xmem_data[65][5] ), .ZN(n24893) );
  AOI22_X1 U28478 ( .A1(n27710), .A2(\xmem_data[88][5] ), .B1(n29697), .B2(
        \xmem_data[89][5] ), .ZN(n24892) );
  AOI22_X1 U28479 ( .A1(n29580), .A2(\xmem_data[80][5] ), .B1(n29579), .B2(
        \xmem_data[81][5] ), .ZN(n24887) );
  AOI22_X1 U28480 ( .A1(n29581), .A2(\xmem_data[82][5] ), .B1(n29725), .B2(
        \xmem_data[83][5] ), .ZN(n24886) );
  AOI22_X1 U28481 ( .A1(n29619), .A2(\xmem_data[84][5] ), .B1(n29618), .B2(
        \xmem_data[85][5] ), .ZN(n24885) );
  AOI22_X1 U28482 ( .A1(n29621), .A2(\xmem_data[86][5] ), .B1(n3142), .B2(
        \xmem_data[87][5] ), .ZN(n24884) );
  NAND4_X1 U28483 ( .A1(n24887), .A2(n24886), .A3(n24885), .A4(n24884), .ZN(
        n24890) );
  AOI22_X1 U28484 ( .A1(n27713), .A2(\xmem_data[76][5] ), .B1(n30170), .B2(
        \xmem_data[77][5] ), .ZN(n24888) );
  INV_X1 U28485 ( .A(n24888), .ZN(n24889) );
  NOR2_X1 U28486 ( .A1(n24890), .A2(n24889), .ZN(n24891) );
  OAI21_X1 U28487 ( .B1(n24895), .B2(n24894), .A(n29600), .ZN(n24946) );
  AOI22_X1 U28488 ( .A1(n27710), .A2(\xmem_data[24][5] ), .B1(n30100), .B2(
        \xmem_data[25][5] ), .ZN(n24899) );
  AOI22_X1 U28489 ( .A1(n29423), .A2(\xmem_data[26][5] ), .B1(n30278), .B2(
        \xmem_data[27][5] ), .ZN(n24898) );
  AOI22_X1 U28490 ( .A1(n29674), .A2(\xmem_data[28][5] ), .B1(n29761), .B2(
        \xmem_data[29][5] ), .ZN(n24897) );
  AOI22_X1 U28491 ( .A1(n29667), .A2(\xmem_data[30][5] ), .B1(n30295), .B2(
        \xmem_data[31][5] ), .ZN(n24896) );
  NAND4_X1 U28492 ( .A1(n24899), .A2(n24898), .A3(n24897), .A4(n24896), .ZN(
        n24915) );
  AOI22_X1 U28493 ( .A1(n28739), .A2(\xmem_data[0][5] ), .B1(n3369), .B2(
        \xmem_data[1][5] ), .ZN(n24903) );
  AOI22_X1 U28494 ( .A1(n3239), .A2(\xmem_data[2][5] ), .B1(n30663), .B2(
        \xmem_data[3][5] ), .ZN(n24902) );
  AOI22_X1 U28495 ( .A1(n27754), .A2(\xmem_data[4][5] ), .B1(n26884), .B2(
        \xmem_data[5][5] ), .ZN(n24901) );
  AOI22_X1 U28496 ( .A1(n29649), .A2(\xmem_data[6][5] ), .B1(n28231), .B2(
        \xmem_data[7][5] ), .ZN(n24900) );
  NAND4_X1 U28497 ( .A1(n24903), .A2(n24902), .A3(n24901), .A4(n24900), .ZN(
        n24914) );
  AOI22_X1 U28498 ( .A1(n3167), .A2(\xmem_data[8][5] ), .B1(n3184), .B2(
        \xmem_data[9][5] ), .ZN(n24907) );
  AOI22_X1 U28499 ( .A1(n28755), .A2(\xmem_data[10][5] ), .B1(n27855), .B2(
        \xmem_data[11][5] ), .ZN(n24906) );
  AOI22_X1 U28500 ( .A1(n30063), .A2(\xmem_data[12][5] ), .B1(n30765), .B2(
        \xmem_data[13][5] ), .ZN(n24905) );
  AOI22_X1 U28501 ( .A1(n29641), .A2(\xmem_data[14][5] ), .B1(n3301), .B2(
        \xmem_data[15][5] ), .ZN(n24904) );
  NAND4_X1 U28502 ( .A1(n24907), .A2(n24906), .A3(n24905), .A4(n24904), .ZN(
        n24913) );
  AOI22_X1 U28503 ( .A1(n29656), .A2(\xmem_data[16][5] ), .B1(n29579), .B2(
        \xmem_data[17][5] ), .ZN(n24911) );
  AOI22_X1 U28504 ( .A1(n29658), .A2(\xmem_data[18][5] ), .B1(n29657), .B2(
        \xmem_data[19][5] ), .ZN(n24910) );
  AOI22_X1 U28505 ( .A1(n29660), .A2(\xmem_data[20][5] ), .B1(n29659), .B2(
        \xmem_data[21][5] ), .ZN(n24909) );
  AOI22_X1 U28506 ( .A1(n29662), .A2(\xmem_data[22][5] ), .B1(n29661), .B2(
        \xmem_data[23][5] ), .ZN(n24908) );
  NAND4_X1 U28507 ( .A1(n24911), .A2(n24910), .A3(n24909), .A4(n24908), .ZN(
        n24912) );
  NAND2_X1 U28508 ( .A1(n24916), .A2(n29681), .ZN(n24945) );
  AOI22_X1 U28509 ( .A1(n28700), .A2(\xmem_data[58][5] ), .B1(n29627), .B2(
        \xmem_data[59][5] ), .ZN(n24917) );
  INV_X1 U28510 ( .A(n24917), .ZN(n24921) );
  AOI22_X1 U28511 ( .A1(n29436), .A2(\xmem_data[36][5] ), .B1(n30634), .B2(
        \xmem_data[37][5] ), .ZN(n24919) );
  AOI22_X1 U28512 ( .A1(n29667), .A2(\xmem_data[62][5] ), .B1(n3135), .B2(
        \xmem_data[63][5] ), .ZN(n24918) );
  NAND2_X1 U28513 ( .A1(n24919), .A2(n24918), .ZN(n24920) );
  NOR2_X1 U28514 ( .A1(n24921), .A2(n24920), .ZN(n24934) );
  AOI22_X1 U28515 ( .A1(n29476), .A2(\xmem_data[42][5] ), .B1(n22717), .B2(
        \xmem_data[43][5] ), .ZN(n24933) );
  AOI22_X1 U28516 ( .A1(n29566), .A2(\xmem_data[60][5] ), .B1(n27833), .B2(
        \xmem_data[61][5] ), .ZN(n24932) );
  AOI22_X1 U28517 ( .A1(n29580), .A2(\xmem_data[48][5] ), .B1(n29579), .B2(
        \xmem_data[49][5] ), .ZN(n24925) );
  AOI22_X1 U28518 ( .A1(n29581), .A2(\xmem_data[50][5] ), .B1(n20577), .B2(
        \xmem_data[51][5] ), .ZN(n24924) );
  AOI22_X1 U28519 ( .A1(n29619), .A2(\xmem_data[52][5] ), .B1(n29618), .B2(
        \xmem_data[53][5] ), .ZN(n24923) );
  AOI22_X1 U28520 ( .A1(n29621), .A2(\xmem_data[54][5] ), .B1(n3142), .B2(
        \xmem_data[55][5] ), .ZN(n24922) );
  NAND4_X1 U28521 ( .A1(n24925), .A2(n24924), .A3(n24923), .A4(n24922), .ZN(
        n24930) );
  AOI22_X1 U28522 ( .A1(n29641), .A2(\xmem_data[46][5] ), .B1(n3270), .B2(
        \xmem_data[47][5] ), .ZN(n24928) );
  AOI22_X1 U28523 ( .A1(n29649), .A2(\xmem_data[38][5] ), .B1(n27455), .B2(
        \xmem_data[39][5] ), .ZN(n24927) );
  AOI22_X1 U28524 ( .A1(n29603), .A2(\xmem_data[34][5] ), .B1(n24640), .B2(
        \xmem_data[35][5] ), .ZN(n24926) );
  NOR2_X1 U28525 ( .A1(n24930), .A2(n24929), .ZN(n24931) );
  NAND4_X1 U28526 ( .A1(n24934), .A2(n24933), .A3(n24932), .A4(n24931), .ZN(
        n24943) );
  AOI22_X1 U28527 ( .A1(n29390), .A2(\xmem_data[32][5] ), .B1(n30730), .B2(
        \xmem_data[33][5] ), .ZN(n24941) );
  AOI22_X1 U28528 ( .A1(n30223), .A2(\xmem_data[56][5] ), .B1(n27832), .B2(
        \xmem_data[57][5] ), .ZN(n24935) );
  INV_X1 U28529 ( .A(n24935), .ZN(n24939) );
  AOI22_X1 U28530 ( .A1(n29815), .A2(\xmem_data[44][5] ), .B1(n29640), .B2(
        \xmem_data[45][5] ), .ZN(n24937) );
  AOI22_X1 U28531 ( .A1(n3161), .A2(\xmem_data[40][5] ), .B1(n3186), .B2(
        \xmem_data[41][5] ), .ZN(n24936) );
  NAND2_X1 U28532 ( .A1(n24937), .A2(n24936), .ZN(n24938) );
  NOR2_X1 U28533 ( .A1(n24939), .A2(n24938), .ZN(n24940) );
  NAND2_X1 U28534 ( .A1(n24941), .A2(n24940), .ZN(n24942) );
  OAI21_X1 U28535 ( .B1(n24943), .B2(n24942), .A(n29683), .ZN(n24944) );
  NAND4_X2 U28536 ( .A1(n24945), .A2(n24946), .A3(n24947), .A4(n24944), .ZN(
        n33027) );
  XNOR2_X1 U28537 ( .A(n33027), .B(\fmem_data[7][7] ), .ZN(n35141) );
  AOI22_X1 U28538 ( .A1(n3165), .A2(\xmem_data[72][4] ), .B1(n3188), .B2(
        \xmem_data[73][4] ), .ZN(n24951) );
  AOI22_X1 U28539 ( .A1(n30075), .A2(\xmem_data[74][4] ), .B1(n16990), .B2(
        \xmem_data[75][4] ), .ZN(n24950) );
  AOI22_X1 U28540 ( .A1(n30063), .A2(\xmem_data[76][4] ), .B1(n29721), .B2(
        \xmem_data[77][4] ), .ZN(n24949) );
  AOI22_X1 U28541 ( .A1(n29641), .A2(\xmem_data[78][4] ), .B1(n21056), .B2(
        \xmem_data[79][4] ), .ZN(n24948) );
  AOI22_X1 U28542 ( .A1(n29630), .A2(\xmem_data[92][4] ), .B1(n30293), .B2(
        \xmem_data[93][4] ), .ZN(n24955) );
  AOI22_X1 U28543 ( .A1(n3392), .A2(\xmem_data[90][4] ), .B1(n29627), .B2(
        \xmem_data[91][4] ), .ZN(n24954) );
  AOI22_X1 U28544 ( .A1(n29421), .A2(\xmem_data[88][4] ), .B1(n26616), .B2(
        \xmem_data[89][4] ), .ZN(n24953) );
  AOI22_X1 U28545 ( .A1(n29667), .A2(\xmem_data[94][4] ), .B1(n3140), .B2(
        \xmem_data[95][4] ), .ZN(n24952) );
  AOI22_X1 U28546 ( .A1(n28739), .A2(\xmem_data[64][4] ), .B1(n30190), .B2(
        \xmem_data[65][4] ), .ZN(n24966) );
  AOI22_X1 U28547 ( .A1(n29616), .A2(\xmem_data[80][4] ), .B1(n29579), .B2(
        \xmem_data[81][4] ), .ZN(n24959) );
  AOI22_X1 U28548 ( .A1(n29617), .A2(\xmem_data[82][4] ), .B1(n31308), .B2(
        \xmem_data[83][4] ), .ZN(n24958) );
  AOI22_X1 U28549 ( .A1(n29619), .A2(\xmem_data[84][4] ), .B1(n29618), .B2(
        \xmem_data[85][4] ), .ZN(n24957) );
  AOI22_X1 U28550 ( .A1(n29621), .A2(\xmem_data[86][4] ), .B1(n3142), .B2(
        \xmem_data[87][4] ), .ZN(n24956) );
  NAND4_X1 U28551 ( .A1(n24959), .A2(n24958), .A3(n24957), .A4(n24956), .ZN(
        n24964) );
  AOI22_X1 U28552 ( .A1(n29714), .A2(\xmem_data[68][4] ), .B1(n30084), .B2(
        \xmem_data[69][4] ), .ZN(n24962) );
  AOI22_X1 U28553 ( .A1(n29649), .A2(\xmem_data[70][4] ), .B1(n28053), .B2(
        \xmem_data[71][4] ), .ZN(n24961) );
  AOI22_X1 U28554 ( .A1(n29603), .A2(\xmem_data[66][4] ), .B1(n30744), .B2(
        \xmem_data[67][4] ), .ZN(n24960) );
  NOR2_X1 U28555 ( .A1(n24964), .A2(n24963), .ZN(n24965) );
  NAND4_X1 U28556 ( .A1(n3855), .A2(n24967), .A3(n24966), .A4(n24965), .ZN(
        n24968) );
  NAND2_X1 U28557 ( .A1(n24968), .A2(n29600), .ZN(n25047) );
  AOI22_X1 U28558 ( .A1(n29433), .A2(\xmem_data[24][4] ), .B1(n26616), .B2(
        \xmem_data[25][4] ), .ZN(n24985) );
  AOI22_X1 U28559 ( .A1(n29656), .A2(\xmem_data[16][4] ), .B1(n29615), .B2(
        \xmem_data[17][4] ), .ZN(n24972) );
  AOI22_X1 U28560 ( .A1(n29658), .A2(\xmem_data[18][4] ), .B1(n29657), .B2(
        \xmem_data[19][4] ), .ZN(n24971) );
  AOI22_X1 U28561 ( .A1(n29660), .A2(\xmem_data[20][4] ), .B1(n29659), .B2(
        \xmem_data[21][4] ), .ZN(n24970) );
  AOI22_X1 U28562 ( .A1(n29662), .A2(\xmem_data[22][4] ), .B1(n29661), .B2(
        \xmem_data[23][4] ), .ZN(n24969) );
  NAND4_X1 U28563 ( .A1(n24972), .A2(n24971), .A3(n24970), .A4(n24969), .ZN(
        n24977) );
  AOI22_X1 U28564 ( .A1(n28755), .A2(\xmem_data[10][4] ), .B1(n29639), .B2(
        \xmem_data[11][4] ), .ZN(n24973) );
  INV_X1 U28565 ( .A(n24973), .ZN(n24976) );
  AOI22_X1 U28566 ( .A1(n29641), .A2(\xmem_data[14][4] ), .B1(n30600), .B2(
        \xmem_data[15][4] ), .ZN(n24974) );
  INV_X1 U28567 ( .A(n24974), .ZN(n24975) );
  NOR3_X1 U28568 ( .A1(n24977), .A2(n24976), .A3(n24975), .ZN(n24984) );
  AOI22_X1 U28569 ( .A1(n29446), .A2(\xmem_data[0][4] ), .B1(n3117), .B2(
        \xmem_data[1][4] ), .ZN(n24983) );
  AOI22_X1 U28570 ( .A1(n3161), .A2(\xmem_data[8][4] ), .B1(n3183), .B2(
        \xmem_data[9][4] ), .ZN(n24978) );
  INV_X1 U28571 ( .A(n24978), .ZN(n24981) );
  AOI22_X1 U28572 ( .A1(n28680), .A2(\xmem_data[12][4] ), .B1(n29487), .B2(
        \xmem_data[13][4] ), .ZN(n24979) );
  INV_X1 U28573 ( .A(n24979), .ZN(n24980) );
  NOR2_X1 U28574 ( .A1(n24981), .A2(n24980), .ZN(n24982) );
  NAND4_X1 U28575 ( .A1(n24985), .A2(n24984), .A3(n24983), .A4(n24982), .ZN(
        n24996) );
  AOI22_X1 U28576 ( .A1(n29674), .A2(\xmem_data[28][4] ), .B1(n29556), .B2(
        \xmem_data[29][4] ), .ZN(n24994) );
  AOI22_X1 U28577 ( .A1(n29790), .A2(\xmem_data[26][4] ), .B1(n29565), .B2(
        \xmem_data[27][4] ), .ZN(n24993) );
  AOI22_X1 U28578 ( .A1(n29667), .A2(\xmem_data[30][4] ), .B1(n30295), .B2(
        \xmem_data[31][4] ), .ZN(n24986) );
  INV_X1 U28579 ( .A(n24986), .ZN(n24991) );
  AOI22_X1 U28580 ( .A1(n28751), .A2(\xmem_data[4][4] ), .B1(n28778), .B2(
        \xmem_data[5][4] ), .ZN(n24989) );
  AOI22_X1 U28581 ( .A1(n29649), .A2(\xmem_data[6][4] ), .B1(n28516), .B2(
        \xmem_data[7][4] ), .ZN(n24988) );
  AOI22_X1 U28582 ( .A1(n3239), .A2(\xmem_data[2][4] ), .B1(n25457), .B2(
        \xmem_data[3][4] ), .ZN(n24987) );
  NOR2_X1 U28583 ( .A1(n24991), .A2(n24990), .ZN(n24992) );
  OAI21_X1 U28584 ( .B1(n24996), .B2(n24995), .A(n29681), .ZN(n25046) );
  AOI22_X1 U28585 ( .A1(n3163), .A2(\xmem_data[40][4] ), .B1(n3186), .B2(
        \xmem_data[41][4] ), .ZN(n25000) );
  AOI22_X1 U28586 ( .A1(n29716), .A2(\xmem_data[42][4] ), .B1(n29410), .B2(
        \xmem_data[43][4] ), .ZN(n24999) );
  AOI22_X1 U28587 ( .A1(n30766), .A2(\xmem_data[44][4] ), .B1(n30644), .B2(
        \xmem_data[45][4] ), .ZN(n24998) );
  AOI22_X1 U28588 ( .A1(n29641), .A2(\xmem_data[46][4] ), .B1(n3307), .B2(
        \xmem_data[47][4] ), .ZN(n24997) );
  NAND4_X1 U28589 ( .A1(n25000), .A2(n24999), .A3(n24998), .A4(n24997), .ZN(
        n25018) );
  AOI22_X1 U28590 ( .A1(n30633), .A2(\xmem_data[32][4] ), .B1(n29589), .B2(
        \xmem_data[33][4] ), .ZN(n25016) );
  AOI22_X1 U28591 ( .A1(n29616), .A2(\xmem_data[48][4] ), .B1(n29615), .B2(
        \xmem_data[49][4] ), .ZN(n25004) );
  AOI22_X1 U28592 ( .A1(n29617), .A2(\xmem_data[50][4] ), .B1(n28772), .B2(
        \xmem_data[51][4] ), .ZN(n25003) );
  AOI22_X1 U28593 ( .A1(n29619), .A2(\xmem_data[52][4] ), .B1(n29618), .B2(
        \xmem_data[53][4] ), .ZN(n25002) );
  AOI22_X1 U28594 ( .A1(n29621), .A2(\xmem_data[54][4] ), .B1(n3142), .B2(
        \xmem_data[55][4] ), .ZN(n25001) );
  AOI22_X1 U28595 ( .A1(n28700), .A2(\xmem_data[58][4] ), .B1(n29627), .B2(
        \xmem_data[59][4] ), .ZN(n25005) );
  AOI22_X1 U28596 ( .A1(n28779), .A2(\xmem_data[36][4] ), .B1(n29592), .B2(
        \xmem_data[37][4] ), .ZN(n25006) );
  AOI22_X1 U28597 ( .A1(n29626), .A2(\xmem_data[56][4] ), .B1(n30222), .B2(
        \xmem_data[57][4] ), .ZN(n25007) );
  INV_X1 U28598 ( .A(n25007), .ZN(n25012) );
  AOI22_X1 U28599 ( .A1(n29667), .A2(\xmem_data[62][4] ), .B1(n28344), .B2(
        \xmem_data[63][4] ), .ZN(n25010) );
  AOI22_X1 U28600 ( .A1(n29649), .A2(\xmem_data[38][4] ), .B1(n3121), .B2(
        \xmem_data[39][4] ), .ZN(n25009) );
  AOI22_X1 U28601 ( .A1(n29603), .A2(\xmem_data[34][4] ), .B1(n22738), .B2(
        \xmem_data[35][4] ), .ZN(n25008) );
  NOR2_X1 U28602 ( .A1(n25012), .A2(n25011), .ZN(n25014) );
  AOI22_X1 U28603 ( .A1(n29630), .A2(\xmem_data[60][4] ), .B1(n29761), .B2(
        \xmem_data[61][4] ), .ZN(n25013) );
  NAND4_X1 U28604 ( .A1(n25016), .A2(n25015), .A3(n25014), .A4(n25013), .ZN(
        n25017) );
  OAI21_X1 U28605 ( .B1(n25018), .B2(n25017), .A(n29683), .ZN(n25045) );
  AOI22_X1 U28606 ( .A1(n29580), .A2(\xmem_data[112][4] ), .B1(n29579), .B2(
        \xmem_data[113][4] ), .ZN(n25022) );
  AOI22_X1 U28607 ( .A1(n29581), .A2(\xmem_data[114][4] ), .B1(n23730), .B2(
        \xmem_data[115][4] ), .ZN(n25021) );
  AOI22_X1 U28608 ( .A1(n29583), .A2(\xmem_data[116][4] ), .B1(n29582), .B2(
        \xmem_data[117][4] ), .ZN(n25020) );
  AOI22_X1 U28609 ( .A1(n29584), .A2(\xmem_data[118][4] ), .B1(n3348), .B2(
        \xmem_data[119][4] ), .ZN(n25019) );
  NAND4_X1 U28610 ( .A1(n25022), .A2(n25021), .A3(n25020), .A4(n25019), .ZN(
        n25027) );
  AOI22_X1 U28611 ( .A1(n28755), .A2(\xmem_data[106][4] ), .B1(n29639), .B2(
        \xmem_data[107][4] ), .ZN(n25023) );
  INV_X1 U28612 ( .A(n25023), .ZN(n25026) );
  AOI22_X1 U28613 ( .A1(n3165), .A2(\xmem_data[104][4] ), .B1(n3185), .B2(
        \xmem_data[105][4] ), .ZN(n25024) );
  INV_X1 U28614 ( .A(n25024), .ZN(n25025) );
  NOR3_X1 U28615 ( .A1(n25027), .A2(n25026), .A3(n25025), .ZN(n25037) );
  AOI22_X1 U28616 ( .A1(n28700), .A2(\xmem_data[122][4] ), .B1(n29565), .B2(
        \xmem_data[123][4] ), .ZN(n25036) );
  AOI22_X1 U28617 ( .A1(n29566), .A2(\xmem_data[124][4] ), .B1(n30696), .B2(
        \xmem_data[125][4] ), .ZN(n25035) );
  AOI22_X1 U28618 ( .A1(n30291), .A2(\xmem_data[120][4] ), .B1(n29697), .B2(
        \xmem_data[121][4] ), .ZN(n25028) );
  INV_X1 U28619 ( .A(n25028), .ZN(n25033) );
  AOI22_X1 U28620 ( .A1(n30717), .A2(\xmem_data[108][4] ), .B1(n30685), .B2(
        \xmem_data[109][4] ), .ZN(n25031) );
  AOI22_X1 U28621 ( .A1(n29574), .A2(\xmem_data[110][4] ), .B1(n29573), .B2(
        \xmem_data[111][4] ), .ZN(n25030) );
  AOI22_X1 U28622 ( .A1(n29568), .A2(\xmem_data[126][4] ), .B1(n3345), .B2(
        \xmem_data[127][4] ), .ZN(n25029) );
  NOR2_X1 U28623 ( .A1(n25033), .A2(n25032), .ZN(n25034) );
  NAND4_X1 U28624 ( .A1(n25037), .A2(n25036), .A3(n25035), .A4(n25034), .ZN(
        n25043) );
  AOI22_X1 U28625 ( .A1(n27703), .A2(\xmem_data[96][4] ), .B1(n3368), .B2(
        \xmem_data[97][4] ), .ZN(n25041) );
  AOI22_X1 U28626 ( .A1(n3239), .A2(\xmem_data[98][4] ), .B1(n29591), .B2(
        \xmem_data[99][4] ), .ZN(n25040) );
  AOI22_X1 U28627 ( .A1(n3174), .A2(\xmem_data[100][4] ), .B1(n30249), .B2(
        \xmem_data[101][4] ), .ZN(n25039) );
  AOI22_X1 U28628 ( .A1(n29593), .A2(\xmem_data[102][4] ), .B1(n25461), .B2(
        \xmem_data[103][4] ), .ZN(n25038) );
  NAND4_X1 U28629 ( .A1(n25041), .A2(n25040), .A3(n25039), .A4(n25038), .ZN(
        n25042) );
  OAI21_X1 U28630 ( .B1(n25043), .B2(n25042), .A(n29598), .ZN(n25044) );
  XNOR2_X1 U28631 ( .A(n32174), .B(\fmem_data[7][7] ), .ZN(n31938) );
  OAI22_X1 U28632 ( .A1(n35141), .A2(n35619), .B1(n31938), .B2(n35618), .ZN(
        n31796) );
  XNOR2_X1 U28633 ( .A(n35242), .B(\fmem_data[27][5] ), .ZN(n34902) );
  XNOR2_X1 U28634 ( .A(n35145), .B(\fmem_data[27][5] ), .ZN(n31981) );
  XOR2_X1 U28635 ( .A(\fmem_data[27][4] ), .B(\fmem_data[27][5] ), .Z(n25048)
         );
  OAI22_X1 U28636 ( .A1(n34902), .A2(n34903), .B1(n31981), .B2(n34904), .ZN(
        n31795) );
  XNOR2_X1 U28637 ( .A(n34859), .B(\fmem_data[25][5] ), .ZN(n33042) );
  XNOR2_X1 U28638 ( .A(n34982), .B(\fmem_data[25][5] ), .ZN(n31825) );
  OAI22_X1 U28639 ( .A1(n33042), .A2(n34985), .B1(n31825), .B2(n34986), .ZN(
        n31644) );
  AOI22_X1 U28640 ( .A1(n28355), .A2(\xmem_data[68][7] ), .B1(n3219), .B2(
        \xmem_data[69][7] ), .ZN(n25056) );
  AOI22_X1 U28641 ( .A1(n28354), .A2(\xmem_data[64][7] ), .B1(n27499), .B2(
        \xmem_data[65][7] ), .ZN(n25055) );
  AOI22_X1 U28642 ( .A1(n20805), .A2(\xmem_data[70][7] ), .B1(n28356), .B2(
        \xmem_data[71][7] ), .ZN(n25050) );
  INV_X1 U28643 ( .A(n25050), .ZN(n25053) );
  AOI22_X1 U28644 ( .A1(n3386), .A2(\xmem_data[66][7] ), .B1(n27437), .B2(
        \xmem_data[67][7] ), .ZN(n25051) );
  INV_X1 U28645 ( .A(n25051), .ZN(n25052) );
  NOR2_X1 U28646 ( .A1(n25053), .A2(n25052), .ZN(n25054) );
  NAND3_X1 U28647 ( .A1(n25054), .A2(n25055), .A3(n25056), .ZN(n25072) );
  AOI22_X1 U28648 ( .A1(n28428), .A2(\xmem_data[88][7] ), .B1(n21009), .B2(
        \xmem_data[89][7] ), .ZN(n25060) );
  AOI22_X1 U28649 ( .A1(n24623), .A2(\xmem_data[90][7] ), .B1(n27975), .B2(
        \xmem_data[91][7] ), .ZN(n25059) );
  AOI22_X1 U28650 ( .A1(n3179), .A2(\xmem_data[92][7] ), .B1(n28328), .B2(
        \xmem_data[93][7] ), .ZN(n25058) );
  AOI22_X1 U28651 ( .A1(n28241), .A2(\xmem_data[94][7] ), .B1(n28329), .B2(
        \xmem_data[95][7] ), .ZN(n25057) );
  NAND4_X1 U28652 ( .A1(n25060), .A2(n25059), .A3(n25058), .A4(n25057), .ZN(
        n25071) );
  AOI22_X1 U28653 ( .A1(n28336), .A2(\xmem_data[82][7] ), .B1(n28335), .B2(
        \xmem_data[83][7] ), .ZN(n25064) );
  AOI22_X1 U28654 ( .A1(n28334), .A2(\xmem_data[80][7] ), .B1(n27536), .B2(
        \xmem_data[81][7] ), .ZN(n25063) );
  AOI22_X1 U28655 ( .A1(n28337), .A2(\xmem_data[84][7] ), .B1(n29048), .B2(
        \xmem_data[85][7] ), .ZN(n25062) );
  AOI22_X1 U28656 ( .A1(n30893), .A2(\xmem_data[86][7] ), .B1(n29318), .B2(
        \xmem_data[87][7] ), .ZN(n25061) );
  NAND4_X1 U28657 ( .A1(n25064), .A2(n25063), .A3(n25062), .A4(n25061), .ZN(
        n25070) );
  AOI22_X1 U28658 ( .A1(n17010), .A2(\xmem_data[72][7] ), .B1(n28342), .B2(
        \xmem_data[73][7] ), .ZN(n25068) );
  AOI22_X1 U28659 ( .A1(n28344), .A2(\xmem_data[74][7] ), .B1(n3231), .B2(
        \xmem_data[75][7] ), .ZN(n25067) );
  AOI22_X1 U28660 ( .A1(n30885), .A2(\xmem_data[76][7] ), .B1(n29180), .B2(
        \xmem_data[77][7] ), .ZN(n25066) );
  AOI22_X1 U28661 ( .A1(n28346), .A2(\xmem_data[78][7] ), .B1(n28345), .B2(
        \xmem_data[79][7] ), .ZN(n25065) );
  NAND4_X1 U28662 ( .A1(n25068), .A2(n25067), .A3(n25066), .A4(n25065), .ZN(
        n25069) );
  OR4_X1 U28663 ( .A1(n25072), .A2(n25071), .A3(n25070), .A4(n25069), .ZN(
        n25073) );
  NAND2_X1 U28664 ( .A1(n25073), .A2(n28324), .ZN(n25144) );
  AND2_X1 U28665 ( .A1(n3221), .A2(\xmem_data[37][7] ), .ZN(n25074) );
  AOI21_X1 U28666 ( .B1(n28355), .B2(\xmem_data[36][7] ), .A(n25074), .ZN(
        n25081) );
  AOI22_X1 U28667 ( .A1(n28354), .A2(\xmem_data[32][7] ), .B1(n25357), .B2(
        \xmem_data[33][7] ), .ZN(n25080) );
  AOI22_X1 U28668 ( .A1(n24533), .A2(\xmem_data[38][7] ), .B1(n28356), .B2(
        \xmem_data[39][7] ), .ZN(n25075) );
  INV_X1 U28669 ( .A(n25075), .ZN(n25078) );
  AOI22_X1 U28670 ( .A1(n3245), .A2(\xmem_data[34][7] ), .B1(n28501), .B2(
        \xmem_data[35][7] ), .ZN(n25076) );
  INV_X1 U28671 ( .A(n25076), .ZN(n25077) );
  NOR2_X1 U28672 ( .A1(n25078), .A2(n25077), .ZN(n25079) );
  NAND3_X1 U28673 ( .A1(n25081), .A2(n25080), .A3(n25079), .ZN(n25097) );
  AOI22_X1 U28674 ( .A1(n22683), .A2(\xmem_data[56][7] ), .B1(n23778), .B2(
        \xmem_data[57][7] ), .ZN(n25085) );
  AOI22_X1 U28675 ( .A1(n28202), .A2(\xmem_data[58][7] ), .B1(n29245), .B2(
        \xmem_data[59][7] ), .ZN(n25084) );
  AOI22_X1 U28676 ( .A1(n3179), .A2(\xmem_data[60][7] ), .B1(n28328), .B2(
        \xmem_data[61][7] ), .ZN(n25083) );
  AOI22_X1 U28677 ( .A1(n28467), .A2(\xmem_data[62][7] ), .B1(n28329), .B2(
        \xmem_data[63][7] ), .ZN(n25082) );
  NAND4_X1 U28678 ( .A1(n25085), .A2(n25084), .A3(n25083), .A4(n25082), .ZN(
        n25096) );
  AOI22_X1 U28679 ( .A1(n28334), .A2(\xmem_data[48][7] ), .B1(n29309), .B2(
        \xmem_data[49][7] ), .ZN(n25089) );
  AOI22_X1 U28680 ( .A1(n28336), .A2(\xmem_data[50][7] ), .B1(n28335), .B2(
        \xmem_data[51][7] ), .ZN(n25088) );
  AOI22_X1 U28681 ( .A1(n28337), .A2(\xmem_data[52][7] ), .B1(n29048), .B2(
        \xmem_data[53][7] ), .ZN(n25087) );
  AOI22_X1 U28682 ( .A1(n24710), .A2(\xmem_data[54][7] ), .B1(n29280), .B2(
        \xmem_data[55][7] ), .ZN(n25086) );
  NAND4_X1 U28683 ( .A1(n25089), .A2(n25088), .A3(n25087), .A4(n25086), .ZN(
        n25095) );
  AOI22_X1 U28684 ( .A1(n24565), .A2(\xmem_data[40][7] ), .B1(n28342), .B2(
        \xmem_data[41][7] ), .ZN(n25093) );
  AOI22_X1 U28685 ( .A1(n28344), .A2(\xmem_data[42][7] ), .B1(n23771), .B2(
        \xmem_data[43][7] ), .ZN(n25092) );
  AOI22_X1 U28686 ( .A1(n25422), .A2(\xmem_data[44][7] ), .B1(n3357), .B2(
        \xmem_data[45][7] ), .ZN(n25091) );
  AOI22_X1 U28687 ( .A1(n28346), .A2(\xmem_data[46][7] ), .B1(n28345), .B2(
        \xmem_data[47][7] ), .ZN(n25090) );
  NAND4_X1 U28688 ( .A1(n25093), .A2(n25092), .A3(n25091), .A4(n25090), .ZN(
        n25094) );
  OR4_X1 U28689 ( .A1(n25097), .A2(n25096), .A3(n25095), .A4(n25094), .ZN(
        n25098) );
  NAND2_X1 U28690 ( .A1(n25098), .A2(n28361), .ZN(n25143) );
  AOI22_X1 U28691 ( .A1(n24548), .A2(\xmem_data[120][7] ), .B1(n28291), .B2(
        \xmem_data[121][7] ), .ZN(n25102) );
  AOI22_X1 U28692 ( .A1(n30269), .A2(\xmem_data[122][7] ), .B1(n27975), .B2(
        \xmem_data[123][7] ), .ZN(n25101) );
  AOI22_X1 U28693 ( .A1(n28293), .A2(\xmem_data[124][7] ), .B1(n28292), .B2(
        \xmem_data[125][7] ), .ZN(n25100) );
  AOI22_X1 U28694 ( .A1(n20577), .A2(\xmem_data[126][7] ), .B1(n28035), .B2(
        \xmem_data[127][7] ), .ZN(n25099) );
  NAND4_X1 U28695 ( .A1(n25102), .A2(n25101), .A3(n25100), .A4(n25099), .ZN(
        n25113) );
  AOI22_X1 U28696 ( .A1(n28298), .A2(\xmem_data[112][7] ), .B1(n23793), .B2(
        \xmem_data[113][7] ), .ZN(n25106) );
  AOI22_X1 U28697 ( .A1(n3158), .A2(\xmem_data[114][7] ), .B1(n28299), .B2(
        \xmem_data[115][7] ), .ZN(n25105) );
  AOI22_X1 U28698 ( .A1(n23717), .A2(\xmem_data[116][7] ), .B1(n29316), .B2(
        \xmem_data[117][7] ), .ZN(n25104) );
  AOI22_X1 U28699 ( .A1(n28302), .A2(\xmem_data[118][7] ), .B1(n28301), .B2(
        \xmem_data[119][7] ), .ZN(n25103) );
  NAND4_X1 U28700 ( .A1(n25106), .A2(n25105), .A3(n25104), .A4(n25103), .ZN(
        n25112) );
  AOI22_X1 U28701 ( .A1(n25490), .A2(\xmem_data[104][7] ), .B1(n31275), .B2(
        \xmem_data[105][7] ), .ZN(n25110) );
  AOI22_X1 U28702 ( .A1(n28308), .A2(\xmem_data[106][7] ), .B1(n28307), .B2(
        \xmem_data[107][7] ), .ZN(n25109) );
  AOI22_X1 U28703 ( .A1(n30885), .A2(\xmem_data[108][7] ), .B1(n28481), .B2(
        \xmem_data[109][7] ), .ZN(n25108) );
  AOI22_X1 U28704 ( .A1(n28309), .A2(\xmem_data[110][7] ), .B1(n21015), .B2(
        \xmem_data[111][7] ), .ZN(n25107) );
  NAND4_X1 U28705 ( .A1(n25110), .A2(n25109), .A3(n25108), .A4(n25107), .ZN(
        n25111) );
  OR3_X1 U28706 ( .A1(n25113), .A2(n25112), .A3(n25111), .ZN(n25119) );
  AOI22_X1 U28707 ( .A1(n28318), .A2(\xmem_data[100][7] ), .B1(n3222), .B2(
        \xmem_data[101][7] ), .ZN(n25117) );
  AOI22_X1 U28708 ( .A1(n3245), .A2(\xmem_data[98][7] ), .B1(n29286), .B2(
        \xmem_data[99][7] ), .ZN(n25116) );
  AOI22_X1 U28709 ( .A1(n25724), .A2(\xmem_data[96][7] ), .B1(n28317), .B2(
        \xmem_data[97][7] ), .ZN(n25115) );
  AOI22_X1 U28710 ( .A1(n20724), .A2(\xmem_data[102][7] ), .B1(n28319), .B2(
        \xmem_data[103][7] ), .ZN(n25114) );
  NAND4_X1 U28711 ( .A1(n25117), .A2(n25116), .A3(n25115), .A4(n25114), .ZN(
        n25118) );
  OAI21_X1 U28712 ( .B1(n25119), .B2(n25118), .A(n28288), .ZN(n25142) );
  AOI22_X1 U28713 ( .A1(n28038), .A2(\xmem_data[0][7] ), .B1(n28366), .B2(
        \xmem_data[1][7] ), .ZN(n25123) );
  AOI22_X1 U28714 ( .A1(n3305), .A2(\xmem_data[2][7] ), .B1(n25687), .B2(
        \xmem_data[3][7] ), .ZN(n25122) );
  AOI22_X1 U28715 ( .A1(n28364), .A2(\xmem_data[4][7] ), .B1(n3218), .B2(
        \xmem_data[5][7] ), .ZN(n25121) );
  AOI22_X1 U28716 ( .A1(n28367), .A2(\xmem_data[6][7] ), .B1(n28508), .B2(
        \xmem_data[7][7] ), .ZN(n25120) );
  NAND4_X1 U28717 ( .A1(n25123), .A2(n25122), .A3(n25121), .A4(n25120), .ZN(
        n25139) );
  AOI22_X1 U28718 ( .A1(n28083), .A2(\xmem_data[8][7] ), .B1(n28372), .B2(
        \xmem_data[9][7] ), .ZN(n25127) );
  AOI22_X1 U28719 ( .A1(n28084), .A2(\xmem_data[10][7] ), .B1(n3231), .B2(
        \xmem_data[11][7] ), .ZN(n25126) );
  AOI22_X1 U28720 ( .A1(n28374), .A2(\xmem_data[12][7] ), .B1(n3357), .B2(
        \xmem_data[13][7] ), .ZN(n25125) );
  AOI22_X1 U28721 ( .A1(n27944), .A2(\xmem_data[14][7] ), .B1(n28375), .B2(
        \xmem_data[15][7] ), .ZN(n25124) );
  NAND4_X1 U28722 ( .A1(n25127), .A2(n25126), .A3(n25125), .A4(n25124), .ZN(
        n25138) );
  AOI22_X1 U28723 ( .A1(n25710), .A2(\xmem_data[16][7] ), .B1(n22741), .B2(
        \xmem_data[17][7] ), .ZN(n25131) );
  AOI22_X1 U28724 ( .A1(n24458), .A2(\xmem_data[18][7] ), .B1(n28993), .B2(
        \xmem_data[19][7] ), .ZN(n25130) );
  AOI22_X1 U28725 ( .A1(n24593), .A2(\xmem_data[20][7] ), .B1(n23796), .B2(
        \xmem_data[21][7] ), .ZN(n25129) );
  AOI22_X1 U28726 ( .A1(n21008), .A2(\xmem_data[22][7] ), .B1(n28380), .B2(
        \xmem_data[23][7] ), .ZN(n25128) );
  NAND4_X1 U28727 ( .A1(n25131), .A2(n25130), .A3(n25129), .A4(n25128), .ZN(
        n25137) );
  AOI22_X1 U28728 ( .A1(n28385), .A2(\xmem_data[24][7] ), .B1(n29281), .B2(
        \xmem_data[25][7] ), .ZN(n25135) );
  AOI22_X1 U28729 ( .A1(n3337), .A2(\xmem_data[26][7] ), .B1(n20983), .B2(
        \xmem_data[27][7] ), .ZN(n25134) );
  AOI22_X1 U28730 ( .A1(n3179), .A2(\xmem_data[28][7] ), .B1(n22751), .B2(
        \xmem_data[29][7] ), .ZN(n25133) );
  AOI22_X1 U28731 ( .A1(n13420), .A2(\xmem_data[30][7] ), .B1(n24624), .B2(
        \xmem_data[31][7] ), .ZN(n25132) );
  NAND4_X1 U28732 ( .A1(n25135), .A2(n25134), .A3(n25133), .A4(n25132), .ZN(
        n25136) );
  OR4_X1 U28733 ( .A1(n25139), .A2(n25138), .A3(n25137), .A4(n25136), .ZN(
        n25140) );
  NAND2_X1 U28734 ( .A1(n25140), .A2(n28395), .ZN(n25141) );
  NAND4_X2 U28735 ( .A1(n25144), .A2(n25143), .A3(n25142), .A4(n25141), .ZN(
        n35108) );
  XNOR2_X1 U28736 ( .A(n35108), .B(\fmem_data[18][3] ), .ZN(n33036) );
  XNOR2_X1 U28737 ( .A(n31644), .B(n31645), .ZN(n25147) );
  XNOR2_X1 U28738 ( .A(n31219), .B(\fmem_data[26][7] ), .ZN(n32022) );
  XNOR2_X1 U28739 ( .A(n25147), .B(n31646), .ZN(n30155) );
  XNOR2_X1 U28740 ( .A(n35280), .B(\fmem_data[1][3] ), .ZN(n33190) );
  XOR2_X1 U28741 ( .A(\fmem_data[1][2] ), .B(\fmem_data[1][3] ), .Z(n25148) );
  AOI22_X1 U28742 ( .A1(n3341), .A2(\xmem_data[12][7] ), .B1(n27994), .B2(
        \xmem_data[13][7] ), .ZN(n25150) );
  INV_X1 U28743 ( .A(n25150), .ZN(n25154) );
  AOI22_X1 U28744 ( .A1(n28137), .A2(\xmem_data[10][7] ), .B1(n28356), .B2(
        \xmem_data[11][7] ), .ZN(n25152) );
  NAND2_X1 U28745 ( .A1(n27905), .A2(\xmem_data[14][7] ), .ZN(n25151) );
  NAND2_X1 U28746 ( .A1(n25152), .A2(n25151), .ZN(n25153) );
  NOR2_X1 U28747 ( .A1(n25154), .A2(n25153), .ZN(n25164) );
  AND2_X1 U28748 ( .A1(n29125), .A2(\xmem_data[3][7] ), .ZN(n25155) );
  AOI21_X1 U28749 ( .B1(n28036), .B2(\xmem_data[2][7] ), .A(n25155), .ZN(
        n25163) );
  AOI22_X1 U28750 ( .A1(n30588), .A2(\xmem_data[4][7] ), .B1(n28366), .B2(
        \xmem_data[5][7] ), .ZN(n25156) );
  INV_X1 U28751 ( .A(n25156), .ZN(n25160) );
  AOI22_X1 U28752 ( .A1(n27542), .A2(\xmem_data[0][7] ), .B1(n27981), .B2(
        \xmem_data[1][7] ), .ZN(n25158) );
  AOI22_X1 U28753 ( .A1(n3228), .A2(\xmem_data[6][7] ), .B1(n3247), .B2(
        \xmem_data[7][7] ), .ZN(n25157) );
  NAND2_X1 U28754 ( .A1(n25158), .A2(n25157), .ZN(n25159) );
  NOR2_X1 U28755 ( .A1(n25160), .A2(n25159), .ZN(n25162) );
  AOI22_X1 U28756 ( .A1(n28318), .A2(\xmem_data[8][7] ), .B1(n3220), .B2(
        \xmem_data[9][7] ), .ZN(n25161) );
  NAND4_X1 U28757 ( .A1(n25164), .A2(n25163), .A3(n25162), .A4(n25161), .ZN(
        n25176) );
  AOI22_X1 U28758 ( .A1(n24554), .A2(\xmem_data[16][7] ), .B1(n27988), .B2(
        \xmem_data[17][7] ), .ZN(n25168) );
  AOI22_X1 U28759 ( .A1(n30508), .A2(\xmem_data[18][7] ), .B1(n13168), .B2(
        \xmem_data[19][7] ), .ZN(n25167) );
  AOI22_X1 U28760 ( .A1(n27515), .A2(\xmem_data[20][7] ), .B1(n25458), .B2(
        \xmem_data[21][7] ), .ZN(n25166) );
  AOI22_X1 U28761 ( .A1(n28231), .A2(\xmem_data[22][7] ), .B1(n27989), .B2(
        \xmem_data[23][7] ), .ZN(n25165) );
  NAND4_X1 U28762 ( .A1(n25168), .A2(n25167), .A3(n25166), .A4(n25165), .ZN(
        n25174) );
  AOI22_X1 U28763 ( .A1(n17020), .A2(\xmem_data[24][7] ), .B1(n25398), .B2(
        \xmem_data[25][7] ), .ZN(n25172) );
  AOI22_X1 U28764 ( .A1(n25400), .A2(\xmem_data[26][7] ), .B1(n24221), .B2(
        \xmem_data[27][7] ), .ZN(n25171) );
  AOI22_X1 U28765 ( .A1(n27974), .A2(\xmem_data[28][7] ), .B1(n3372), .B2(
        \xmem_data[29][7] ), .ZN(n25170) );
  AOI22_X1 U28766 ( .A1(n3329), .A2(\xmem_data[30][7] ), .B1(n27975), .B2(
        \xmem_data[31][7] ), .ZN(n25169) );
  NAND4_X1 U28767 ( .A1(n25172), .A2(n25171), .A3(n25170), .A4(n25169), .ZN(
        n25173) );
  NOR2_X1 U28768 ( .A1(n25176), .A2(n25175), .ZN(n25178) );
  NAND2_X1 U28769 ( .A1(n28007), .A2(\xmem_data[15][7] ), .ZN(n25177) );
  AOI21_X1 U28770 ( .B1(n25178), .B2(n25177), .A(n24043), .ZN(n25179) );
  INV_X1 U28771 ( .A(n25179), .ZN(n25245) );
  AOI22_X1 U28772 ( .A1(n24572), .A2(\xmem_data[96][7] ), .B1(n20733), .B2(
        \xmem_data[97][7] ), .ZN(n25183) );
  AOI22_X1 U28773 ( .A1(n28036), .A2(\xmem_data[98][7] ), .B1(n28035), .B2(
        \xmem_data[99][7] ), .ZN(n25182) );
  AOI22_X1 U28774 ( .A1(n28038), .A2(\xmem_data[100][7] ), .B1(n28037), .B2(
        \xmem_data[101][7] ), .ZN(n25181) );
  AOI22_X1 U28775 ( .A1(n28039), .A2(\xmem_data[102][7] ), .B1(n31347), .B2(
        \xmem_data[103][7] ), .ZN(n25180) );
  NAND4_X1 U28776 ( .A1(n25183), .A2(n25182), .A3(n25181), .A4(n25180), .ZN(
        n25199) );
  AOI22_X1 U28777 ( .A1(n28044), .A2(\xmem_data[104][7] ), .B1(n3221), .B2(
        \xmem_data[105][7] ), .ZN(n25187) );
  AOI22_X1 U28778 ( .A1(n24632), .A2(\xmem_data[106][7] ), .B1(n25491), .B2(
        \xmem_data[107][7] ), .ZN(n25186) );
  AOI22_X1 U28779 ( .A1(n24141), .A2(\xmem_data[108][7] ), .B1(n23811), .B2(
        \xmem_data[109][7] ), .ZN(n25185) );
  AOI22_X1 U28780 ( .A1(n23742), .A2(\xmem_data[110][7] ), .B1(n3231), .B2(
        \xmem_data[111][7] ), .ZN(n25184) );
  NAND4_X1 U28781 ( .A1(n25187), .A2(n25186), .A3(n25185), .A4(n25184), .ZN(
        n25198) );
  AOI22_X1 U28782 ( .A1(n28050), .A2(\xmem_data[112][7] ), .B1(n28373), .B2(
        \xmem_data[113][7] ), .ZN(n25191) );
  AOI22_X1 U28783 ( .A1(n28051), .A2(\xmem_data[114][7] ), .B1(n24159), .B2(
        \xmem_data[115][7] ), .ZN(n25190) );
  AOI22_X1 U28784 ( .A1(n17041), .A2(\xmem_data[116][7] ), .B1(n28052), .B2(
        \xmem_data[117][7] ), .ZN(n25189) );
  AOI22_X1 U28785 ( .A1(n20718), .A2(\xmem_data[118][7] ), .B1(n27516), .B2(
        \xmem_data[119][7] ), .ZN(n25188) );
  NAND4_X1 U28786 ( .A1(n25191), .A2(n25190), .A3(n25189), .A4(n25188), .ZN(
        n25197) );
  AOI22_X1 U28787 ( .A1(n28059), .A2(\xmem_data[120][7] ), .B1(n28058), .B2(
        \xmem_data[121][7] ), .ZN(n25195) );
  AOI22_X1 U28788 ( .A1(n20815), .A2(\xmem_data[122][7] ), .B1(n24221), .B2(
        \xmem_data[123][7] ), .ZN(n25194) );
  AOI22_X1 U28789 ( .A1(n28061), .A2(\xmem_data[124][7] ), .B1(n28060), .B2(
        \xmem_data[125][7] ), .ZN(n25193) );
  AOI22_X1 U28790 ( .A1(n3271), .A2(\xmem_data[126][7] ), .B1(n28062), .B2(
        \xmem_data[127][7] ), .ZN(n25192) );
  NAND4_X1 U28791 ( .A1(n25195), .A2(n25194), .A3(n25193), .A4(n25192), .ZN(
        n25196) );
  OR4_X1 U28792 ( .A1(n25199), .A2(n25198), .A3(n25197), .A4(n25196), .ZN(
        n25221) );
  AOI22_X1 U28793 ( .A1(n25582), .A2(\xmem_data[64][7] ), .B1(n20488), .B2(
        \xmem_data[65][7] ), .ZN(n25203) );
  AOI22_X1 U28794 ( .A1(n30901), .A2(\xmem_data[66][7] ), .B1(n30524), .B2(
        \xmem_data[67][7] ), .ZN(n25202) );
  AOI22_X1 U28795 ( .A1(n28076), .A2(\xmem_data[68][7] ), .B1(n28075), .B2(
        \xmem_data[69][7] ), .ZN(n25201) );
  AOI22_X1 U28796 ( .A1(n3434), .A2(\xmem_data[70][7] ), .B1(n3247), .B2(
        \xmem_data[71][7] ), .ZN(n25200) );
  NAND4_X1 U28797 ( .A1(n25203), .A2(n25202), .A3(n25201), .A4(n25200), .ZN(
        n25219) );
  AOI22_X1 U28798 ( .A1(n28082), .A2(\xmem_data[72][7] ), .B1(n3217), .B2(
        \xmem_data[73][7] ), .ZN(n25207) );
  AOI22_X1 U28799 ( .A1(n29494), .A2(\xmem_data[74][7] ), .B1(n22710), .B2(
        \xmem_data[75][7] ), .ZN(n25206) );
  AOI22_X1 U28800 ( .A1(n28083), .A2(\xmem_data[76][7] ), .B1(n3256), .B2(
        \xmem_data[77][7] ), .ZN(n25205) );
  AOI22_X1 U28801 ( .A1(n28084), .A2(\xmem_data[78][7] ), .B1(n25492), .B2(
        \xmem_data[79][7] ), .ZN(n25204) );
  NAND4_X1 U28802 ( .A1(n25207), .A2(n25206), .A3(n25205), .A4(n25204), .ZN(
        n25218) );
  AOI22_X1 U28803 ( .A1(n27551), .A2(\xmem_data[80][7] ), .B1(n13475), .B2(
        \xmem_data[81][7] ), .ZN(n25211) );
  AOI22_X1 U28804 ( .A1(n28089), .A2(\xmem_data[82][7] ), .B1(n24212), .B2(
        \xmem_data[83][7] ), .ZN(n25210) );
  AOI22_X1 U28805 ( .A1(n23763), .A2(\xmem_data[84][7] ), .B1(n28090), .B2(
        \xmem_data[85][7] ), .ZN(n25209) );
  AOI22_X1 U28806 ( .A1(n27517), .A2(\xmem_data[86][7] ), .B1(n3208), .B2(
        \xmem_data[87][7] ), .ZN(n25208) );
  NAND4_X1 U28807 ( .A1(n25211), .A2(n25210), .A3(n25209), .A4(n25208), .ZN(
        n25217) );
  AOI22_X1 U28808 ( .A1(n28096), .A2(\xmem_data[88][7] ), .B1(n29316), .B2(
        \xmem_data[89][7] ), .ZN(n25215) );
  AOI22_X1 U28809 ( .A1(n27825), .A2(\xmem_data[90][7] ), .B1(n28097), .B2(
        \xmem_data[91][7] ), .ZN(n25214) );
  AOI22_X1 U28810 ( .A1(n28460), .A2(\xmem_data[92][7] ), .B1(n23778), .B2(
        \xmem_data[93][7] ), .ZN(n25213) );
  AOI22_X1 U28811 ( .A1(n29297), .A2(\xmem_data[94][7] ), .B1(n28098), .B2(
        \xmem_data[95][7] ), .ZN(n25212) );
  NAND4_X1 U28812 ( .A1(n25215), .A2(n25214), .A3(n25213), .A4(n25212), .ZN(
        n25216) );
  OR4_X1 U28813 ( .A1(n25219), .A2(n25218), .A3(n25217), .A4(n25216), .ZN(
        n25220) );
  AOI22_X1 U28814 ( .A1(n28071), .A2(n25221), .B1(n28033), .B2(n25220), .ZN(
        n25244) );
  AOI22_X1 U28815 ( .A1(n3171), .A2(\xmem_data[32][7] ), .B1(n20488), .B2(
        \xmem_data[33][7] ), .ZN(n25225) );
  AOI22_X1 U28816 ( .A1(n25407), .A2(\xmem_data[34][7] ), .B1(n25528), .B2(
        \xmem_data[35][7] ), .ZN(n25224) );
  AOI22_X1 U28817 ( .A1(n28076), .A2(\xmem_data[36][7] ), .B1(n28075), .B2(
        \xmem_data[37][7] ), .ZN(n25223) );
  AOI22_X1 U28818 ( .A1(n3434), .A2(\xmem_data[38][7] ), .B1(n3247), .B2(
        \xmem_data[39][7] ), .ZN(n25222) );
  NAND4_X1 U28819 ( .A1(n25225), .A2(n25224), .A3(n25223), .A4(n25222), .ZN(
        n25241) );
  AOI22_X1 U28820 ( .A1(n28082), .A2(\xmem_data[40][7] ), .B1(n3219), .B2(
        \xmem_data[41][7] ), .ZN(n25229) );
  AOI22_X1 U28821 ( .A1(n23740), .A2(\xmem_data[42][7] ), .B1(n24695), .B2(
        \xmem_data[43][7] ), .ZN(n25228) );
  AOI22_X1 U28822 ( .A1(n28083), .A2(\xmem_data[44][7] ), .B1(n27994), .B2(
        \xmem_data[45][7] ), .ZN(n25227) );
  AOI22_X1 U28823 ( .A1(n28084), .A2(\xmem_data[46][7] ), .B1(n25514), .B2(
        \xmem_data[47][7] ), .ZN(n25226) );
  NAND4_X1 U28824 ( .A1(n25229), .A2(n25228), .A3(n25227), .A4(n25226), .ZN(
        n25240) );
  AOI22_X1 U28825 ( .A1(n27551), .A2(\xmem_data[48][7] ), .B1(n13475), .B2(
        \xmem_data[49][7] ), .ZN(n25233) );
  AOI22_X1 U28826 ( .A1(n28089), .A2(\xmem_data[50][7] ), .B1(n24212), .B2(
        \xmem_data[51][7] ), .ZN(n25232) );
  AOI22_X1 U28827 ( .A1(n25567), .A2(\xmem_data[52][7] ), .B1(n28090), .B2(
        \xmem_data[53][7] ), .ZN(n25231) );
  AOI22_X1 U28828 ( .A1(n29437), .A2(\xmem_data[54][7] ), .B1(n23716), .B2(
        \xmem_data[55][7] ), .ZN(n25230) );
  NAND4_X1 U28829 ( .A1(n25233), .A2(n25232), .A3(n25231), .A4(n25230), .ZN(
        n25239) );
  AOI22_X1 U28830 ( .A1(n28096), .A2(\xmem_data[56][7] ), .B1(n27918), .B2(
        \xmem_data[57][7] ), .ZN(n25237) );
  AOI22_X1 U28831 ( .A1(n28687), .A2(\xmem_data[58][7] ), .B1(n28097), .B2(
        \xmem_data[59][7] ), .ZN(n25236) );
  AOI22_X1 U28832 ( .A1(n28428), .A2(\xmem_data[60][7] ), .B1(n25581), .B2(
        \xmem_data[61][7] ), .ZN(n25235) );
  AOI22_X1 U28833 ( .A1(n20817), .A2(\xmem_data[62][7] ), .B1(n28098), .B2(
        \xmem_data[63][7] ), .ZN(n25234) );
  NAND4_X1 U28834 ( .A1(n25237), .A2(n25236), .A3(n25235), .A4(n25234), .ZN(
        n25238) );
  OR4_X1 U28835 ( .A1(n25241), .A2(n25240), .A3(n25239), .A4(n25238), .ZN(
        n25242) );
  NAND2_X1 U28836 ( .A1(n25242), .A2(n28107), .ZN(n25243) );
  XNOR2_X1 U28837 ( .A(n35072), .B(\fmem_data[22][3] ), .ZN(n33050) );
  AOI22_X1 U28838 ( .A1(n24685), .A2(\xmem_data[32][6] ), .B1(n28468), .B2(
        \xmem_data[33][6] ), .ZN(n25249) );
  AOI22_X1 U28839 ( .A1(n30901), .A2(\xmem_data[34][6] ), .B1(n29125), .B2(
        \xmem_data[35][6] ), .ZN(n25248) );
  AOI22_X1 U28840 ( .A1(n28076), .A2(\xmem_data[36][6] ), .B1(n28075), .B2(
        \xmem_data[37][6] ), .ZN(n25247) );
  AOI22_X1 U28841 ( .A1(n3434), .A2(\xmem_data[38][6] ), .B1(n3247), .B2(
        \xmem_data[39][6] ), .ZN(n25246) );
  NAND4_X1 U28842 ( .A1(n25249), .A2(n25248), .A3(n25247), .A4(n25246), .ZN(
        n25265) );
  AOI22_X1 U28843 ( .A1(n28082), .A2(\xmem_data[40][6] ), .B1(n3220), .B2(
        \xmem_data[41][6] ), .ZN(n25253) );
  AOI22_X1 U28844 ( .A1(n20724), .A2(\xmem_data[42][6] ), .B1(n29255), .B2(
        \xmem_data[43][6] ), .ZN(n25252) );
  AOI22_X1 U28845 ( .A1(n28083), .A2(\xmem_data[44][6] ), .B1(n3256), .B2(
        \xmem_data[45][6] ), .ZN(n25251) );
  AOI22_X1 U28846 ( .A1(n28084), .A2(\xmem_data[46][6] ), .B1(n24553), .B2(
        \xmem_data[47][6] ), .ZN(n25250) );
  NAND4_X1 U28847 ( .A1(n25253), .A2(n25252), .A3(n25251), .A4(n25250), .ZN(
        n25264) );
  AOI22_X1 U28848 ( .A1(n27551), .A2(\xmem_data[48][6] ), .B1(n13475), .B2(
        \xmem_data[49][6] ), .ZN(n25257) );
  AOI22_X1 U28849 ( .A1(n28089), .A2(\xmem_data[50][6] ), .B1(n24212), .B2(
        \xmem_data[51][6] ), .ZN(n25256) );
  AOI22_X1 U28850 ( .A1(n30891), .A2(\xmem_data[52][6] ), .B1(n28090), .B2(
        \xmem_data[53][6] ), .ZN(n25255) );
  AOI22_X1 U28851 ( .A1(n30746), .A2(\xmem_data[54][6] ), .B1(n29279), .B2(
        \xmem_data[55][6] ), .ZN(n25254) );
  NAND4_X1 U28852 ( .A1(n25257), .A2(n25256), .A3(n25255), .A4(n25254), .ZN(
        n25263) );
  AOI22_X1 U28853 ( .A1(n28096), .A2(\xmem_data[56][6] ), .B1(n28492), .B2(
        \xmem_data[57][6] ), .ZN(n25261) );
  AOI22_X1 U28854 ( .A1(n29047), .A2(\xmem_data[58][6] ), .B1(n28097), .B2(
        \xmem_data[59][6] ), .ZN(n25260) );
  AOI22_X1 U28855 ( .A1(n25632), .A2(\xmem_data[60][6] ), .B1(n30898), .B2(
        \xmem_data[61][6] ), .ZN(n25259) );
  AOI22_X1 U28856 ( .A1(n23724), .A2(\xmem_data[62][6] ), .B1(n28098), .B2(
        \xmem_data[63][6] ), .ZN(n25258) );
  NAND4_X1 U28857 ( .A1(n25261), .A2(n25260), .A3(n25259), .A4(n25258), .ZN(
        n25262) );
  OR4_X1 U28858 ( .A1(n25265), .A2(n25264), .A3(n25263), .A4(n25262), .ZN(
        n25288) );
  AOI22_X1 U28859 ( .A1(n20782), .A2(\xmem_data[0][6] ), .B1(n27981), .B2(
        \xmem_data[1][6] ), .ZN(n25269) );
  AOI22_X1 U28860 ( .A1(n29820), .A2(\xmem_data[2][6] ), .B1(n24468), .B2(
        \xmem_data[3][6] ), .ZN(n25268) );
  AOI22_X1 U28861 ( .A1(n30862), .A2(\xmem_data[4][6] ), .B1(n25561), .B2(
        \xmem_data[5][6] ), .ZN(n25267) );
  AOI22_X1 U28862 ( .A1(n3449), .A2(\xmem_data[6][6] ), .B1(n28501), .B2(
        \xmem_data[7][6] ), .ZN(n25266) );
  NAND4_X1 U28863 ( .A1(n25269), .A2(n25268), .A3(n25267), .A4(n25266), .ZN(
        n25285) );
  AOI22_X1 U28864 ( .A1(n28318), .A2(\xmem_data[8][6] ), .B1(n3218), .B2(
        \xmem_data[9][6] ), .ZN(n25273) );
  AOI22_X1 U28865 ( .A1(n29627), .A2(\xmem_data[10][6] ), .B1(n24695), .B2(
        \xmem_data[11][6] ), .ZN(n25272) );
  AOI22_X1 U28866 ( .A1(n24565), .A2(\xmem_data[12][6] ), .B1(n27994), .B2(
        \xmem_data[13][6] ), .ZN(n25271) );
  AOI22_X1 U28867 ( .A1(n3137), .A2(\xmem_data[14][6] ), .B1(n30877), .B2(
        \xmem_data[15][6] ), .ZN(n25270) );
  NAND4_X1 U28868 ( .A1(n25273), .A2(n25272), .A3(n25271), .A4(n25270), .ZN(
        n25284) );
  AOI22_X1 U28869 ( .A1(n25422), .A2(\xmem_data[16][6] ), .B1(n27988), .B2(
        \xmem_data[17][6] ), .ZN(n25277) );
  AOI22_X1 U28870 ( .A1(n27514), .A2(\xmem_data[18][6] ), .B1(n28416), .B2(
        \xmem_data[19][6] ), .ZN(n25276) );
  AOI22_X1 U28871 ( .A1(n17041), .A2(\xmem_data[20][6] ), .B1(n24160), .B2(
        \xmem_data[21][6] ), .ZN(n25275) );
  AOI22_X1 U28872 ( .A1(n27945), .A2(\xmem_data[22][6] ), .B1(n27989), .B2(
        \xmem_data[23][6] ), .ZN(n25274) );
  NAND4_X1 U28873 ( .A1(n25277), .A2(n25276), .A3(n25275), .A4(n25274), .ZN(
        n25283) );
  AOI22_X1 U28874 ( .A1(n25434), .A2(\xmem_data[24][6] ), .B1(n25398), .B2(
        \xmem_data[25][6] ), .ZN(n25281) );
  AOI22_X1 U28875 ( .A1(n28781), .A2(\xmem_data[26][6] ), .B1(n31254), .B2(
        \xmem_data[27][6] ), .ZN(n25280) );
  AOI22_X1 U28876 ( .A1(n27974), .A2(\xmem_data[28][6] ), .B1(n25716), .B2(
        \xmem_data[29][6] ), .ZN(n25279) );
  AOI22_X1 U28877 ( .A1(n3330), .A2(\xmem_data[30][6] ), .B1(n27975), .B2(
        \xmem_data[31][6] ), .ZN(n25278) );
  NAND4_X1 U28878 ( .A1(n25281), .A2(n25280), .A3(n25279), .A4(n25278), .ZN(
        n25282) );
  OR4_X1 U28879 ( .A1(n25285), .A2(n25284), .A3(n25283), .A4(n25282), .ZN(
        n25286) );
  AOI22_X1 U28880 ( .A1(n28107), .A2(n25288), .B1(n25287), .B2(n25286), .ZN(
        n25332) );
  AOI22_X1 U28881 ( .A1(n24572), .A2(\xmem_data[96][6] ), .B1(n20733), .B2(
        \xmem_data[97][6] ), .ZN(n25292) );
  AOI22_X1 U28882 ( .A1(n28036), .A2(\xmem_data[98][6] ), .B1(n28035), .B2(
        \xmem_data[99][6] ), .ZN(n25291) );
  AOI22_X1 U28883 ( .A1(n28038), .A2(\xmem_data[100][6] ), .B1(n28037), .B2(
        \xmem_data[101][6] ), .ZN(n25290) );
  AOI22_X1 U28884 ( .A1(n28039), .A2(\xmem_data[102][6] ), .B1(n28501), .B2(
        \xmem_data[103][6] ), .ZN(n25289) );
  NAND4_X1 U28885 ( .A1(n25292), .A2(n25291), .A3(n25290), .A4(n25289), .ZN(
        n25308) );
  AOI22_X1 U28886 ( .A1(n28044), .A2(\xmem_data[104][6] ), .B1(n3217), .B2(
        \xmem_data[105][6] ), .ZN(n25296) );
  AOI22_X1 U28887 ( .A1(n23770), .A2(\xmem_data[106][6] ), .B1(n29095), .B2(
        \xmem_data[107][6] ), .ZN(n25295) );
  AOI22_X1 U28888 ( .A1(n28475), .A2(\xmem_data[108][6] ), .B1(n29181), .B2(
        \xmem_data[109][6] ), .ZN(n25294) );
  AOI22_X1 U28889 ( .A1(n17063), .A2(\xmem_data[110][6] ), .B1(n25450), .B2(
        \xmem_data[111][6] ), .ZN(n25293) );
  NAND4_X1 U28890 ( .A1(n25296), .A2(n25295), .A3(n25294), .A4(n25293), .ZN(
        n25307) );
  AOI22_X1 U28891 ( .A1(n28050), .A2(\xmem_data[112][6] ), .B1(n24590), .B2(
        \xmem_data[113][6] ), .ZN(n25300) );
  AOI22_X1 U28892 ( .A1(n28051), .A2(\xmem_data[114][6] ), .B1(n24212), .B2(
        \xmem_data[115][6] ), .ZN(n25299) );
  AOI22_X1 U28893 ( .A1(n20495), .A2(\xmem_data[116][6] ), .B1(n28052), .B2(
        \xmem_data[117][6] ), .ZN(n25298) );
  AOI22_X1 U28894 ( .A1(n29315), .A2(\xmem_data[118][6] ), .B1(n29279), .B2(
        \xmem_data[119][6] ), .ZN(n25297) );
  NAND4_X1 U28895 ( .A1(n25300), .A2(n25299), .A3(n25298), .A4(n25297), .ZN(
        n25306) );
  AOI22_X1 U28896 ( .A1(n28059), .A2(\xmem_data[120][6] ), .B1(n28058), .B2(
        \xmem_data[121][6] ), .ZN(n25304) );
  AOI22_X1 U28897 ( .A1(n25678), .A2(\xmem_data[122][6] ), .B1(n31254), .B2(
        \xmem_data[123][6] ), .ZN(n25303) );
  AOI22_X1 U28898 ( .A1(n28061), .A2(\xmem_data[124][6] ), .B1(n28060), .B2(
        \xmem_data[125][6] ), .ZN(n25302) );
  AOI22_X1 U28899 ( .A1(n3338), .A2(\xmem_data[126][6] ), .B1(n28062), .B2(
        \xmem_data[127][6] ), .ZN(n25301) );
  NAND4_X1 U28900 ( .A1(n25304), .A2(n25303), .A3(n25302), .A4(n25301), .ZN(
        n25305) );
  OR4_X1 U28901 ( .A1(n25308), .A2(n25307), .A3(n25306), .A4(n25305), .ZN(
        n25330) );
  AOI22_X1 U28902 ( .A1(n30497), .A2(\xmem_data[64][6] ), .B1(n27981), .B2(
        \xmem_data[65][6] ), .ZN(n25312) );
  AOI22_X1 U28903 ( .A1(n25407), .A2(\xmem_data[66][6] ), .B1(n20769), .B2(
        \xmem_data[67][6] ), .ZN(n25311) );
  AOI22_X1 U28904 ( .A1(n28076), .A2(\xmem_data[68][6] ), .B1(n28075), .B2(
        \xmem_data[69][6] ), .ZN(n25310) );
  AOI22_X1 U28905 ( .A1(n3434), .A2(\xmem_data[70][6] ), .B1(n3247), .B2(
        \xmem_data[71][6] ), .ZN(n25309) );
  NAND4_X1 U28906 ( .A1(n25312), .A2(n25311), .A3(n25310), .A4(n25309), .ZN(
        n25328) );
  AOI22_X1 U28907 ( .A1(n28082), .A2(\xmem_data[72][6] ), .B1(n3218), .B2(
        \xmem_data[73][6] ), .ZN(n25316) );
  AOI22_X1 U28908 ( .A1(n24696), .A2(\xmem_data[74][6] ), .B1(n27869), .B2(
        \xmem_data[75][6] ), .ZN(n25315) );
  AOI22_X1 U28909 ( .A1(n28083), .A2(\xmem_data[76][6] ), .B1(n24564), .B2(
        \xmem_data[77][6] ), .ZN(n25314) );
  AOI22_X1 U28910 ( .A1(n28084), .A2(\xmem_data[78][6] ), .B1(n28307), .B2(
        \xmem_data[79][6] ), .ZN(n25313) );
  NAND4_X1 U28911 ( .A1(n25316), .A2(n25315), .A3(n25314), .A4(n25313), .ZN(
        n25327) );
  AOI22_X1 U28912 ( .A1(n27551), .A2(\xmem_data[80][6] ), .B1(n13475), .B2(
        \xmem_data[81][6] ), .ZN(n25320) );
  AOI22_X1 U28913 ( .A1(n28089), .A2(\xmem_data[82][6] ), .B1(n24159), .B2(
        \xmem_data[83][6] ), .ZN(n25319) );
  AOI22_X1 U28914 ( .A1(n29109), .A2(\xmem_data[84][6] ), .B1(n28090), .B2(
        \xmem_data[85][6] ), .ZN(n25318) );
  AOI22_X1 U28915 ( .A1(n21048), .A2(\xmem_data[86][6] ), .B1(n29279), .B2(
        \xmem_data[87][6] ), .ZN(n25317) );
  NAND4_X1 U28916 ( .A1(n25320), .A2(n25319), .A3(n25318), .A4(n25317), .ZN(
        n25326) );
  AOI22_X1 U28917 ( .A1(n28096), .A2(\xmem_data[88][6] ), .B1(n25677), .B2(
        \xmem_data[89][6] ), .ZN(n25324) );
  AOI22_X1 U28918 ( .A1(n30309), .A2(\xmem_data[90][6] ), .B1(n28097), .B2(
        \xmem_data[91][6] ), .ZN(n25323) );
  AOI22_X1 U28919 ( .A1(n3206), .A2(\xmem_data[92][6] ), .B1(n25581), .B2(
        \xmem_data[93][6] ), .ZN(n25322) );
  AOI22_X1 U28920 ( .A1(n20817), .A2(\xmem_data[94][6] ), .B1(n28098), .B2(
        \xmem_data[95][6] ), .ZN(n25321) );
  NAND4_X1 U28921 ( .A1(n25324), .A2(n25323), .A3(n25322), .A4(n25321), .ZN(
        n25325) );
  OR4_X1 U28922 ( .A1(n25328), .A2(n25327), .A3(n25326), .A4(n25325), .ZN(
        n25329) );
  AOI22_X1 U28923 ( .A1(n28071), .A2(n25330), .B1(n28033), .B2(n25329), .ZN(
        n25331) );
  NAND2_X1 U28924 ( .A1(n25332), .A2(n25331), .ZN(n35073) );
  XOR2_X1 U28925 ( .A(\fmem_data[22][3] ), .B(\fmem_data[22][2] ), .Z(n25333)
         );
  OAI22_X1 U28926 ( .A1(n33050), .A2(n34414), .B1(n30370), .B2(n34416), .ZN(
        n28934) );
  AOI22_X1 U28927 ( .A1(n25434), .A2(\xmem_data[32][7] ), .B1(n28427), .B2(
        \xmem_data[33][7] ), .ZN(n25337) );
  AOI22_X1 U28928 ( .A1(n24115), .A2(\xmem_data[34][7] ), .B1(n25435), .B2(
        \xmem_data[35][7] ), .ZN(n25336) );
  AOI22_X1 U28929 ( .A1(n28428), .A2(\xmem_data[36][7] ), .B1(n23778), .B2(
        \xmem_data[37][7] ), .ZN(n25335) );
  AOI22_X1 U28930 ( .A1(n3308), .A2(\xmem_data[38][7] ), .B1(n24223), .B2(
        \xmem_data[39][7] ), .ZN(n25334) );
  NAND4_X1 U28931 ( .A1(n25337), .A2(n25336), .A3(n25335), .A4(n25334), .ZN(
        n25353) );
  AOI22_X1 U28932 ( .A1(n21058), .A2(\xmem_data[40][7] ), .B1(n28328), .B2(
        \xmem_data[41][7] ), .ZN(n25341) );
  AOI22_X1 U28933 ( .A1(n30901), .A2(\xmem_data[42][7] ), .B1(n25440), .B2(
        \xmem_data[43][7] ), .ZN(n25340) );
  AOI22_X1 U28934 ( .A1(n25441), .A2(\xmem_data[44][7] ), .B1(n29118), .B2(
        \xmem_data[45][7] ), .ZN(n25339) );
  AOI22_X1 U28935 ( .A1(n25443), .A2(\xmem_data[46][7] ), .B1(n25442), .B2(
        \xmem_data[47][7] ), .ZN(n25338) );
  NAND4_X1 U28936 ( .A1(n25341), .A2(n25340), .A3(n25339), .A4(n25338), .ZN(
        n25352) );
  AOI22_X1 U28937 ( .A1(n25413), .A2(\xmem_data[48][7] ), .B1(n3218), .B2(
        \xmem_data[49][7] ), .ZN(n25345) );
  AOI22_X1 U28938 ( .A1(n25448), .A2(\xmem_data[50][7] ), .B1(n20558), .B2(
        \xmem_data[51][7] ), .ZN(n25344) );
  AOI22_X1 U28939 ( .A1(n25449), .A2(\xmem_data[52][7] ), .B1(n28372), .B2(
        \xmem_data[53][7] ), .ZN(n25343) );
  AOI22_X1 U28940 ( .A1(n25451), .A2(\xmem_data[54][7] ), .B1(n30877), .B2(
        \xmem_data[55][7] ), .ZN(n25342) );
  NAND4_X1 U28941 ( .A1(n25345), .A2(n25344), .A3(n25343), .A4(n25342), .ZN(
        n25351) );
  AOI22_X1 U28942 ( .A1(n25670), .A2(\xmem_data[56][7] ), .B1(n27943), .B2(
        \xmem_data[57][7] ), .ZN(n25349) );
  AOI22_X1 U28943 ( .A1(n25457), .A2(\xmem_data[58][7] ), .B1(n27452), .B2(
        \xmem_data[59][7] ), .ZN(n25348) );
  AOI22_X1 U28944 ( .A1(n25459), .A2(\xmem_data[60][7] ), .B1(n25458), .B2(
        \xmem_data[61][7] ), .ZN(n25347) );
  AOI22_X1 U28945 ( .A1(n20718), .A2(\xmem_data[62][7] ), .B1(n25460), .B2(
        \xmem_data[63][7] ), .ZN(n25346) );
  NAND4_X1 U28946 ( .A1(n25349), .A2(n25348), .A3(n25347), .A4(n25346), .ZN(
        n25350) );
  OR4_X1 U28947 ( .A1(n25353), .A2(n25352), .A3(n25351), .A4(n25350), .ZN(
        n25397) );
  NAND2_X1 U28948 ( .A1(n25354), .A2(\xmem_data[16][7] ), .ZN(n25356) );
  NAND2_X1 U28949 ( .A1(n3217), .A2(\xmem_data[17][7] ), .ZN(n25355) );
  NAND2_X1 U28950 ( .A1(n25356), .A2(n25355), .ZN(n25375) );
  AOI22_X1 U28951 ( .A1(n25358), .A2(\xmem_data[12][7] ), .B1(n25357), .B2(
        \xmem_data[13][7] ), .ZN(n25373) );
  AOI22_X1 U28952 ( .A1(n29151), .A2(\xmem_data[8][7] ), .B1(n25359), .B2(
        \xmem_data[9][7] ), .ZN(n25363) );
  AOI22_X1 U28953 ( .A1(n30864), .A2(\xmem_data[14][7] ), .B1(n25360), .B2(
        \xmem_data[15][7] ), .ZN(n25362) );
  NAND2_X1 U28954 ( .A1(n25514), .A2(\xmem_data[23][7] ), .ZN(n25361) );
  AOI22_X1 U28955 ( .A1(n30849), .A2(\xmem_data[4][7] ), .B1(n25364), .B2(
        \xmem_data[5][7] ), .ZN(n25372) );
  AOI22_X1 U28956 ( .A1(n29010), .A2(\xmem_data[0][7] ), .B1(n24645), .B2(
        \xmem_data[1][7] ), .ZN(n25366) );
  AOI22_X1 U28957 ( .A1(n25718), .A2(\xmem_data[6][7] ), .B1(n27975), .B2(
        \xmem_data[7][7] ), .ZN(n25365) );
  NAND2_X1 U28958 ( .A1(n25366), .A2(n25365), .ZN(n25370) );
  AOI22_X1 U28959 ( .A1(n17021), .A2(\xmem_data[2][7] ), .B1(n25367), .B2(
        \xmem_data[3][7] ), .ZN(n25368) );
  INV_X1 U28960 ( .A(n25368), .ZN(n25369) );
  NOR2_X1 U28961 ( .A1(n25370), .A2(n25369), .ZN(n25371) );
  NAND4_X1 U28962 ( .A1(n25373), .A2(n3910), .A3(n25372), .A4(n25371), .ZN(
        n25374) );
  NOR2_X1 U28963 ( .A1(n25375), .A2(n25374), .ZN(n25394) );
  AOI22_X1 U28964 ( .A1(n27904), .A2(\xmem_data[20][7] ), .B1(n24140), .B2(
        \xmem_data[21][7] ), .ZN(n25376) );
  INV_X1 U28965 ( .A(n25376), .ZN(n25381) );
  AOI22_X1 U28966 ( .A1(n24696), .A2(\xmem_data[18][7] ), .B1(n20598), .B2(
        \xmem_data[19][7] ), .ZN(n25379) );
  NAND2_X1 U28967 ( .A1(n25377), .A2(\xmem_data[22][7] ), .ZN(n25378) );
  NAND2_X1 U28968 ( .A1(n25379), .A2(n25378), .ZN(n25380) );
  AOI22_X1 U28969 ( .A1(n24638), .A2(\xmem_data[24][7] ), .B1(n13475), .B2(
        \xmem_data[25][7] ), .ZN(n25387) );
  AOI22_X1 U28970 ( .A1(n30744), .A2(\xmem_data[26][7] ), .B1(n17012), .B2(
        \xmem_data[27][7] ), .ZN(n25386) );
  AOI22_X1 U28971 ( .A1(n30514), .A2(\xmem_data[28][7] ), .B1(n25382), .B2(
        \xmem_data[29][7] ), .ZN(n25385) );
  AOI22_X1 U28972 ( .A1(n29807), .A2(\xmem_data[30][7] ), .B1(n25383), .B2(
        \xmem_data[31][7] ), .ZN(n25384) );
  NAND4_X1 U28973 ( .A1(n25387), .A2(n25386), .A3(n25385), .A4(n25384), .ZN(
        n25391) );
  AOI22_X1 U28974 ( .A1(n27568), .A2(\xmem_data[10][7] ), .B1(n25388), .B2(
        \xmem_data[11][7] ), .ZN(n25389) );
  INV_X1 U28975 ( .A(n25389), .ZN(n25390) );
  NOR3_X1 U28976 ( .A1(n3959), .A2(n25391), .A3(n25390), .ZN(n25393) );
  AOI21_X1 U28977 ( .B1(n25394), .B2(n25393), .A(n25392), .ZN(n25395) );
  AOI21_X1 U28978 ( .B1(n25397), .B2(n25396), .A(n25395), .ZN(n25475) );
  AOI22_X1 U28979 ( .A1(n23717), .A2(\xmem_data[96][7] ), .B1(n25398), .B2(
        \xmem_data[97][7] ), .ZN(n25405) );
  AOI22_X1 U28980 ( .A1(n25400), .A2(\xmem_data[98][7] ), .B1(n25399), .B2(
        \xmem_data[99][7] ), .ZN(n25404) );
  AOI22_X1 U28981 ( .A1(n21010), .A2(\xmem_data[100][7] ), .B1(n28327), .B2(
        \xmem_data[101][7] ), .ZN(n25403) );
  AOI22_X1 U28982 ( .A1(n25401), .A2(\xmem_data[102][7] ), .B1(n14975), .B2(
        \xmem_data[103][7] ), .ZN(n25402) );
  NAND4_X1 U28983 ( .A1(n25405), .A2(n25404), .A3(n25403), .A4(n25402), .ZN(
        n25433) );
  AOI22_X1 U28984 ( .A1(n20818), .A2(\xmem_data[104][7] ), .B1(n25406), .B2(
        \xmem_data[105][7] ), .ZN(n25412) );
  AOI22_X1 U28985 ( .A1(n25407), .A2(\xmem_data[106][7] ), .B1(n31344), .B2(
        \xmem_data[107][7] ), .ZN(n25411) );
  AOI22_X1 U28986 ( .A1(n25408), .A2(\xmem_data[108][7] ), .B1(n20578), .B2(
        \xmem_data[109][7] ), .ZN(n25410) );
  AOI22_X1 U28987 ( .A1(n3318), .A2(\xmem_data[110][7] ), .B1(n25485), .B2(
        \xmem_data[111][7] ), .ZN(n25409) );
  NAND4_X1 U28988 ( .A1(n25412), .A2(n25411), .A3(n25410), .A4(n25409), .ZN(
        n25432) );
  AOI22_X1 U28989 ( .A1(n25413), .A2(\xmem_data[112][7] ), .B1(n3222), .B2(
        \xmem_data[113][7] ), .ZN(n25421) );
  AOI22_X1 U28990 ( .A1(n25414), .A2(\xmem_data[114][7] ), .B1(n22667), .B2(
        \xmem_data[115][7] ), .ZN(n25420) );
  AOI22_X1 U28991 ( .A1(n25416), .A2(\xmem_data[116][7] ), .B1(n25415), .B2(
        \xmem_data[117][7] ), .ZN(n25419) );
  AOI22_X1 U28992 ( .A1(n25417), .A2(\xmem_data[118][7] ), .B1(n25492), .B2(
        \xmem_data[119][7] ), .ZN(n25418) );
  NAND4_X1 U28993 ( .A1(n25421), .A2(n25420), .A3(n25419), .A4(n25418), .ZN(
        n25431) );
  AOI22_X1 U28994 ( .A1(n25422), .A2(\xmem_data[120][7] ), .B1(n20588), .B2(
        \xmem_data[121][7] ), .ZN(n25429) );
  AOI22_X1 U28995 ( .A1(n25424), .A2(\xmem_data[122][7] ), .B1(n25423), .B2(
        \xmem_data[123][7] ), .ZN(n25428) );
  AOI22_X1 U28996 ( .A1(n25425), .A2(\xmem_data[124][7] ), .B1(n28052), .B2(
        \xmem_data[125][7] ), .ZN(n25427) );
  AOI22_X1 U28997 ( .A1(n17018), .A2(\xmem_data[126][7] ), .B1(n3213), .B2(
        \xmem_data[127][7] ), .ZN(n25426) );
  NAND4_X1 U28998 ( .A1(n25429), .A2(n25428), .A3(n25427), .A4(n25426), .ZN(
        n25430) );
  OR4_X1 U28999 ( .A1(n25433), .A2(n25432), .A3(n25431), .A4(n25430), .ZN(
        n25472) );
  AOI22_X1 U29000 ( .A1(n25434), .A2(\xmem_data[64][7] ), .B1(n23796), .B2(
        \xmem_data[65][7] ), .ZN(n25439) );
  AOI22_X1 U29001 ( .A1(n28994), .A2(\xmem_data[66][7] ), .B1(n25435), .B2(
        \xmem_data[67][7] ), .ZN(n25438) );
  AOI22_X1 U29002 ( .A1(n24461), .A2(\xmem_data[68][7] ), .B1(n25581), .B2(
        \xmem_data[69][7] ), .ZN(n25437) );
  AOI22_X1 U29003 ( .A1(n3308), .A2(\xmem_data[70][7] ), .B1(n22685), .B2(
        \xmem_data[71][7] ), .ZN(n25436) );
  NAND4_X1 U29004 ( .A1(n25439), .A2(n25438), .A3(n25437), .A4(n25436), .ZN(
        n25469) );
  AOI22_X1 U29005 ( .A1(n20734), .A2(\xmem_data[72][7] ), .B1(n28468), .B2(
        \xmem_data[73][7] ), .ZN(n25447) );
  AOI22_X1 U29006 ( .A1(n25407), .A2(\xmem_data[74][7] ), .B1(n25440), .B2(
        \xmem_data[75][7] ), .ZN(n25446) );
  AOI22_X1 U29007 ( .A1(n25441), .A2(\xmem_data[76][7] ), .B1(n29118), .B2(
        \xmem_data[77][7] ), .ZN(n25445) );
  AOI22_X1 U29008 ( .A1(n25443), .A2(\xmem_data[78][7] ), .B1(n25442), .B2(
        \xmem_data[79][7] ), .ZN(n25444) );
  NAND4_X1 U29009 ( .A1(n25447), .A2(n25446), .A3(n25445), .A4(n25444), .ZN(
        n25468) );
  AOI22_X1 U29010 ( .A1(n30592), .A2(\xmem_data[80][7] ), .B1(n3217), .B2(
        \xmem_data[81][7] ), .ZN(n25455) );
  AOI22_X1 U29011 ( .A1(n25448), .A2(\xmem_data[82][7] ), .B1(n24695), .B2(
        \xmem_data[83][7] ), .ZN(n25454) );
  AOI22_X1 U29012 ( .A1(n25449), .A2(\xmem_data[84][7] ), .B1(n13444), .B2(
        \xmem_data[85][7] ), .ZN(n25453) );
  AOI22_X1 U29013 ( .A1(n25451), .A2(\xmem_data[86][7] ), .B1(n28510), .B2(
        \xmem_data[87][7] ), .ZN(n25452) );
  NAND4_X1 U29014 ( .A1(n25455), .A2(n25454), .A3(n25453), .A4(n25452), .ZN(
        n25467) );
  AOI22_X1 U29015 ( .A1(n27508), .A2(\xmem_data[88][7] ), .B1(n27943), .B2(
        \xmem_data[89][7] ), .ZN(n25465) );
  AOI22_X1 U29016 ( .A1(n25457), .A2(\xmem_data[90][7] ), .B1(n13168), .B2(
        \xmem_data[91][7] ), .ZN(n25464) );
  AOI22_X1 U29017 ( .A1(n25459), .A2(\xmem_data[92][7] ), .B1(n25458), .B2(
        \xmem_data[93][7] ), .ZN(n25463) );
  AOI22_X1 U29018 ( .A1(n25461), .A2(\xmem_data[94][7] ), .B1(n25460), .B2(
        \xmem_data[95][7] ), .ZN(n25462) );
  NAND4_X1 U29019 ( .A1(n25465), .A2(n25464), .A3(n25463), .A4(n25462), .ZN(
        n25466) );
  OR4_X1 U29020 ( .A1(n25469), .A2(n25468), .A3(n25467), .A4(n25466), .ZN(
        n25470) );
  AOI22_X1 U29021 ( .A1(n25473), .A2(n25472), .B1(n25471), .B2(n25470), .ZN(
        n25474) );
  XNOR2_X1 U29022 ( .A(n35076), .B(\fmem_data[30][3] ), .ZN(n33232) );
  OAI22_X1 U29023 ( .A1(n33232), .A2(n34435), .B1(n31997), .B2(n34437), .ZN(
        n28933) );
  AOI22_X1 U29024 ( .A1(n14999), .A2(\xmem_data[16][7] ), .B1(n29008), .B2(
        \xmem_data[17][7] ), .ZN(n25479) );
  AOI22_X1 U29025 ( .A1(n22742), .A2(\xmem_data[18][7] ), .B1(n30949), .B2(
        \xmem_data[19][7] ), .ZN(n25478) );
  AOI22_X1 U29026 ( .A1(n29048), .A2(\xmem_data[20][7] ), .B1(n29239), .B2(
        \xmem_data[21][7] ), .ZN(n25477) );
  AOI22_X1 U29027 ( .A1(n20814), .A2(\xmem_data[22][7] ), .B1(n25521), .B2(
        \xmem_data[23][7] ), .ZN(n25476) );
  AOI22_X1 U29028 ( .A1(n29118), .A2(\xmem_data[0][7] ), .B1(n27813), .B2(
        \xmem_data[1][7] ), .ZN(n25480) );
  AOI22_X1 U29029 ( .A1(n25481), .A2(\xmem_data[12][7] ), .B1(n28233), .B2(
        \xmem_data[13][7] ), .ZN(n25482) );
  INV_X1 U29030 ( .A(n25482), .ZN(n25483) );
  AOI22_X1 U29031 ( .A1(n25485), .A2(\xmem_data[2][7] ), .B1(n24443), .B2(
        \xmem_data[3][7] ), .ZN(n25499) );
  AOI22_X1 U29032 ( .A1(n25486), .A2(\xmem_data[8][7] ), .B1(n3375), .B2(
        \xmem_data[9][7] ), .ZN(n25489) );
  AOI22_X1 U29033 ( .A1(n29232), .A2(\xmem_data[14][7] ), .B1(n27913), .B2(
        \xmem_data[15][7] ), .ZN(n25488) );
  NAND2_X1 U29034 ( .A1(n30885), .A2(\xmem_data[11][7] ), .ZN(n25487) );
  NAND3_X1 U29035 ( .A1(n25489), .A2(n25488), .A3(n25487), .ZN(n25497) );
  AOI22_X1 U29036 ( .A1(n25491), .A2(\xmem_data[6][7] ), .B1(n25490), .B2(
        \xmem_data[7][7] ), .ZN(n25495) );
  AOI22_X1 U29037 ( .A1(n3219), .A2(\xmem_data[4][7] ), .B1(n29422), .B2(
        \xmem_data[5][7] ), .ZN(n25494) );
  NAND2_X1 U29038 ( .A1(n25492), .A2(\xmem_data[10][7] ), .ZN(n25493) );
  NAND3_X1 U29039 ( .A1(n25495), .A2(n25494), .A3(n25493), .ZN(n25496) );
  AOI22_X1 U29040 ( .A1(n28327), .A2(\xmem_data[24][7] ), .B1(n29573), .B2(
        \xmem_data[25][7] ), .ZN(n25504) );
  AOI22_X1 U29041 ( .A1(n24167), .A2(\xmem_data[26][7] ), .B1(n3209), .B2(
        \xmem_data[27][7] ), .ZN(n25503) );
  AOI22_X1 U29042 ( .A1(n20733), .A2(\xmem_data[28][7] ), .B1(n20708), .B2(
        \xmem_data[29][7] ), .ZN(n25502) );
  AOI22_X1 U29043 ( .A1(n25528), .A2(\xmem_data[30][7] ), .B1(n30862), .B2(
        \xmem_data[31][7] ), .ZN(n25501) );
  NAND4_X1 U29044 ( .A1(n25504), .A2(n25503), .A3(n25502), .A4(n25501), .ZN(
        n25506) );
  AOI22_X1 U29045 ( .A1(n3203), .A2(\xmem_data[96][7] ), .B1(n3434), .B2(
        \xmem_data[97][7] ), .ZN(n25513) );
  AOI22_X1 U29046 ( .A1(n30589), .A2(\xmem_data[98][7] ), .B1(n25508), .B2(
        \xmem_data[99][7] ), .ZN(n25512) );
  AOI22_X1 U29047 ( .A1(n3217), .A2(\xmem_data[100][7] ), .B1(n27831), .B2(
        \xmem_data[101][7] ), .ZN(n25511) );
  AOI22_X1 U29048 ( .A1(n25509), .A2(\xmem_data[102][7] ), .B1(n25449), .B2(
        \xmem_data[103][7] ), .ZN(n25510) );
  NAND4_X1 U29049 ( .A1(n25513), .A2(n25512), .A3(n25511), .A4(n25510), .ZN(
        n25536) );
  AOI22_X1 U29050 ( .A1(n24564), .A2(\xmem_data[104][7] ), .B1(n30295), .B2(
        \xmem_data[105][7] ), .ZN(n25518) );
  AOI22_X1 U29051 ( .A1(n25514), .A2(\xmem_data[106][7] ), .B1(n28972), .B2(
        \xmem_data[107][7] ), .ZN(n25517) );
  AOI22_X1 U29052 ( .A1(n25481), .A2(\xmem_data[108][7] ), .B1(n30744), .B2(
        \xmem_data[109][7] ), .ZN(n25516) );
  AOI22_X1 U29053 ( .A1(n24516), .A2(\xmem_data[110][7] ), .B1(n30514), .B2(
        \xmem_data[111][7] ), .ZN(n25515) );
  NAND4_X1 U29054 ( .A1(n25518), .A2(n25517), .A3(n25516), .A4(n25515), .ZN(
        n25535) );
  AOI22_X1 U29055 ( .A1(n25671), .A2(\xmem_data[112][7] ), .B1(n25519), .B2(
        \xmem_data[113][7] ), .ZN(n25525) );
  AOI22_X1 U29056 ( .A1(n25460), .A2(\xmem_data[114][7] ), .B1(n25635), .B2(
        \xmem_data[115][7] ), .ZN(n25524) );
  AOI22_X1 U29057 ( .A1(n25520), .A2(\xmem_data[116][7] ), .B1(n28781), .B2(
        \xmem_data[117][7] ), .ZN(n25523) );
  AOI22_X1 U29058 ( .A1(n30871), .A2(\xmem_data[118][7] ), .B1(n25521), .B2(
        \xmem_data[119][7] ), .ZN(n25522) );
  NAND4_X1 U29059 ( .A1(n25525), .A2(n25524), .A3(n25523), .A4(n25522), .ZN(
        n25534) );
  AOI22_X1 U29060 ( .A1(n20943), .A2(\xmem_data[120][7] ), .B1(n24571), .B2(
        \xmem_data[121][7] ), .ZN(n25532) );
  AOI22_X1 U29061 ( .A1(n20553), .A2(\xmem_data[122][7] ), .B1(n25526), .B2(
        \xmem_data[123][7] ), .ZN(n25531) );
  AOI22_X1 U29062 ( .A1(n25527), .A2(\xmem_data[124][7] ), .B1(n20567), .B2(
        \xmem_data[125][7] ), .ZN(n25530) );
  AOI22_X1 U29063 ( .A1(n25528), .A2(\xmem_data[126][7] ), .B1(n27564), .B2(
        \xmem_data[127][7] ), .ZN(n25529) );
  NAND4_X1 U29064 ( .A1(n25532), .A2(n25531), .A3(n25530), .A4(n25529), .ZN(
        n25533) );
  OR4_X1 U29065 ( .A1(n25536), .A2(n25535), .A3(n25534), .A4(n25533), .ZN(
        n25559) );
  AOI22_X1 U29066 ( .A1(n25561), .A2(\xmem_data[64][7] ), .B1(n23732), .B2(
        \xmem_data[65][7] ), .ZN(n25540) );
  AOI22_X1 U29067 ( .A1(n27501), .A2(\xmem_data[66][7] ), .B1(n20518), .B2(
        \xmem_data[67][7] ), .ZN(n25539) );
  AOI22_X1 U29068 ( .A1(n3218), .A2(\xmem_data[68][7] ), .B1(n29627), .B2(
        \xmem_data[69][7] ), .ZN(n25538) );
  AOI22_X1 U29069 ( .A1(n25562), .A2(\xmem_data[70][7] ), .B1(n3341), .B2(
        \xmem_data[71][7] ), .ZN(n25537) );
  NAND4_X1 U29070 ( .A1(n25540), .A2(n25539), .A3(n25538), .A4(n25537), .ZN(
        n25556) );
  AOI22_X1 U29071 ( .A1(n30882), .A2(\xmem_data[72][7] ), .B1(n3138), .B2(
        \xmem_data[73][7] ), .ZN(n25544) );
  AOI22_X1 U29072 ( .A1(n27446), .A2(\xmem_data[74][7] ), .B1(n16974), .B2(
        \xmem_data[75][7] ), .ZN(n25543) );
  AOI22_X1 U29073 ( .A1(n20546), .A2(\xmem_data[76][7] ), .B1(n27944), .B2(
        \xmem_data[77][7] ), .ZN(n25542) );
  AOI22_X1 U29074 ( .A1(n14998), .A2(\xmem_data[78][7] ), .B1(n25567), .B2(
        \xmem_data[79][7] ), .ZN(n25541) );
  NAND4_X1 U29075 ( .A1(n25544), .A2(n25543), .A3(n25542), .A4(n25541), .ZN(
        n25555) );
  AOI22_X1 U29076 ( .A1(n23715), .A2(\xmem_data[80][7] ), .B1(n24213), .B2(
        \xmem_data[81][7] ), .ZN(n25548) );
  AOI22_X1 U29077 ( .A1(n25574), .A2(\xmem_data[82][7] ), .B1(n25573), .B2(
        \xmem_data[83][7] ), .ZN(n25547) );
  AOI22_X1 U29078 ( .A1(n31270), .A2(\xmem_data[84][7] ), .B1(n17044), .B2(
        \xmem_data[85][7] ), .ZN(n25546) );
  AOI22_X1 U29079 ( .A1(n25576), .A2(\xmem_data[86][7] ), .B1(n25575), .B2(
        \xmem_data[87][7] ), .ZN(n25545) );
  NAND4_X1 U29080 ( .A1(n25548), .A2(n25547), .A3(n25546), .A4(n25545), .ZN(
        n25554) );
  AOI22_X1 U29081 ( .A1(n25679), .A2(\xmem_data[88][7] ), .B1(n3307), .B2(
        \xmem_data[89][7] ), .ZN(n25552) );
  AOI22_X1 U29082 ( .A1(n25583), .A2(\xmem_data[90][7] ), .B1(n25582), .B2(
        \xmem_data[91][7] ), .ZN(n25551) );
  AOI22_X1 U29083 ( .A1(n28500), .A2(\xmem_data[92][7] ), .B1(n25584), .B2(
        \xmem_data[93][7] ), .ZN(n25550) );
  AOI22_X1 U29084 ( .A1(n30601), .A2(\xmem_data[94][7] ), .B1(n30909), .B2(
        \xmem_data[95][7] ), .ZN(n25549) );
  NAND4_X1 U29085 ( .A1(n25552), .A2(n25551), .A3(n25550), .A4(n25549), .ZN(
        n25553) );
  OR4_X1 U29086 ( .A1(n25556), .A2(n25555), .A3(n25554), .A4(n25553), .ZN(
        n25557) );
  AOI22_X1 U29087 ( .A1(n25560), .A2(n25559), .B1(n25558), .B2(n25557), .ZN(
        n25596) );
  AOI22_X1 U29088 ( .A1(n25561), .A2(\xmem_data[32][7] ), .B1(n3352), .B2(
        \xmem_data[33][7] ), .ZN(n25566) );
  AOI22_X1 U29089 ( .A1(n25687), .A2(\xmem_data[34][7] ), .B1(n24694), .B2(
        \xmem_data[35][7] ), .ZN(n25565) );
  AOI22_X1 U29090 ( .A1(n3220), .A2(\xmem_data[36][7] ), .B1(n31368), .B2(
        \xmem_data[37][7] ), .ZN(n25564) );
  AOI22_X1 U29091 ( .A1(n25562), .A2(\xmem_data[38][7] ), .B1(n3341), .B2(
        \xmem_data[39][7] ), .ZN(n25563) );
  NAND4_X1 U29092 ( .A1(n25566), .A2(n25565), .A3(n25564), .A4(n25563), .ZN(
        n25592) );
  AOI22_X1 U29093 ( .A1(n23811), .A2(\xmem_data[40][7] ), .B1(n30698), .B2(
        \xmem_data[41][7] ), .ZN(n25571) );
  AOI22_X1 U29094 ( .A1(n31252), .A2(\xmem_data[42][7] ), .B1(n23813), .B2(
        \xmem_data[43][7] ), .ZN(n25570) );
  AOI22_X1 U29095 ( .A1(n29180), .A2(\xmem_data[44][7] ), .B1(n24157), .B2(
        \xmem_data[45][7] ), .ZN(n25569) );
  AOI22_X1 U29096 ( .A1(n24555), .A2(\xmem_data[46][7] ), .B1(n25567), .B2(
        \xmem_data[47][7] ), .ZN(n25568) );
  NAND4_X1 U29097 ( .A1(n25571), .A2(n25570), .A3(n25569), .A4(n25568), .ZN(
        n25591) );
  AOI22_X1 U29098 ( .A1(n25572), .A2(\xmem_data[48][7] ), .B1(n30892), .B2(
        \xmem_data[49][7] ), .ZN(n25580) );
  AOI22_X1 U29099 ( .A1(n25574), .A2(\xmem_data[50][7] ), .B1(n25573), .B2(
        \xmem_data[51][7] ), .ZN(n25579) );
  AOI22_X1 U29100 ( .A1(n30544), .A2(\xmem_data[52][7] ), .B1(n31255), .B2(
        \xmem_data[53][7] ), .ZN(n25578) );
  AOI22_X1 U29101 ( .A1(n25576), .A2(\xmem_data[54][7] ), .B1(n25575), .B2(
        \xmem_data[55][7] ), .ZN(n25577) );
  NAND4_X1 U29102 ( .A1(n25580), .A2(n25579), .A3(n25578), .A4(n25577), .ZN(
        n25590) );
  AOI22_X1 U29103 ( .A1(n28429), .A2(\xmem_data[56][7] ), .B1(n28701), .B2(
        \xmem_data[57][7] ), .ZN(n25588) );
  AOI22_X1 U29104 ( .A1(n25583), .A2(\xmem_data[58][7] ), .B1(n25582), .B2(
        \xmem_data[59][7] ), .ZN(n25587) );
  AOI22_X1 U29105 ( .A1(n21057), .A2(\xmem_data[60][7] ), .B1(n25584), .B2(
        \xmem_data[61][7] ), .ZN(n25586) );
  AOI22_X1 U29106 ( .A1(n29125), .A2(\xmem_data[62][7] ), .B1(n24607), .B2(
        \xmem_data[63][7] ), .ZN(n25585) );
  NAND4_X1 U29107 ( .A1(n25588), .A2(n25587), .A3(n25586), .A4(n25585), .ZN(
        n25589) );
  OR4_X1 U29108 ( .A1(n25592), .A2(n25591), .A3(n25590), .A4(n25589), .ZN(
        n25594) );
  NAND2_X1 U29109 ( .A1(n25594), .A2(n25593), .ZN(n25595) );
  XNOR2_X1 U29110 ( .A(n35074), .B(\fmem_data[17][3] ), .ZN(n33248) );
  XNOR2_X1 U29111 ( .A(n31705), .B(\fmem_data[17][3] ), .ZN(n32645) );
  OAI22_X1 U29112 ( .A1(n33250), .A2(n33248), .B1(n32645), .B2(n33249), .ZN(
        n28932) );
  XNOR2_X1 U29113 ( .A(n3367), .B(\fmem_data[3][7] ), .ZN(n31815) );
  XNOR2_X1 U29114 ( .A(n3262), .B(\fmem_data[3][7] ), .ZN(n31982) );
  OAI22_X1 U29115 ( .A1(n31815), .A2(n35638), .B1(n31982), .B2(n35637), .ZN(
        n31779) );
  XNOR2_X1 U29116 ( .A(n35258), .B(\fmem_data[23][5] ), .ZN(n34907) );
  XNOR2_X1 U29117 ( .A(n35114), .B(\fmem_data[23][5] ), .ZN(n31941) );
  XOR2_X1 U29118 ( .A(\fmem_data[23][4] ), .B(\fmem_data[23][5] ), .Z(n25598)
         );
  OAI22_X1 U29119 ( .A1(n34907), .A2(n34909), .B1(n31941), .B2(n34908), .ZN(
        n31778) );
  XNOR2_X1 U29120 ( .A(n35110), .B(\fmem_data[31][5] ), .ZN(n31970) );
  XNOR2_X1 U29121 ( .A(n35256), .B(\fmem_data[31][5] ), .ZN(n34947) );
  OAI22_X1 U29122 ( .A1(n31970), .A2(n34945), .B1(n34947), .B2(n34944), .ZN(
        n31777) );
  FA_X1 U29123 ( .A(n25601), .B(n25600), .CI(n25599), .CO(n31784), .S(n26036)
         );
  XNOR2_X1 U29124 ( .A(n31799), .B(\fmem_data[14][3] ), .ZN(n31944) );
  OAI22_X1 U29125 ( .A1(n25602), .A2(n33741), .B1(n31944), .B2(n33603), .ZN(
        n29541) );
  XNOR2_X1 U29126 ( .A(n31663), .B(\fmem_data[12][3] ), .ZN(n33273) );
  OAI22_X1 U29127 ( .A1(n25603), .A2(n34340), .B1(n33273), .B2(n33582), .ZN(
        n29540) );
  AOI22_X1 U29128 ( .A1(n25604), .A2(\xmem_data[0][2] ), .B1(n3357), .B2(
        \xmem_data[1][2] ), .ZN(n25611) );
  AOI22_X1 U29129 ( .A1(n20716), .A2(\xmem_data[2][2] ), .B1(n25605), .B2(
        \xmem_data[3][2] ), .ZN(n25610) );
  AOI22_X1 U29130 ( .A1(n28980), .A2(\xmem_data[4][2] ), .B1(n25606), .B2(
        \xmem_data[5][2] ), .ZN(n25609) );
  AOI22_X1 U29131 ( .A1(n28516), .A2(\xmem_data[6][2] ), .B1(n28335), .B2(
        \xmem_data[7][2] ), .ZN(n25608) );
  AND4_X1 U29132 ( .A1(n25611), .A2(n25610), .A3(n25609), .A4(n25608), .ZN(
        n25615) );
  NAND2_X1 U29133 ( .A1(n28476), .A2(\xmem_data[27][2] ), .ZN(n25614) );
  NAND2_X1 U29134 ( .A1(n25612), .A2(\xmem_data[26][2] ), .ZN(n25613) );
  NAND2_X1 U29135 ( .A1(n25615), .A2(n4015), .ZN(n25622) );
  AOI22_X1 U29136 ( .A1(n24562), .A2(\xmem_data[24][2] ), .B1(n3221), .B2(
        \xmem_data[25][2] ), .ZN(n25620) );
  AOI22_X1 U29137 ( .A1(n25617), .A2(\xmem_data[28][2] ), .B1(n25616), .B2(
        \xmem_data[29][2] ), .ZN(n25619) );
  NAND2_X1 U29138 ( .A1(n30698), .A2(\xmem_data[30][2] ), .ZN(n25618) );
  NAND3_X1 U29139 ( .A1(n25620), .A2(n25619), .A3(n25618), .ZN(n25621) );
  AOI22_X1 U29140 ( .A1(n21058), .A2(\xmem_data[16][2] ), .B1(n27526), .B2(
        \xmem_data[17][2] ), .ZN(n25623) );
  AOI22_X1 U29141 ( .A1(n25624), .A2(\xmem_data[22][2] ), .B1(n30589), .B2(
        \xmem_data[23][2] ), .ZN(n25625) );
  AOI22_X1 U29142 ( .A1(n25628), .A2(\xmem_data[18][2] ), .B1(n10456), .B2(
        \xmem_data[19][2] ), .ZN(n25644) );
  AOI22_X1 U29143 ( .A1(n25630), .A2(\xmem_data[20][2] ), .B1(n25629), .B2(
        \xmem_data[21][2] ), .ZN(n25643) );
  AOI22_X1 U29144 ( .A1(n28781), .A2(\xmem_data[10][2] ), .B1(n27950), .B2(
        \xmem_data[11][2] ), .ZN(n25631) );
  INV_X1 U29145 ( .A(n25631), .ZN(n25641) );
  NAND2_X1 U29146 ( .A1(n25632), .A2(\xmem_data[12][2] ), .ZN(n25634) );
  NAND2_X1 U29147 ( .A1(n3372), .A2(\xmem_data[13][2] ), .ZN(n25633) );
  NAND2_X1 U29148 ( .A1(n25634), .A2(n25633), .ZN(n25640) );
  AOI22_X1 U29149 ( .A1(n25635), .A2(\xmem_data[8][2] ), .B1(n17043), .B2(
        \xmem_data[9][2] ), .ZN(n25638) );
  AOI22_X1 U29150 ( .A1(n25636), .A2(\xmem_data[14][2] ), .B1(n28062), .B2(
        \xmem_data[15][2] ), .ZN(n25637) );
  NAND2_X1 U29151 ( .A1(n25638), .A2(n25637), .ZN(n25639) );
  NOR3_X1 U29152 ( .A1(n25641), .A2(n25640), .A3(n25639), .ZN(n25642) );
  NAND4_X1 U29153 ( .A1(n25645), .A2(n25644), .A3(n25643), .A4(n25642), .ZN(
        n25646) );
  NOR2_X1 U29154 ( .A1(n25646), .A2(n3885), .ZN(n25648) );
  AOI21_X1 U29155 ( .B1(n3940), .B2(n25648), .A(n25647), .ZN(n25649) );
  INV_X1 U29156 ( .A(n25649), .ZN(n25745) );
  AOI22_X1 U29157 ( .A1(n25670), .A2(\xmem_data[96][2] ), .B1(n24130), .B2(
        \xmem_data[97][2] ), .ZN(n25653) );
  AOI22_X1 U29158 ( .A1(n17064), .A2(\xmem_data[98][2] ), .B1(n21075), .B2(
        \xmem_data[99][2] ), .ZN(n25652) );
  AOI22_X1 U29159 ( .A1(n20959), .A2(\xmem_data[100][2] ), .B1(n25671), .B2(
        \xmem_data[101][2] ), .ZN(n25651) );
  AOI22_X1 U29160 ( .A1(n25672), .A2(\xmem_data[102][2] ), .B1(n30615), .B2(
        \xmem_data[103][2] ), .ZN(n25650) );
  NAND4_X1 U29161 ( .A1(n25653), .A2(n25652), .A3(n25651), .A4(n25650), .ZN(
        n25669) );
  AOI22_X1 U29162 ( .A1(n23764), .A2(\xmem_data[104][2] ), .B1(n25677), .B2(
        \xmem_data[105][2] ), .ZN(n25657) );
  AOI22_X1 U29163 ( .A1(n25678), .A2(\xmem_data[106][2] ), .B1(n30616), .B2(
        \xmem_data[107][2] ), .ZN(n25656) );
  AOI22_X1 U29164 ( .A1(n28385), .A2(\xmem_data[108][2] ), .B1(n25679), .B2(
        \xmem_data[109][2] ), .ZN(n25655) );
  AOI22_X1 U29165 ( .A1(n3307), .A2(\xmem_data[110][2] ), .B1(n28495), .B2(
        \xmem_data[111][2] ), .ZN(n25654) );
  NAND4_X1 U29166 ( .A1(n25657), .A2(n25656), .A3(n25655), .A4(n25654), .ZN(
        n25668) );
  AOI22_X1 U29167 ( .A1(n25526), .A2(\xmem_data[112][2] ), .B1(n27526), .B2(
        \xmem_data[113][2] ), .ZN(n25661) );
  AOI22_X1 U29168 ( .A1(n25684), .A2(\xmem_data[114][2] ), .B1(n29125), .B2(
        \xmem_data[115][2] ), .ZN(n25660) );
  AOI22_X1 U29169 ( .A1(n25686), .A2(\xmem_data[116][2] ), .B1(n25685), .B2(
        \xmem_data[117][2] ), .ZN(n25659) );
  AOI22_X1 U29170 ( .A1(n3228), .A2(\xmem_data[118][2] ), .B1(n25687), .B2(
        \xmem_data[119][2] ), .ZN(n25658) );
  NAND4_X1 U29171 ( .A1(n25661), .A2(n25660), .A3(n25659), .A4(n25658), .ZN(
        n25667) );
  AOI22_X1 U29172 ( .A1(n25692), .A2(\xmem_data[120][2] ), .B1(n3221), .B2(
        \xmem_data[121][2] ), .ZN(n25665) );
  AOI22_X1 U29173 ( .A1(n25693), .A2(\xmem_data[122][2] ), .B1(n25509), .B2(
        \xmem_data[123][2] ), .ZN(n25664) );
  AOI22_X1 U29174 ( .A1(n25694), .A2(\xmem_data[124][2] ), .B1(n13444), .B2(
        \xmem_data[125][2] ), .ZN(n25663) );
  AOI22_X1 U29175 ( .A1(n3374), .A2(\xmem_data[126][2] ), .B1(n13474), .B2(
        \xmem_data[127][2] ), .ZN(n25662) );
  NAND4_X1 U29176 ( .A1(n25665), .A2(n25664), .A3(n25663), .A4(n25662), .ZN(
        n25666) );
  AOI22_X1 U29177 ( .A1(n25670), .A2(\xmem_data[64][2] ), .B1(n27988), .B2(
        \xmem_data[65][2] ), .ZN(n25676) );
  AOI22_X1 U29178 ( .A1(n24157), .A2(\xmem_data[66][2] ), .B1(n23761), .B2(
        \xmem_data[67][2] ), .ZN(n25675) );
  AOI22_X1 U29179 ( .A1(n25425), .A2(\xmem_data[68][2] ), .B1(n25671), .B2(
        \xmem_data[69][2] ), .ZN(n25674) );
  AOI22_X1 U29180 ( .A1(n25672), .A2(\xmem_data[70][2] ), .B1(n22677), .B2(
        \xmem_data[71][2] ), .ZN(n25673) );
  NAND4_X1 U29181 ( .A1(n25676), .A2(n25675), .A3(n25674), .A4(n25673), .ZN(
        n25702) );
  AOI22_X1 U29182 ( .A1(n17020), .A2(\xmem_data[72][2] ), .B1(n25677), .B2(
        \xmem_data[73][2] ), .ZN(n25683) );
  AOI22_X1 U29183 ( .A1(n25678), .A2(\xmem_data[74][2] ), .B1(n24116), .B2(
        \xmem_data[75][2] ), .ZN(n25682) );
  AOI22_X1 U29184 ( .A1(n25632), .A2(\xmem_data[76][2] ), .B1(n28327), .B2(
        \xmem_data[77][2] ), .ZN(n25681) );
  AOI22_X1 U29185 ( .A1(n3307), .A2(\xmem_data[78][2] ), .B1(n24622), .B2(
        \xmem_data[79][2] ), .ZN(n25680) );
  NAND4_X1 U29186 ( .A1(n25683), .A2(n25682), .A3(n25681), .A4(n25680), .ZN(
        n25701) );
  AOI22_X1 U29187 ( .A1(n25582), .A2(\xmem_data[80][2] ), .B1(n29017), .B2(
        \xmem_data[81][2] ), .ZN(n25691) );
  AOI22_X1 U29188 ( .A1(n25684), .A2(\xmem_data[82][2] ), .B1(n16999), .B2(
        \xmem_data[83][2] ), .ZN(n25690) );
  AOI22_X1 U29189 ( .A1(n25686), .A2(\xmem_data[84][2] ), .B1(n25685), .B2(
        \xmem_data[85][2] ), .ZN(n25689) );
  AOI22_X1 U29190 ( .A1(n3433), .A2(\xmem_data[86][2] ), .B1(n25687), .B2(
        \xmem_data[87][2] ), .ZN(n25688) );
  NAND4_X1 U29191 ( .A1(n25691), .A2(n25690), .A3(n25689), .A4(n25688), .ZN(
        n25700) );
  AOI22_X1 U29192 ( .A1(n25692), .A2(\xmem_data[88][2] ), .B1(n3217), .B2(
        \xmem_data[89][2] ), .ZN(n25698) );
  AOI22_X1 U29193 ( .A1(n25693), .A2(\xmem_data[90][2] ), .B1(n20723), .B2(
        \xmem_data[91][2] ), .ZN(n25697) );
  AOI22_X1 U29194 ( .A1(n25694), .A2(\xmem_data[92][2] ), .B1(n13444), .B2(
        \xmem_data[93][2] ), .ZN(n25696) );
  AOI22_X1 U29195 ( .A1(n25417), .A2(\xmem_data[94][2] ), .B1(n13474), .B2(
        \xmem_data[95][2] ), .ZN(n25695) );
  NAND4_X1 U29196 ( .A1(n25698), .A2(n25697), .A3(n25696), .A4(n25695), .ZN(
        n25699) );
  OR4_X1 U29197 ( .A1(n25702), .A2(n25701), .A3(n25700), .A4(n25699), .ZN(
        n25703) );
  AOI22_X1 U29198 ( .A1(n25706), .A2(n25705), .B1(n25704), .B2(n25703), .ZN(
        n25744) );
  AOI22_X1 U29199 ( .A1(n25707), .A2(\xmem_data[32][2] ), .B1(n28373), .B2(
        \xmem_data[33][2] ), .ZN(n25714) );
  AOI22_X1 U29200 ( .A1(n25708), .A2(\xmem_data[34][2] ), .B1(n28375), .B2(
        \xmem_data[35][2] ), .ZN(n25713) );
  AOI22_X1 U29201 ( .A1(n20495), .A2(\xmem_data[36][2] ), .B1(n25709), .B2(
        \xmem_data[37][2] ), .ZN(n25712) );
  AOI22_X1 U29202 ( .A1(n3466), .A2(\xmem_data[38][2] ), .B1(n25383), .B2(
        \xmem_data[39][2] ), .ZN(n25711) );
  NAND4_X1 U29203 ( .A1(n25714), .A2(n25713), .A3(n25712), .A4(n25711), .ZN(
        n25740) );
  AOI22_X1 U29204 ( .A1(n25573), .A2(\xmem_data[40][2] ), .B1(n25715), .B2(
        \xmem_data[41][2] ), .ZN(n25722) );
  AOI22_X1 U29205 ( .A1(n28302), .A2(\xmem_data[42][2] ), .B1(n30871), .B2(
        \xmem_data[43][2] ), .ZN(n25721) );
  AOI22_X1 U29206 ( .A1(n17002), .A2(\xmem_data[44][2] ), .B1(n21009), .B2(
        \xmem_data[45][2] ), .ZN(n25720) );
  AOI22_X1 U29207 ( .A1(n25718), .A2(\xmem_data[46][2] ), .B1(n27365), .B2(
        \xmem_data[47][2] ), .ZN(n25719) );
  NAND4_X1 U29208 ( .A1(n25722), .A2(n25721), .A3(n25720), .A4(n25719), .ZN(
        n25739) );
  AOI22_X1 U29209 ( .A1(n25582), .A2(\xmem_data[48][2] ), .B1(n25723), .B2(
        \xmem_data[49][2] ), .ZN(n25729) );
  AOI22_X1 U29210 ( .A1(n27498), .A2(\xmem_data[50][2] ), .B1(n31344), .B2(
        \xmem_data[51][2] ), .ZN(n25728) );
  AOI22_X1 U29211 ( .A1(n25724), .A2(\xmem_data[52][2] ), .B1(n28366), .B2(
        \xmem_data[53][2] ), .ZN(n25727) );
  AOI22_X1 U29212 ( .A1(n25725), .A2(\xmem_data[54][2] ), .B1(n27501), .B2(
        \xmem_data[55][2] ), .ZN(n25726) );
  NAND4_X1 U29213 ( .A1(n25729), .A2(n25728), .A3(n25727), .A4(n25726), .ZN(
        n25738) );
  AOI22_X1 U29214 ( .A1(n25730), .A2(\xmem_data[56][2] ), .B1(n3220), .B2(
        \xmem_data[57][2] ), .ZN(n25736) );
  AOI22_X1 U29215 ( .A1(n25731), .A2(\xmem_data[58][2] ), .B1(n29095), .B2(
        \xmem_data[59][2] ), .ZN(n25735) );
  AOI22_X1 U29216 ( .A1(n20725), .A2(\xmem_data[60][2] ), .B1(n20993), .B2(
        \xmem_data[61][2] ), .ZN(n25734) );
  AOI22_X1 U29217 ( .A1(n25732), .A2(\xmem_data[62][2] ), .B1(n3231), .B2(
        \xmem_data[63][2] ), .ZN(n25733) );
  NAND4_X1 U29218 ( .A1(n25736), .A2(n25735), .A3(n25734), .A4(n25733), .ZN(
        n25737) );
  OR4_X1 U29219 ( .A1(n25740), .A2(n25739), .A3(n25738), .A4(n25737), .ZN(
        n25742) );
  NAND2_X1 U29220 ( .A1(n25742), .A2(n25741), .ZN(n25743) );
  XNOR2_X1 U29221 ( .A(n32117), .B(\fmem_data[6][7] ), .ZN(n32001) );
  OAI22_X1 U29222 ( .A1(n25746), .A2(n35512), .B1(n35511), .B2(n32001), .ZN(
        n29539) );
  XNOR2_X1 U29223 ( .A(n35106), .B(\fmem_data[26][3] ), .ZN(n32021) );
  OAI22_X1 U29224 ( .A1(n30381), .A2(n35507), .B1(n25747), .B2(n35508), .ZN(
        n26031) );
  AOI22_X1 U29225 ( .A1(n30295), .A2(\xmem_data[32][7] ), .B1(n28007), .B2(
        \xmem_data[33][7] ), .ZN(n25751) );
  AOI22_X1 U29226 ( .A1(n30885), .A2(\xmem_data[34][7] ), .B1(n29307), .B2(
        \xmem_data[35][7] ), .ZN(n25750) );
  AOI22_X1 U29227 ( .A1(n29308), .A2(\xmem_data[36][7] ), .B1(n31326), .B2(
        \xmem_data[37][7] ), .ZN(n25749) );
  AOI22_X1 U29228 ( .A1(n29310), .A2(\xmem_data[38][7] ), .B1(n29309), .B2(
        \xmem_data[39][7] ), .ZN(n25748) );
  NAND4_X1 U29229 ( .A1(n25751), .A2(n25750), .A3(n25749), .A4(n25748), .ZN(
        n25768) );
  AOI22_X1 U29230 ( .A1(n30746), .A2(\xmem_data[40][7] ), .B1(n3207), .B2(
        \xmem_data[41][7] ), .ZN(n25755) );
  AOI22_X1 U29231 ( .A1(n29317), .A2(\xmem_data[42][7] ), .B1(n29316), .B2(
        \xmem_data[43][7] ), .ZN(n25754) );
  AOI22_X1 U29232 ( .A1(n29319), .A2(\xmem_data[44][7] ), .B1(n29318), .B2(
        \xmem_data[45][7] ), .ZN(n25753) );
  AOI22_X1 U29233 ( .A1(n28385), .A2(\xmem_data[46][7] ), .B1(n23778), .B2(
        \xmem_data[47][7] ), .ZN(n25752) );
  NAND4_X1 U29234 ( .A1(n25755), .A2(n25754), .A3(n25753), .A4(n25752), .ZN(
        n25767) );
  AOI22_X1 U29235 ( .A1(n29324), .A2(\xmem_data[48][7] ), .B1(n14975), .B2(
        \xmem_data[49][7] ), .ZN(n25760) );
  AOI22_X1 U29236 ( .A1(n29325), .A2(\xmem_data[50][7] ), .B1(n20733), .B2(
        \xmem_data[51][7] ), .ZN(n25759) );
  AND2_X1 U29237 ( .A1(n29326), .A2(\xmem_data[53][7] ), .ZN(n25756) );
  AOI21_X1 U29238 ( .B1(n29327), .B2(\xmem_data[52][7] ), .A(n25756), .ZN(
        n25758) );
  AOI22_X1 U29239 ( .A1(n20953), .A2(\xmem_data[54][7] ), .B1(n29328), .B2(
        \xmem_data[55][7] ), .ZN(n25757) );
  NAND4_X1 U29240 ( .A1(n25760), .A2(n25759), .A3(n25758), .A4(n25757), .ZN(
        n25766) );
  AOI22_X1 U29241 ( .A1(n3382), .A2(\xmem_data[56][7] ), .B1(n25360), .B2(
        \xmem_data[57][7] ), .ZN(n25764) );
  AOI22_X1 U29242 ( .A1(n24532), .A2(\xmem_data[58][7] ), .B1(n3218), .B2(
        \xmem_data[59][7] ), .ZN(n25763) );
  AOI22_X1 U29243 ( .A1(n24139), .A2(\xmem_data[60][7] ), .B1(n30534), .B2(
        \xmem_data[61][7] ), .ZN(n25762) );
  AOI22_X1 U29244 ( .A1(n29027), .A2(\xmem_data[62][7] ), .B1(n29104), .B2(
        \xmem_data[63][7] ), .ZN(n25761) );
  NAND4_X1 U29245 ( .A1(n25764), .A2(n25763), .A3(n25762), .A4(n25761), .ZN(
        n25765) );
  OR4_X1 U29246 ( .A1(n25768), .A2(n25767), .A3(n25766), .A4(n25765), .ZN(
        n25791) );
  AOI22_X1 U29247 ( .A1(n3135), .A2(\xmem_data[0][7] ), .B1(n29103), .B2(
        \xmem_data[1][7] ), .ZN(n25772) );
  AOI22_X1 U29248 ( .A1(n25422), .A2(\xmem_data[2][7] ), .B1(n3358), .B2(
        \xmem_data[3][7] ), .ZN(n25771) );
  AOI22_X1 U29249 ( .A1(n27911), .A2(\xmem_data[4][7] ), .B1(n25605), .B2(
        \xmem_data[5][7] ), .ZN(n25770) );
  AOI22_X1 U29250 ( .A1(n29272), .A2(\xmem_data[6][7] ), .B1(n29271), .B2(
        \xmem_data[7][7] ), .ZN(n25769) );
  NAND4_X1 U29251 ( .A1(n25772), .A2(n25771), .A3(n25770), .A4(n25769), .ZN(
        n25788) );
  AOI22_X1 U29252 ( .A1(n30543), .A2(\xmem_data[8][7] ), .B1(n29279), .B2(
        \xmem_data[9][7] ), .ZN(n25776) );
  AOI22_X1 U29253 ( .A1(n25573), .A2(\xmem_data[10][7] ), .B1(n25715), .B2(
        \xmem_data[11][7] ), .ZN(n25775) );
  AOI22_X1 U29254 ( .A1(n29047), .A2(\xmem_data[12][7] ), .B1(n29280), .B2(
        \xmem_data[13][7] ), .ZN(n25774) );
  AOI22_X1 U29255 ( .A1(n28385), .A2(\xmem_data[14][7] ), .B1(n29281), .B2(
        \xmem_data[15][7] ), .ZN(n25773) );
  NAND4_X1 U29256 ( .A1(n25776), .A2(n25775), .A3(n25774), .A4(n25773), .ZN(
        n25787) );
  AOI22_X1 U29257 ( .A1(n29297), .A2(\xmem_data[16][7] ), .B1(n20983), .B2(
        \xmem_data[17][7] ), .ZN(n25780) );
  AOI22_X1 U29258 ( .A1(n24572), .A2(\xmem_data[18][7] ), .B1(n28328), .B2(
        \xmem_data[19][7] ), .ZN(n25779) );
  AOI22_X1 U29259 ( .A1(n29298), .A2(\xmem_data[20][7] ), .B1(n29326), .B2(
        \xmem_data[21][7] ), .ZN(n25778) );
  AOI22_X1 U29260 ( .A1(n29057), .A2(\xmem_data[22][7] ), .B1(n28037), .B2(
        \xmem_data[23][7] ), .ZN(n25777) );
  NAND4_X1 U29261 ( .A1(n25780), .A2(n25779), .A3(n25778), .A4(n25777), .ZN(
        n25786) );
  AOI22_X1 U29262 ( .A1(n3335), .A2(\xmem_data[24][7] ), .B1(n29286), .B2(
        \xmem_data[25][7] ), .ZN(n25784) );
  AOI22_X1 U29263 ( .A1(n29064), .A2(\xmem_data[26][7] ), .B1(n3221), .B2(
        \xmem_data[27][7] ), .ZN(n25783) );
  AOI22_X1 U29264 ( .A1(n29288), .A2(\xmem_data[28][7] ), .B1(n27869), .B2(
        \xmem_data[29][7] ), .ZN(n25782) );
  AOI22_X1 U29265 ( .A1(n29289), .A2(\xmem_data[30][7] ), .B1(n3255), .B2(
        \xmem_data[31][7] ), .ZN(n25781) );
  NAND4_X1 U29266 ( .A1(n25784), .A2(n25783), .A3(n25782), .A4(n25781), .ZN(
        n25785) );
  OR4_X1 U29267 ( .A1(n25788), .A2(n25787), .A3(n25786), .A4(n25785), .ZN(
        n25789) );
  AOI22_X1 U29268 ( .A1(n29343), .A2(n25791), .B1(n25790), .B2(n25789), .ZN(
        n25837) );
  AOI22_X1 U29269 ( .A1(n29762), .A2(\xmem_data[64][7] ), .B1(n3231), .B2(
        \xmem_data[65][7] ), .ZN(n25795) );
  AOI22_X1 U29270 ( .A1(n27508), .A2(\xmem_data[66][7] ), .B1(n29307), .B2(
        \xmem_data[67][7] ), .ZN(n25794) );
  AOI22_X1 U29271 ( .A1(n29308), .A2(\xmem_data[68][7] ), .B1(n27535), .B2(
        \xmem_data[69][7] ), .ZN(n25793) );
  AOI22_X1 U29272 ( .A1(n29310), .A2(\xmem_data[70][7] ), .B1(n29309), .B2(
        \xmem_data[71][7] ), .ZN(n25792) );
  NAND4_X1 U29273 ( .A1(n25795), .A2(n25794), .A3(n25793), .A4(n25792), .ZN(
        n25812) );
  AOI22_X1 U29274 ( .A1(n29237), .A2(\xmem_data[72][7] ), .B1(n24134), .B2(
        \xmem_data[73][7] ), .ZN(n25799) );
  AOI22_X1 U29275 ( .A1(n29317), .A2(\xmem_data[74][7] ), .B1(n29316), .B2(
        \xmem_data[75][7] ), .ZN(n25798) );
  AOI22_X1 U29276 ( .A1(n29319), .A2(\xmem_data[76][7] ), .B1(n29318), .B2(
        \xmem_data[77][7] ), .ZN(n25797) );
  AOI22_X1 U29277 ( .A1(n27974), .A2(\xmem_data[78][7] ), .B1(n30598), .B2(
        \xmem_data[79][7] ), .ZN(n25796) );
  NAND4_X1 U29278 ( .A1(n25799), .A2(n25798), .A3(n25797), .A4(n25796), .ZN(
        n25811) );
  AOI22_X1 U29279 ( .A1(n29324), .A2(\xmem_data[80][7] ), .B1(n14975), .B2(
        \xmem_data[81][7] ), .ZN(n25804) );
  AOI22_X1 U29280 ( .A1(n29325), .A2(\xmem_data[82][7] ), .B1(n28979), .B2(
        \xmem_data[83][7] ), .ZN(n25803) );
  AOI22_X1 U29281 ( .A1(n29327), .A2(\xmem_data[84][7] ), .B1(n29326), .B2(
        \xmem_data[85][7] ), .ZN(n25802) );
  AND2_X1 U29282 ( .A1(n29124), .A2(\xmem_data[86][7] ), .ZN(n25800) );
  AOI21_X1 U29283 ( .B1(n29328), .B2(\xmem_data[87][7] ), .A(n25800), .ZN(
        n25801) );
  NAND4_X1 U29284 ( .A1(n25804), .A2(n25803), .A3(n25802), .A4(n25801), .ZN(
        n25810) );
  AOI22_X1 U29285 ( .A1(n3383), .A2(\xmem_data[88][7] ), .B1(n31347), .B2(
        \xmem_data[89][7] ), .ZN(n25808) );
  AOI22_X1 U29286 ( .A1(n20576), .A2(\xmem_data[90][7] ), .B1(n3222), .B2(
        \xmem_data[91][7] ), .ZN(n25807) );
  AOI22_X1 U29287 ( .A1(n25693), .A2(\xmem_data[92][7] ), .B1(n25509), .B2(
        \xmem_data[93][7] ), .ZN(n25806) );
  AOI22_X1 U29288 ( .A1(n20994), .A2(\xmem_data[94][7] ), .B1(n20806), .B2(
        \xmem_data[95][7] ), .ZN(n25805) );
  NAND4_X1 U29289 ( .A1(n25808), .A2(n25807), .A3(n25806), .A4(n25805), .ZN(
        n25809) );
  OR4_X1 U29290 ( .A1(n25812), .A2(n25811), .A3(n25810), .A4(n25809), .ZN(
        n25813) );
  NAND2_X1 U29291 ( .A1(n25813), .A2(n29267), .ZN(n25836) );
  AOI22_X1 U29292 ( .A1(n28973), .A2(\xmem_data[120][7] ), .B1(n29253), .B2(
        \xmem_data[121][7] ), .ZN(n25817) );
  AOI22_X1 U29293 ( .A1(n29254), .A2(\xmem_data[122][7] ), .B1(n3220), .B2(
        \xmem_data[123][7] ), .ZN(n25816) );
  AOI22_X1 U29294 ( .A1(n29256), .A2(\xmem_data[124][7] ), .B1(n29255), .B2(
        \xmem_data[125][7] ), .ZN(n25815) );
  AOI22_X1 U29295 ( .A1(n29257), .A2(\xmem_data[126][7] ), .B1(n25616), .B2(
        \xmem_data[127][7] ), .ZN(n25814) );
  NAND4_X1 U29296 ( .A1(n25817), .A2(n25816), .A3(n25815), .A4(n25814), .ZN(
        n25833) );
  AOI22_X1 U29297 ( .A1(n29246), .A2(\xmem_data[112][7] ), .B1(n29245), .B2(
        \xmem_data[113][7] ), .ZN(n25821) );
  AOI22_X1 U29298 ( .A1(n29325), .A2(\xmem_data[114][7] ), .B1(n29247), .B2(
        \xmem_data[115][7] ), .ZN(n25820) );
  AOI22_X1 U29299 ( .A1(n30674), .A2(\xmem_data[116][7] ), .B1(n29248), .B2(
        \xmem_data[117][7] ), .ZN(n25819) );
  AOI22_X1 U29300 ( .A1(n27564), .A2(\xmem_data[118][7] ), .B1(n31262), .B2(
        \xmem_data[119][7] ), .ZN(n25818) );
  NAND4_X1 U29301 ( .A1(n25821), .A2(n25820), .A3(n25819), .A4(n25818), .ZN(
        n25832) );
  AOI22_X1 U29302 ( .A1(n29231), .A2(\xmem_data[96][7] ), .B1(n25450), .B2(
        \xmem_data[97][7] ), .ZN(n25825) );
  AOI22_X1 U29303 ( .A1(n27447), .A2(\xmem_data[98][7] ), .B1(n3357), .B2(
        \xmem_data[99][7] ), .ZN(n25824) );
  AOI22_X1 U29304 ( .A1(n22738), .A2(\xmem_data[100][7] ), .B1(n29232), .B2(
        \xmem_data[101][7] ), .ZN(n25823) );
  AOI22_X1 U29305 ( .A1(n25710), .A2(\xmem_data[102][7] ), .B1(n22703), .B2(
        \xmem_data[103][7] ), .ZN(n25822) );
  NAND4_X1 U29306 ( .A1(n25825), .A2(n25824), .A3(n25823), .A4(n25822), .ZN(
        n25831) );
  AOI22_X1 U29307 ( .A1(n23795), .A2(\xmem_data[104][7] ), .B1(n24457), .B2(
        \xmem_data[105][7] ), .ZN(n25829) );
  AOI22_X1 U29308 ( .A1(n23717), .A2(\xmem_data[106][7] ), .B1(n17043), .B2(
        \xmem_data[107][7] ), .ZN(n25828) );
  AOI22_X1 U29309 ( .A1(n29239), .A2(\xmem_data[108][7] ), .B1(n29238), .B2(
        \xmem_data[109][7] ), .ZN(n25827) );
  AOI22_X1 U29310 ( .A1(n29240), .A2(\xmem_data[110][7] ), .B1(n20551), .B2(
        \xmem_data[111][7] ), .ZN(n25826) );
  NAND4_X1 U29311 ( .A1(n25829), .A2(n25828), .A3(n25827), .A4(n25826), .ZN(
        n25830) );
  OR4_X1 U29312 ( .A1(n25833), .A2(n25832), .A3(n25831), .A4(n25830), .ZN(
        n25834) );
  NAND2_X1 U29313 ( .A1(n25834), .A2(n29269), .ZN(n25835) );
  XNOR2_X1 U29314 ( .A(n35328), .B(\fmem_data[8][3] ), .ZN(n33062) );
  XOR2_X1 U29315 ( .A(\fmem_data[8][2] ), .B(\fmem_data[8][3] ), .Z(n25838) );
  AND2_X1 U29316 ( .A1(n34208), .A2(n34206), .ZN(n25839) );
  XNOR2_X1 U29317 ( .A(n3272), .B(\fmem_data[31][7] ), .ZN(n35111) );
  XNOR2_X1 U29318 ( .A(n3320), .B(\fmem_data[31][7] ), .ZN(n31974) );
  AOI22_X1 U29319 ( .A1(n28700), .A2(\xmem_data[106][5] ), .B1(n28733), .B2(
        \xmem_data[107][5] ), .ZN(n25841) );
  AOI22_X1 U29320 ( .A1(n29433), .A2(\xmem_data[104][5] ), .B1(n30100), .B2(
        \xmem_data[105][5] ), .ZN(n25840) );
  NAND2_X1 U29321 ( .A1(n25841), .A2(n25840), .ZN(n25847) );
  AOI22_X1 U29322 ( .A1(n29390), .A2(\xmem_data[112][5] ), .B1(n30662), .B2(
        \xmem_data[113][5] ), .ZN(n25845) );
  AOI22_X1 U29323 ( .A1(n30664), .A2(\xmem_data[114][5] ), .B1(n30663), .B2(
        \xmem_data[115][5] ), .ZN(n25844) );
  AOI22_X1 U29324 ( .A1(n27754), .A2(\xmem_data[116][5] ), .B1(n26884), .B2(
        \xmem_data[117][5] ), .ZN(n25843) );
  AOI22_X1 U29325 ( .A1(n30667), .A2(\xmem_data[118][5] ), .B1(n29396), .B2(
        \xmem_data[119][5] ), .ZN(n25842) );
  NAND4_X1 U29326 ( .A1(n25845), .A2(n25844), .A3(n25843), .A4(n25842), .ZN(
        n25846) );
  OR2_X1 U29327 ( .A1(n25847), .A2(n25846), .ZN(n25861) );
  AOI22_X1 U29328 ( .A1(n30673), .A2(\xmem_data[96][5] ), .B1(n30672), .B2(
        \xmem_data[97][5] ), .ZN(n25851) );
  AOI22_X1 U29329 ( .A1(n30675), .A2(\xmem_data[98][5] ), .B1(n30674), .B2(
        \xmem_data[99][5] ), .ZN(n25850) );
  AOI22_X1 U29330 ( .A1(n30677), .A2(\xmem_data[100][5] ), .B1(n30676), .B2(
        \xmem_data[101][5] ), .ZN(n25849) );
  AOI22_X1 U29331 ( .A1(n30678), .A2(\xmem_data[102][5] ), .B1(n28164), .B2(
        \xmem_data[103][5] ), .ZN(n25848) );
  AOI22_X1 U29332 ( .A1(n3162), .A2(\xmem_data[120][5] ), .B1(n3182), .B2(
        \xmem_data[121][5] ), .ZN(n25854) );
  AOI22_X1 U29333 ( .A1(n30687), .A2(\xmem_data[126][5] ), .B1(n30686), .B2(
        \xmem_data[127][5] ), .ZN(n25853) );
  AOI22_X1 U29334 ( .A1(n30699), .A2(\xmem_data[110][5] ), .B1(n30698), .B2(
        \xmem_data[111][5] ), .ZN(n25852) );
  NOR2_X1 U29335 ( .A1(n3970), .A2(n25855), .ZN(n25859) );
  AOI22_X1 U29336 ( .A1(n30697), .A2(\xmem_data[108][5] ), .B1(n30696), .B2(
        \xmem_data[109][5] ), .ZN(n25858) );
  AOI22_X1 U29337 ( .A1(n30764), .A2(\xmem_data[122][5] ), .B1(n28232), .B2(
        \xmem_data[123][5] ), .ZN(n25857) );
  AOI22_X1 U29338 ( .A1(n29488), .A2(\xmem_data[124][5] ), .B1(n29487), .B2(
        \xmem_data[125][5] ), .ZN(n25856) );
  NAND4_X1 U29339 ( .A1(n25859), .A2(n25858), .A3(n25857), .A4(n25856), .ZN(
        n25860) );
  OAI21_X1 U29340 ( .B1(n25861), .B2(n25860), .A(n30659), .ZN(n25936) );
  AOI22_X1 U29341 ( .A1(n30777), .A2(\xmem_data[76][5] ), .B1(n27833), .B2(
        \xmem_data[77][5] ), .ZN(n25882) );
  AOI22_X1 U29342 ( .A1(n30753), .A2(\xmem_data[64][5] ), .B1(n30752), .B2(
        \xmem_data[65][5] ), .ZN(n25865) );
  AOI22_X1 U29343 ( .A1(n30755), .A2(\xmem_data[66][5] ), .B1(n30754), .B2(
        \xmem_data[67][5] ), .ZN(n25864) );
  AOI22_X1 U29344 ( .A1(n30757), .A2(\xmem_data[68][5] ), .B1(n30756), .B2(
        \xmem_data[69][5] ), .ZN(n25863) );
  AOI22_X1 U29345 ( .A1(n30759), .A2(\xmem_data[70][5] ), .B1(n3144), .B2(
        \xmem_data[71][5] ), .ZN(n25862) );
  NAND4_X1 U29346 ( .A1(n25865), .A2(n25864), .A3(n25863), .A4(n25862), .ZN(
        n25870) );
  AOI22_X1 U29347 ( .A1(n28689), .A2(\xmem_data[90][5] ), .B1(n22717), .B2(
        \xmem_data[91][5] ), .ZN(n25866) );
  INV_X1 U29348 ( .A(n25866), .ZN(n25869) );
  AOI22_X1 U29349 ( .A1(n29801), .A2(\xmem_data[80][5] ), .B1(n29704), .B2(
        \xmem_data[81][5] ), .ZN(n25867) );
  INV_X1 U29350 ( .A(n25867), .ZN(n25868) );
  NOR3_X1 U29351 ( .A1(n25870), .A2(n25869), .A3(n25868), .ZN(n25881) );
  AOI22_X1 U29352 ( .A1(n3224), .A2(\xmem_data[78][5] ), .B1(n30710), .B2(
        \xmem_data[79][5] ), .ZN(n25874) );
  AOI22_X1 U29353 ( .A1(n30747), .A2(\xmem_data[86][5] ), .B1(n30543), .B2(
        \xmem_data[87][5] ), .ZN(n25873) );
  AOI22_X1 U29354 ( .A1(n26543), .A2(\xmem_data[82][5] ), .B1(n30744), .B2(
        \xmem_data[83][5] ), .ZN(n25872) );
  AOI22_X1 U29355 ( .A1(n30767), .A2(\xmem_data[94][5] ), .B1(n3269), .B2(
        \xmem_data[95][5] ), .ZN(n25871) );
  AOI22_X1 U29356 ( .A1(n3166), .A2(\xmem_data[88][5] ), .B1(n3189), .B2(
        \xmem_data[89][5] ), .ZN(n25875) );
  NAND2_X1 U29357 ( .A1(n3802), .A2(n25875), .ZN(n25878) );
  AOI22_X1 U29358 ( .A1(n30665), .A2(\xmem_data[84][5] ), .B1(n29739), .B2(
        \xmem_data[85][5] ), .ZN(n25876) );
  INV_X1 U29359 ( .A(n25876), .ZN(n25877) );
  NOR2_X1 U29360 ( .A1(n25878), .A2(n25877), .ZN(n25880) );
  AOI22_X1 U29361 ( .A1(n29815), .A2(\xmem_data[92][5] ), .B1(n30765), .B2(
        \xmem_data[93][5] ), .ZN(n25879) );
  NAND4_X1 U29362 ( .A1(n25882), .A2(n25881), .A3(n25880), .A4(n25879), .ZN(
        n25886) );
  AOI22_X1 U29363 ( .A1(n30279), .A2(\xmem_data[74][5] ), .B1(n28218), .B2(
        \xmem_data[75][5] ), .ZN(n25884) );
  AOI22_X1 U29364 ( .A1(n29421), .A2(\xmem_data[72][5] ), .B1(n29753), .B2(
        \xmem_data[73][5] ), .ZN(n25883) );
  NAND2_X1 U29365 ( .A1(n25884), .A2(n25883), .ZN(n25885) );
  OAI21_X1 U29366 ( .B1(n25886), .B2(n25885), .A(n30704), .ZN(n25935) );
  AOI22_X1 U29367 ( .A1(n30764), .A2(\xmem_data[26][5] ), .B1(n29639), .B2(
        \xmem_data[27][5] ), .ZN(n25897) );
  AOI22_X1 U29368 ( .A1(n29488), .A2(\xmem_data[28][5] ), .B1(n30266), .B2(
        \xmem_data[29][5] ), .ZN(n25896) );
  AOI22_X1 U29369 ( .A1(n3161), .A2(\xmem_data[24][5] ), .B1(n3188), .B2(
        \xmem_data[25][5] ), .ZN(n25895) );
  AOI22_X1 U29370 ( .A1(n7041), .A2(\xmem_data[0][5] ), .B1(n7042), .B2(
        \xmem_data[1][5] ), .ZN(n25890) );
  AOI22_X1 U29371 ( .A1(n30722), .A2(\xmem_data[2][5] ), .B1(n31345), .B2(
        \xmem_data[3][5] ), .ZN(n25889) );
  AOI22_X1 U29372 ( .A1(n30724), .A2(\xmem_data[4][5] ), .B1(n30723), .B2(
        \xmem_data[5][5] ), .ZN(n25888) );
  AOI22_X1 U29373 ( .A1(n30725), .A2(\xmem_data[6][5] ), .B1(n3414), .B2(
        \xmem_data[7][5] ), .ZN(n25887) );
  NAND4_X1 U29374 ( .A1(n25890), .A2(n25889), .A3(n25888), .A4(n25887), .ZN(
        n25893) );
  AOI22_X1 U29375 ( .A1(n30767), .A2(\xmem_data[30][5] ), .B1(n30686), .B2(
        \xmem_data[31][5] ), .ZN(n25891) );
  INV_X1 U29376 ( .A(n25891), .ZN(n25892) );
  NOR2_X1 U29377 ( .A1(n25893), .A2(n25892), .ZN(n25894) );
  NAND4_X1 U29378 ( .A1(n25897), .A2(n25896), .A3(n25895), .A4(n25894), .ZN(
        n25903) );
  AOI22_X1 U29379 ( .A1(n28739), .A2(\xmem_data[16][5] ), .B1(n3368), .B2(
        \xmem_data[17][5] ), .ZN(n25901) );
  AOI22_X1 U29380 ( .A1(n30731), .A2(\xmem_data[18][5] ), .B1(n28152), .B2(
        \xmem_data[19][5] ), .ZN(n25900) );
  AOI22_X1 U29381 ( .A1(n28779), .A2(\xmem_data[20][5] ), .B1(n26884), .B2(
        \xmem_data[21][5] ), .ZN(n25899) );
  AOI22_X1 U29382 ( .A1(n30732), .A2(\xmem_data[22][5] ), .B1(n30746), .B2(
        \xmem_data[23][5] ), .ZN(n25898) );
  NAND4_X1 U29383 ( .A1(n25901), .A2(n25900), .A3(n25899), .A4(n25898), .ZN(
        n25902) );
  OR2_X1 U29384 ( .A1(n25903), .A2(n25902), .ZN(n25909) );
  AOI22_X1 U29385 ( .A1(n28136), .A2(\xmem_data[8][5] ), .B1(n28766), .B2(
        \xmem_data[9][5] ), .ZN(n25907) );
  AOI22_X1 U29386 ( .A1(n28700), .A2(\xmem_data[10][5] ), .B1(n27445), .B2(
        \xmem_data[11][5] ), .ZN(n25906) );
  AOI22_X1 U29387 ( .A1(n30280), .A2(\xmem_data[12][5] ), .B1(n30217), .B2(
        \xmem_data[13][5] ), .ZN(n25905) );
  AOI22_X1 U29388 ( .A1(n3224), .A2(\xmem_data[14][5] ), .B1(n30710), .B2(
        \xmem_data[15][5] ), .ZN(n25904) );
  NAND4_X1 U29389 ( .A1(n25907), .A2(n25906), .A3(n25905), .A4(n25904), .ZN(
        n25908) );
  OAI21_X1 U29390 ( .B1(n25909), .B2(n25908), .A(n30741), .ZN(n25934) );
  AOI22_X1 U29391 ( .A1(n29801), .A2(\xmem_data[48][5] ), .B1(n28238), .B2(
        \xmem_data[49][5] ), .ZN(n25913) );
  AOI22_X1 U29392 ( .A1(n26543), .A2(\xmem_data[50][5] ), .B1(n30744), .B2(
        \xmem_data[51][5] ), .ZN(n25912) );
  AOI22_X1 U29393 ( .A1(n30665), .A2(\xmem_data[52][5] ), .B1(n30193), .B2(
        \xmem_data[53][5] ), .ZN(n25911) );
  AOI22_X1 U29394 ( .A1(n30747), .A2(\xmem_data[54][5] ), .B1(n20718), .B2(
        \xmem_data[55][5] ), .ZN(n25910) );
  NAND4_X1 U29395 ( .A1(n25913), .A2(n25912), .A3(n25911), .A4(n25910), .ZN(
        n25919) );
  AOI22_X1 U29396 ( .A1(n3168), .A2(\xmem_data[56][5] ), .B1(n3185), .B2(
        \xmem_data[57][5] ), .ZN(n25917) );
  AOI22_X1 U29397 ( .A1(n30310), .A2(\xmem_data[58][5] ), .B1(n28781), .B2(
        \xmem_data[59][5] ), .ZN(n25916) );
  AOI22_X1 U29398 ( .A1(n30717), .A2(\xmem_data[60][5] ), .B1(n30716), .B2(
        \xmem_data[61][5] ), .ZN(n25915) );
  AOI22_X1 U29399 ( .A1(n30646), .A2(\xmem_data[62][5] ), .B1(n30645), .B2(
        \xmem_data[63][5] ), .ZN(n25914) );
  NAND4_X1 U29400 ( .A1(n25917), .A2(n25916), .A3(n25915), .A4(n25914), .ZN(
        n25918) );
  OR2_X1 U29401 ( .A1(n25919), .A2(n25918), .ZN(n25932) );
  AOI22_X1 U29402 ( .A1(n30777), .A2(\xmem_data[44][5] ), .B1(n30293), .B2(
        \xmem_data[45][5] ), .ZN(n25930) );
  AOI22_X1 U29403 ( .A1(n27740), .A2(\xmem_data[42][5] ), .B1(n29565), .B2(
        \xmem_data[43][5] ), .ZN(n25929) );
  AOI22_X1 U29404 ( .A1(n28734), .A2(\xmem_data[40][5] ), .B1(n30654), .B2(
        \xmem_data[41][5] ), .ZN(n25928) );
  AOI22_X1 U29405 ( .A1(n30753), .A2(\xmem_data[32][5] ), .B1(n30752), .B2(
        \xmem_data[33][5] ), .ZN(n25923) );
  AOI22_X1 U29406 ( .A1(n30755), .A2(\xmem_data[34][5] ), .B1(n30754), .B2(
        \xmem_data[35][5] ), .ZN(n25922) );
  AOI22_X1 U29407 ( .A1(n30757), .A2(\xmem_data[36][5] ), .B1(n30756), .B2(
        \xmem_data[37][5] ), .ZN(n25921) );
  AOI22_X1 U29408 ( .A1(n30759), .A2(\xmem_data[38][5] ), .B1(n3144), .B2(
        \xmem_data[39][5] ), .ZN(n25920) );
  NAND4_X1 U29409 ( .A1(n25923), .A2(n25922), .A3(n25921), .A4(n25920), .ZN(
        n25926) );
  AOI22_X1 U29410 ( .A1(n3224), .A2(\xmem_data[46][5] ), .B1(n30295), .B2(
        \xmem_data[47][5] ), .ZN(n25924) );
  INV_X1 U29411 ( .A(n25924), .ZN(n25925) );
  NOR2_X1 U29412 ( .A1(n25926), .A2(n25925), .ZN(n25927) );
  NAND4_X1 U29413 ( .A1(n25930), .A2(n25929), .A3(n25928), .A4(n25927), .ZN(
        n25931) );
  OAI21_X1 U29414 ( .B1(n25932), .B2(n25931), .A(n30782), .ZN(n25933) );
  AOI22_X1 U29415 ( .A1(n30753), .A2(\xmem_data[32][4] ), .B1(n30752), .B2(
        \xmem_data[33][4] ), .ZN(n25940) );
  AOI22_X1 U29416 ( .A1(n30755), .A2(\xmem_data[34][4] ), .B1(n30754), .B2(
        \xmem_data[35][4] ), .ZN(n25939) );
  AOI22_X1 U29417 ( .A1(n30757), .A2(\xmem_data[36][4] ), .B1(n30756), .B2(
        \xmem_data[37][4] ), .ZN(n25938) );
  AOI22_X1 U29418 ( .A1(n30759), .A2(\xmem_data[38][4] ), .B1(n3144), .B2(
        \xmem_data[39][4] ), .ZN(n25937) );
  NAND4_X1 U29419 ( .A1(n25940), .A2(n25939), .A3(n25938), .A4(n25937), .ZN(
        n25956) );
  AOI22_X1 U29420 ( .A1(n29433), .A2(\xmem_data[40][4] ), .B1(n29753), .B2(
        \xmem_data[41][4] ), .ZN(n25944) );
  AOI22_X1 U29421 ( .A1(n29790), .A2(\xmem_data[42][4] ), .B1(n30292), .B2(
        \xmem_data[43][4] ), .ZN(n25943) );
  AOI22_X1 U29422 ( .A1(n30777), .A2(\xmem_data[44][4] ), .B1(n29798), .B2(
        \xmem_data[45][4] ), .ZN(n25942) );
  AOI22_X1 U29423 ( .A1(n3224), .A2(\xmem_data[46][4] ), .B1(n30295), .B2(
        \xmem_data[47][4] ), .ZN(n25941) );
  NAND4_X1 U29424 ( .A1(n25944), .A2(n25943), .A3(n25942), .A4(n25941), .ZN(
        n25955) );
  AOI22_X1 U29425 ( .A1(n3249), .A2(\xmem_data[48][4] ), .B1(n30662), .B2(
        \xmem_data[49][4] ), .ZN(n25948) );
  AOI22_X1 U29426 ( .A1(n30664), .A2(\xmem_data[50][4] ), .B1(n30744), .B2(
        \xmem_data[51][4] ), .ZN(n25947) );
  AOI22_X1 U29427 ( .A1(n27754), .A2(\xmem_data[52][4] ), .B1(n30090), .B2(
        \xmem_data[53][4] ), .ZN(n25946) );
  AOI22_X1 U29428 ( .A1(n30747), .A2(\xmem_data[54][4] ), .B1(n30543), .B2(
        \xmem_data[55][4] ), .ZN(n25945) );
  NAND4_X1 U29429 ( .A1(n25948), .A2(n25947), .A3(n25946), .A4(n25945), .ZN(
        n25954) );
  AOI22_X1 U29430 ( .A1(n3162), .A2(\xmem_data[56][4] ), .B1(n3187), .B2(
        \xmem_data[57][4] ), .ZN(n25952) );
  AOI22_X1 U29431 ( .A1(n30062), .A2(\xmem_data[58][4] ), .B1(n24710), .B2(
        \xmem_data[59][4] ), .ZN(n25951) );
  AOI22_X1 U29432 ( .A1(n29488), .A2(\xmem_data[60][4] ), .B1(n30716), .B2(
        \xmem_data[61][4] ), .ZN(n25950) );
  AOI22_X1 U29433 ( .A1(n30687), .A2(\xmem_data[62][4] ), .B1(n30686), .B2(
        \xmem_data[63][4] ), .ZN(n25949) );
  NAND4_X1 U29434 ( .A1(n25951), .A2(n25952), .A3(n25950), .A4(n25949), .ZN(
        n25953) );
  OR4_X1 U29435 ( .A1(n25956), .A2(n25955), .A3(n25954), .A4(n25953), .ZN(
        n25978) );
  AOI22_X1 U29436 ( .A1(n30673), .A2(\xmem_data[0][4] ), .B1(n7042), .B2(
        \xmem_data[1][4] ), .ZN(n25960) );
  AOI22_X1 U29437 ( .A1(n30722), .A2(\xmem_data[2][4] ), .B1(n29383), .B2(
        \xmem_data[3][4] ), .ZN(n25959) );
  AOI22_X1 U29438 ( .A1(n30724), .A2(\xmem_data[4][4] ), .B1(n30723), .B2(
        \xmem_data[5][4] ), .ZN(n25958) );
  AOI22_X1 U29439 ( .A1(n30725), .A2(\xmem_data[6][4] ), .B1(n3414), .B2(
        \xmem_data[7][4] ), .ZN(n25957) );
  NAND4_X1 U29440 ( .A1(n25960), .A2(n25959), .A3(n25958), .A4(n25957), .ZN(
        n25976) );
  AOI22_X1 U29441 ( .A1(n29788), .A2(\xmem_data[8][4] ), .B1(n27832), .B2(
        \xmem_data[9][4] ), .ZN(n25964) );
  AOI22_X1 U29442 ( .A1(n30215), .A2(\xmem_data[10][4] ), .B1(n29431), .B2(
        \xmem_data[11][4] ), .ZN(n25963) );
  AOI22_X1 U29443 ( .A1(n28209), .A2(\xmem_data[12][4] ), .B1(n28667), .B2(
        \xmem_data[13][4] ), .ZN(n25962) );
  AOI22_X1 U29444 ( .A1(n3224), .A2(\xmem_data[14][4] ), .B1(n30710), .B2(
        \xmem_data[15][4] ), .ZN(n25961) );
  NAND4_X1 U29445 ( .A1(n25964), .A2(n25963), .A3(n25962), .A4(n25961), .ZN(
        n25975) );
  AOI22_X1 U29446 ( .A1(n28739), .A2(\xmem_data[16][4] ), .B1(n30730), .B2(
        \xmem_data[17][4] ), .ZN(n25968) );
  AOI22_X1 U29447 ( .A1(n30731), .A2(\xmem_data[18][4] ), .B1(n30083), .B2(
        \xmem_data[19][4] ), .ZN(n25967) );
  AOI22_X1 U29448 ( .A1(n29714), .A2(\xmem_data[20][4] ), .B1(n30084), .B2(
        \xmem_data[21][4] ), .ZN(n25966) );
  AOI22_X1 U29449 ( .A1(n30732), .A2(\xmem_data[22][4] ), .B1(n30303), .B2(
        \xmem_data[23][4] ), .ZN(n25965) );
  NAND4_X1 U29450 ( .A1(n25968), .A2(n25967), .A3(n25966), .A4(n25965), .ZN(
        n25974) );
  AOI22_X1 U29451 ( .A1(n29476), .A2(\xmem_data[26][4] ), .B1(n28754), .B2(
        \xmem_data[27][4] ), .ZN(n25972) );
  AOI22_X1 U29452 ( .A1(n27713), .A2(\xmem_data[28][4] ), .B1(n30716), .B2(
        \xmem_data[29][4] ), .ZN(n25971) );
  AOI22_X1 U29453 ( .A1(n3165), .A2(\xmem_data[24][4] ), .B1(n3191), .B2(
        \xmem_data[25][4] ), .ZN(n25970) );
  AOI22_X1 U29454 ( .A1(n30687), .A2(\xmem_data[30][4] ), .B1(n30686), .B2(
        \xmem_data[31][4] ), .ZN(n25969) );
  NAND4_X1 U29455 ( .A1(n25972), .A2(n25971), .A3(n25970), .A4(n25969), .ZN(
        n25973) );
  AOI22_X1 U29456 ( .A1(n30782), .A2(n25978), .B1(n30741), .B2(n25977), .ZN(
        n26022) );
  AOI22_X1 U29457 ( .A1(n30673), .A2(\xmem_data[96][4] ), .B1(n30672), .B2(
        \xmem_data[97][4] ), .ZN(n25982) );
  AOI22_X1 U29458 ( .A1(n30675), .A2(\xmem_data[98][4] ), .B1(n30674), .B2(
        \xmem_data[99][4] ), .ZN(n25981) );
  AOI22_X1 U29459 ( .A1(n30677), .A2(\xmem_data[100][4] ), .B1(n30676), .B2(
        \xmem_data[101][4] ), .ZN(n25980) );
  AOI22_X1 U29460 ( .A1(n30678), .A2(\xmem_data[102][4] ), .B1(n28245), .B2(
        \xmem_data[103][4] ), .ZN(n25979) );
  NAND4_X1 U29461 ( .A1(n25982), .A2(n25981), .A3(n25980), .A4(n25979), .ZN(
        n25998) );
  AOI22_X1 U29462 ( .A1(n30291), .A2(\xmem_data[104][4] ), .B1(n30100), .B2(
        \xmem_data[105][4] ), .ZN(n25986) );
  AOI22_X1 U29463 ( .A1(n28700), .A2(\xmem_data[106][4] ), .B1(n28367), .B2(
        \xmem_data[107][4] ), .ZN(n25985) );
  AOI22_X1 U29464 ( .A1(n30697), .A2(\xmem_data[108][4] ), .B1(n30293), .B2(
        \xmem_data[109][4] ), .ZN(n25984) );
  AOI22_X1 U29465 ( .A1(n30699), .A2(\xmem_data[110][4] ), .B1(n30698), .B2(
        \xmem_data[111][4] ), .ZN(n25983) );
  NAND4_X1 U29466 ( .A1(n25986), .A2(n25985), .A3(n25984), .A4(n25983), .ZN(
        n25997) );
  AOI22_X1 U29467 ( .A1(n28146), .A2(\xmem_data[112][4] ), .B1(n29589), .B2(
        \xmem_data[113][4] ), .ZN(n25990) );
  AOI22_X1 U29468 ( .A1(n30664), .A2(\xmem_data[114][4] ), .B1(n30663), .B2(
        \xmem_data[115][4] ), .ZN(n25989) );
  AOI22_X1 U29469 ( .A1(n29714), .A2(\xmem_data[116][4] ), .B1(n29768), .B2(
        \xmem_data[117][4] ), .ZN(n25988) );
  AOI22_X1 U29470 ( .A1(n30667), .A2(\xmem_data[118][4] ), .B1(n29237), .B2(
        \xmem_data[119][4] ), .ZN(n25987) );
  NAND4_X1 U29471 ( .A1(n25990), .A2(n25989), .A3(n25988), .A4(n25987), .ZN(
        n25996) );
  AOI22_X1 U29472 ( .A1(n3166), .A2(\xmem_data[120][4] ), .B1(n3183), .B2(
        \xmem_data[121][4] ), .ZN(n25994) );
  AOI22_X1 U29473 ( .A1(n30075), .A2(\xmem_data[122][4] ), .B1(n30950), .B2(
        \xmem_data[123][4] ), .ZN(n25993) );
  AOI22_X1 U29474 ( .A1(n29722), .A2(\xmem_data[124][4] ), .B1(n30765), .B2(
        \xmem_data[125][4] ), .ZN(n25992) );
  AOI22_X1 U29475 ( .A1(n30767), .A2(\xmem_data[126][4] ), .B1(n3328), .B2(
        \xmem_data[127][4] ), .ZN(n25991) );
  NAND4_X1 U29476 ( .A1(n25994), .A2(n25993), .A3(n25992), .A4(n25991), .ZN(
        n25995) );
  OR4_X1 U29477 ( .A1(n25998), .A2(n25997), .A3(n25996), .A4(n25995), .ZN(
        n26020) );
  AOI22_X1 U29478 ( .A1(n29433), .A2(\xmem_data[72][4] ), .B1(n29697), .B2(
        \xmem_data[73][4] ), .ZN(n26002) );
  AOI22_X1 U29479 ( .A1(n29790), .A2(\xmem_data[74][4] ), .B1(n28218), .B2(
        \xmem_data[75][4] ), .ZN(n26001) );
  AOI22_X1 U29480 ( .A1(n30777), .A2(\xmem_data[76][4] ), .B1(n29708), .B2(
        \xmem_data[77][4] ), .ZN(n26000) );
  AOI22_X1 U29481 ( .A1(n3224), .A2(\xmem_data[78][4] ), .B1(n3131), .B2(
        \xmem_data[79][4] ), .ZN(n25999) );
  NAND4_X1 U29482 ( .A1(n26002), .A2(n26001), .A3(n26000), .A4(n25999), .ZN(
        n26018) );
  AOI22_X1 U29483 ( .A1(n30743), .A2(\xmem_data[80][4] ), .B1(n30662), .B2(
        \xmem_data[81][4] ), .ZN(n26006) );
  AOI22_X1 U29484 ( .A1(n30664), .A2(\xmem_data[82][4] ), .B1(n30744), .B2(
        \xmem_data[83][4] ), .ZN(n26005) );
  AOI22_X1 U29485 ( .A1(n28779), .A2(\xmem_data[84][4] ), .B1(n27728), .B2(
        \xmem_data[85][4] ), .ZN(n26004) );
  AOI22_X1 U29486 ( .A1(n30747), .A2(\xmem_data[86][4] ), .B1(n28516), .B2(
        \xmem_data[87][4] ), .ZN(n26003) );
  NAND4_X1 U29487 ( .A1(n26006), .A2(n26005), .A3(n26004), .A4(n26003), .ZN(
        n26017) );
  AOI22_X1 U29488 ( .A1(n3161), .A2(\xmem_data[88][4] ), .B1(n3182), .B2(
        \xmem_data[89][4] ), .ZN(n26010) );
  AOI22_X1 U29489 ( .A1(n30684), .A2(\xmem_data[90][4] ), .B1(n20942), .B2(
        \xmem_data[91][4] ), .ZN(n26009) );
  AOI22_X1 U29490 ( .A1(n30717), .A2(\xmem_data[92][4] ), .B1(n30644), .B2(
        \xmem_data[93][4] ), .ZN(n26008) );
  AOI22_X1 U29491 ( .A1(n30767), .A2(\xmem_data[94][4] ), .B1(n30311), .B2(
        \xmem_data[95][4] ), .ZN(n26007) );
  NAND4_X1 U29492 ( .A1(n26010), .A2(n26009), .A3(n26008), .A4(n26007), .ZN(
        n26016) );
  AOI22_X1 U29493 ( .A1(n30753), .A2(\xmem_data[64][4] ), .B1(n30752), .B2(
        \xmem_data[65][4] ), .ZN(n26014) );
  AOI22_X1 U29494 ( .A1(n30755), .A2(\xmem_data[66][4] ), .B1(n30754), .B2(
        \xmem_data[67][4] ), .ZN(n26013) );
  AOI22_X1 U29495 ( .A1(n30757), .A2(\xmem_data[68][4] ), .B1(n30756), .B2(
        \xmem_data[69][4] ), .ZN(n26012) );
  AOI22_X1 U29496 ( .A1(n30759), .A2(\xmem_data[70][4] ), .B1(n3144), .B2(
        \xmem_data[71][4] ), .ZN(n26011) );
  NAND4_X1 U29497 ( .A1(n26014), .A2(n26013), .A3(n26012), .A4(n26011), .ZN(
        n26015) );
  AOI22_X1 U29498 ( .A1(n26020), .A2(n30659), .B1(n30704), .B2(n26019), .ZN(
        n26021) );
  NAND2_X1 U29499 ( .A1(n26022), .A2(n26021), .ZN(n32256) );
  XNOR2_X1 U29500 ( .A(n32256), .B(\fmem_data[23][7] ), .ZN(n33020) );
  XOR2_X1 U29501 ( .A(\fmem_data[23][6] ), .B(\fmem_data[23][7] ), .Z(n26023)
         );
  OAI22_X1 U29502 ( .A1(n35115), .A2(n35652), .B1(n33020), .B2(n35651), .ZN(
        n31678) );
  FA_X1 U29503 ( .A(n26026), .B(n26025), .CI(n26024), .CO(n31677), .S(n26038)
         );
  FA_X1 U29504 ( .A(n26028), .B(n3495), .CI(n26027), .CO(n31838), .S(n16356)
         );
  FA_X1 U29505 ( .A(n3491), .B(n26030), .CI(n26029), .CO(n31837), .S(n24839)
         );
  XNOR2_X1 U29506 ( .A(n31838), .B(n31837), .ZN(n26033) );
  FA_X1 U29507 ( .A(n26032), .B(n26031), .CI(n3730), .CO(n31836), .S(n26034)
         );
  XNOR2_X1 U29508 ( .A(n26033), .B(n31836), .ZN(n31789) );
  FA_X1 U29509 ( .A(n26036), .B(n26035), .CI(n26034), .CO(n31791), .S(n30135)
         );
  XNOR2_X1 U29510 ( .A(n26038), .B(n26037), .ZN(n26040) );
  XNOR2_X1 U29511 ( .A(n26040), .B(n26039), .ZN(n30134) );
  NOR2_X1 U29512 ( .A1(n30135), .A2(n30134), .ZN(n26259) );
  FA_X1 U29513 ( .A(n26043), .B(n26042), .CI(n26041), .CO(n30138), .S(n27322)
         );
  AOI22_X1 U29514 ( .A1(n29628), .A2(\xmem_data[82][1] ), .B1(n28218), .B2(
        \xmem_data[83][1] ), .ZN(n26047) );
  AOI22_X1 U29515 ( .A1(n27741), .A2(\xmem_data[80][1] ), .B1(n30654), .B2(
        \xmem_data[81][1] ), .ZN(n26046) );
  AOI22_X1 U29516 ( .A1(n28219), .A2(\xmem_data[84][1] ), .B1(n29798), .B2(
        \xmem_data[85][1] ), .ZN(n26045) );
  AOI22_X1 U29517 ( .A1(n28220), .A2(\xmem_data[86][1] ), .B1(n25451), .B2(
        \xmem_data[87][1] ), .ZN(n26044) );
  NAND4_X1 U29518 ( .A1(n26047), .A2(n26046), .A3(n26045), .A4(n26044), .ZN(
        n26048) );
  NAND2_X1 U29519 ( .A1(n26048), .A2(n28258), .ZN(n26094) );
  AOI22_X1 U29520 ( .A1(n29433), .A2(\xmem_data[112][1] ), .B1(n29831), .B2(
        \xmem_data[113][1] ), .ZN(n26052) );
  AOI22_X1 U29521 ( .A1(n27740), .A2(\xmem_data[114][1] ), .B1(n28218), .B2(
        \xmem_data[115][1] ), .ZN(n26051) );
  AOI22_X1 U29522 ( .A1(n28219), .A2(\xmem_data[116][1] ), .B1(n29629), .B2(
        \xmem_data[117][1] ), .ZN(n26050) );
  AOI22_X1 U29523 ( .A1(n28220), .A2(\xmem_data[118][1] ), .B1(n29231), .B2(
        \xmem_data[119][1] ), .ZN(n26049) );
  NAND4_X1 U29524 ( .A1(n26052), .A2(n26051), .A3(n26050), .A4(n26049), .ZN(
        n26053) );
  NAND2_X1 U29525 ( .A1(n26053), .A2(n28133), .ZN(n26093) );
  AOI22_X1 U29526 ( .A1(n30633), .A2(\xmem_data[88][1] ), .B1(n28145), .B2(
        \xmem_data[89][1] ), .ZN(n26060) );
  AOI22_X1 U29527 ( .A1(n29769), .A2(\xmem_data[92][1] ), .B1(n27728), .B2(
        \xmem_data[93][1] ), .ZN(n26054) );
  INV_X1 U29528 ( .A(n26054), .ZN(n26058) );
  AOI22_X1 U29529 ( .A1(n3240), .A2(\xmem_data[94][1] ), .B1(n28231), .B2(
        \xmem_data[95][1] ), .ZN(n26056) );
  AOI22_X1 U29530 ( .A1(n3241), .A2(\xmem_data[90][1] ), .B1(n28233), .B2(
        \xmem_data[91][1] ), .ZN(n26055) );
  NAND2_X1 U29531 ( .A1(n26056), .A2(n26055), .ZN(n26057) );
  NOR2_X1 U29532 ( .A1(n26058), .A2(n26057), .ZN(n26059) );
  NAND2_X1 U29533 ( .A1(n26060), .A2(n26059), .ZN(n26073) );
  AOI22_X1 U29534 ( .A1(n30310), .A2(\xmem_data[66][1] ), .B1(n28232), .B2(
        \xmem_data[67][1] ), .ZN(n26071) );
  AOI22_X1 U29535 ( .A1(n29722), .A2(\xmem_data[68][1] ), .B1(n30716), .B2(
        \xmem_data[69][1] ), .ZN(n26070) );
  AOI22_X1 U29536 ( .A1(n3166), .A2(\xmem_data[64][1] ), .B1(n3186), .B2(
        \xmem_data[65][1] ), .ZN(n26069) );
  AOI22_X1 U29537 ( .A1(n28240), .A2(\xmem_data[72][1] ), .B1(n28239), .B2(
        \xmem_data[73][1] ), .ZN(n26064) );
  AOI22_X1 U29538 ( .A1(n28242), .A2(\xmem_data[74][1] ), .B1(n28241), .B2(
        \xmem_data[75][1] ), .ZN(n26063) );
  AOI22_X1 U29539 ( .A1(n28244), .A2(\xmem_data[76][1] ), .B1(n28243), .B2(
        \xmem_data[77][1] ), .ZN(n26062) );
  AOI22_X1 U29540 ( .A1(n28246), .A2(\xmem_data[78][1] ), .B1(n28245), .B2(
        \xmem_data[79][1] ), .ZN(n26061) );
  NAND4_X1 U29541 ( .A1(n26064), .A2(n26063), .A3(n26062), .A4(n26061), .ZN(
        n26067) );
  AOI22_X1 U29542 ( .A1(n3233), .A2(\xmem_data[70][1] ), .B1(n28226), .B2(
        \xmem_data[71][1] ), .ZN(n26065) );
  INV_X1 U29543 ( .A(n26065), .ZN(n26066) );
  NOR2_X1 U29544 ( .A1(n26067), .A2(n26066), .ZN(n26068) );
  NAND4_X1 U29545 ( .A1(n26071), .A2(n26070), .A3(n26069), .A4(n26068), .ZN(
        n26072) );
  OAI21_X1 U29546 ( .B1(n26073), .B2(n26072), .A(n28258), .ZN(n26092) );
  AOI22_X1 U29547 ( .A1(n30743), .A2(\xmem_data[120][1] ), .B1(n29347), .B2(
        \xmem_data[121][1] ), .ZN(n26077) );
  AOI22_X1 U29548 ( .A1(n3241), .A2(\xmem_data[122][1] ), .B1(n28233), .B2(
        \xmem_data[123][1] ), .ZN(n26076) );
  AOI22_X1 U29549 ( .A1(n29436), .A2(\xmem_data[124][1] ), .B1(n30634), .B2(
        \xmem_data[125][1] ), .ZN(n26075) );
  AOI22_X1 U29550 ( .A1(n3240), .A2(\xmem_data[126][1] ), .B1(n28231), .B2(
        \xmem_data[127][1] ), .ZN(n26074) );
  NAND4_X1 U29551 ( .A1(n26077), .A2(n26076), .A3(n26075), .A4(n26074), .ZN(
        n26090) );
  AOI22_X1 U29552 ( .A1(n28755), .A2(\xmem_data[98][1] ), .B1(n28232), .B2(
        \xmem_data[99][1] ), .ZN(n26088) );
  AOI22_X1 U29553 ( .A1(n29547), .A2(\xmem_data[100][1] ), .B1(n30716), .B2(
        \xmem_data[101][1] ), .ZN(n26087) );
  AOI22_X1 U29554 ( .A1(n3164), .A2(\xmem_data[96][1] ), .B1(n3187), .B2(
        \xmem_data[97][1] ), .ZN(n26086) );
  AOI22_X1 U29555 ( .A1(n28240), .A2(\xmem_data[104][1] ), .B1(n28239), .B2(
        \xmem_data[105][1] ), .ZN(n26081) );
  AOI22_X1 U29556 ( .A1(n28242), .A2(\xmem_data[106][1] ), .B1(n28241), .B2(
        \xmem_data[107][1] ), .ZN(n26080) );
  AOI22_X1 U29557 ( .A1(n28244), .A2(\xmem_data[108][1] ), .B1(n28243), .B2(
        \xmem_data[109][1] ), .ZN(n26079) );
  AOI22_X1 U29558 ( .A1(n28246), .A2(\xmem_data[110][1] ), .B1(n28245), .B2(
        \xmem_data[111][1] ), .ZN(n26078) );
  NAND4_X1 U29559 ( .A1(n26081), .A2(n26080), .A3(n26079), .A4(n26078), .ZN(
        n26084) );
  AOI22_X1 U29560 ( .A1(n3233), .A2(\xmem_data[102][1] ), .B1(n28226), .B2(
        \xmem_data[103][1] ), .ZN(n26082) );
  INV_X1 U29561 ( .A(n26082), .ZN(n26083) );
  NOR2_X1 U29562 ( .A1(n26084), .A2(n26083), .ZN(n26085) );
  NAND4_X1 U29563 ( .A1(n26088), .A2(n26087), .A3(n26086), .A4(n26085), .ZN(
        n26089) );
  OAI21_X1 U29564 ( .B1(n26090), .B2(n26089), .A(n28133), .ZN(n26091) );
  AND4_X1 U29565 ( .A1(n26094), .A2(n26093), .A3(n26092), .A4(n26091), .ZN(
        n26147) );
  AOI22_X1 U29566 ( .A1(n11444), .A2(\xmem_data[32][1] ), .B1(n3190), .B2(
        \xmem_data[33][1] ), .ZN(n26098) );
  AOI22_X1 U29567 ( .A1(n29610), .A2(\xmem_data[34][1] ), .B1(n28147), .B2(
        \xmem_data[35][1] ), .ZN(n26097) );
  AOI22_X1 U29568 ( .A1(n30766), .A2(\xmem_data[36][1] ), .B1(n30716), .B2(
        \xmem_data[37][1] ), .ZN(n26096) );
  AOI22_X1 U29569 ( .A1(n28151), .A2(\xmem_data[38][1] ), .B1(n30311), .B2(
        \xmem_data[39][1] ), .ZN(n26095) );
  AOI22_X1 U29570 ( .A1(n28138), .A2(\xmem_data[50][1] ), .B1(n28137), .B2(
        \xmem_data[51][1] ), .ZN(n26099) );
  INV_X1 U29571 ( .A(n26099), .ZN(n26113) );
  AOI22_X1 U29572 ( .A1(n28180), .A2(\xmem_data[56][1] ), .B1(n29482), .B2(
        \xmem_data[57][1] ), .ZN(n26111) );
  AOI22_X1 U29573 ( .A1(n3174), .A2(\xmem_data[60][1] ), .B1(n30249), .B2(
        \xmem_data[61][1] ), .ZN(n26110) );
  AOI22_X1 U29574 ( .A1(n28160), .A2(\xmem_data[40][1] ), .B1(n28159), .B2(
        \xmem_data[41][1] ), .ZN(n26103) );
  AOI22_X1 U29575 ( .A1(n28161), .A2(\xmem_data[42][1] ), .B1(n24687), .B2(
        \xmem_data[43][1] ), .ZN(n26102) );
  AOI22_X1 U29576 ( .A1(n28163), .A2(\xmem_data[44][1] ), .B1(n28162), .B2(
        \xmem_data[45][1] ), .ZN(n26101) );
  AOI22_X1 U29577 ( .A1(n28165), .A2(\xmem_data[46][1] ), .B1(n28164), .B2(
        \xmem_data[47][1] ), .ZN(n26100) );
  NAND4_X1 U29578 ( .A1(n26103), .A2(n26102), .A3(n26101), .A4(n26100), .ZN(
        n26108) );
  AOI22_X1 U29579 ( .A1(n28155), .A2(\xmem_data[62][1] ), .B1(n28154), .B2(
        \xmem_data[63][1] ), .ZN(n26106) );
  AOI22_X1 U29580 ( .A1(n28153), .A2(\xmem_data[58][1] ), .B1(n28152), .B2(
        \xmem_data[59][1] ), .ZN(n26105) );
  AOI22_X1 U29581 ( .A1(n28140), .A2(\xmem_data[54][1] ), .B1(n28308), .B2(
        \xmem_data[55][1] ), .ZN(n26104) );
  NAND3_X1 U29582 ( .A1(n26106), .A2(n26105), .A3(n26104), .ZN(n26107) );
  NOR2_X1 U29583 ( .A1(n26108), .A2(n26107), .ZN(n26109) );
  NAND3_X1 U29584 ( .A1(n26111), .A2(n26110), .A3(n26109), .ZN(n26112) );
  NOR2_X1 U29585 ( .A1(n26113), .A2(n26112), .ZN(n26116) );
  AOI22_X1 U29586 ( .A1(n28139), .A2(\xmem_data[52][1] ), .B1(n28667), .B2(
        \xmem_data[53][1] ), .ZN(n26115) );
  AOI22_X1 U29587 ( .A1(n29433), .A2(\xmem_data[48][1] ), .B1(n30222), .B2(
        \xmem_data[49][1] ), .ZN(n26114) );
  NAND4_X1 U29588 ( .A1(n3863), .A2(n26116), .A3(n26115), .A4(n26114), .ZN(
        n26117) );
  NAND2_X1 U29589 ( .A1(n26117), .A2(n28177), .ZN(n26146) );
  AOI22_X1 U29590 ( .A1(n27710), .A2(\xmem_data[16][1] ), .B1(n27013), .B2(
        \xmem_data[17][1] ), .ZN(n26121) );
  AOI22_X1 U29591 ( .A1(n29699), .A2(\xmem_data[18][1] ), .B1(n25414), .B2(
        \xmem_data[19][1] ), .ZN(n26120) );
  AOI22_X1 U29592 ( .A1(n28209), .A2(\xmem_data[20][1] ), .B1(n29629), .B2(
        \xmem_data[21][1] ), .ZN(n26119) );
  AOI22_X1 U29593 ( .A1(n28210), .A2(\xmem_data[22][1] ), .B1(n3147), .B2(
        \xmem_data[23][1] ), .ZN(n26118) );
  NAND4_X1 U29594 ( .A1(n26121), .A2(n26120), .A3(n26119), .A4(n26118), .ZN(
        n26131) );
  NAND2_X1 U29595 ( .A1(n30266), .A2(\xmem_data[5][1] ), .ZN(n26129) );
  AOI22_X1 U29596 ( .A1(n30715), .A2(\xmem_data[2][1] ), .B1(n28754), .B2(
        \xmem_data[3][1] ), .ZN(n26128) );
  AOI22_X1 U29597 ( .A1(n3241), .A2(\xmem_data[26][1] ), .B1(n29591), .B2(
        \xmem_data[27][1] ), .ZN(n26124) );
  AOI22_X1 U29598 ( .A1(n3240), .A2(\xmem_data[30][1] ), .B1(n17018), .B2(
        \xmem_data[31][1] ), .ZN(n26123) );
  NAND2_X1 U29599 ( .A1(n28684), .A2(\xmem_data[29][1] ), .ZN(n26122) );
  NAND3_X1 U29600 ( .A1(n26124), .A2(n26123), .A3(n26122), .ZN(n26125) );
  AOI21_X1 U29601 ( .B1(n29714), .B2(\xmem_data[28][1] ), .A(n26125), .ZN(
        n26127) );
  AOI22_X1 U29602 ( .A1(n29801), .A2(\xmem_data[24][1] ), .B1(n29589), .B2(
        \xmem_data[25][1] ), .ZN(n26126) );
  NAND4_X1 U29603 ( .A1(n26129), .A2(n26128), .A3(n26127), .A4(n26126), .ZN(
        n26130) );
  NOR2_X1 U29604 ( .A1(n26131), .A2(n26130), .ZN(n26143) );
  AOI22_X1 U29605 ( .A1(n28191), .A2(\xmem_data[8][1] ), .B1(n28190), .B2(
        \xmem_data[9][1] ), .ZN(n26135) );
  AOI22_X1 U29606 ( .A1(n28193), .A2(\xmem_data[10][1] ), .B1(n28192), .B2(
        \xmem_data[11][1] ), .ZN(n26134) );
  AOI22_X1 U29607 ( .A1(n28195), .A2(\xmem_data[12][1] ), .B1(n28194), .B2(
        \xmem_data[13][1] ), .ZN(n26133) );
  AOI22_X1 U29608 ( .A1(n28196), .A2(\xmem_data[14][1] ), .B1(n3144), .B2(
        \xmem_data[15][1] ), .ZN(n26132) );
  AND4_X1 U29609 ( .A1(n26135), .A2(n26134), .A3(n26133), .A4(n26132), .ZN(
        n26140) );
  AOI22_X1 U29610 ( .A1(n3161), .A2(\xmem_data[0][1] ), .B1(n3188), .B2(
        \xmem_data[1][1] ), .ZN(n26139) );
  AOI22_X1 U29611 ( .A1(n3233), .A2(\xmem_data[6][1] ), .B1(n28202), .B2(
        \xmem_data[7][1] ), .ZN(n26137) );
  NAND2_X1 U29612 ( .A1(n30717), .A2(\xmem_data[4][1] ), .ZN(n26136) );
  AND2_X1 U29613 ( .A1(n26137), .A2(n26136), .ZN(n26138) );
  AND3_X1 U29614 ( .A1(n26140), .A2(n26139), .A3(n26138), .ZN(n26142) );
  INV_X1 U29615 ( .A(n28215), .ZN(n26141) );
  AOI21_X1 U29616 ( .B1(n26143), .B2(n26142), .A(n26141), .ZN(n26144) );
  INV_X1 U29617 ( .A(n26144), .ZN(n26145) );
  XNOR2_X1 U29618 ( .A(n33483), .B(\fmem_data[31][7] ), .ZN(n32258) );
  OAI22_X1 U29619 ( .A1(n26148), .A2(n35663), .B1(n35662), .B2(n32258), .ZN(
        n29526) );
  OR2_X1 U29620 ( .A1(n33751), .A2(n3653), .ZN(n26149) );
  OAI22_X1 U29621 ( .A1(n26149), .A2(n35581), .B1(n35580), .B2(n3653), .ZN(
        n31012) );
  OR2_X1 U29622 ( .A1(n36296), .A2(n3637), .ZN(n26150) );
  OAI22_X1 U29623 ( .A1(n26150), .A2(n35494), .B1(n35493), .B2(n3637), .ZN(
        n31011) );
  XNOR2_X1 U29624 ( .A(n3276), .B(\fmem_data[26][3] ), .ZN(n32143) );
  OAI22_X1 U29625 ( .A1(n26151), .A2(n32780), .B1(n32143), .B2(n32779), .ZN(
        n31010) );
  XNOR2_X1 U29626 ( .A(n3452), .B(\fmem_data[11][3] ), .ZN(n32261) );
  OAI22_X1 U29627 ( .A1(n32261), .A2(n34429), .B1(n26152), .B2(n34533), .ZN(
        n29524) );
  AOI22_X1 U29628 ( .A1(n30753), .A2(\xmem_data[32][3] ), .B1(n30752), .B2(
        \xmem_data[33][3] ), .ZN(n26156) );
  AOI22_X1 U29629 ( .A1(n30755), .A2(\xmem_data[34][3] ), .B1(n30754), .B2(
        \xmem_data[35][3] ), .ZN(n26155) );
  AOI22_X1 U29630 ( .A1(n30757), .A2(\xmem_data[36][3] ), .B1(n30756), .B2(
        \xmem_data[37][3] ), .ZN(n26154) );
  AOI22_X1 U29631 ( .A1(n30759), .A2(\xmem_data[38][3] ), .B1(n3144), .B2(
        \xmem_data[39][3] ), .ZN(n26153) );
  NAND4_X1 U29632 ( .A1(n26156), .A2(n26155), .A3(n26154), .A4(n26153), .ZN(
        n26172) );
  AOI22_X1 U29633 ( .A1(n29626), .A2(\xmem_data[40][3] ), .B1(n30290), .B2(
        \xmem_data[41][3] ), .ZN(n26160) );
  AOI22_X1 U29634 ( .A1(n29628), .A2(\xmem_data[42][3] ), .B1(n29565), .B2(
        \xmem_data[43][3] ), .ZN(n26159) );
  AOI22_X1 U29635 ( .A1(n30777), .A2(\xmem_data[44][3] ), .B1(n30293), .B2(
        \xmem_data[45][3] ), .ZN(n26158) );
  AOI22_X1 U29636 ( .A1(n3224), .A2(\xmem_data[46][3] ), .B1(n3345), .B2(
        \xmem_data[47][3] ), .ZN(n26157) );
  NAND4_X1 U29637 ( .A1(n26160), .A2(n26159), .A3(n26158), .A4(n26157), .ZN(
        n26171) );
  AOI22_X1 U29638 ( .A1(n29705), .A2(\xmem_data[48][3] ), .B1(n27761), .B2(
        \xmem_data[49][3] ), .ZN(n26164) );
  AOI22_X1 U29639 ( .A1(n30731), .A2(\xmem_data[50][3] ), .B1(n30744), .B2(
        \xmem_data[51][3] ), .ZN(n26163) );
  AOI22_X1 U29640 ( .A1(n29436), .A2(\xmem_data[52][3] ), .B1(n29648), .B2(
        \xmem_data[53][3] ), .ZN(n26162) );
  AOI22_X1 U29641 ( .A1(n30747), .A2(\xmem_data[54][3] ), .B1(n25461), .B2(
        \xmem_data[55][3] ), .ZN(n26161) );
  NAND4_X1 U29642 ( .A1(n26164), .A2(n26163), .A3(n26162), .A4(n26161), .ZN(
        n26170) );
  AOI22_X1 U29643 ( .A1(n3166), .A2(\xmem_data[56][3] ), .B1(n3190), .B2(
        \xmem_data[57][3] ), .ZN(n26168) );
  AOI22_X1 U29644 ( .A1(n27031), .A2(\xmem_data[58][3] ), .B1(n25400), .B2(
        \xmem_data[59][3] ), .ZN(n26167) );
  AOI22_X1 U29645 ( .A1(n29547), .A2(\xmem_data[60][3] ), .B1(n30266), .B2(
        \xmem_data[61][3] ), .ZN(n26166) );
  AOI22_X1 U29646 ( .A1(n30767), .A2(\xmem_data[62][3] ), .B1(n3151), .B2(
        \xmem_data[63][3] ), .ZN(n26165) );
  NAND4_X1 U29647 ( .A1(n26168), .A2(n26167), .A3(n26166), .A4(n26165), .ZN(
        n26169) );
  OR4_X1 U29648 ( .A1(n26172), .A2(n26171), .A3(n26170), .A4(n26169), .ZN(
        n26206) );
  AOI22_X1 U29649 ( .A1(n28180), .A2(\xmem_data[16][3] ), .B1(n29389), .B2(
        \xmem_data[17][3] ), .ZN(n26173) );
  INV_X1 U29650 ( .A(n26173), .ZN(n26178) );
  AOI22_X1 U29651 ( .A1(n29714), .A2(\xmem_data[20][3] ), .B1(n28778), .B2(
        \xmem_data[21][3] ), .ZN(n26176) );
  AOI22_X1 U29652 ( .A1(n30732), .A2(\xmem_data[22][3] ), .B1(n30892), .B2(
        \xmem_data[23][3] ), .ZN(n26175) );
  AOI22_X1 U29653 ( .A1(n30731), .A2(\xmem_data[18][3] ), .B1(n29591), .B2(
        \xmem_data[19][3] ), .ZN(n26174) );
  NAND3_X1 U29654 ( .A1(n26176), .A2(n26175), .A3(n26174), .ZN(n26177) );
  INV_X1 U29655 ( .A(n30741), .ZN(n26179) );
  OAI21_X1 U29656 ( .B1(n26178), .B2(n26177), .A(n30741), .ZN(n26183) );
  NOR2_X1 U29657 ( .A1(n26179), .A2(n39011), .ZN(n26181) );
  NOR2_X1 U29658 ( .A1(n26179), .A2(n39018), .ZN(n26180) );
  AOI22_X1 U29659 ( .A1(n28209), .A2(n26181), .B1(n30776), .B2(n26180), .ZN(
        n26182) );
  NAND2_X1 U29660 ( .A1(n26183), .A2(n26182), .ZN(n26190) );
  AOI22_X1 U29661 ( .A1(n3167), .A2(\xmem_data[24][3] ), .B1(n3185), .B2(
        \xmem_data[25][3] ), .ZN(n26187) );
  AOI22_X1 U29662 ( .A1(n29476), .A2(\xmem_data[26][3] ), .B1(n28147), .B2(
        \xmem_data[27][3] ), .ZN(n26186) );
  AOI22_X1 U29663 ( .A1(n30198), .A2(\xmem_data[28][3] ), .B1(n30685), .B2(
        \xmem_data[29][3] ), .ZN(n26185) );
  AOI22_X1 U29664 ( .A1(n30646), .A2(\xmem_data[30][3] ), .B1(n30645), .B2(
        \xmem_data[31][3] ), .ZN(n26184) );
  NAND4_X1 U29665 ( .A1(n26187), .A2(n26186), .A3(n26185), .A4(n26184), .ZN(
        n26188) );
  AND2_X1 U29666 ( .A1(n26188), .A2(n30741), .ZN(n26189) );
  NOR2_X1 U29667 ( .A1(n26190), .A2(n26189), .ZN(n26204) );
  AOI22_X1 U29668 ( .A1(n7041), .A2(\xmem_data[0][3] ), .B1(n7042), .B2(
        \xmem_data[1][3] ), .ZN(n26194) );
  AOI22_X1 U29669 ( .A1(n30722), .A2(\xmem_data[2][3] ), .B1(n21060), .B2(
        \xmem_data[3][3] ), .ZN(n26193) );
  AOI22_X1 U29670 ( .A1(n30724), .A2(\xmem_data[4][3] ), .B1(n30723), .B2(
        \xmem_data[5][3] ), .ZN(n26192) );
  AOI22_X1 U29671 ( .A1(n30725), .A2(\xmem_data[6][3] ), .B1(n3413), .B2(
        \xmem_data[7][3] ), .ZN(n26191) );
  NAND2_X1 U29672 ( .A1(n29753), .A2(\xmem_data[9][3] ), .ZN(n26196) );
  AOI22_X1 U29673 ( .A1(n3224), .A2(\xmem_data[14][3] ), .B1(n30710), .B2(
        \xmem_data[15][3] ), .ZN(n26195) );
  AOI22_X1 U29674 ( .A1(n30215), .A2(\xmem_data[10][3] ), .B1(n29565), .B2(
        \xmem_data[11][3] ), .ZN(n26200) );
  INV_X1 U29675 ( .A(n26200), .ZN(n26201) );
  OAI21_X1 U29676 ( .B1(n26202), .B2(n26201), .A(n30741), .ZN(n26203) );
  NAND2_X1 U29677 ( .A1(n26204), .A2(n26203), .ZN(n26205) );
  AOI21_X1 U29678 ( .B1(n26206), .B2(n30782), .A(n26205), .ZN(n26251) );
  AOI22_X1 U29679 ( .A1(n30673), .A2(\xmem_data[96][3] ), .B1(n30672), .B2(
        \xmem_data[97][3] ), .ZN(n26210) );
  AOI22_X1 U29680 ( .A1(n30675), .A2(\xmem_data[98][3] ), .B1(n30674), .B2(
        \xmem_data[99][3] ), .ZN(n26209) );
  AOI22_X1 U29681 ( .A1(n30677), .A2(\xmem_data[100][3] ), .B1(n30676), .B2(
        \xmem_data[101][3] ), .ZN(n26208) );
  AOI22_X1 U29682 ( .A1(n30678), .A2(\xmem_data[102][3] ), .B1(n3153), .B2(
        \xmem_data[103][3] ), .ZN(n26207) );
  NAND4_X1 U29683 ( .A1(n26210), .A2(n26209), .A3(n26208), .A4(n26207), .ZN(
        n26226) );
  AOI22_X1 U29684 ( .A1(n28136), .A2(\xmem_data[104][3] ), .B1(n30290), .B2(
        \xmem_data[105][3] ), .ZN(n26214) );
  AOI22_X1 U29685 ( .A1(n29628), .A2(\xmem_data[106][3] ), .B1(n29256), .B2(
        \xmem_data[107][3] ), .ZN(n26213) );
  AOI22_X1 U29686 ( .A1(n30697), .A2(\xmem_data[108][3] ), .B1(n28208), .B2(
        \xmem_data[109][3] ), .ZN(n26212) );
  AOI22_X1 U29687 ( .A1(n30699), .A2(\xmem_data[110][3] ), .B1(n30698), .B2(
        \xmem_data[111][3] ), .ZN(n26211) );
  NAND4_X1 U29688 ( .A1(n26214), .A2(n26213), .A3(n26212), .A4(n26211), .ZN(
        n26225) );
  AOI22_X1 U29689 ( .A1(n28146), .A2(\xmem_data[112][3] ), .B1(n29389), .B2(
        \xmem_data[113][3] ), .ZN(n26218) );
  AOI22_X1 U29690 ( .A1(n30664), .A2(\xmem_data[114][3] ), .B1(n30663), .B2(
        \xmem_data[115][3] ), .ZN(n26217) );
  AOI22_X1 U29691 ( .A1(n29436), .A2(\xmem_data[116][3] ), .B1(n28110), .B2(
        \xmem_data[117][3] ), .ZN(n26216) );
  AOI22_X1 U29692 ( .A1(n30667), .A2(\xmem_data[118][3] ), .B1(n17018), .B2(
        \xmem_data[119][3] ), .ZN(n26215) );
  NAND4_X1 U29693 ( .A1(n26218), .A2(n26217), .A3(n26216), .A4(n26215), .ZN(
        n26224) );
  AOI22_X1 U29694 ( .A1(n3166), .A2(\xmem_data[120][3] ), .B1(n3187), .B2(
        \xmem_data[121][3] ), .ZN(n26222) );
  AOI22_X1 U29695 ( .A1(n30684), .A2(\xmem_data[122][3] ), .B1(n28147), .B2(
        \xmem_data[123][3] ), .ZN(n26221) );
  AOI22_X1 U29696 ( .A1(n30076), .A2(\xmem_data[124][3] ), .B1(n29721), .B2(
        \xmem_data[125][3] ), .ZN(n26220) );
  AOI22_X1 U29697 ( .A1(n30646), .A2(\xmem_data[126][3] ), .B1(n30645), .B2(
        \xmem_data[127][3] ), .ZN(n26219) );
  NAND4_X1 U29698 ( .A1(n26222), .A2(n26221), .A3(n26220), .A4(n26219), .ZN(
        n26223) );
  OR4_X1 U29699 ( .A1(n26226), .A2(n26225), .A3(n26224), .A4(n26223), .ZN(
        n26249) );
  AOI22_X1 U29700 ( .A1(n30673), .A2(\xmem_data[64][3] ), .B1(n30672), .B2(
        \xmem_data[65][3] ), .ZN(n26230) );
  AOI22_X1 U29701 ( .A1(n30675), .A2(\xmem_data[66][3] ), .B1(n30674), .B2(
        \xmem_data[67][3] ), .ZN(n26229) );
  AOI22_X1 U29702 ( .A1(n30677), .A2(\xmem_data[68][3] ), .B1(n30676), .B2(
        \xmem_data[69][3] ), .ZN(n26228) );
  AOI22_X1 U29703 ( .A1(n30678), .A2(\xmem_data[70][3] ), .B1(n3144), .B2(
        \xmem_data[71][3] ), .ZN(n26227) );
  NAND4_X1 U29704 ( .A1(n26230), .A2(n26229), .A3(n26228), .A4(n26227), .ZN(
        n26247) );
  AOI22_X1 U29705 ( .A1(n28734), .A2(\xmem_data[72][3] ), .B1(n29432), .B2(
        \xmem_data[73][3] ), .ZN(n26234) );
  AOI22_X1 U29706 ( .A1(n28207), .A2(\xmem_data[74][3] ), .B1(n29422), .B2(
        \xmem_data[75][3] ), .ZN(n26233) );
  AOI22_X1 U29707 ( .A1(n30697), .A2(\xmem_data[76][3] ), .B1(n28208), .B2(
        \xmem_data[77][3] ), .ZN(n26232) );
  AOI22_X1 U29708 ( .A1(n30699), .A2(\xmem_data[78][3] ), .B1(n30698), .B2(
        \xmem_data[79][3] ), .ZN(n26231) );
  NAND4_X1 U29709 ( .A1(n26234), .A2(n26233), .A3(n26232), .A4(n26231), .ZN(
        n26246) );
  AOI22_X1 U29710 ( .A1(n28739), .A2(\xmem_data[80][3] ), .B1(n28145), .B2(
        \xmem_data[81][3] ), .ZN(n26238) );
  AOI22_X1 U29711 ( .A1(n30664), .A2(\xmem_data[82][3] ), .B1(n30663), .B2(
        \xmem_data[83][3] ), .ZN(n26237) );
  AOI22_X1 U29712 ( .A1(n3174), .A2(\xmem_data[84][3] ), .B1(n29648), .B2(
        \xmem_data[85][3] ), .ZN(n26236) );
  AOI22_X1 U29713 ( .A1(n30667), .A2(\xmem_data[86][3] ), .B1(n30303), .B2(
        \xmem_data[87][3] ), .ZN(n26235) );
  NAND4_X1 U29714 ( .A1(n26238), .A2(n26237), .A3(n26236), .A4(n26235), .ZN(
        n26245) );
  AND2_X1 U29715 ( .A1(n28232), .A2(\xmem_data[91][3] ), .ZN(n26239) );
  AOI21_X1 U29716 ( .B1(n30310), .B2(\xmem_data[90][3] ), .A(n26239), .ZN(
        n26243) );
  AOI22_X1 U29717 ( .A1(n3164), .A2(\xmem_data[88][3] ), .B1(n3189), .B2(
        \xmem_data[89][3] ), .ZN(n26242) );
  AOI22_X1 U29718 ( .A1(n27713), .A2(\xmem_data[92][3] ), .B1(n30266), .B2(
        \xmem_data[93][3] ), .ZN(n26241) );
  AOI22_X1 U29719 ( .A1(n30687), .A2(\xmem_data[94][3] ), .B1(n3151), .B2(
        \xmem_data[95][3] ), .ZN(n26240) );
  NAND4_X1 U29720 ( .A1(n26243), .A2(n26242), .A3(n26241), .A4(n26240), .ZN(
        n26244) );
  AOI22_X1 U29721 ( .A1(n30659), .A2(n26249), .B1(n30704), .B2(n26248), .ZN(
        n26250) );
  XNOR2_X1 U29722 ( .A(n33019), .B(\fmem_data[23][5] ), .ZN(n32150) );
  XNOR2_X1 U29723 ( .A(n32256), .B(\fmem_data[23][5] ), .ZN(n34234) );
  XNOR2_X1 U29724 ( .A(n3365), .B(\fmem_data[9][7] ), .ZN(n26253) );
  OAI22_X1 U29725 ( .A1(n26254), .A2(n35726), .B1(n26253), .B2(n35725), .ZN(
        n29531) );
  XNOR2_X1 U29726 ( .A(n35397), .B(\fmem_data[16][1] ), .ZN(n31990) );
  XNOR2_X1 U29727 ( .A(n34980), .B(\fmem_data[16][1] ), .ZN(n32167) );
  XNOR2_X1 U29728 ( .A(n34929), .B(\fmem_data[6][3] ), .ZN(n30445) );
  OAI22_X1 U29729 ( .A1(n31881), .A2(n33598), .B1(n30445), .B2(n33596), .ZN(
        n28904) );
  OAI21_X1 U29730 ( .B1(n28905), .B2(n28906), .A(n28904), .ZN(n26256) );
  NAND2_X1 U29731 ( .A1(n26256), .A2(n26255), .ZN(n27320) );
  INV_X1 U29732 ( .A(n30136), .ZN(n26258) );
  NAND2_X1 U29733 ( .A1(n30135), .A2(n30134), .ZN(n26257) );
  OAI21_X1 U29734 ( .B1(n26259), .B2(n26258), .A(n26257), .ZN(n31810) );
  XNOR2_X1 U29735 ( .A(n31774), .B(n31773), .ZN(n27308) );
  FA_X1 U29736 ( .A(n26262), .B(n26261), .CI(n26260), .CO(n31851), .S(n27309)
         );
  XNOR2_X1 U29737 ( .A(n26264), .B(n26263), .ZN(n26265) );
  XNOR2_X1 U29738 ( .A(n26265), .B(n26266), .ZN(n27310) );
  FA_X1 U29739 ( .A(n26269), .B(n26268), .CI(n26267), .CO(n26377), .S(n28916)
         );
  XNOR2_X1 U29740 ( .A(n31511), .B(\fmem_data[16][3] ), .ZN(n31163) );
  XNOR2_X1 U29741 ( .A(n32600), .B(\fmem_data[14][3] ), .ZN(n31122) );
  FA_X1 U29742 ( .A(n26274), .B(n26273), .CI(n26272), .CO(n23584), .S(n31483)
         );
  AOI22_X1 U29743 ( .A1(n28492), .A2(\xmem_data[96][1] ), .B1(n23802), .B2(
        \xmem_data[97][1] ), .ZN(n26278) );
  AOI22_X1 U29744 ( .A1(n30515), .A2(\xmem_data[98][1] ), .B1(n28493), .B2(
        \xmem_data[99][1] ), .ZN(n26277) );
  AOI22_X1 U29745 ( .A1(n28494), .A2(\xmem_data[100][1] ), .B1(n28202), .B2(
        \xmem_data[101][1] ), .ZN(n26276) );
  AOI22_X1 U29746 ( .A1(n28495), .A2(\xmem_data[102][1] ), .B1(n20734), .B2(
        \xmem_data[103][1] ), .ZN(n26275) );
  NAND4_X1 U29747 ( .A1(n26278), .A2(n26277), .A3(n26276), .A4(n26275), .ZN(
        n26294) );
  AOI22_X1 U29748 ( .A1(n28500), .A2(\xmem_data[104][1] ), .B1(n30901), .B2(
        \xmem_data[105][1] ), .ZN(n26282) );
  AOI22_X1 U29749 ( .A1(n20951), .A2(\xmem_data[106][1] ), .B1(n27564), .B2(
        \xmem_data[107][1] ), .ZN(n26281) );
  AOI22_X1 U29750 ( .A1(n31262), .A2(\xmem_data[108][1] ), .B1(n16980), .B2(
        \xmem_data[109][1] ), .ZN(n26280) );
  AOI22_X1 U29751 ( .A1(n28501), .A2(\xmem_data[110][1] ), .B1(n28503), .B2(
        \xmem_data[111][1] ), .ZN(n26279) );
  NAND4_X1 U29752 ( .A1(n26282), .A2(n26281), .A3(n26280), .A4(n26279), .ZN(
        n26293) );
  AOI22_X1 U29753 ( .A1(n3221), .A2(\xmem_data[112][1] ), .B1(n24563), .B2(
        \xmem_data[113][1] ), .ZN(n26286) );
  AOI22_X1 U29754 ( .A1(n28508), .A2(\xmem_data[114][1] ), .B1(n3342), .B2(
        \xmem_data[115][1] ), .ZN(n26285) );
  AOI22_X1 U29755 ( .A1(n28509), .A2(\xmem_data[116][1] ), .B1(n3345), .B2(
        \xmem_data[117][1] ), .ZN(n26284) );
  AOI22_X1 U29756 ( .A1(n25450), .A2(\xmem_data[118][1] ), .B1(n28374), .B2(
        \xmem_data[119][1] ), .ZN(n26283) );
  NAND4_X1 U29757 ( .A1(n26286), .A2(n26285), .A3(n26284), .A4(n26283), .ZN(
        n26292) );
  AOI22_X1 U29758 ( .A1(n14933), .A2(\xmem_data[120][1] ), .B1(n20545), .B2(
        \xmem_data[121][1] ), .ZN(n26290) );
  AOI22_X1 U29759 ( .A1(n28515), .A2(\xmem_data[122][1] ), .B1(n31268), .B2(
        \xmem_data[123][1] ), .ZN(n26289) );
  AOI22_X1 U29760 ( .A1(n28517), .A2(\xmem_data[124][1] ), .B1(n31354), .B2(
        \xmem_data[125][1] ), .ZN(n26288) );
  AOI22_X1 U29761 ( .A1(n20586), .A2(\xmem_data[126][1] ), .B1(n25573), .B2(
        \xmem_data[127][1] ), .ZN(n26287) );
  NAND4_X1 U29762 ( .A1(n26290), .A2(n26289), .A3(n26288), .A4(n26287), .ZN(
        n26291) );
  OR4_X1 U29763 ( .A1(n26294), .A2(n26293), .A3(n26292), .A4(n26291), .ZN(
        n26316) );
  AOI22_X1 U29764 ( .A1(n28492), .A2(\xmem_data[64][1] ), .B1(n29319), .B2(
        \xmem_data[65][1] ), .ZN(n26298) );
  AOI22_X1 U29765 ( .A1(n24460), .A2(\xmem_data[66][1] ), .B1(n28493), .B2(
        \xmem_data[67][1] ), .ZN(n26297) );
  AOI22_X1 U29766 ( .A1(n28494), .A2(\xmem_data[68][1] ), .B1(n30600), .B2(
        \xmem_data[69][1] ), .ZN(n26296) );
  AOI22_X1 U29767 ( .A1(n28495), .A2(\xmem_data[70][1] ), .B1(n3171), .B2(
        \xmem_data[71][1] ), .ZN(n26295) );
  NAND4_X1 U29768 ( .A1(n26298), .A2(n26297), .A3(n26296), .A4(n26295), .ZN(
        n26314) );
  AOI22_X1 U29769 ( .A1(n28500), .A2(\xmem_data[72][1] ), .B1(n30754), .B2(
        \xmem_data[73][1] ), .ZN(n26302) );
  AOI22_X1 U29770 ( .A1(n27957), .A2(\xmem_data[74][1] ), .B1(n27500), .B2(
        \xmem_data[75][1] ), .ZN(n26301) );
  AOI22_X1 U29771 ( .A1(n28037), .A2(\xmem_data[76][1] ), .B1(n25725), .B2(
        \xmem_data[77][1] ), .ZN(n26300) );
  AOI22_X1 U29772 ( .A1(n28501), .A2(\xmem_data[78][1] ), .B1(n28503), .B2(
        \xmem_data[79][1] ), .ZN(n26299) );
  NAND4_X1 U29773 ( .A1(n26302), .A2(n26301), .A3(n26300), .A4(n26299), .ZN(
        n26313) );
  AOI22_X1 U29774 ( .A1(n3218), .A2(\xmem_data[80][1] ), .B1(n29431), .B2(
        \xmem_data[81][1] ), .ZN(n26306) );
  AOI22_X1 U29775 ( .A1(n28508), .A2(\xmem_data[82][1] ), .B1(n3342), .B2(
        \xmem_data[83][1] ), .ZN(n26305) );
  AOI22_X1 U29776 ( .A1(n28509), .A2(\xmem_data[84][1] ), .B1(n30698), .B2(
        \xmem_data[85][1] ), .ZN(n26304) );
  AOI22_X1 U29777 ( .A1(n31252), .A2(\xmem_data[86][1] ), .B1(n28374), .B2(
        \xmem_data[87][1] ), .ZN(n26303) );
  NAND4_X1 U29778 ( .A1(n26306), .A2(n26305), .A3(n26304), .A4(n26303), .ZN(
        n26312) );
  AOI22_X1 U29779 ( .A1(n14933), .A2(\xmem_data[88][1] ), .B1(n28051), .B2(
        \xmem_data[89][1] ), .ZN(n26310) );
  AOI22_X1 U29780 ( .A1(n28515), .A2(\xmem_data[90][1] ), .B1(n25710), .B2(
        \xmem_data[91][1] ), .ZN(n26309) );
  AOI22_X1 U29781 ( .A1(n28517), .A2(\xmem_data[92][1] ), .B1(n30543), .B2(
        \xmem_data[93][1] ), .ZN(n26308) );
  AOI22_X1 U29782 ( .A1(n31269), .A2(\xmem_data[94][1] ), .B1(n25635), .B2(
        \xmem_data[95][1] ), .ZN(n26307) );
  NAND4_X1 U29783 ( .A1(n26310), .A2(n26309), .A3(n26308), .A4(n26307), .ZN(
        n26311) );
  OR4_X1 U29784 ( .A1(n26314), .A2(n26313), .A3(n26312), .A4(n26311), .ZN(
        n26315) );
  AOI22_X1 U29785 ( .A1(n28458), .A2(n26316), .B1(n28526), .B2(n26315), .ZN(
        n26369) );
  NOR2_X1 U29786 ( .A1(n15043), .A2(n39002), .ZN(n26317) );
  NAND2_X1 U29787 ( .A1(n27547), .A2(n26317), .ZN(n26368) );
  AOI22_X1 U29788 ( .A1(n27918), .A2(\xmem_data[32][1] ), .B1(n28781), .B2(
        \xmem_data[33][1] ), .ZN(n26321) );
  AOI22_X1 U29789 ( .A1(n24460), .A2(\xmem_data[34][1] ), .B1(n25717), .B2(
        \xmem_data[35][1] ), .ZN(n26320) );
  AOI22_X1 U29790 ( .A1(n28462), .A2(\xmem_data[36][1] ), .B1(n28461), .B2(
        \xmem_data[37][1] ), .ZN(n26319) );
  AOI22_X1 U29791 ( .A1(n24521), .A2(\xmem_data[38][1] ), .B1(n3172), .B2(
        \xmem_data[39][1] ), .ZN(n26318) );
  NAND4_X1 U29792 ( .A1(n26321), .A2(n26320), .A3(n26319), .A4(n26318), .ZN(
        n26337) );
  AOI22_X1 U29793 ( .A1(n28468), .A2(\xmem_data[40][1] ), .B1(n28467), .B2(
        \xmem_data[41][1] ), .ZN(n26325) );
  AOI22_X1 U29794 ( .A1(n20579), .A2(\xmem_data[42][1] ), .B1(n24526), .B2(
        \xmem_data[43][1] ), .ZN(n26324) );
  AOI22_X1 U29795 ( .A1(n3203), .A2(\xmem_data[44][1] ), .B1(n25443), .B2(
        \xmem_data[45][1] ), .ZN(n26323) );
  AOI22_X1 U29796 ( .A1(n29173), .A2(\xmem_data[46][1] ), .B1(n28470), .B2(
        \xmem_data[47][1] ), .ZN(n26322) );
  NAND4_X1 U29797 ( .A1(n26325), .A2(n26324), .A3(n26323), .A4(n26322), .ZN(
        n26336) );
  AOI22_X1 U29798 ( .A1(n3217), .A2(\xmem_data[48][1] ), .B1(n29789), .B2(
        \xmem_data[49][1] ), .ZN(n26329) );
  AOI22_X1 U29799 ( .A1(n28476), .A2(\xmem_data[50][1] ), .B1(n28475), .B2(
        \xmem_data[51][1] ), .ZN(n26328) );
  AOI22_X1 U29800 ( .A1(n22711), .A2(\xmem_data[52][1] ), .B1(n27905), .B2(
        \xmem_data[53][1] ), .ZN(n26327) );
  AOI22_X1 U29801 ( .A1(n30877), .A2(\xmem_data[54][1] ), .B1(n27551), .B2(
        \xmem_data[55][1] ), .ZN(n26326) );
  NAND4_X1 U29802 ( .A1(n26329), .A2(n26328), .A3(n26327), .A4(n26326), .ZN(
        n26335) );
  AOI22_X1 U29803 ( .A1(n28481), .A2(\xmem_data[56][1] ), .B1(n27763), .B2(
        \xmem_data[57][1] ), .ZN(n26333) );
  AOI22_X1 U29804 ( .A1(n22702), .A2(\xmem_data[58][1] ), .B1(n16986), .B2(
        \xmem_data[59][1] ), .ZN(n26332) );
  AOI22_X1 U29805 ( .A1(n25572), .A2(\xmem_data[60][1] ), .B1(n27455), .B2(
        \xmem_data[61][1] ), .ZN(n26331) );
  AOI22_X1 U29806 ( .A1(n27454), .A2(\xmem_data[62][1] ), .B1(n21007), .B2(
        \xmem_data[63][1] ), .ZN(n26330) );
  NAND4_X1 U29807 ( .A1(n26333), .A2(n26332), .A3(n26331), .A4(n26330), .ZN(
        n26334) );
  OR4_X1 U29808 ( .A1(n26337), .A2(n26336), .A3(n26335), .A4(n26334), .ZN(
        n26366) );
  AOI22_X1 U29809 ( .A1(n27437), .A2(\xmem_data[14][1] ), .B1(n20991), .B2(
        \xmem_data[15][1] ), .ZN(n26348) );
  AOI22_X1 U29810 ( .A1(n30571), .A2(\xmem_data[12][1] ), .B1(n29661), .B2(
        \xmem_data[13][1] ), .ZN(n26338) );
  INV_X1 U29811 ( .A(n26338), .ZN(n26341) );
  AOI22_X1 U29812 ( .A1(n22727), .A2(\xmem_data[10][1] ), .B1(n30862), .B2(
        \xmem_data[11][1] ), .ZN(n26339) );
  INV_X1 U29813 ( .A(n26339), .ZN(n26340) );
  NOR2_X1 U29814 ( .A1(n26341), .A2(n26340), .ZN(n26347) );
  AOI22_X1 U29815 ( .A1(n28468), .A2(\xmem_data[8][1] ), .B1(n27717), .B2(
        \xmem_data[9][1] ), .ZN(n26346) );
  AOI22_X1 U29816 ( .A1(n28427), .A2(\xmem_data[0][1] ), .B1(n28302), .B2(
        \xmem_data[1][1] ), .ZN(n26345) );
  AOI22_X1 U29817 ( .A1(n25435), .A2(\xmem_data[2][1] ), .B1(n28428), .B2(
        \xmem_data[3][1] ), .ZN(n26344) );
  AOI22_X1 U29818 ( .A1(n3372), .A2(\xmem_data[4][1] ), .B1(n3308), .B2(
        \xmem_data[5][1] ), .ZN(n26343) );
  AOI22_X1 U29819 ( .A1(n20781), .A2(\xmem_data[6][1] ), .B1(n21058), .B2(
        \xmem_data[7][1] ), .ZN(n26342) );
  NAND4_X1 U29820 ( .A1(n26348), .A2(n26347), .A3(n26346), .A4(n3785), .ZN(
        n26363) );
  AOI22_X1 U29821 ( .A1(n3221), .A2(\xmem_data[16][1] ), .B1(n29627), .B2(
        \xmem_data[17][1] ), .ZN(n26355) );
  AOI22_X1 U29822 ( .A1(n24140), .A2(\xmem_data[20][1] ), .B1(n3375), .B2(
        \xmem_data[21][1] ), .ZN(n26349) );
  INV_X1 U29823 ( .A(n26349), .ZN(n26353) );
  AOI22_X1 U29824 ( .A1(n22710), .A2(\xmem_data[18][1] ), .B1(n25416), .B2(
        \xmem_data[19][1] ), .ZN(n26351) );
  NAND2_X1 U29825 ( .A1(n25422), .A2(\xmem_data[23][1] ), .ZN(n26350) );
  NAND2_X1 U29826 ( .A1(n26351), .A2(n26350), .ZN(n26352) );
  NOR2_X1 U29827 ( .A1(n26353), .A2(n26352), .ZN(n26354) );
  NAND2_X1 U29828 ( .A1(n26355), .A2(n26354), .ZN(n26361) );
  AOI22_X1 U29829 ( .A1(n3358), .A2(\xmem_data[24][1] ), .B1(n28233), .B2(
        \xmem_data[25][1] ), .ZN(n26359) );
  AOI22_X1 U29830 ( .A1(n28416), .A2(\xmem_data[26][1] ), .B1(n16986), .B2(
        \xmem_data[27][1] ), .ZN(n26358) );
  AOI22_X1 U29831 ( .A1(n21076), .A2(\xmem_data[28][1] ), .B1(n23795), .B2(
        \xmem_data[29][1] ), .ZN(n26357) );
  AOI22_X1 U29832 ( .A1(n24457), .A2(\xmem_data[30][1] ), .B1(n23764), .B2(
        \xmem_data[31][1] ), .ZN(n26356) );
  NAND4_X1 U29833 ( .A1(n26359), .A2(n26358), .A3(n26357), .A4(n26356), .ZN(
        n26360) );
  OR2_X1 U29834 ( .A1(n26361), .A2(n26360), .ZN(n26362) );
  NOR2_X1 U29835 ( .A1(n26363), .A2(n26362), .ZN(n26364) );
  NOR2_X1 U29836 ( .A1(n26364), .A2(n15043), .ZN(n26365) );
  AOI21_X1 U29837 ( .B1(n26366), .B2(n28490), .A(n26365), .ZN(n26367) );
  OAI22_X1 U29838 ( .A1(n31173), .A2(n35084), .B1(n26370), .B2(n35083), .ZN(
        n31481) );
  XNOR2_X1 U29839 ( .A(n3425), .B(\fmem_data[15][3] ), .ZN(n32205) );
  XNOR2_X1 U29840 ( .A(n32597), .B(\fmem_data[15][3] ), .ZN(n26805) );
  OAI22_X1 U29841 ( .A1(n32205), .A2(n34363), .B1(n26805), .B2(n34364), .ZN(
        n31482) );
  OAI21_X1 U29842 ( .B1(n31483), .B2(n31481), .A(n31482), .ZN(n26372) );
  NAND2_X1 U29843 ( .A1(n31483), .A2(n31481), .ZN(n26371) );
  NAND2_X1 U29844 ( .A1(n26372), .A2(n26371), .ZN(n28918) );
  OAI21_X1 U29845 ( .B1(n28916), .B2(n28917), .A(n28918), .ZN(n26374) );
  NAND2_X1 U29846 ( .A1(n26374), .A2(n26373), .ZN(n34168) );
  XNOR2_X1 U29847 ( .A(n26376), .B(n26375), .ZN(n26378) );
  XNOR2_X1 U29848 ( .A(n26378), .B(n26377), .ZN(n34167) );
  FA_X1 U29849 ( .A(n26381), .B(n26380), .CI(n26379), .CO(n26376), .S(n28408)
         );
  FA_X1 U29850 ( .A(n26384), .B(n26383), .CI(n26382), .CO(n26803), .S(n28407)
         );
  OR2_X1 U29851 ( .A1(n34615), .A2(n3665), .ZN(n26385) );
  OAI22_X1 U29852 ( .A1(n26385), .A2(n34195), .B1(n34194), .B2(n3665), .ZN(
        n31472) );
  AOI22_X1 U29853 ( .A1(n25358), .A2(\xmem_data[8][0] ), .B1(n30571), .B2(
        \xmem_data[9][0] ), .ZN(n26390) );
  AOI22_X1 U29854 ( .A1(n24630), .A2(\xmem_data[10][0] ), .B1(n25360), .B2(
        \xmem_data[11][0] ), .ZN(n26389) );
  AND2_X1 U29855 ( .A1(n3217), .A2(\xmem_data[13][0] ), .ZN(n26386) );
  AOI21_X1 U29856 ( .B1(n30503), .B2(\xmem_data[12][0] ), .A(n26386), .ZN(
        n26388) );
  AOI22_X1 U29857 ( .A1(n24696), .A2(\xmem_data[14][0] ), .B1(n30534), .B2(
        \xmem_data[15][0] ), .ZN(n26387) );
  NAND4_X1 U29858 ( .A1(n26390), .A2(n26389), .A3(n26388), .A4(n26387), .ZN(
        n26406) );
  AOI22_X1 U29859 ( .A1(n30557), .A2(\xmem_data[0][0] ), .B1(n20816), .B2(
        \xmem_data[1][0] ), .ZN(n26394) );
  AOI22_X1 U29860 ( .A1(n24623), .A2(\xmem_data[2][0] ), .B1(n31314), .B2(
        \xmem_data[3][0] ), .ZN(n26393) );
  AOI22_X1 U29861 ( .A1(n3172), .A2(\xmem_data[4][0] ), .B1(n11008), .B2(
        \xmem_data[5][0] ), .ZN(n26392) );
  AOI22_X1 U29862 ( .A1(n27852), .A2(\xmem_data[6][0] ), .B1(n30524), .B2(
        \xmem_data[7][0] ), .ZN(n26391) );
  NAND4_X1 U29863 ( .A1(n26394), .A2(n26393), .A3(n26392), .A4(n26391), .ZN(
        n26405) );
  AOI22_X1 U29864 ( .A1(n20807), .A2(\xmem_data[16][0] ), .B1(n30550), .B2(
        \xmem_data[17][0] ), .ZN(n26398) );
  AOI22_X1 U29865 ( .A1(n28952), .A2(\xmem_data[18][0] ), .B1(n29306), .B2(
        \xmem_data[19][0] ), .ZN(n26397) );
  AOI22_X1 U29866 ( .A1(n30551), .A2(\xmem_data[20][0] ), .B1(n24130), .B2(
        \xmem_data[21][0] ), .ZN(n26396) );
  AOI22_X1 U29867 ( .A1(n20799), .A2(\xmem_data[22][0] ), .B1(n30552), .B2(
        \xmem_data[23][0] ), .ZN(n26395) );
  NAND4_X1 U29868 ( .A1(n26398), .A2(n26397), .A3(n26396), .A4(n26395), .ZN(
        n26404) );
  AOI22_X1 U29869 ( .A1(n30891), .A2(\xmem_data[24][0] ), .B1(n30541), .B2(
        \xmem_data[25][0] ), .ZN(n26402) );
  AOI22_X1 U29870 ( .A1(n25461), .A2(\xmem_data[26][0] ), .B1(n30542), .B2(
        \xmem_data[27][0] ), .ZN(n26401) );
  AOI22_X1 U29871 ( .A1(n24593), .A2(\xmem_data[28][0] ), .B1(n30544), .B2(
        \xmem_data[29][0] ), .ZN(n26400) );
  AOI22_X1 U29872 ( .A1(n27855), .A2(\xmem_data[30][0] ), .B1(n30545), .B2(
        \xmem_data[31][0] ), .ZN(n26399) );
  NAND4_X1 U29873 ( .A1(n26402), .A2(n26401), .A3(n26400), .A4(n26399), .ZN(
        n26403) );
  OR4_X1 U29874 ( .A1(n26406), .A2(n26405), .A3(n26404), .A4(n26403), .ZN(
        n26407) );
  NAND2_X1 U29875 ( .A1(n26407), .A2(n30563), .ZN(n26481) );
  AOI22_X1 U29876 ( .A1(n30588), .A2(\xmem_data[40][0] ), .B1(n30571), .B2(
        \xmem_data[41][0] ), .ZN(n26411) );
  AOI22_X1 U29877 ( .A1(n3306), .A2(\xmem_data[42][0] ), .B1(n27437), .B2(
        \xmem_data[43][0] ), .ZN(n26410) );
  AOI22_X1 U29878 ( .A1(n30503), .A2(\xmem_data[44][0] ), .B1(n3219), .B2(
        \xmem_data[45][0] ), .ZN(n26409) );
  AOI22_X1 U29879 ( .A1(n25693), .A2(\xmem_data[46][0] ), .B1(n20723), .B2(
        \xmem_data[47][0] ), .ZN(n26408) );
  NAND4_X1 U29880 ( .A1(n26411), .A2(n26410), .A3(n26409), .A4(n26408), .ZN(
        n26429) );
  AOI22_X1 U29881 ( .A1(n22683), .A2(\xmem_data[32][0] ), .B1(n30495), .B2(
        \xmem_data[33][0] ), .ZN(n26412) );
  INV_X1 U29882 ( .A(n26412), .ZN(n26416) );
  AOI22_X1 U29883 ( .A1(n30497), .A2(\xmem_data[36][0] ), .B1(n30496), .B2(
        \xmem_data[37][0] ), .ZN(n26414) );
  AOI22_X1 U29884 ( .A1(n24522), .A2(\xmem_data[34][0] ), .B1(n20949), .B2(
        \xmem_data[35][0] ), .ZN(n26413) );
  NAND2_X1 U29885 ( .A1(n26414), .A2(n26413), .ZN(n26415) );
  NOR2_X1 U29886 ( .A1(n26416), .A2(n26415), .ZN(n26427) );
  AOI22_X1 U29887 ( .A1(n24438), .A2(\xmem_data[48][0] ), .B1(n3256), .B2(
        \xmem_data[49][0] ), .ZN(n26420) );
  AOI22_X1 U29888 ( .A1(n25451), .A2(\xmem_data[50][0] ), .B1(n28510), .B2(
        \xmem_data[51][0] ), .ZN(n26419) );
  AOI22_X1 U29889 ( .A1(n30607), .A2(\xmem_data[52][0] ), .B1(n20588), .B2(
        \xmem_data[53][0] ), .ZN(n26418) );
  AOI22_X1 U29890 ( .A1(n30508), .A2(\xmem_data[54][0] ), .B1(n22740), .B2(
        \xmem_data[55][0] ), .ZN(n26417) );
  AOI22_X1 U29891 ( .A1(n3207), .A2(\xmem_data[59][0] ), .B1(
        \xmem_data[58][0] ), .B2(n24213), .ZN(n26424) );
  AOI22_X1 U29892 ( .A1(n28781), .A2(\xmem_data[62][0] ), .B1(n30515), .B2(
        \xmem_data[63][0] ), .ZN(n26423) );
  AOI22_X1 U29893 ( .A1(n30514), .A2(\xmem_data[56][0] ), .B1(n30513), .B2(
        \xmem_data[57][0] ), .ZN(n26422) );
  AOI22_X1 U29894 ( .A1(n20542), .A2(\xmem_data[60][0] ), .B1(n24645), .B2(
        \xmem_data[61][0] ), .ZN(n26421) );
  AOI22_X1 U29895 ( .A1(n23730), .A2(\xmem_data[38][0] ), .B1(n30498), .B2(
        \xmem_data[39][0] ), .ZN(n26425) );
  NAND4_X1 U29896 ( .A1(n26427), .A2(n3823), .A3(n26426), .A4(n26425), .ZN(
        n26428) );
  OAI21_X1 U29897 ( .B1(n26429), .B2(n26428), .A(n30565), .ZN(n26480) );
  AOI22_X1 U29898 ( .A1(n30588), .A2(\xmem_data[72][0] ), .B1(n21309), .B2(
        \xmem_data[73][0] ), .ZN(n26433) );
  AOI22_X1 U29899 ( .A1(n3229), .A2(\xmem_data[74][0] ), .B1(n30589), .B2(
        \xmem_data[75][0] ), .ZN(n26432) );
  AOI22_X1 U29900 ( .A1(n30592), .A2(\xmem_data[76][0] ), .B1(n3220), .B2(
        \xmem_data[77][0] ), .ZN(n26431) );
  AOI22_X1 U29901 ( .A1(n30593), .A2(\xmem_data[78][0] ), .B1(n27444), .B2(
        \xmem_data[79][0] ), .ZN(n26430) );
  NAND4_X1 U29902 ( .A1(n26433), .A2(n26432), .A3(n26431), .A4(n26430), .ZN(
        n26455) );
  NAND2_X1 U29903 ( .A1(n27974), .A2(\xmem_data[64][0] ), .ZN(n26435) );
  NAND2_X1 U29904 ( .A1(n29281), .A2(\xmem_data[65][0] ), .ZN(n26434) );
  NAND2_X1 U29905 ( .A1(n26435), .A2(n26434), .ZN(n26439) );
  AOI22_X1 U29906 ( .A1(n20782), .A2(\xmem_data[68][0] ), .B1(n17003), .B2(
        \xmem_data[69][0] ), .ZN(n26437) );
  AOI22_X1 U29907 ( .A1(n30600), .A2(\xmem_data[66][0] ), .B1(n30599), .B2(
        \xmem_data[67][0] ), .ZN(n26436) );
  NAND2_X1 U29908 ( .A1(n26437), .A2(n26436), .ZN(n26438) );
  NOR2_X1 U29909 ( .A1(n26439), .A2(n26438), .ZN(n26453) );
  AOI22_X1 U29910 ( .A1(n30607), .A2(\xmem_data[84][0] ), .B1(n28415), .B2(
        \xmem_data[85][0] ), .ZN(n26440) );
  INV_X1 U29911 ( .A(n26440), .ZN(n26446) );
  AOI22_X1 U29912 ( .A1(n30608), .A2(\xmem_data[86][0] ), .B1(n21075), .B2(
        \xmem_data[87][0] ), .ZN(n26442) );
  AOI22_X1 U29913 ( .A1(n21074), .A2(\xmem_data[82][0] ), .B1(n28343), .B2(
        \xmem_data[83][0] ), .ZN(n26441) );
  NAND2_X1 U29914 ( .A1(n26442), .A2(n26441), .ZN(n26445) );
  AOI22_X1 U29915 ( .A1(n30606), .A2(\xmem_data[80][0] ), .B1(n20559), .B2(
        \xmem_data[81][0] ), .ZN(n26443) );
  INV_X1 U29916 ( .A(n26443), .ZN(n26444) );
  NOR3_X1 U29917 ( .A1(n26446), .A2(n26445), .A3(n26444), .ZN(n26452) );
  AOI22_X1 U29918 ( .A1(n21005), .A2(\xmem_data[90][0] ), .B1(n30615), .B2(
        \xmem_data[91][0] ), .ZN(n26450) );
  AOI22_X1 U29919 ( .A1(n30614), .A2(\xmem_data[88][0] ), .B1(n30613), .B2(
        \xmem_data[89][0] ), .ZN(n26449) );
  AOI22_X1 U29920 ( .A1(n21007), .A2(\xmem_data[92][0] ), .B1(n21006), .B2(
        \xmem_data[93][0] ), .ZN(n26448) );
  AOI22_X1 U29921 ( .A1(n30617), .A2(\xmem_data[94][0] ), .B1(n30616), .B2(
        \xmem_data[95][0] ), .ZN(n26447) );
  AOI22_X1 U29922 ( .A1(n27717), .A2(\xmem_data[70][0] ), .B1(n30601), .B2(
        \xmem_data[71][0] ), .ZN(n26451) );
  NAND4_X1 U29923 ( .A1(n26453), .A2(n26452), .A3(n3765), .A4(n26451), .ZN(
        n26454) );
  OAI21_X1 U29924 ( .B1(n26455), .B2(n26454), .A(n30628), .ZN(n26479) );
  AOI22_X1 U29925 ( .A1(n30588), .A2(\xmem_data[104][0] ), .B1(n24525), .B2(
        \xmem_data[105][0] ), .ZN(n26459) );
  AOI22_X1 U29926 ( .A1(n3229), .A2(\xmem_data[106][0] ), .B1(n30589), .B2(
        \xmem_data[107][0] ), .ZN(n26458) );
  AOI22_X1 U29927 ( .A1(n30592), .A2(\xmem_data[108][0] ), .B1(n3217), .B2(
        \xmem_data[109][0] ), .ZN(n26457) );
  AOI22_X1 U29928 ( .A1(n30593), .A2(\xmem_data[110][0] ), .B1(n31367), .B2(
        \xmem_data[111][0] ), .ZN(n26456) );
  NAND4_X1 U29929 ( .A1(n26459), .A2(n26458), .A3(n26457), .A4(n26456), .ZN(
        n26477) );
  AOI22_X1 U29930 ( .A1(n24647), .A2(\xmem_data[96][0] ), .B1(n20506), .B2(
        \xmem_data[97][0] ), .ZN(n26464) );
  AOI22_X1 U29931 ( .A1(n30600), .A2(\xmem_data[98][0] ), .B1(n30599), .B2(
        \xmem_data[99][0] ), .ZN(n26463) );
  AOI22_X1 U29932 ( .A1(n20782), .A2(\xmem_data[100][0] ), .B1(n28468), .B2(
        \xmem_data[101][0] ), .ZN(n26462) );
  AND2_X1 U29933 ( .A1(n30601), .A2(\xmem_data[103][0] ), .ZN(n26460) );
  AOI21_X1 U29934 ( .B1(n30901), .B2(\xmem_data[102][0] ), .A(n26460), .ZN(
        n26461) );
  NAND4_X1 U29935 ( .A1(n26464), .A2(n26463), .A3(n26462), .A4(n26461), .ZN(
        n26475) );
  AOI22_X1 U29936 ( .A1(n20939), .A2(\xmem_data[122][0] ), .B1(n30615), .B2(
        \xmem_data[123][0] ), .ZN(n26468) );
  AOI22_X1 U29937 ( .A1(n30614), .A2(\xmem_data[120][0] ), .B1(n30613), .B2(
        \xmem_data[121][0] ), .ZN(n26467) );
  AOI22_X1 U29938 ( .A1(n23764), .A2(\xmem_data[124][0] ), .B1(n25715), .B2(
        \xmem_data[125][0] ), .ZN(n26466) );
  AOI22_X1 U29939 ( .A1(n30617), .A2(\xmem_data[126][0] ), .B1(n30616), .B2(
        \xmem_data[127][0] ), .ZN(n26465) );
  NAND4_X1 U29940 ( .A1(n26468), .A2(n26467), .A3(n26466), .A4(n26465), .ZN(
        n26474) );
  AOI22_X1 U29941 ( .A1(n30606), .A2(\xmem_data[112][0] ), .B1(n17061), .B2(
        \xmem_data[113][0] ), .ZN(n26472) );
  AOI22_X1 U29942 ( .A1(n29567), .A2(\xmem_data[114][0] ), .B1(n28007), .B2(
        \xmem_data[115][0] ), .ZN(n26471) );
  AOI22_X1 U29943 ( .A1(n30607), .A2(\xmem_data[116][0] ), .B1(n14996), .B2(
        \xmem_data[117][0] ), .ZN(n26470) );
  AOI22_X1 U29944 ( .A1(n30608), .A2(\xmem_data[118][0] ), .B1(n28375), .B2(
        \xmem_data[119][0] ), .ZN(n26469) );
  NAND4_X1 U29945 ( .A1(n26472), .A2(n26471), .A3(n26470), .A4(n26469), .ZN(
        n26473) );
  OR3_X1 U29946 ( .A1(n26475), .A2(n26474), .A3(n26473), .ZN(n26476) );
  OAI21_X1 U29947 ( .B1(n26477), .B2(n26476), .A(n30626), .ZN(n26478) );
  NAND4_X2 U29948 ( .A1(n26481), .A2(n26480), .A3(n26479), .A4(n26478), .ZN(
        n36111) );
  OR2_X1 U29949 ( .A1(n36111), .A2(n3677), .ZN(n26482) );
  OAI22_X1 U29950 ( .A1(n26482), .A2(n35034), .B1(n35033), .B2(n3677), .ZN(
        n31471) );
  INV_X1 U29951 ( .A(n33956), .ZN(n26483) );
  INV_X1 U29952 ( .A(n34195), .ZN(n26484) );
  NAND2_X1 U29953 ( .A1(n34615), .A2(n26484), .ZN(n28533) );
  INV_X1 U29954 ( .A(n28533), .ZN(n26485) );
  NAND2_X1 U29955 ( .A1(n29629), .A2(\xmem_data[45][2] ), .ZN(n26487) );
  NAND2_X1 U29956 ( .A1(n30777), .A2(\xmem_data[44][2] ), .ZN(n26486) );
  NAND2_X1 U29957 ( .A1(n26487), .A2(n26486), .ZN(n26490) );
  AOI22_X1 U29958 ( .A1(n30076), .A2(\xmem_data[60][2] ), .B1(n30685), .B2(
        \xmem_data[61][2] ), .ZN(n26488) );
  INV_X1 U29959 ( .A(n26488), .ZN(n26489) );
  NOR2_X1 U29960 ( .A1(n26490), .A2(n26489), .ZN(n26509) );
  NAND2_X1 U29961 ( .A1(n29704), .A2(\xmem_data[49][2] ), .ZN(n26498) );
  NAND2_X1 U29962 ( .A1(n28180), .A2(\xmem_data[48][2] ), .ZN(n26497) );
  NAND2_X1 U29963 ( .A1(n28755), .A2(\xmem_data[58][2] ), .ZN(n26496) );
  AOI22_X1 U29964 ( .A1(n26491), .A2(\xmem_data[46][2] ), .B1(n3137), .B2(
        \xmem_data[47][2] ), .ZN(n26493) );
  AOI22_X1 U29965 ( .A1(n29639), .A2(\xmem_data[59][2] ), .B1(n29627), .B2(
        \xmem_data[43][2] ), .ZN(n26492) );
  NAND2_X1 U29966 ( .A1(n26493), .A2(n26492), .ZN(n26494) );
  AOI21_X1 U29967 ( .B1(n29769), .B2(\xmem_data[52][2] ), .A(n26494), .ZN(
        n26495) );
  AOI22_X1 U29968 ( .A1(n30753), .A2(\xmem_data[32][2] ), .B1(n30752), .B2(
        \xmem_data[33][2] ), .ZN(n26502) );
  AOI22_X1 U29969 ( .A1(n30755), .A2(\xmem_data[34][2] ), .B1(n30754), .B2(
        \xmem_data[35][2] ), .ZN(n26501) );
  AOI22_X1 U29970 ( .A1(n30757), .A2(\xmem_data[36][2] ), .B1(n30756), .B2(
        \xmem_data[37][2] ), .ZN(n26500) );
  AOI22_X1 U29971 ( .A1(n30759), .A2(\xmem_data[38][2] ), .B1(n3144), .B2(
        \xmem_data[39][2] ), .ZN(n26499) );
  NAND4_X1 U29972 ( .A1(n26502), .A2(n26501), .A3(n26500), .A4(n26499), .ZN(
        n26507) );
  AOI22_X1 U29973 ( .A1(n30731), .A2(\xmem_data[50][2] ), .B1(n30744), .B2(
        \xmem_data[51][2] ), .ZN(n26505) );
  NAND2_X1 U29974 ( .A1(n3188), .A2(\xmem_data[57][2] ), .ZN(n26504) );
  NAND2_X1 U29975 ( .A1(n3168), .A2(\xmem_data[56][2] ), .ZN(n26503) );
  NOR2_X1 U29976 ( .A1(n26507), .A2(n26506), .ZN(n26508) );
  NAND3_X1 U29977 ( .A1(n26509), .A2(n3869), .A3(n26508), .ZN(n26518) );
  AOI22_X1 U29978 ( .A1(n30223), .A2(\xmem_data[40][2] ), .B1(n30695), .B2(
        \xmem_data[41][2] ), .ZN(n26516) );
  AOI22_X1 U29979 ( .A1(n30747), .A2(\xmem_data[54][2] ), .B1(n29315), .B2(
        \xmem_data[55][2] ), .ZN(n26513) );
  AOI22_X1 U29980 ( .A1(n30646), .A2(\xmem_data[62][2] ), .B1(n30645), .B2(
        \xmem_data[63][2] ), .ZN(n26512) );
  NAND2_X1 U29981 ( .A1(n28110), .A2(\xmem_data[53][2] ), .ZN(n26511) );
  AOI21_X1 U29982 ( .B1(\xmem_data[42][2] ), .B2(n28207), .A(n26514), .ZN(
        n26515) );
  NAND2_X1 U29983 ( .A1(n26516), .A2(n26515), .ZN(n26517) );
  OAI21_X1 U29984 ( .B1(n26518), .B2(n26517), .A(n30782), .ZN(n26594) );
  AOI22_X1 U29985 ( .A1(n29801), .A2(\xmem_data[80][2] ), .B1(n29589), .B2(
        \xmem_data[81][2] ), .ZN(n26522) );
  AOI22_X1 U29986 ( .A1(n30664), .A2(\xmem_data[82][2] ), .B1(n30663), .B2(
        \xmem_data[83][2] ), .ZN(n26521) );
  AOI22_X1 U29987 ( .A1(n30302), .A2(\xmem_data[84][2] ), .B1(n29768), .B2(
        \xmem_data[85][2] ), .ZN(n26520) );
  AOI22_X1 U29988 ( .A1(n30667), .A2(\xmem_data[86][2] ), .B1(n3158), .B2(
        \xmem_data[87][2] ), .ZN(n26519) );
  NAND4_X1 U29989 ( .A1(n26522), .A2(n26521), .A3(n26520), .A4(n26519), .ZN(
        n26534) );
  AND2_X1 U29990 ( .A1(n30309), .A2(\xmem_data[91][2] ), .ZN(n26523) );
  AOI21_X1 U29991 ( .B1(n30075), .B2(\xmem_data[90][2] ), .A(n26523), .ZN(
        n26527) );
  AOI22_X1 U29992 ( .A1(n3166), .A2(\xmem_data[88][2] ), .B1(n3182), .B2(
        \xmem_data[89][2] ), .ZN(n26526) );
  AOI22_X1 U29993 ( .A1(n29547), .A2(\xmem_data[92][2] ), .B1(n30644), .B2(
        \xmem_data[93][2] ), .ZN(n26525) );
  AOI22_X1 U29994 ( .A1(n30646), .A2(\xmem_data[94][2] ), .B1(n30645), .B2(
        \xmem_data[95][2] ), .ZN(n26524) );
  NAND4_X1 U29995 ( .A1(n26527), .A2(n26526), .A3(n26525), .A4(n26524), .ZN(
        n26533) );
  AOI22_X1 U29996 ( .A1(n30673), .A2(\xmem_data[64][2] ), .B1(n30672), .B2(
        \xmem_data[65][2] ), .ZN(n26531) );
  AOI22_X1 U29997 ( .A1(n30675), .A2(\xmem_data[66][2] ), .B1(n30674), .B2(
        \xmem_data[67][2] ), .ZN(n26530) );
  AOI22_X1 U29998 ( .A1(n30677), .A2(\xmem_data[68][2] ), .B1(n30676), .B2(
        \xmem_data[69][2] ), .ZN(n26529) );
  AOI22_X1 U29999 ( .A1(n30678), .A2(\xmem_data[70][2] ), .B1(n27813), .B2(
        \xmem_data[71][2] ), .ZN(n26528) );
  NAND4_X1 U30000 ( .A1(n26531), .A2(n26530), .A3(n26529), .A4(n26528), .ZN(
        n26532) );
  OR3_X1 U30001 ( .A1(n26534), .A2(n26533), .A3(n26532), .ZN(n26540) );
  AOI22_X1 U30002 ( .A1(n27710), .A2(\xmem_data[72][2] ), .B1(n28766), .B2(
        \xmem_data[73][2] ), .ZN(n26538) );
  AOI22_X1 U30003 ( .A1(n30215), .A2(\xmem_data[74][2] ), .B1(n27708), .B2(
        \xmem_data[75][2] ), .ZN(n26537) );
  AOI22_X1 U30004 ( .A1(n30697), .A2(\xmem_data[76][2] ), .B1(n27833), .B2(
        \xmem_data[77][2] ), .ZN(n26536) );
  AOI22_X1 U30005 ( .A1(n30699), .A2(\xmem_data[78][2] ), .B1(n30698), .B2(
        \xmem_data[79][2] ), .ZN(n26535) );
  NAND4_X1 U30006 ( .A1(n26538), .A2(n26537), .A3(n26536), .A4(n26535), .ZN(
        n26539) );
  OAI21_X1 U30007 ( .B1(n26540), .B2(n26539), .A(n30704), .ZN(n26593) );
  AOI22_X1 U30008 ( .A1(n29481), .A2(\xmem_data[112][2] ), .B1(n27761), .B2(
        \xmem_data[113][2] ), .ZN(n26549) );
  NAND2_X1 U30009 ( .A1(n29592), .A2(\xmem_data[117][2] ), .ZN(n26542) );
  NAND2_X1 U30010 ( .A1(n29769), .A2(\xmem_data[116][2] ), .ZN(n26541) );
  NAND2_X1 U30011 ( .A1(n26542), .A2(n26541), .ZN(n26547) );
  AOI22_X1 U30012 ( .A1(n30667), .A2(\xmem_data[118][2] ), .B1(n29315), .B2(
        \xmem_data[119][2] ), .ZN(n26545) );
  AOI22_X1 U30013 ( .A1(n26543), .A2(\xmem_data[114][2] ), .B1(n30663), .B2(
        \xmem_data[115][2] ), .ZN(n26544) );
  NAND2_X1 U30014 ( .A1(n26545), .A2(n26544), .ZN(n26546) );
  NOR2_X1 U30015 ( .A1(n26547), .A2(n26546), .ZN(n26548) );
  NAND2_X1 U30016 ( .A1(n26549), .A2(n26548), .ZN(n26561) );
  AND2_X1 U30017 ( .A1(n28147), .A2(\xmem_data[123][2] ), .ZN(n26550) );
  AOI21_X1 U30018 ( .B1(n30070), .B2(\xmem_data[122][2] ), .A(n26550), .ZN(
        n26554) );
  AOI22_X1 U30019 ( .A1(n3165), .A2(\xmem_data[120][2] ), .B1(n3185), .B2(
        \xmem_data[121][2] ), .ZN(n26553) );
  AOI22_X1 U30020 ( .A1(n28680), .A2(\xmem_data[124][2] ), .B1(n29487), .B2(
        \xmem_data[125][2] ), .ZN(n26552) );
  AOI22_X1 U30021 ( .A1(n30687), .A2(\xmem_data[126][2] ), .B1(n30686), .B2(
        \xmem_data[127][2] ), .ZN(n26551) );
  NAND4_X1 U30022 ( .A1(n26554), .A2(n26553), .A3(n26552), .A4(n26551), .ZN(
        n26560) );
  AOI22_X1 U30023 ( .A1(n30673), .A2(\xmem_data[96][2] ), .B1(n30672), .B2(
        \xmem_data[97][2] ), .ZN(n26558) );
  AOI22_X1 U30024 ( .A1(n30675), .A2(\xmem_data[98][2] ), .B1(n30674), .B2(
        \xmem_data[99][2] ), .ZN(n26557) );
  AOI22_X1 U30025 ( .A1(n30677), .A2(\xmem_data[100][2] ), .B1(n30676), .B2(
        \xmem_data[101][2] ), .ZN(n26556) );
  AOI22_X1 U30026 ( .A1(n30678), .A2(\xmem_data[102][2] ), .B1(n3149), .B2(
        \xmem_data[103][2] ), .ZN(n26555) );
  NAND4_X1 U30027 ( .A1(n26558), .A2(n26557), .A3(n26556), .A4(n26555), .ZN(
        n26559) );
  AOI22_X1 U30028 ( .A1(n27710), .A2(\xmem_data[104][2] ), .B1(n27013), .B2(
        \xmem_data[105][2] ), .ZN(n26565) );
  AOI22_X1 U30029 ( .A1(n29628), .A2(\xmem_data[106][2] ), .B1(n28137), .B2(
        \xmem_data[107][2] ), .ZN(n26564) );
  AOI22_X1 U30030 ( .A1(n30697), .A2(\xmem_data[108][2] ), .B1(n30776), .B2(
        \xmem_data[109][2] ), .ZN(n26563) );
  AOI22_X1 U30031 ( .A1(n30699), .A2(\xmem_data[110][2] ), .B1(n30698), .B2(
        \xmem_data[111][2] ), .ZN(n26562) );
  NAND4_X1 U30032 ( .A1(n26565), .A2(n26564), .A3(n26563), .A4(n26562), .ZN(
        n26566) );
  OAI21_X1 U30033 ( .B1(n26567), .B2(n26566), .A(n30659), .ZN(n26592) );
  AOI22_X1 U30034 ( .A1(n27703), .A2(\xmem_data[16][2] ), .B1(n28145), .B2(
        \xmem_data[17][2] ), .ZN(n26578) );
  AOI22_X1 U30035 ( .A1(n30745), .A2(\xmem_data[20][2] ), .B1(n28110), .B2(
        \xmem_data[21][2] ), .ZN(n26577) );
  AOI22_X1 U30036 ( .A1(n7041), .A2(\xmem_data[0][2] ), .B1(n7042), .B2(
        \xmem_data[1][2] ), .ZN(n26571) );
  AOI22_X1 U30037 ( .A1(n30722), .A2(\xmem_data[2][2] ), .B1(n25407), .B2(
        \xmem_data[3][2] ), .ZN(n26570) );
  AOI22_X1 U30038 ( .A1(n30724), .A2(\xmem_data[4][2] ), .B1(n30723), .B2(
        \xmem_data[5][2] ), .ZN(n26569) );
  AOI22_X1 U30039 ( .A1(n30725), .A2(\xmem_data[6][2] ), .B1(n3413), .B2(
        \xmem_data[7][2] ), .ZN(n26568) );
  AOI22_X1 U30040 ( .A1(n30732), .A2(\xmem_data[22][2] ), .B1(n27818), .B2(
        \xmem_data[23][2] ), .ZN(n26572) );
  INV_X1 U30041 ( .A(n26572), .ZN(n26575) );
  AOI22_X1 U30042 ( .A1(n30731), .A2(\xmem_data[18][2] ), .B1(n28152), .B2(
        \xmem_data[19][2] ), .ZN(n26573) );
  INV_X1 U30043 ( .A(n26573), .ZN(n26574) );
  NOR2_X1 U30044 ( .A1(n26575), .A2(n26574), .ZN(n26576) );
  NAND4_X1 U30045 ( .A1(n26578), .A2(n26577), .A3(n3770), .A4(n26576), .ZN(
        n26589) );
  AOI22_X1 U30046 ( .A1(n29423), .A2(\xmem_data[10][2] ), .B1(n28218), .B2(
        \xmem_data[11][2] ), .ZN(n26582) );
  AOI22_X1 U30047 ( .A1(n29421), .A2(\xmem_data[8][2] ), .B1(n27013), .B2(
        \xmem_data[9][2] ), .ZN(n26581) );
  AOI22_X1 U30048 ( .A1(n29674), .A2(\xmem_data[12][2] ), .B1(n30217), .B2(
        \xmem_data[13][2] ), .ZN(n26580) );
  AOI22_X1 U30049 ( .A1(n3224), .A2(\xmem_data[14][2] ), .B1(n30710), .B2(
        \xmem_data[15][2] ), .ZN(n26579) );
  NAND4_X1 U30050 ( .A1(n26582), .A2(n26581), .A3(n26580), .A4(n26579), .ZN(
        n26588) );
  AOI22_X1 U30051 ( .A1(n3161), .A2(\xmem_data[24][2] ), .B1(n3188), .B2(
        \xmem_data[25][2] ), .ZN(n26586) );
  AOI22_X1 U30052 ( .A1(n29610), .A2(\xmem_data[26][2] ), .B1(n28147), .B2(
        \xmem_data[27][2] ), .ZN(n26585) );
  AOI22_X1 U30053 ( .A1(n29547), .A2(\xmem_data[28][2] ), .B1(n30685), .B2(
        \xmem_data[29][2] ), .ZN(n26584) );
  AOI22_X1 U30054 ( .A1(n30687), .A2(\xmem_data[30][2] ), .B1(n30311), .B2(
        \xmem_data[31][2] ), .ZN(n26583) );
  NAND4_X1 U30055 ( .A1(n26586), .A2(n26585), .A3(n26584), .A4(n26583), .ZN(
        n26587) );
  OR3_X1 U30056 ( .A1(n26589), .A2(n26588), .A3(n26587), .ZN(n26590) );
  NAND2_X1 U30057 ( .A1(n26590), .A2(n30741), .ZN(n26591) );
  NAND4_X1 U30058 ( .A1(n26594), .A2(n26593), .A3(n26592), .A4(n26591), .ZN(
        n32929) );
  XNOR2_X1 U30059 ( .A(n32929), .B(\fmem_data[23][5] ), .ZN(n32149) );
  AOI22_X1 U30060 ( .A1(n29788), .A2(\xmem_data[72][1] ), .B1(n30775), .B2(
        \xmem_data[73][1] ), .ZN(n26598) );
  AOI22_X1 U30061 ( .A1(n29790), .A2(\xmem_data[74][1] ), .B1(n29494), .B2(
        \xmem_data[75][1] ), .ZN(n26597) );
  AOI22_X1 U30062 ( .A1(n30697), .A2(\xmem_data[76][1] ), .B1(n3198), .B2(
        \xmem_data[77][1] ), .ZN(n26596) );
  AOI22_X1 U30063 ( .A1(n30699), .A2(\xmem_data[78][1] ), .B1(n30698), .B2(
        \xmem_data[79][1] ), .ZN(n26595) );
  NAND4_X1 U30064 ( .A1(n26598), .A2(n26597), .A3(n26596), .A4(n26595), .ZN(
        n26615) );
  AOI22_X1 U30065 ( .A1(n29481), .A2(\xmem_data[80][1] ), .B1(n28738), .B2(
        \xmem_data[81][1] ), .ZN(n26602) );
  AOI22_X1 U30066 ( .A1(n30664), .A2(\xmem_data[82][1] ), .B1(n30663), .B2(
        \xmem_data[83][1] ), .ZN(n26601) );
  AOI22_X1 U30067 ( .A1(n30302), .A2(\xmem_data[84][1] ), .B1(n30237), .B2(
        \xmem_data[85][1] ), .ZN(n26600) );
  AOI22_X1 U30068 ( .A1(n30667), .A2(\xmem_data[86][1] ), .B1(n28154), .B2(
        \xmem_data[87][1] ), .ZN(n26599) );
  NAND4_X1 U30069 ( .A1(n26602), .A2(n26601), .A3(n26600), .A4(n26599), .ZN(
        n26613) );
  AOI22_X1 U30070 ( .A1(n30075), .A2(\xmem_data[90][1] ), .B1(n14971), .B2(
        \xmem_data[91][1] ), .ZN(n26606) );
  AOI22_X1 U30071 ( .A1(n3164), .A2(\xmem_data[88][1] ), .B1(n3184), .B2(
        \xmem_data[89][1] ), .ZN(n26605) );
  AOI22_X1 U30072 ( .A1(n30717), .A2(\xmem_data[92][1] ), .B1(n30716), .B2(
        \xmem_data[93][1] ), .ZN(n26604) );
  AOI22_X1 U30073 ( .A1(n30687), .A2(\xmem_data[94][1] ), .B1(n30686), .B2(
        \xmem_data[95][1] ), .ZN(n26603) );
  NAND4_X1 U30074 ( .A1(n26606), .A2(n26605), .A3(n26604), .A4(n26603), .ZN(
        n26612) );
  AOI22_X1 U30075 ( .A1(n30673), .A2(\xmem_data[64][1] ), .B1(n30672), .B2(
        \xmem_data[65][1] ), .ZN(n26610) );
  AOI22_X1 U30076 ( .A1(n30675), .A2(\xmem_data[66][1] ), .B1(n30674), .B2(
        \xmem_data[67][1] ), .ZN(n26609) );
  AOI22_X1 U30077 ( .A1(n30677), .A2(\xmem_data[68][1] ), .B1(n30676), .B2(
        \xmem_data[69][1] ), .ZN(n26608) );
  AOI22_X1 U30078 ( .A1(n30678), .A2(\xmem_data[70][1] ), .B1(n3149), .B2(
        \xmem_data[71][1] ), .ZN(n26607) );
  NAND4_X1 U30079 ( .A1(n26610), .A2(n26609), .A3(n26608), .A4(n26607), .ZN(
        n26611) );
  OAI21_X1 U30080 ( .B1(n26615), .B2(n26614), .A(n30704), .ZN(n26687) );
  AOI22_X1 U30081 ( .A1(n27710), .A2(\xmem_data[104][1] ), .B1(n29753), .B2(
        \xmem_data[105][1] ), .ZN(n26620) );
  AOI22_X1 U30082 ( .A1(n3392), .A2(\xmem_data[106][1] ), .B1(n29431), .B2(
        \xmem_data[107][1] ), .ZN(n26619) );
  AOI22_X1 U30083 ( .A1(n30697), .A2(\xmem_data[108][1] ), .B1(n3198), .B2(
        \xmem_data[109][1] ), .ZN(n26618) );
  AOI22_X1 U30084 ( .A1(n30699), .A2(\xmem_data[110][1] ), .B1(n30698), .B2(
        \xmem_data[111][1] ), .ZN(n26617) );
  NAND4_X1 U30085 ( .A1(n26620), .A2(n26619), .A3(n26618), .A4(n26617), .ZN(
        n26638) );
  AOI22_X1 U30086 ( .A1(n3249), .A2(\xmem_data[112][1] ), .B1(n29646), .B2(
        \xmem_data[113][1] ), .ZN(n26624) );
  AOI22_X1 U30087 ( .A1(n30664), .A2(\xmem_data[114][1] ), .B1(n30663), .B2(
        \xmem_data[115][1] ), .ZN(n26623) );
  AOI22_X1 U30088 ( .A1(n30250), .A2(\xmem_data[116][1] ), .B1(n30193), .B2(
        \xmem_data[117][1] ), .ZN(n26622) );
  AOI22_X1 U30089 ( .A1(n30667), .A2(\xmem_data[118][1] ), .B1(n29396), .B2(
        \xmem_data[119][1] ), .ZN(n26621) );
  NAND4_X1 U30090 ( .A1(n26624), .A2(n26623), .A3(n26622), .A4(n26621), .ZN(
        n26636) );
  AND2_X1 U30091 ( .A1(n29639), .A2(\xmem_data[123][1] ), .ZN(n26625) );
  AOI21_X1 U30092 ( .B1(n30062), .B2(\xmem_data[122][1] ), .A(n26625), .ZN(
        n26629) );
  AOI22_X1 U30093 ( .A1(n3162), .A2(\xmem_data[120][1] ), .B1(n3189), .B2(
        \xmem_data[121][1] ), .ZN(n26628) );
  AOI22_X1 U30094 ( .A1(n28173), .A2(\xmem_data[124][1] ), .B1(n30685), .B2(
        \xmem_data[125][1] ), .ZN(n26627) );
  AOI22_X1 U30095 ( .A1(n30767), .A2(\xmem_data[126][1] ), .B1(n29379), .B2(
        \xmem_data[127][1] ), .ZN(n26626) );
  NAND4_X1 U30096 ( .A1(n26629), .A2(n26628), .A3(n26627), .A4(n26626), .ZN(
        n26635) );
  AOI22_X1 U30097 ( .A1(n30673), .A2(\xmem_data[96][1] ), .B1(n30672), .B2(
        \xmem_data[97][1] ), .ZN(n26633) );
  AOI22_X1 U30098 ( .A1(n30675), .A2(\xmem_data[98][1] ), .B1(n30674), .B2(
        \xmem_data[99][1] ), .ZN(n26632) );
  AOI22_X1 U30099 ( .A1(n30677), .A2(\xmem_data[100][1] ), .B1(n30676), .B2(
        \xmem_data[101][1] ), .ZN(n26631) );
  AOI22_X1 U30100 ( .A1(n30678), .A2(\xmem_data[102][1] ), .B1(n3149), .B2(
        \xmem_data[103][1] ), .ZN(n26630) );
  NAND4_X1 U30101 ( .A1(n26633), .A2(n26632), .A3(n26631), .A4(n26630), .ZN(
        n26634) );
  OR3_X1 U30102 ( .A1(n26636), .A2(n26635), .A3(n26634), .ZN(n26637) );
  OAI21_X1 U30103 ( .B1(n26638), .B2(n26637), .A(n30659), .ZN(n26686) );
  AOI22_X1 U30104 ( .A1(n7041), .A2(\xmem_data[0][1] ), .B1(n7042), .B2(
        \xmem_data[1][1] ), .ZN(n26642) );
  AOI22_X1 U30105 ( .A1(n30722), .A2(\xmem_data[2][1] ), .B1(n20577), .B2(
        \xmem_data[3][1] ), .ZN(n26641) );
  AOI22_X1 U30106 ( .A1(n30724), .A2(\xmem_data[4][1] ), .B1(n30723), .B2(
        \xmem_data[5][1] ), .ZN(n26640) );
  AOI22_X1 U30107 ( .A1(n30725), .A2(\xmem_data[6][1] ), .B1(n3413), .B2(
        \xmem_data[7][1] ), .ZN(n26639) );
  NAND4_X1 U30108 ( .A1(n26642), .A2(n26641), .A3(n26640), .A4(n26639), .ZN(
        n26645) );
  AOI22_X1 U30109 ( .A1(n30646), .A2(\xmem_data[30][1] ), .B1(n30645), .B2(
        \xmem_data[31][1] ), .ZN(n26643) );
  INV_X1 U30110 ( .A(n26643), .ZN(n26644) );
  NOR2_X1 U30111 ( .A1(n26645), .A2(n26644), .ZN(n26649) );
  AOI22_X1 U30112 ( .A1(n30062), .A2(\xmem_data[26][1] ), .B1(n28754), .B2(
        \xmem_data[27][1] ), .ZN(n26648) );
  AOI22_X1 U30113 ( .A1(n3165), .A2(\xmem_data[24][1] ), .B1(n3188), .B2(
        \xmem_data[25][1] ), .ZN(n26647) );
  AOI22_X1 U30114 ( .A1(n30266), .A2(\xmem_data[29][1] ), .B1(n29722), .B2(
        \xmem_data[28][1] ), .ZN(n26646) );
  NAND4_X1 U30115 ( .A1(n26649), .A2(n26648), .A3(n26647), .A4(n26646), .ZN(
        n26655) );
  AOI22_X1 U30116 ( .A1(n29602), .A2(\xmem_data[16][1] ), .B1(n29589), .B2(
        \xmem_data[17][1] ), .ZN(n26653) );
  AOI22_X1 U30117 ( .A1(n30731), .A2(\xmem_data[18][1] ), .B1(n30083), .B2(
        \xmem_data[19][1] ), .ZN(n26652) );
  AOI22_X1 U30118 ( .A1(n30745), .A2(\xmem_data[20][1] ), .B1(n29592), .B2(
        \xmem_data[21][1] ), .ZN(n26651) );
  AOI22_X1 U30119 ( .A1(n30732), .A2(\xmem_data[22][1] ), .B1(n29605), .B2(
        \xmem_data[23][1] ), .ZN(n26650) );
  NAND4_X1 U30120 ( .A1(n26653), .A2(n26652), .A3(n26651), .A4(n26650), .ZN(
        n26654) );
  NOR2_X1 U30121 ( .A1(n26655), .A2(n26654), .ZN(n26661) );
  AOI22_X1 U30122 ( .A1(n3392), .A2(\xmem_data[10][1] ), .B1(n29832), .B2(
        \xmem_data[11][1] ), .ZN(n26659) );
  AOI22_X1 U30123 ( .A1(n28734), .A2(\xmem_data[8][1] ), .B1(n28206), .B2(
        \xmem_data[9][1] ), .ZN(n26658) );
  AOI22_X1 U30124 ( .A1(n28209), .A2(\xmem_data[12][1] ), .B1(n3198), .B2(
        \xmem_data[13][1] ), .ZN(n26657) );
  AOI22_X1 U30125 ( .A1(n3224), .A2(\xmem_data[14][1] ), .B1(n30710), .B2(
        \xmem_data[15][1] ), .ZN(n26656) );
  NAND2_X1 U30126 ( .A1(n26661), .A2(n26660), .ZN(n26662) );
  NAND2_X1 U30127 ( .A1(n26662), .A2(n30741), .ZN(n26685) );
  AOI22_X1 U30128 ( .A1(n27741), .A2(\xmem_data[40][1] ), .B1(n26510), .B2(
        \xmem_data[41][1] ), .ZN(n26666) );
  AOI22_X1 U30129 ( .A1(n3392), .A2(\xmem_data[42][1] ), .B1(n29422), .B2(
        \xmem_data[43][1] ), .ZN(n26665) );
  AOI22_X1 U30130 ( .A1(n30777), .A2(\xmem_data[44][1] ), .B1(n3170), .B2(
        \xmem_data[45][1] ), .ZN(n26664) );
  AOI22_X1 U30131 ( .A1(n3224), .A2(\xmem_data[46][1] ), .B1(n3132), .B2(
        \xmem_data[47][1] ), .ZN(n26663) );
  NAND4_X1 U30132 ( .A1(n26666), .A2(n26665), .A3(n26664), .A4(n26663), .ZN(
        n26683) );
  AOI22_X1 U30133 ( .A1(n30664), .A2(\xmem_data[50][1] ), .B1(n30744), .B2(
        \xmem_data[51][1] ), .ZN(n26669) );
  AOI22_X1 U30134 ( .A1(n30665), .A2(\xmem_data[52][1] ), .B1(n30084), .B2(
        \xmem_data[53][1] ), .ZN(n26668) );
  AOI22_X1 U30135 ( .A1(n30747), .A2(\xmem_data[54][1] ), .B1(n30746), .B2(
        \xmem_data[55][1] ), .ZN(n26667) );
  NAND4_X1 U30136 ( .A1(n26670), .A2(n26669), .A3(n26668), .A4(n26667), .ZN(
        n26681) );
  AOI22_X1 U30137 ( .A1(n3161), .A2(\xmem_data[56][1] ), .B1(n3184), .B2(
        \xmem_data[57][1] ), .ZN(n26674) );
  AOI22_X1 U30138 ( .A1(n26812), .A2(\xmem_data[58][1] ), .B1(n28147), .B2(
        \xmem_data[59][1] ), .ZN(n26673) );
  AOI22_X1 U30139 ( .A1(n30198), .A2(\xmem_data[60][1] ), .B1(n30170), .B2(
        \xmem_data[61][1] ), .ZN(n26672) );
  AOI22_X1 U30140 ( .A1(n30687), .A2(\xmem_data[62][1] ), .B1(n30686), .B2(
        \xmem_data[63][1] ), .ZN(n26671) );
  NAND4_X1 U30141 ( .A1(n26674), .A2(n26673), .A3(n26672), .A4(n26671), .ZN(
        n26680) );
  AOI22_X1 U30142 ( .A1(n30753), .A2(\xmem_data[32][1] ), .B1(n30752), .B2(
        \xmem_data[33][1] ), .ZN(n26678) );
  AOI22_X1 U30143 ( .A1(n30755), .A2(\xmem_data[34][1] ), .B1(n30754), .B2(
        \xmem_data[35][1] ), .ZN(n26677) );
  AOI22_X1 U30144 ( .A1(n30757), .A2(\xmem_data[36][1] ), .B1(n30756), .B2(
        \xmem_data[37][1] ), .ZN(n26676) );
  AOI22_X1 U30145 ( .A1(n30759), .A2(\xmem_data[38][1] ), .B1(n3144), .B2(
        \xmem_data[39][1] ), .ZN(n26675) );
  NAND4_X1 U30146 ( .A1(n26678), .A2(n26677), .A3(n26676), .A4(n26675), .ZN(
        n26679) );
  OAI21_X1 U30147 ( .B1(n26683), .B2(n26682), .A(n30782), .ZN(n26684) );
  XNOR2_X1 U30148 ( .A(n34361), .B(n3687), .ZN(n31196) );
  OAI22_X1 U30149 ( .A1(n32149), .A2(n34909), .B1(n34908), .B2(n31196), .ZN(
        n31479) );
  AOI22_X1 U30150 ( .A1(n29363), .A2(\xmem_data[80][1] ), .B1(n30765), .B2(
        \xmem_data[81][1] ), .ZN(n26691) );
  AOI22_X1 U30151 ( .A1(n28720), .A2(\xmem_data[82][1] ), .B1(n30311), .B2(
        \xmem_data[83][1] ), .ZN(n26690) );
  AOI22_X1 U30152 ( .A1(n28725), .A2(\xmem_data[84][1] ), .B1(n28724), .B2(
        \xmem_data[85][1] ), .ZN(n26689) );
  AOI22_X1 U30153 ( .A1(n28727), .A2(\xmem_data[86][1] ), .B1(n29298), .B2(
        \xmem_data[87][1] ), .ZN(n26688) );
  NAND4_X1 U30154 ( .A1(n26691), .A2(n26690), .A3(n26689), .A4(n26688), .ZN(
        n26694) );
  AOI22_X1 U30155 ( .A1(n27031), .A2(\xmem_data[78][1] ), .B1(n28754), .B2(
        \xmem_data[79][1] ), .ZN(n26692) );
  INV_X1 U30156 ( .A(n26692), .ZN(n26693) );
  NOR2_X1 U30157 ( .A1(n26694), .A2(n26693), .ZN(n26706) );
  AOI22_X1 U30158 ( .A1(n28740), .A2(\xmem_data[64][1] ), .B1(n30293), .B2(
        \xmem_data[65][1] ), .ZN(n26705) );
  AOI22_X1 U30159 ( .A1(n29705), .A2(\xmem_data[68][1] ), .B1(n29347), .B2(
        \xmem_data[69][1] ), .ZN(n26704) );
  AOI22_X1 U30160 ( .A1(n28753), .A2(\xmem_data[74][1] ), .B1(n30948), .B2(
        \xmem_data[75][1] ), .ZN(n26695) );
  INV_X1 U30161 ( .A(n26695), .ZN(n26702) );
  AOI22_X1 U30162 ( .A1(n28751), .A2(\xmem_data[72][1] ), .B1(n26884), .B2(
        \xmem_data[73][1] ), .ZN(n26696) );
  INV_X1 U30163 ( .A(n26696), .ZN(n26701) );
  AOI22_X1 U30164 ( .A1(n3167), .A2(\xmem_data[76][1] ), .B1(n3183), .B2(
        \xmem_data[77][1] ), .ZN(n26699) );
  AOI22_X1 U30165 ( .A1(n3244), .A2(\xmem_data[66][1] ), .B1(n3126), .B2(
        \xmem_data[67][1] ), .ZN(n26698) );
  AOI22_X1 U30166 ( .A1(n28744), .A2(\xmem_data[70][1] ), .B1(n28743), .B2(
        \xmem_data[71][1] ), .ZN(n26697) );
  NAND2_X1 U30167 ( .A1(n26699), .A2(n3926), .ZN(n26700) );
  NOR3_X1 U30168 ( .A1(n26702), .A2(n26701), .A3(n26700), .ZN(n26703) );
  NAND4_X1 U30169 ( .A1(n26706), .A2(n26705), .A3(n26704), .A4(n26703), .ZN(
        n26712) );
  AOI22_X1 U30170 ( .A1(n29786), .A2(\xmem_data[88][1] ), .B1(n29418), .B2(
        \xmem_data[89][1] ), .ZN(n26710) );
  AOI22_X1 U30171 ( .A1(n28719), .A2(\xmem_data[90][1] ), .B1(n28718), .B2(
        \xmem_data[91][1] ), .ZN(n26709) );
  AOI22_X1 U30172 ( .A1(n29788), .A2(\xmem_data[92][1] ), .B1(n26616), .B2(
        \xmem_data[93][1] ), .ZN(n26708) );
  AOI22_X1 U30173 ( .A1(n29699), .A2(\xmem_data[94][1] ), .B1(n28733), .B2(
        \xmem_data[95][1] ), .ZN(n26707) );
  NAND4_X1 U30174 ( .A1(n26710), .A2(n26709), .A3(n26708), .A4(n26707), .ZN(
        n26711) );
  OAI21_X1 U30175 ( .B1(n26712), .B2(n26711), .A(n28662), .ZN(n26793) );
  AOI22_X1 U30176 ( .A1(n30198), .A2(\xmem_data[112][1] ), .B1(n30765), .B2(
        \xmem_data[113][1] ), .ZN(n26716) );
  AOI22_X1 U30177 ( .A1(n28720), .A2(\xmem_data[114][1] ), .B1(n29573), .B2(
        \xmem_data[115][1] ), .ZN(n26715) );
  AOI22_X1 U30178 ( .A1(n28725), .A2(\xmem_data[116][1] ), .B1(n28724), .B2(
        \xmem_data[117][1] ), .ZN(n26714) );
  AOI22_X1 U30179 ( .A1(n28727), .A2(\xmem_data[118][1] ), .B1(n21060), .B2(
        \xmem_data[119][1] ), .ZN(n26713) );
  NAND4_X1 U30180 ( .A1(n26716), .A2(n26715), .A3(n26714), .A4(n26713), .ZN(
        n26720) );
  AND2_X1 U30181 ( .A1(n28687), .A2(\xmem_data[111][1] ), .ZN(n26717) );
  AOI21_X1 U30182 ( .B1(n28755), .B2(\xmem_data[110][1] ), .A(n26717), .ZN(
        n26718) );
  INV_X1 U30183 ( .A(n26718), .ZN(n26719) );
  NOR2_X1 U30184 ( .A1(n26720), .A2(n26719), .ZN(n26733) );
  AOI22_X1 U30185 ( .A1(n28740), .A2(\xmem_data[96][1] ), .B1(n28786), .B2(
        \xmem_data[97][1] ), .ZN(n26732) );
  AOI22_X1 U30186 ( .A1(n30743), .A2(\xmem_data[100][1] ), .B1(n29704), .B2(
        \xmem_data[101][1] ), .ZN(n26731) );
  AOI22_X1 U30187 ( .A1(n28779), .A2(\xmem_data[104][1] ), .B1(n30090), .B2(
        \xmem_data[105][1] ), .ZN(n26724) );
  AOI22_X1 U30188 ( .A1(n3244), .A2(\xmem_data[98][1] ), .B1(n3126), .B2(
        \xmem_data[99][1] ), .ZN(n26722) );
  AOI22_X1 U30189 ( .A1(n28744), .A2(\xmem_data[102][1] ), .B1(n28743), .B2(
        \xmem_data[103][1] ), .ZN(n26721) );
  NAND2_X1 U30190 ( .A1(n26724), .A2(n26723), .ZN(n26729) );
  AOI22_X1 U30191 ( .A1(n28753), .A2(\xmem_data[106][1] ), .B1(n28091), .B2(
        \xmem_data[107][1] ), .ZN(n26725) );
  INV_X1 U30192 ( .A(n26725), .ZN(n26728) );
  AOI22_X1 U30193 ( .A1(n3167), .A2(\xmem_data[108][1] ), .B1(n3187), .B2(
        \xmem_data[109][1] ), .ZN(n26726) );
  INV_X1 U30194 ( .A(n26726), .ZN(n26727) );
  NOR3_X1 U30195 ( .A1(n26729), .A2(n26728), .A3(n26727), .ZN(n26730) );
  NAND4_X1 U30196 ( .A1(n26733), .A2(n26732), .A3(n26731), .A4(n26730), .ZN(
        n26740) );
  AOI22_X1 U30197 ( .A1(n29829), .A2(\xmem_data[120][1] ), .B1(n29497), .B2(
        \xmem_data[121][1] ), .ZN(n26738) );
  AOI22_X1 U30198 ( .A1(n28719), .A2(\xmem_data[122][1] ), .B1(n28718), .B2(
        \xmem_data[123][1] ), .ZN(n26737) );
  AOI22_X1 U30199 ( .A1(n29788), .A2(\xmem_data[124][1] ), .B1(n30182), .B2(
        \xmem_data[125][1] ), .ZN(n26736) );
  AND2_X1 U30200 ( .A1(n28733), .A2(\xmem_data[127][1] ), .ZN(n26734) );
  AOI21_X1 U30201 ( .B1(n29628), .B2(\xmem_data[126][1] ), .A(n26734), .ZN(
        n26735) );
  NAND4_X1 U30202 ( .A1(n26738), .A2(n26737), .A3(n26736), .A4(n26735), .ZN(
        n26739) );
  OAI21_X1 U30203 ( .B1(n26740), .B2(n26739), .A(n28762), .ZN(n26792) );
  AOI22_X1 U30204 ( .A1(n3167), .A2(\xmem_data[44][1] ), .B1(n3183), .B2(
        \xmem_data[45][1] ), .ZN(n26745) );
  AOI22_X1 U30205 ( .A1(n30635), .A2(\xmem_data[40][1] ), .B1(n30237), .B2(
        \xmem_data[41][1] ), .ZN(n26744) );
  AOI22_X1 U30206 ( .A1(n28686), .A2(\xmem_data[42][1] ), .B1(n20776), .B2(
        \xmem_data[43][1] ), .ZN(n26743) );
  AND2_X1 U30207 ( .A1(n28754), .A2(\xmem_data[47][1] ), .ZN(n26741) );
  AOI21_X1 U30208 ( .B1(n29810), .B2(\xmem_data[46][1] ), .A(n26741), .ZN(
        n26742) );
  NAND4_X1 U30209 ( .A1(n26745), .A2(n26744), .A3(n26743), .A4(n26742), .ZN(
        n26751) );
  AOI22_X1 U30210 ( .A1(n28765), .A2(\xmem_data[56][1] ), .B1(n27723), .B2(
        \xmem_data[57][1] ), .ZN(n26749) );
  AOI22_X1 U30211 ( .A1(n3227), .A2(\xmem_data[58][1] ), .B1(n28677), .B2(
        \xmem_data[59][1] ), .ZN(n26748) );
  AOI22_X1 U30212 ( .A1(n29433), .A2(\xmem_data[60][1] ), .B1(n29831), .B2(
        \xmem_data[61][1] ), .ZN(n26747) );
  AOI22_X1 U30213 ( .A1(n3392), .A2(\xmem_data[62][1] ), .B1(n29832), .B2(
        \xmem_data[63][1] ), .ZN(n26746) );
  NAND4_X1 U30214 ( .A1(n26749), .A2(n26748), .A3(n26747), .A4(n26746), .ZN(
        n26750) );
  OR2_X1 U30215 ( .A1(n26751), .A2(n26750), .ZN(n26764) );
  AOI22_X1 U30216 ( .A1(n29722), .A2(\xmem_data[48][1] ), .B1(n29487), .B2(
        \xmem_data[49][1] ), .ZN(n26755) );
  AOI22_X1 U30217 ( .A1(n28702), .A2(\xmem_data[50][1] ), .B1(n28701), .B2(
        \xmem_data[51][1] ), .ZN(n26754) );
  AOI22_X1 U30218 ( .A1(n28725), .A2(\xmem_data[52][1] ), .B1(n28696), .B2(
        \xmem_data[53][1] ), .ZN(n26753) );
  AOI22_X1 U30219 ( .A1(n28681), .A2(\xmem_data[54][1] ), .B1(n25684), .B2(
        \xmem_data[55][1] ), .ZN(n26752) );
  AOI22_X1 U30220 ( .A1(n29799), .A2(\xmem_data[32][1] ), .B1(n29495), .B2(
        \xmem_data[33][1] ), .ZN(n26762) );
  AOI22_X1 U30221 ( .A1(n29481), .A2(\xmem_data[36][1] ), .B1(n30662), .B2(
        \xmem_data[37][1] ), .ZN(n26761) );
  AOI22_X1 U30222 ( .A1(n28670), .A2(\xmem_data[34][1] ), .B1(n29706), .B2(
        \xmem_data[35][1] ), .ZN(n26756) );
  INV_X1 U30223 ( .A(n26756), .ZN(n26759) );
  AOI22_X1 U30224 ( .A1(n28744), .A2(\xmem_data[38][1] ), .B1(n28671), .B2(
        \xmem_data[39][1] ), .ZN(n26757) );
  INV_X1 U30225 ( .A(n26757), .ZN(n26758) );
  NOR2_X1 U30226 ( .A1(n26759), .A2(n26758), .ZN(n26760) );
  NAND4_X1 U30227 ( .A1(n3856), .A2(n26762), .A3(n26761), .A4(n26760), .ZN(
        n26763) );
  OAI21_X1 U30228 ( .B1(n26764), .B2(n26763), .A(n28713), .ZN(n26791) );
  AOI22_X1 U30229 ( .A1(n28787), .A2(\xmem_data[0][1] ), .B1(n30293), .B2(
        \xmem_data[1][1] ), .ZN(n26768) );
  AOI22_X1 U30230 ( .A1(n3244), .A2(\xmem_data[2][1] ), .B1(n3131), .B2(
        \xmem_data[3][1] ), .ZN(n26767) );
  AOI22_X1 U30231 ( .A1(n29602), .A2(\xmem_data[4][1] ), .B1(n3368), .B2(
        \xmem_data[5][1] ), .ZN(n26766) );
  AOI22_X1 U30232 ( .A1(n28788), .A2(\xmem_data[6][1] ), .B1(n30663), .B2(
        \xmem_data[7][1] ), .ZN(n26765) );
  AND4_X1 U30233 ( .A1(n26768), .A2(n26767), .A3(n26766), .A4(n26765), .ZN(
        n26774) );
  AOI22_X1 U30234 ( .A1(n28779), .A2(\xmem_data[8][1] ), .B1(n29648), .B2(
        \xmem_data[9][1] ), .ZN(n26772) );
  AOI22_X1 U30235 ( .A1(n28753), .A2(\xmem_data[10][1] ), .B1(n27517), .B2(
        \xmem_data[11][1] ), .ZN(n26771) );
  AOI22_X1 U30236 ( .A1(n11444), .A2(\xmem_data[12][1] ), .B1(n3188), .B2(
        \xmem_data[13][1] ), .ZN(n26770) );
  AOI22_X1 U30237 ( .A1(n30062), .A2(\xmem_data[14][1] ), .B1(n28781), .B2(
        \xmem_data[15][1] ), .ZN(n26769) );
  AND4_X1 U30238 ( .A1(n26772), .A2(n26771), .A3(n26770), .A4(n26769), .ZN(
        n26773) );
  NAND2_X1 U30239 ( .A1(n26774), .A2(n26773), .ZN(n26789) );
  AOI22_X1 U30240 ( .A1(n29421), .A2(\xmem_data[28][1] ), .B1(n26510), .B2(
        \xmem_data[29][1] ), .ZN(n26775) );
  INV_X1 U30241 ( .A(n26775), .ZN(n26781) );
  AOI22_X1 U30242 ( .A1(n28700), .A2(\xmem_data[30][1] ), .B1(n30278), .B2(
        \xmem_data[31][1] ), .ZN(n26776) );
  INV_X1 U30243 ( .A(n26776), .ZN(n26780) );
  AOI22_X1 U30244 ( .A1(n28765), .A2(\xmem_data[24][1] ), .B1(n27723), .B2(
        \xmem_data[25][1] ), .ZN(n26778) );
  AOI22_X1 U30245 ( .A1(n3227), .A2(\xmem_data[26][1] ), .B1(n3149), .B2(
        \xmem_data[27][1] ), .ZN(n26777) );
  NAND2_X1 U30246 ( .A1(n26778), .A2(n26777), .ZN(n26779) );
  NOR3_X1 U30247 ( .A1(n26781), .A2(n26780), .A3(n26779), .ZN(n26787) );
  AOI22_X1 U30248 ( .A1(n29363), .A2(\xmem_data[16][1] ), .B1(n30266), .B2(
        \xmem_data[17][1] ), .ZN(n26785) );
  AOI22_X1 U30249 ( .A1(n28720), .A2(\xmem_data[18][1] ), .B1(n30311), .B2(
        \xmem_data[19][1] ), .ZN(n26784) );
  AOI22_X1 U30250 ( .A1(n29819), .A2(\xmem_data[20][1] ), .B1(n28696), .B2(
        \xmem_data[21][1] ), .ZN(n26783) );
  AOI22_X1 U30251 ( .A1(n27806), .A2(\xmem_data[22][1] ), .B1(n28772), .B2(
        \xmem_data[23][1] ), .ZN(n26782) );
  AND4_X1 U30252 ( .A1(n26785), .A2(n26784), .A3(n26783), .A4(n26782), .ZN(
        n26786) );
  NAND2_X1 U30253 ( .A1(n26787), .A2(n26786), .ZN(n26788) );
  OAI21_X1 U30254 ( .B1(n26789), .B2(n26788), .A(n28794), .ZN(n26790) );
  NAND4_X1 U30255 ( .A1(n26793), .A2(n26792), .A3(n26791), .A4(n26790), .ZN(
        n33733) );
  XNOR2_X1 U30256 ( .A(n33733), .B(\fmem_data[11][5] ), .ZN(n31231) );
  XNOR2_X1 U30257 ( .A(n32233), .B(\fmem_data[11][5] ), .ZN(n33972) );
  OAI22_X1 U30258 ( .A1(n31231), .A2(n34933), .B1(n33972), .B2(n34932), .ZN(
        n31478) );
  XNOR2_X1 U30259 ( .A(n26795), .B(n26794), .ZN(n26796) );
  XNOR2_X1 U30260 ( .A(n26797), .B(n26796), .ZN(n34179) );
  FA_X1 U30261 ( .A(n26804), .B(n26803), .CI(n26802), .CO(n26797), .S(n34152)
         );
  XNOR2_X1 U30262 ( .A(n31817), .B(\fmem_data[19][1] ), .ZN(n32151) );
  XNOR2_X1 U30263 ( .A(n31818), .B(\fmem_data[19][1] ), .ZN(n31171) );
  OAI22_X1 U30264 ( .A1(n32151), .A2(n3633), .B1(n31171), .B2(n36226), .ZN(
        n28899) );
  AOI22_X1 U30265 ( .A1(n29390), .A2(\xmem_data[116][1] ), .B1(n29389), .B2(
        \xmem_data[117][1] ), .ZN(n26807) );
  INV_X1 U30266 ( .A(n26807), .ZN(n26811) );
  AOI22_X1 U30267 ( .A1(n3223), .A2(\xmem_data[114][1] ), .B1(n3140), .B2(
        \xmem_data[115][1] ), .ZN(n26809) );
  AOI22_X1 U30268 ( .A1(n29709), .A2(\xmem_data[118][1] ), .B1(n27763), .B2(
        \xmem_data[119][1] ), .ZN(n26808) );
  NAND2_X1 U30269 ( .A1(n26809), .A2(n26808), .ZN(n26810) );
  NOR2_X1 U30270 ( .A1(n26811), .A2(n26810), .ZN(n26822) );
  AOI22_X1 U30271 ( .A1(n27834), .A2(\xmem_data[112][1] ), .B1(n28786), .B2(
        \xmem_data[113][1] ), .ZN(n26821) );
  AOI22_X1 U30272 ( .A1(n3168), .A2(\xmem_data[124][1] ), .B1(n3189), .B2(
        \xmem_data[125][1] ), .ZN(n26816) );
  AOI22_X1 U30273 ( .A1(n27819), .A2(\xmem_data[122][1] ), .B1(n3158), .B2(
        \xmem_data[123][1] ), .ZN(n26815) );
  AOI22_X1 U30274 ( .A1(n29714), .A2(\xmem_data[120][1] ), .B1(n29739), .B2(
        \xmem_data[121][1] ), .ZN(n26814) );
  AOI22_X1 U30275 ( .A1(n26812), .A2(\xmem_data[126][1] ), .B1(n29410), .B2(
        \xmem_data[127][1] ), .ZN(n26813) );
  AOI22_X1 U30276 ( .A1(n28680), .A2(\xmem_data[96][1] ), .B1(n30765), .B2(
        \xmem_data[97][1] ), .ZN(n26820) );
  AOI22_X1 U30277 ( .A1(n27804), .A2(\xmem_data[98][1] ), .B1(n20817), .B2(
        \xmem_data[99][1] ), .ZN(n26819) );
  AOI22_X1 U30278 ( .A1(n29463), .A2(\xmem_data[100][1] ), .B1(n27805), .B2(
        \xmem_data[101][1] ), .ZN(n26818) );
  AOI22_X1 U30279 ( .A1(n27806), .A2(\xmem_data[102][1] ), .B1(n30674), .B2(
        \xmem_data[103][1] ), .ZN(n26817) );
  NAND4_X1 U30280 ( .A1(n26822), .A2(n26821), .A3(n3800), .A4(n3529), .ZN(
        n26828) );
  AOI22_X1 U30281 ( .A1(n7451), .A2(\xmem_data[104][1] ), .B1(n27812), .B2(
        \xmem_data[105][1] ), .ZN(n26826) );
  AOI22_X1 U30282 ( .A1(n27814), .A2(\xmem_data[106][1] ), .B1(n27813), .B2(
        \xmem_data[107][1] ), .ZN(n26825) );
  AOI22_X1 U30283 ( .A1(n28734), .A2(\xmem_data[108][1] ), .B1(n30222), .B2(
        \xmem_data[109][1] ), .ZN(n26824) );
  AOI22_X1 U30284 ( .A1(n28138), .A2(\xmem_data[110][1] ), .B1(n27831), .B2(
        \xmem_data[111][1] ), .ZN(n26823) );
  NAND4_X1 U30285 ( .A1(n26826), .A2(n26825), .A3(n26824), .A4(n26823), .ZN(
        n26827) );
  OAI21_X1 U30286 ( .B1(n26828), .B2(n26827), .A(n27801), .ZN(n26905) );
  AOI22_X1 U30287 ( .A1(n27701), .A2(\xmem_data[48][1] ), .B1(n29761), .B2(
        \xmem_data[49][1] ), .ZN(n26829) );
  AOI22_X1 U30288 ( .A1(n29481), .A2(\xmem_data[52][1] ), .B1(n30190), .B2(
        \xmem_data[53][1] ), .ZN(n26830) );
  AOI22_X1 U30289 ( .A1(n29363), .A2(\xmem_data[32][1] ), .B1(n30266), .B2(
        \xmem_data[33][1] ), .ZN(n26834) );
  AOI22_X1 U30290 ( .A1(n27714), .A2(\xmem_data[34][1] ), .B1(n3270), .B2(
        \xmem_data[35][1] ), .ZN(n26833) );
  AOI22_X1 U30291 ( .A1(n27716), .A2(\xmem_data[36][1] ), .B1(n27715), .B2(
        \xmem_data[37][1] ), .ZN(n26832) );
  AOI22_X1 U30292 ( .A1(n27718), .A2(\xmem_data[38][1] ), .B1(n27717), .B2(
        \xmem_data[39][1] ), .ZN(n26831) );
  AOI22_X1 U30293 ( .A1(n27702), .A2(\xmem_data[50][1] ), .B1(n3147), .B2(
        \xmem_data[51][1] ), .ZN(n26838) );
  AOI22_X1 U30294 ( .A1(n27729), .A2(\xmem_data[58][1] ), .B1(n3158), .B2(
        \xmem_data[59][1] ), .ZN(n26837) );
  NAND2_X1 U30295 ( .A1(n29714), .A2(\xmem_data[56][1] ), .ZN(n26836) );
  NAND2_X1 U30296 ( .A1(n3187), .A2(\xmem_data[61][1] ), .ZN(n26835) );
  NAND4_X1 U30297 ( .A1(n26838), .A2(n26837), .A3(n26836), .A4(n26835), .ZN(
        n26845) );
  NAND2_X1 U30298 ( .A1(n28689), .A2(\xmem_data[62][1] ), .ZN(n26843) );
  AOI22_X1 U30299 ( .A1(n30237), .A2(\xmem_data[57][1] ), .B1(n3168), .B2(
        \xmem_data[60][1] ), .ZN(n26842) );
  AOI22_X1 U30300 ( .A1(n26879), .A2(\xmem_data[54][1] ), .B1(n27763), .B2(
        \xmem_data[55][1] ), .ZN(n26840) );
  NAND2_X1 U30301 ( .A1(n27825), .A2(\xmem_data[63][1] ), .ZN(n26839) );
  NAND3_X1 U30302 ( .A1(n26843), .A2(n26842), .A3(n26841), .ZN(n26844) );
  NOR2_X1 U30303 ( .A1(n26845), .A2(n26844), .ZN(n26846) );
  NAND4_X1 U30304 ( .A1(n26829), .A2(n26830), .A3(n3477), .A4(n26846), .ZN(
        n26852) );
  AOI22_X1 U30305 ( .A1(n29829), .A2(\xmem_data[40][1] ), .B1(n27723), .B2(
        \xmem_data[41][1] ), .ZN(n26850) );
  AOI22_X1 U30306 ( .A1(n11850), .A2(\xmem_data[42][1] ), .B1(n3149), .B2(
        \xmem_data[43][1] ), .ZN(n26849) );
  AOI22_X1 U30307 ( .A1(n28136), .A2(\xmem_data[44][1] ), .B1(n26616), .B2(
        \xmem_data[45][1] ), .ZN(n26848) );
  AOI22_X1 U30308 ( .A1(n29699), .A2(\xmem_data[46][1] ), .B1(n27708), .B2(
        \xmem_data[47][1] ), .ZN(n26847) );
  NAND4_X1 U30309 ( .A1(n26850), .A2(n26849), .A3(n26848), .A4(n26847), .ZN(
        n26851) );
  OAI21_X1 U30310 ( .B1(n26852), .B2(n26851), .A(n27737), .ZN(n26904) );
  AOI22_X1 U30311 ( .A1(n30191), .A2(\xmem_data[20][1] ), .B1(n27761), .B2(
        \xmem_data[21][1] ), .ZN(n26856) );
  AOI22_X1 U30312 ( .A1(n3223), .A2(\xmem_data[18][1] ), .B1(n30295), .B2(
        \xmem_data[19][1] ), .ZN(n26855) );
  AOI22_X1 U30313 ( .A1(n27771), .A2(\xmem_data[16][1] ), .B1(n30696), .B2(
        \xmem_data[17][1] ), .ZN(n26854) );
  AOI22_X1 U30314 ( .A1(n29709), .A2(\xmem_data[22][1] ), .B1(n30083), .B2(
        \xmem_data[23][1] ), .ZN(n26853) );
  NAND4_X1 U30315 ( .A1(n26856), .A2(n26855), .A3(n26854), .A4(n26853), .ZN(
        n26862) );
  AOI22_X1 U30316 ( .A1(n3164), .A2(\xmem_data[28][1] ), .B1(n3183), .B2(
        \xmem_data[29][1] ), .ZN(n26860) );
  AOI22_X1 U30317 ( .A1(n30715), .A2(\xmem_data[30][1] ), .B1(n25400), .B2(
        \xmem_data[31][1] ), .ZN(n26859) );
  AOI22_X1 U30318 ( .A1(n27756), .A2(\xmem_data[26][1] ), .B1(n20718), .B2(
        \xmem_data[27][1] ), .ZN(n26858) );
  AOI22_X1 U30319 ( .A1(n30635), .A2(\xmem_data[24][1] ), .B1(n27753), .B2(
        \xmem_data[25][1] ), .ZN(n26857) );
  NAND4_X1 U30320 ( .A1(n26860), .A2(n26859), .A3(n26858), .A4(n26857), .ZN(
        n26861) );
  NOR2_X1 U30321 ( .A1(n26862), .A2(n26861), .ZN(n26867) );
  AOI22_X1 U30322 ( .A1(n30717), .A2(\xmem_data[0][1] ), .B1(n29721), .B2(
        \xmem_data[1][1] ), .ZN(n26866) );
  AOI22_X1 U30323 ( .A1(n7446), .A2(\xmem_data[2][1] ), .B1(n20732), .B2(
        \xmem_data[3][1] ), .ZN(n26865) );
  AOI22_X1 U30324 ( .A1(n29777), .A2(\xmem_data[4][1] ), .B1(n27805), .B2(
        \xmem_data[5][1] ), .ZN(n26864) );
  AOI22_X1 U30325 ( .A1(n28681), .A2(\xmem_data[6][1] ), .B1(n20826), .B2(
        \xmem_data[7][1] ), .ZN(n26863) );
  NAND2_X1 U30326 ( .A1(n26867), .A2(n3783), .ZN(n26873) );
  AOI22_X1 U30327 ( .A1(n29829), .A2(\xmem_data[8][1] ), .B1(n27743), .B2(
        \xmem_data[9][1] ), .ZN(n26871) );
  AOI22_X1 U30328 ( .A1(n27742), .A2(\xmem_data[10][1] ), .B1(n3144), .B2(
        \xmem_data[11][1] ), .ZN(n26870) );
  AOI22_X1 U30329 ( .A1(n29433), .A2(\xmem_data[12][1] ), .B1(n30182), .B2(
        \xmem_data[13][1] ), .ZN(n26869) );
  AOI22_X1 U30330 ( .A1(n29628), .A2(\xmem_data[14][1] ), .B1(n28218), .B2(
        \xmem_data[15][1] ), .ZN(n26868) );
  NAND4_X1 U30331 ( .A1(n26871), .A2(n26870), .A3(n26869), .A4(n26868), .ZN(
        n26872) );
  OAI21_X1 U30332 ( .B1(n26873), .B2(n26872), .A(n27778), .ZN(n26903) );
  AOI22_X1 U30333 ( .A1(n30198), .A2(\xmem_data[64][1] ), .B1(n29487), .B2(
        \xmem_data[65][1] ), .ZN(n26877) );
  AOI22_X1 U30334 ( .A1(n27804), .A2(\xmem_data[66][1] ), .B1(n28226), .B2(
        \xmem_data[67][1] ), .ZN(n26876) );
  AOI22_X1 U30335 ( .A1(n29382), .A2(\xmem_data[68][1] ), .B1(n27805), .B2(
        \xmem_data[69][1] ), .ZN(n26875) );
  AOI22_X1 U30336 ( .A1(n27806), .A2(\xmem_data[70][1] ), .B1(n30674), .B2(
        \xmem_data[71][1] ), .ZN(n26874) );
  AOI22_X1 U30337 ( .A1(n29421), .A2(\xmem_data[76][1] ), .B1(n28766), .B2(
        \xmem_data[77][1] ), .ZN(n26900) );
  AOI22_X1 U30338 ( .A1(n30279), .A2(\xmem_data[78][1] ), .B1(n27831), .B2(
        \xmem_data[79][1] ), .ZN(n26899) );
  AOI22_X1 U30339 ( .A1(n26878), .A2(\xmem_data[82][1] ), .B1(n30710), .B2(
        \xmem_data[83][1] ), .ZN(n26881) );
  AOI22_X1 U30340 ( .A1(n26879), .A2(\xmem_data[86][1] ), .B1(n28233), .B2(
        \xmem_data[87][1] ), .ZN(n26880) );
  NAND2_X1 U30341 ( .A1(n26881), .A2(n26880), .ZN(n26882) );
  AOI21_X1 U30342 ( .B1(n27834), .B2(\xmem_data[80][1] ), .A(n26882), .ZN(
        n26888) );
  AND2_X1 U30343 ( .A1(n27825), .A2(\xmem_data[95][1] ), .ZN(n26883) );
  AOI21_X1 U30344 ( .B1(n3184), .B2(\xmem_data[93][1] ), .A(n26883), .ZN(
        n26887) );
  NAND2_X1 U30345 ( .A1(n30301), .A2(\xmem_data[89][1] ), .ZN(n26886) );
  NAND2_X1 U30346 ( .A1(n3197), .A2(\xmem_data[81][1] ), .ZN(n26885) );
  NAND4_X1 U30347 ( .A1(n26888), .A2(n26887), .A3(n26886), .A4(n26885), .ZN(
        n26897) );
  AOI22_X1 U30348 ( .A1(\xmem_data[92][1] ), .A2(n3162), .B1(n30250), .B2(
        \xmem_data[88][1] ), .ZN(n26892) );
  NAND2_X1 U30349 ( .A1(n27031), .A2(\xmem_data[94][1] ), .ZN(n26891) );
  NAND2_X1 U30350 ( .A1(n28739), .A2(\xmem_data[84][1] ), .ZN(n26890) );
  NAND2_X1 U30351 ( .A1(n3368), .A2(\xmem_data[85][1] ), .ZN(n26889) );
  NAND4_X1 U30352 ( .A1(n26892), .A2(n26891), .A3(n26890), .A4(n26889), .ZN(
        n26896) );
  AOI22_X1 U30353 ( .A1(n7451), .A2(\xmem_data[72][1] ), .B1(n27812), .B2(
        \xmem_data[73][1] ), .ZN(n26895) );
  AOI22_X1 U30354 ( .A1(n27819), .A2(\xmem_data[90][1] ), .B1(n20776), .B2(
        \xmem_data[91][1] ), .ZN(n26894) );
  AOI22_X1 U30355 ( .A1(n27814), .A2(\xmem_data[74][1] ), .B1(n27813), .B2(
        \xmem_data[75][1] ), .ZN(n26893) );
  NOR3_X1 U30356 ( .A1(n26897), .A2(n26896), .A3(n3998), .ZN(n26898) );
  NAND4_X1 U30357 ( .A1(n3867), .A2(n26900), .A3(n26899), .A4(n26898), .ZN(
        n26901) );
  NAND2_X1 U30358 ( .A1(n26901), .A2(n27839), .ZN(n26902) );
  NAND4_X1 U30359 ( .A1(n26905), .A2(n26904), .A3(n26903), .A4(n26902), .ZN(
        n34334) );
  XNOR2_X1 U30360 ( .A(n34334), .B(\fmem_data[27][5] ), .ZN(n31248) );
  XNOR2_X1 U30361 ( .A(n32978), .B(\fmem_data[27][5] ), .ZN(n32307) );
  OAI22_X1 U30362 ( .A1(n31248), .A2(n34904), .B1(n34903), .B2(n32307), .ZN(
        n28898) );
  AOI22_X1 U30363 ( .A1(n29849), .A2(\xmem_data[32][1] ), .B1(n29848), .B2(
        \xmem_data[33][1] ), .ZN(n26909) );
  AOI22_X1 U30364 ( .A1(n29851), .A2(\xmem_data[34][1] ), .B1(n29850), .B2(
        \xmem_data[35][1] ), .ZN(n26908) );
  AOI22_X1 U30365 ( .A1(n29853), .A2(\xmem_data[36][1] ), .B1(n29852), .B2(
        \xmem_data[37][1] ), .ZN(n26907) );
  AOI22_X1 U30366 ( .A1(n29855), .A2(\xmem_data[38][1] ), .B1(n29854), .B2(
        \xmem_data[39][1] ), .ZN(n26906) );
  AND4_X1 U30367 ( .A1(n26909), .A2(n26908), .A3(n26907), .A4(n26906), .ZN(
        n26925) );
  AOI22_X1 U30368 ( .A1(n29860), .A2(\xmem_data[40][1] ), .B1(n29976), .B2(
        \xmem_data[41][1] ), .ZN(n26913) );
  AOI22_X1 U30369 ( .A1(n29978), .A2(\xmem_data[42][1] ), .B1(n3194), .B2(
        \xmem_data[43][1] ), .ZN(n26912) );
  AOI22_X1 U30370 ( .A1(n29980), .A2(\xmem_data[44][1] ), .B1(n29944), .B2(
        \xmem_data[45][1] ), .ZN(n26911) );
  AOI22_X1 U30371 ( .A1(n29982), .A2(\xmem_data[46][1] ), .B1(n29946), .B2(
        \xmem_data[47][1] ), .ZN(n26910) );
  AND4_X1 U30372 ( .A1(n26913), .A2(n26912), .A3(n26911), .A4(n26910), .ZN(
        n26924) );
  AOI22_X1 U30373 ( .A1(n29866), .A2(\xmem_data[48][1] ), .B1(n29865), .B2(
        \xmem_data[49][1] ), .ZN(n26917) );
  AOI22_X1 U30374 ( .A1(n29868), .A2(\xmem_data[50][1] ), .B1(n29867), .B2(
        \xmem_data[51][1] ), .ZN(n26916) );
  AOI22_X1 U30375 ( .A1(n29870), .A2(\xmem_data[52][1] ), .B1(n29918), .B2(
        \xmem_data[53][1] ), .ZN(n26915) );
  AOI22_X1 U30376 ( .A1(n29871), .A2(\xmem_data[54][1] ), .B1(n29993), .B2(
        \xmem_data[55][1] ), .ZN(n26914) );
  AND4_X1 U30377 ( .A1(n26917), .A2(n26916), .A3(n26915), .A4(n26914), .ZN(
        n26923) );
  AOI22_X1 U30378 ( .A1(n29877), .A2(\xmem_data[56][1] ), .B1(n29876), .B2(
        \xmem_data[57][1] ), .ZN(n26921) );
  AOI22_X1 U30379 ( .A1(n29879), .A2(\xmem_data[58][1] ), .B1(n29878), .B2(
        \xmem_data[59][1] ), .ZN(n26920) );
  AOI22_X1 U30380 ( .A1(n29881), .A2(\xmem_data[60][1] ), .B1(n29880), .B2(
        \xmem_data[61][1] ), .ZN(n26919) );
  AOI22_X1 U30381 ( .A1(n29883), .A2(\xmem_data[62][1] ), .B1(n29882), .B2(
        \xmem_data[63][1] ), .ZN(n26918) );
  AND4_X1 U30382 ( .A1(n26921), .A2(n26920), .A3(n26919), .A4(n26918), .ZN(
        n26922) );
  NAND4_X1 U30383 ( .A1(n26925), .A2(n26924), .A3(n26923), .A4(n26922), .ZN(
        n26947) );
  AOI22_X1 U30384 ( .A1(n29915), .A2(\xmem_data[16][1] ), .B1(n29914), .B2(
        \xmem_data[17][1] ), .ZN(n26929) );
  AOI22_X1 U30385 ( .A1(n29917), .A2(\xmem_data[18][1] ), .B1(n29916), .B2(
        \xmem_data[19][1] ), .ZN(n26928) );
  AOI22_X1 U30386 ( .A1(n29919), .A2(\xmem_data[20][1] ), .B1(n29918), .B2(
        \xmem_data[21][1] ), .ZN(n26927) );
  AOI22_X1 U30387 ( .A1(n29921), .A2(\xmem_data[22][1] ), .B1(n29920), .B2(
        \xmem_data[23][1] ), .ZN(n26926) );
  AND4_X1 U30388 ( .A1(n26929), .A2(n26928), .A3(n26927), .A4(n26926), .ZN(
        n26945) );
  AOI22_X1 U30389 ( .A1(n29904), .A2(\xmem_data[8][1] ), .B1(n29976), .B2(
        \xmem_data[9][1] ), .ZN(n26933) );
  AOI22_X1 U30390 ( .A1(n29905), .A2(\xmem_data[10][1] ), .B1(n3195), .B2(
        \xmem_data[11][1] ), .ZN(n26932) );
  AOI22_X1 U30391 ( .A1(n29907), .A2(\xmem_data[12][1] ), .B1(n29906), .B2(
        \xmem_data[13][1] ), .ZN(n26931) );
  AOI22_X1 U30392 ( .A1(n29909), .A2(\xmem_data[14][1] ), .B1(n29946), .B2(
        \xmem_data[15][1] ), .ZN(n26930) );
  AND4_X1 U30393 ( .A1(n26933), .A2(n26932), .A3(n26931), .A4(n26930), .ZN(
        n26944) );
  AOI22_X1 U30394 ( .A1(n29893), .A2(\xmem_data[0][1] ), .B1(n29892), .B2(
        \xmem_data[1][1] ), .ZN(n26937) );
  AOI22_X1 U30395 ( .A1(n29895), .A2(\xmem_data[2][1] ), .B1(n29894), .B2(
        \xmem_data[3][1] ), .ZN(n26936) );
  AOI22_X1 U30396 ( .A1(n29897), .A2(\xmem_data[4][1] ), .B1(n29896), .B2(
        \xmem_data[5][1] ), .ZN(n26935) );
  AOI22_X1 U30397 ( .A1(n29899), .A2(\xmem_data[6][1] ), .B1(n29898), .B2(
        \xmem_data[7][1] ), .ZN(n26934) );
  AND4_X1 U30398 ( .A1(n26937), .A2(n26936), .A3(n26935), .A4(n26934), .ZN(
        n26943) );
  AOI22_X1 U30399 ( .A1(n3243), .A2(\xmem_data[24][1] ), .B1(n3242), .B2(
        \xmem_data[25][1] ), .ZN(n26941) );
  AOI22_X1 U30400 ( .A1(n3235), .A2(\xmem_data[26][1] ), .B1(n3238), .B2(
        \xmem_data[27][1] ), .ZN(n26940) );
  AOI22_X1 U30401 ( .A1(n3236), .A2(\xmem_data[28][1] ), .B1(n3225), .B2(
        \xmem_data[29][1] ), .ZN(n26939) );
  AOI22_X1 U30402 ( .A1(n3237), .A2(\xmem_data[30][1] ), .B1(n3234), .B2(
        \xmem_data[31][1] ), .ZN(n26938) );
  AND4_X1 U30403 ( .A1(n26941), .A2(n26940), .A3(n26939), .A4(n26938), .ZN(
        n26942) );
  NAND4_X1 U30404 ( .A1(n26945), .A2(n26944), .A3(n26943), .A4(n26942), .ZN(
        n26946) );
  AOI22_X1 U30405 ( .A1(n26947), .A2(n29937), .B1(n26946), .B2(n29935), .ZN(
        n26991) );
  AOI22_X1 U30406 ( .A1(n29966), .A2(\xmem_data[96][1] ), .B1(n29965), .B2(
        \xmem_data[97][1] ), .ZN(n26951) );
  AOI22_X1 U30407 ( .A1(n29968), .A2(\xmem_data[98][1] ), .B1(n29967), .B2(
        \xmem_data[99][1] ), .ZN(n26950) );
  AOI22_X1 U30408 ( .A1(n29969), .A2(\xmem_data[100][1] ), .B1(n29896), .B2(
        \xmem_data[101][1] ), .ZN(n26949) );
  AOI22_X1 U30409 ( .A1(n29971), .A2(\xmem_data[102][1] ), .B1(n29970), .B2(
        \xmem_data[103][1] ), .ZN(n26948) );
  AND4_X1 U30410 ( .A1(n26951), .A2(n26950), .A3(n26949), .A4(n26948), .ZN(
        n26967) );
  AOI22_X1 U30411 ( .A1(n29977), .A2(\xmem_data[104][1] ), .B1(n29976), .B2(
        \xmem_data[105][1] ), .ZN(n26955) );
  AOI22_X1 U30412 ( .A1(n29943), .A2(\xmem_data[106][1] ), .B1(n3196), .B2(
        \xmem_data[107][1] ), .ZN(n26954) );
  AOI22_X1 U30413 ( .A1(n29945), .A2(\xmem_data[108][1] ), .B1(n29944), .B2(
        \xmem_data[109][1] ), .ZN(n26953) );
  AOI22_X1 U30414 ( .A1(n29947), .A2(\xmem_data[110][1] ), .B1(n29946), .B2(
        \xmem_data[111][1] ), .ZN(n26952) );
  AND4_X1 U30415 ( .A1(n26955), .A2(n26954), .A3(n26953), .A4(n26952), .ZN(
        n26966) );
  AOI22_X1 U30416 ( .A1(n29988), .A2(\xmem_data[112][1] ), .B1(n29987), .B2(
        \xmem_data[113][1] ), .ZN(n26959) );
  AOI22_X1 U30417 ( .A1(n29990), .A2(\xmem_data[114][1] ), .B1(n29989), .B2(
        \xmem_data[115][1] ), .ZN(n26958) );
  AOI22_X1 U30418 ( .A1(n29992), .A2(\xmem_data[116][1] ), .B1(n29991), .B2(
        \xmem_data[117][1] ), .ZN(n26957) );
  AOI22_X1 U30419 ( .A1(n29994), .A2(\xmem_data[118][1] ), .B1(n29993), .B2(
        \xmem_data[119][1] ), .ZN(n26956) );
  AND4_X1 U30420 ( .A1(n26959), .A2(n26958), .A3(n26957), .A4(n26956), .ZN(
        n26965) );
  AOI22_X1 U30421 ( .A1(n3243), .A2(\xmem_data[120][1] ), .B1(n3242), .B2(
        \xmem_data[121][1] ), .ZN(n26963) );
  AOI22_X1 U30422 ( .A1(n3235), .A2(\xmem_data[122][1] ), .B1(n3238), .B2(
        \xmem_data[123][1] ), .ZN(n26962) );
  AOI22_X1 U30423 ( .A1(n3236), .A2(\xmem_data[124][1] ), .B1(n3225), .B2(
        \xmem_data[125][1] ), .ZN(n26961) );
  AOI22_X1 U30424 ( .A1(n3237), .A2(\xmem_data[126][1] ), .B1(n3234), .B2(
        \xmem_data[127][1] ), .ZN(n26960) );
  AND4_X1 U30425 ( .A1(n26963), .A2(n26962), .A3(n26961), .A4(n26960), .ZN(
        n26964) );
  NAND4_X1 U30426 ( .A1(n26967), .A2(n26966), .A3(n26965), .A4(n26964), .ZN(
        n26989) );
  AOI22_X1 U30427 ( .A1(n29966), .A2(\xmem_data[64][1] ), .B1(n29965), .B2(
        \xmem_data[65][1] ), .ZN(n26971) );
  AOI22_X1 U30428 ( .A1(n29968), .A2(\xmem_data[66][1] ), .B1(n29967), .B2(
        \xmem_data[67][1] ), .ZN(n26970) );
  AOI22_X1 U30429 ( .A1(n29969), .A2(\xmem_data[68][1] ), .B1(n29896), .B2(
        \xmem_data[69][1] ), .ZN(n26969) );
  AOI22_X1 U30430 ( .A1(n29971), .A2(\xmem_data[70][1] ), .B1(n29970), .B2(
        \xmem_data[71][1] ), .ZN(n26968) );
  AND4_X1 U30431 ( .A1(n26971), .A2(n26970), .A3(n26969), .A4(n26968), .ZN(
        n26987) );
  AOI22_X1 U30432 ( .A1(n29977), .A2(\xmem_data[72][1] ), .B1(n29976), .B2(
        \xmem_data[73][1] ), .ZN(n26975) );
  AOI22_X1 U30433 ( .A1(n29943), .A2(\xmem_data[74][1] ), .B1(n3194), .B2(
        \xmem_data[75][1] ), .ZN(n26974) );
  AOI22_X1 U30434 ( .A1(n29945), .A2(\xmem_data[76][1] ), .B1(n29979), .B2(
        \xmem_data[77][1] ), .ZN(n26973) );
  AOI22_X1 U30435 ( .A1(n29947), .A2(\xmem_data[78][1] ), .B1(n29981), .B2(
        \xmem_data[79][1] ), .ZN(n26972) );
  AND4_X1 U30436 ( .A1(n26975), .A2(n26974), .A3(n26973), .A4(n26972), .ZN(
        n26986) );
  AOI22_X1 U30437 ( .A1(n29988), .A2(\xmem_data[80][1] ), .B1(n29987), .B2(
        \xmem_data[81][1] ), .ZN(n26979) );
  AOI22_X1 U30438 ( .A1(n29990), .A2(\xmem_data[82][1] ), .B1(n29989), .B2(
        \xmem_data[83][1] ), .ZN(n26978) );
  AOI22_X1 U30439 ( .A1(n29992), .A2(\xmem_data[84][1] ), .B1(n29991), .B2(
        \xmem_data[85][1] ), .ZN(n26977) );
  AOI22_X1 U30440 ( .A1(n29994), .A2(\xmem_data[86][1] ), .B1(n29993), .B2(
        \xmem_data[87][1] ), .ZN(n26976) );
  AND4_X1 U30441 ( .A1(n26979), .A2(n26978), .A3(n26977), .A4(n26976), .ZN(
        n26985) );
  AOI22_X1 U30442 ( .A1(n3243), .A2(\xmem_data[88][1] ), .B1(n3242), .B2(
        \xmem_data[89][1] ), .ZN(n26983) );
  AOI22_X1 U30443 ( .A1(n3235), .A2(\xmem_data[90][1] ), .B1(n3238), .B2(
        \xmem_data[91][1] ), .ZN(n26982) );
  AOI22_X1 U30444 ( .A1(n3236), .A2(\xmem_data[92][1] ), .B1(n3225), .B2(
        \xmem_data[93][1] ), .ZN(n26981) );
  AOI22_X1 U30445 ( .A1(n3237), .A2(\xmem_data[94][1] ), .B1(n3234), .B2(
        \xmem_data[95][1] ), .ZN(n26980) );
  AND4_X1 U30446 ( .A1(n26983), .A2(n26982), .A3(n26981), .A4(n26980), .ZN(
        n26984) );
  NAND4_X1 U30447 ( .A1(n26987), .A2(n26986), .A3(n26985), .A4(n26984), .ZN(
        n26988) );
  AOI22_X1 U30448 ( .A1(n30007), .A2(n26989), .B1(n30009), .B2(n26988), .ZN(
        n26990) );
  NAND2_X1 U30449 ( .A1(n26991), .A2(n26990), .ZN(n32939) );
  XNOR2_X1 U30450 ( .A(n32936), .B(\fmem_data[19][5] ), .ZN(n32182) );
  AOI22_X1 U30451 ( .A1(n30191), .A2(\xmem_data[12][1] ), .B1(n28145), .B2(
        \xmem_data[13][1] ), .ZN(n26992) );
  INV_X1 U30452 ( .A(n26992), .ZN(n26997) );
  AOI22_X1 U30453 ( .A1(n29799), .A2(\xmem_data[8][1] ), .B1(n3170), .B2(
        \xmem_data[9][1] ), .ZN(n26995) );
  AOI22_X1 U30454 ( .A1(n29709), .A2(\xmem_data[14][1] ), .B1(n30886), .B2(
        \xmem_data[15][1] ), .ZN(n26994) );
  AOI22_X1 U30455 ( .A1(n29707), .A2(\xmem_data[10][1] ), .B1(n29762), .B2(
        \xmem_data[11][1] ), .ZN(n26993) );
  NOR2_X1 U30456 ( .A1(n26997), .A2(n26996), .ZN(n27012) );
  AOI22_X1 U30457 ( .A1(n28685), .A2(\xmem_data[16][1] ), .B1(n30193), .B2(
        \xmem_data[17][1] ), .ZN(n27001) );
  AOI22_X1 U30458 ( .A1(n29808), .A2(\xmem_data[18][1] ), .B1(n28516), .B2(
        \xmem_data[19][1] ), .ZN(n27000) );
  AOI22_X1 U30459 ( .A1(n3167), .A2(\xmem_data[20][1] ), .B1(n3188), .B2(
        \xmem_data[21][1] ), .ZN(n26999) );
  AOI22_X1 U30460 ( .A1(n30310), .A2(\xmem_data[22][1] ), .B1(n28147), .B2(
        \xmem_data[23][1] ), .ZN(n26998) );
  NAND4_X1 U30461 ( .A1(n27001), .A2(n27000), .A3(n26999), .A4(n26998), .ZN(
        n27010) );
  AOI22_X1 U30462 ( .A1(n30063), .A2(\xmem_data[24][1] ), .B1(n30765), .B2(
        \xmem_data[25][1] ), .ZN(n27008) );
  AOI22_X1 U30463 ( .A1(n29777), .A2(\xmem_data[28][1] ), .B1(n29776), .B2(
        \xmem_data[29][1] ), .ZN(n27002) );
  INV_X1 U30464 ( .A(n27002), .ZN(n27006) );
  AOI22_X1 U30465 ( .A1(n8075), .A2(\xmem_data[30][1] ), .B1(n21060), .B2(
        \xmem_data[31][1] ), .ZN(n27004) );
  AOI22_X1 U30466 ( .A1(n3226), .A2(\xmem_data[26][1] ), .B1(n3338), .B2(
        \xmem_data[27][1] ), .ZN(n27003) );
  NAND2_X1 U30467 ( .A1(n27004), .A2(n27003), .ZN(n27005) );
  NOR2_X1 U30468 ( .A1(n27006), .A2(n27005), .ZN(n27007) );
  NAND2_X1 U30469 ( .A1(n27008), .A2(n27007), .ZN(n27009) );
  NOR2_X1 U30470 ( .A1(n27010), .A2(n27009), .ZN(n27011) );
  NAND2_X1 U30471 ( .A1(n27012), .A2(n27011), .ZN(n27019) );
  AOI22_X1 U30472 ( .A1(n29829), .A2(\xmem_data[0][1] ), .B1(n29695), .B2(
        \xmem_data[1][1] ), .ZN(n27017) );
  AOI22_X1 U30473 ( .A1(n29696), .A2(\xmem_data[2][1] ), .B1(n3142), .B2(
        \xmem_data[3][1] ), .ZN(n27016) );
  AOI22_X1 U30474 ( .A1(n30291), .A2(\xmem_data[4][1] ), .B1(n29432), .B2(
        \xmem_data[5][1] ), .ZN(n27015) );
  AOI22_X1 U30475 ( .A1(n29423), .A2(\xmem_data[6][1] ), .B1(n29698), .B2(
        \xmem_data[7][1] ), .ZN(n27014) );
  NAND4_X1 U30476 ( .A1(n27017), .A2(n27016), .A3(n27015), .A4(n27014), .ZN(
        n27018) );
  OAI21_X1 U30477 ( .B1(n27019), .B2(n27018), .A(n29733), .ZN(n27101) );
  AOI22_X1 U30478 ( .A1(n30766), .A2(\xmem_data[120][1] ), .B1(n29487), .B2(
        \xmem_data[121][1] ), .ZN(n27026) );
  AOI22_X1 U30479 ( .A1(n29819), .A2(\xmem_data[124][1] ), .B1(n29818), .B2(
        \xmem_data[125][1] ), .ZN(n27020) );
  INV_X1 U30480 ( .A(n27020), .ZN(n27024) );
  AOI22_X1 U30481 ( .A1(n29821), .A2(\xmem_data[126][1] ), .B1(n29820), .B2(
        \xmem_data[127][1] ), .ZN(n27022) );
  AOI22_X1 U30482 ( .A1(n29817), .A2(\xmem_data[122][1] ), .B1(n29816), .B2(
        \xmem_data[123][1] ), .ZN(n27021) );
  NAND2_X1 U30483 ( .A1(n27022), .A2(n27021), .ZN(n27023) );
  NOR2_X1 U30484 ( .A1(n27024), .A2(n27023), .ZN(n27025) );
  NAND2_X1 U30485 ( .A1(n27026), .A2(n27025), .ZN(n27038) );
  AOI22_X1 U30486 ( .A1(n29799), .A2(\xmem_data[104][1] ), .B1(n29708), .B2(
        \xmem_data[105][1] ), .ZN(n27030) );
  AOI22_X1 U30487 ( .A1(n29800), .A2(\xmem_data[106][1] ), .B1(n3375), .B2(
        \xmem_data[107][1] ), .ZN(n27029) );
  AOI22_X1 U30488 ( .A1(n3249), .A2(\xmem_data[108][1] ), .B1(n30730), .B2(
        \xmem_data[109][1] ), .ZN(n27028) );
  AOI22_X1 U30489 ( .A1(n29802), .A2(\xmem_data[110][1] ), .B1(n27763), .B2(
        \xmem_data[111][1] ), .ZN(n27027) );
  NAND4_X1 U30490 ( .A1(n27030), .A2(n27029), .A3(n27028), .A4(n27027), .ZN(
        n27037) );
  AOI22_X1 U30491 ( .A1(n28751), .A2(\xmem_data[112][1] ), .B1(n30634), .B2(
        \xmem_data[113][1] ), .ZN(n27035) );
  AOI22_X1 U30492 ( .A1(n29808), .A2(\xmem_data[114][1] ), .B1(n29807), .B2(
        \xmem_data[115][1] ), .ZN(n27034) );
  AOI22_X1 U30493 ( .A1(n3161), .A2(\xmem_data[116][1] ), .B1(n3188), .B2(
        \xmem_data[117][1] ), .ZN(n27033) );
  NAND4_X1 U30494 ( .A1(n27035), .A2(n27034), .A3(n27033), .A4(n27032), .ZN(
        n27036) );
  OR3_X2 U30495 ( .A1(n27038), .A2(n27037), .A3(n27036), .ZN(n27044) );
  AOI22_X1 U30496 ( .A1(n28717), .A2(\xmem_data[96][1] ), .B1(n29785), .B2(
        \xmem_data[97][1] ), .ZN(n27042) );
  AOI22_X1 U30497 ( .A1(n29830), .A2(\xmem_data[98][1] ), .B1(n20828), .B2(
        \xmem_data[99][1] ), .ZN(n27041) );
  AOI22_X1 U30498 ( .A1(n30291), .A2(\xmem_data[100][1] ), .B1(n26510), .B2(
        \xmem_data[101][1] ), .ZN(n27040) );
  AOI22_X1 U30499 ( .A1(n3392), .A2(\xmem_data[102][1] ), .B1(n29832), .B2(
        \xmem_data[103][1] ), .ZN(n27039) );
  NAND4_X1 U30500 ( .A1(n27042), .A2(n27041), .A3(n27040), .A4(n27039), .ZN(
        n27043) );
  OAI21_X1 U30501 ( .B1(n27044), .B2(n27043), .A(n29837), .ZN(n27100) );
  AOI22_X1 U30502 ( .A1(n29707), .A2(\xmem_data[42][1] ), .B1(n29762), .B2(
        \xmem_data[43][1] ), .ZN(n27048) );
  AOI22_X1 U30503 ( .A1(n29763), .A2(\xmem_data[46][1] ), .B1(n28309), .B2(
        \xmem_data[47][1] ), .ZN(n27047) );
  NAND2_X1 U30504 ( .A1(n3186), .A2(\xmem_data[53][1] ), .ZN(n27046) );
  NAND2_X1 U30505 ( .A1(n3168), .A2(\xmem_data[52][1] ), .ZN(n27045) );
  NAND4_X1 U30506 ( .A1(n27048), .A2(n27047), .A3(n27046), .A4(n27045), .ZN(
        n27052) );
  NAND2_X1 U30507 ( .A1(n27833), .A2(\xmem_data[41][1] ), .ZN(n27050) );
  AOI22_X1 U30508 ( .A1(\xmem_data[49][1] ), .A2(n30249), .B1(n30745), .B2(
        \xmem_data[48][1] ), .ZN(n27049) );
  NAND2_X1 U30509 ( .A1(n27050), .A2(n27049), .ZN(n27051) );
  NOR2_X1 U30510 ( .A1(n27052), .A2(n27051), .ZN(n27069) );
  AND2_X1 U30511 ( .A1(n29482), .A2(\xmem_data[45][1] ), .ZN(n27059) );
  AOI22_X1 U30512 ( .A1(n29771), .A2(\xmem_data[50][1] ), .B1(n17018), .B2(
        \xmem_data[51][1] ), .ZN(n27054) );
  NAND2_X1 U30513 ( .A1(n25678), .A2(\xmem_data[55][1] ), .ZN(n27053) );
  NAND2_X1 U30514 ( .A1(n27054), .A2(n27053), .ZN(n27058) );
  NAND2_X1 U30515 ( .A1(n29610), .A2(\xmem_data[54][1] ), .ZN(n27056) );
  NAND2_X1 U30516 ( .A1(n29390), .A2(\xmem_data[44][1] ), .ZN(n27055) );
  NAND2_X1 U30517 ( .A1(n27056), .A2(n27055), .ZN(n27057) );
  NOR3_X1 U30518 ( .A1(n27059), .A2(n27058), .A3(n27057), .ZN(n27068) );
  AOI22_X1 U30519 ( .A1(n28173), .A2(\xmem_data[56][1] ), .B1(n30266), .B2(
        \xmem_data[57][1] ), .ZN(n27066) );
  AOI22_X1 U30520 ( .A1(n29777), .A2(\xmem_data[60][1] ), .B1(n29776), .B2(
        \xmem_data[61][1] ), .ZN(n27060) );
  INV_X1 U30521 ( .A(n27060), .ZN(n27064) );
  AOI22_X1 U30522 ( .A1(n29726), .A2(\xmem_data[62][1] ), .B1(n21060), .B2(
        \xmem_data[63][1] ), .ZN(n27062) );
  AOI22_X1 U30523 ( .A1(n3226), .A2(\xmem_data[58][1] ), .B1(n23724), .B2(
        \xmem_data[59][1] ), .ZN(n27061) );
  NAND2_X1 U30524 ( .A1(n27062), .A2(n27061), .ZN(n27063) );
  NOR2_X1 U30525 ( .A1(n27064), .A2(n27063), .ZN(n27065) );
  AND2_X1 U30526 ( .A1(n27066), .A2(n27065), .ZN(n27067) );
  NAND4_X1 U30527 ( .A1(n27069), .A2(n4006), .A3(n27068), .A4(n27067), .ZN(
        n27075) );
  AOI22_X1 U30528 ( .A1(n29786), .A2(\xmem_data[32][1] ), .B1(n29785), .B2(
        \xmem_data[33][1] ), .ZN(n27073) );
  AOI22_X1 U30529 ( .A1(n29787), .A2(\xmem_data[34][1] ), .B1(n30907), .B2(
        \xmem_data[35][1] ), .ZN(n27072) );
  AOI22_X1 U30530 ( .A1(n29626), .A2(\xmem_data[36][1] ), .B1(n30707), .B2(
        \xmem_data[37][1] ), .ZN(n27071) );
  AOI22_X1 U30531 ( .A1(n28138), .A2(\xmem_data[38][1] ), .B1(n29789), .B2(
        \xmem_data[39][1] ), .ZN(n27070) );
  NAND4_X1 U30532 ( .A1(n27073), .A2(n27072), .A3(n27071), .A4(n27070), .ZN(
        n27074) );
  OAI21_X1 U30533 ( .B1(n27075), .B2(n27074), .A(n29795), .ZN(n27099) );
  AOI22_X1 U30534 ( .A1(n29628), .A2(\xmem_data[70][1] ), .B1(n29832), .B2(
        \xmem_data[71][1] ), .ZN(n27076) );
  AOI22_X1 U30535 ( .A1(n28717), .A2(\xmem_data[64][1] ), .B1(n29785), .B2(
        \xmem_data[65][1] ), .ZN(n27077) );
  AOI22_X1 U30536 ( .A1(n30633), .A2(\xmem_data[76][1] ), .B1(n28238), .B2(
        \xmem_data[77][1] ), .ZN(n27082) );
  AOI22_X1 U30537 ( .A1(n27754), .A2(\xmem_data[80][1] ), .B1(n27728), .B2(
        \xmem_data[81][1] ), .ZN(n27081) );
  AOI22_X1 U30538 ( .A1(n29830), .A2(\xmem_data[66][1] ), .B1(n3142), .B2(
        \xmem_data[67][1] ), .ZN(n27080) );
  AOI22_X1 U30539 ( .A1(n29802), .A2(\xmem_data[78][1] ), .B1(n28051), .B2(
        \xmem_data[79][1] ), .ZN(n27079) );
  AOI22_X1 U30540 ( .A1(n29800), .A2(\xmem_data[74][1] ), .B1(n29706), .B2(
        \xmem_data[75][1] ), .ZN(n27078) );
  AOI22_X1 U30541 ( .A1(n30766), .A2(\xmem_data[88][1] ), .B1(n29487), .B2(
        \xmem_data[89][1] ), .ZN(n27084) );
  AOI22_X1 U30542 ( .A1(n30062), .A2(\xmem_data[86][1] ), .B1(n28687), .B2(
        \xmem_data[87][1] ), .ZN(n27083) );
  NAND3_X1 U30543 ( .A1(n27076), .A2(n3478), .A3(n27085), .ZN(n27097) );
  AOI22_X1 U30544 ( .A1(n30223), .A2(\xmem_data[68][1] ), .B1(n30775), .B2(
        \xmem_data[69][1] ), .ZN(n27095) );
  AOI22_X1 U30545 ( .A1(n3168), .A2(\xmem_data[84][1] ), .B1(n3191), .B2(
        \xmem_data[85][1] ), .ZN(n27086) );
  AOI22_X1 U30546 ( .A1(n29726), .A2(\xmem_data[94][1] ), .B1(n29725), .B2(
        \xmem_data[95][1] ), .ZN(n27089) );
  AOI22_X1 U30547 ( .A1(n29808), .A2(\xmem_data[82][1] ), .B1(n29807), .B2(
        \xmem_data[83][1] ), .ZN(n27088) );
  AOI22_X1 U30548 ( .A1(n29817), .A2(\xmem_data[90][1] ), .B1(n3151), .B2(
        \xmem_data[91][1] ), .ZN(n27087) );
  AOI22_X1 U30549 ( .A1(n29724), .A2(\xmem_data[92][1] ), .B1(n29723), .B2(
        \xmem_data[93][1] ), .ZN(n27090) );
  INV_X1 U30550 ( .A(n27090), .ZN(n27091) );
  NOR2_X1 U30551 ( .A1(n27092), .A2(n27091), .ZN(n27094) );
  AOI22_X1 U30552 ( .A1(n29799), .A2(\xmem_data[72][1] ), .B1(n29798), .B2(
        \xmem_data[73][1] ), .ZN(n27093) );
  NAND4_X1 U30553 ( .A1(n27095), .A2(n27086), .A3(n27094), .A4(n27093), .ZN(
        n27096) );
  OAI21_X1 U30554 ( .B1(n27097), .B2(n27096), .A(n29758), .ZN(n27098) );
  OAI22_X1 U30555 ( .A1(n32182), .A2(n34923), .B1(n31395), .B2(n34922), .ZN(
        n33636) );
  AOI22_X1 U30556 ( .A1(n28309), .A2(\xmem_data[110][1] ), .B1(n24212), .B2(
        \xmem_data[111][1] ), .ZN(n27112) );
  AOI22_X1 U30557 ( .A1(n25632), .A2(\xmem_data[120][1] ), .B1(n28291), .B2(
        \xmem_data[121][1] ), .ZN(n27106) );
  AOI22_X1 U30558 ( .A1(n3302), .A2(\xmem_data[122][1] ), .B1(n24570), .B2(
        \xmem_data[123][1] ), .ZN(n27105) );
  AOI22_X1 U30559 ( .A1(n28293), .A2(\xmem_data[124][1] ), .B1(n28292), .B2(
        \xmem_data[125][1] ), .ZN(n27104) );
  AND2_X1 U30560 ( .A1(n24686), .A2(\xmem_data[127][1] ), .ZN(n27102) );
  AOI21_X1 U30561 ( .B1(n28192), .B2(\xmem_data[126][1] ), .A(n27102), .ZN(
        n27103) );
  NAND4_X1 U30562 ( .A1(n27106), .A2(n27105), .A3(n27104), .A4(n27103), .ZN(
        n27110) );
  AOI22_X1 U30563 ( .A1(n24565), .A2(\xmem_data[104][1] ), .B1(n24564), .B2(
        \xmem_data[105][1] ), .ZN(n27108) );
  AOI22_X1 U30564 ( .A1(n24450), .A2(\xmem_data[108][1] ), .B1(n13475), .B2(
        \xmem_data[109][1] ), .ZN(n27107) );
  NAND2_X1 U30565 ( .A1(n27108), .A2(n27107), .ZN(n27109) );
  NOR2_X1 U30566 ( .A1(n27110), .A2(n27109), .ZN(n27111) );
  NAND2_X1 U30567 ( .A1(n27112), .A2(n27111), .ZN(n27118) );
  AOI22_X1 U30568 ( .A1(n24688), .A2(\xmem_data[96][1] ), .B1(n28317), .B2(
        \xmem_data[97][1] ), .ZN(n27116) );
  AOI22_X1 U30569 ( .A1(n3424), .A2(\xmem_data[98][1] ), .B1(n31347), .B2(
        \xmem_data[99][1] ), .ZN(n27115) );
  AOI22_X1 U30570 ( .A1(n28318), .A2(\xmem_data[100][1] ), .B1(n3219), .B2(
        \xmem_data[101][1] ), .ZN(n27114) );
  AOI22_X1 U30571 ( .A1(n25414), .A2(\xmem_data[102][1] ), .B1(n28319), .B2(
        \xmem_data[103][1] ), .ZN(n27113) );
  NAND4_X1 U30572 ( .A1(n27116), .A2(n27115), .A3(n27114), .A4(n27113), .ZN(
        n27117) );
  AOI22_X1 U30573 ( .A1(n28298), .A2(\xmem_data[112][1] ), .B1(n25606), .B2(
        \xmem_data[113][1] ), .ZN(n27122) );
  AOI22_X1 U30574 ( .A1(n29437), .A2(\xmem_data[114][1] ), .B1(n28299), .B2(
        \xmem_data[115][1] ), .ZN(n27121) );
  AOI22_X1 U30575 ( .A1(n21007), .A2(\xmem_data[116][1] ), .B1(n17043), .B2(
        \xmem_data[117][1] ), .ZN(n27120) );
  AOI22_X1 U30576 ( .A1(n28302), .A2(\xmem_data[118][1] ), .B1(n28301), .B2(
        \xmem_data[119][1] ), .ZN(n27119) );
  NAND4_X1 U30577 ( .A1(n27122), .A2(n27121), .A3(n27120), .A4(n27119), .ZN(
        n27125) );
  AOI22_X1 U30578 ( .A1(n28308), .A2(\xmem_data[106][1] ), .B1(n28307), .B2(
        \xmem_data[107][1] ), .ZN(n27123) );
  INV_X1 U30579 ( .A(n27123), .ZN(n27124) );
  NOR2_X1 U30580 ( .A1(n27125), .A2(n27124), .ZN(n27127) );
  INV_X1 U30581 ( .A(n28288), .ZN(n27126) );
  AOI21_X1 U30582 ( .B1(n27128), .B2(n27127), .A(n27126), .ZN(n27155) );
  AOI22_X1 U30583 ( .A1(n28344), .A2(\xmem_data[42][1] ), .B1(n3231), .B2(
        \xmem_data[43][1] ), .ZN(n27153) );
  AOI22_X1 U30584 ( .A1(n28346), .A2(\xmem_data[46][1] ), .B1(n28345), .B2(
        \xmem_data[47][1] ), .ZN(n27138) );
  AOI22_X1 U30585 ( .A1(n21010), .A2(\xmem_data[56][1] ), .B1(n25581), .B2(
        \xmem_data[57][1] ), .ZN(n27132) );
  AOI22_X1 U30586 ( .A1(n23780), .A2(\xmem_data[58][1] ), .B1(n23723), .B2(
        \xmem_data[59][1] ), .ZN(n27131) );
  AOI22_X1 U30587 ( .A1(n3179), .A2(\xmem_data[60][1] ), .B1(n28328), .B2(
        \xmem_data[61][1] ), .ZN(n27130) );
  AOI22_X1 U30588 ( .A1(n28467), .A2(\xmem_data[62][1] ), .B1(n28329), .B2(
        \xmem_data[63][1] ), .ZN(n27129) );
  NAND4_X1 U30589 ( .A1(n27132), .A2(n27131), .A3(n27130), .A4(n27129), .ZN(
        n27136) );
  AOI22_X1 U30590 ( .A1(n25617), .A2(\xmem_data[40][1] ), .B1(n28342), .B2(
        \xmem_data[41][1] ), .ZN(n27134) );
  AOI22_X1 U30591 ( .A1(n22712), .A2(\xmem_data[44][1] ), .B1(n20982), .B2(
        \xmem_data[45][1] ), .ZN(n27133) );
  NAND2_X1 U30592 ( .A1(n27134), .A2(n27133), .ZN(n27135) );
  NOR2_X1 U30593 ( .A1(n27136), .A2(n27135), .ZN(n27137) );
  NAND2_X1 U30594 ( .A1(n27138), .A2(n27137), .ZN(n27150) );
  AOI22_X1 U30595 ( .A1(n28354), .A2(\xmem_data[32][1] ), .B1(n25629), .B2(
        \xmem_data[33][1] ), .ZN(n27142) );
  AOI22_X1 U30596 ( .A1(n3229), .A2(\xmem_data[34][1] ), .B1(n31347), .B2(
        \xmem_data[35][1] ), .ZN(n27141) );
  AOI22_X1 U30597 ( .A1(n28355), .A2(\xmem_data[36][1] ), .B1(n3218), .B2(
        \xmem_data[37][1] ), .ZN(n27140) );
  AOI22_X1 U30598 ( .A1(n29026), .A2(\xmem_data[38][1] ), .B1(n28356), .B2(
        \xmem_data[39][1] ), .ZN(n27139) );
  NAND4_X1 U30599 ( .A1(n27142), .A2(n27141), .A3(n27140), .A4(n27139), .ZN(
        n27148) );
  AOI22_X1 U30600 ( .A1(n28334), .A2(\xmem_data[48][1] ), .B1(n29009), .B2(
        \xmem_data[49][1] ), .ZN(n27146) );
  AOI22_X1 U30601 ( .A1(n28336), .A2(\xmem_data[50][1] ), .B1(n28335), .B2(
        \xmem_data[51][1] ), .ZN(n27145) );
  AOI22_X1 U30602 ( .A1(n28337), .A2(\xmem_data[52][1] ), .B1(n14912), .B2(
        \xmem_data[53][1] ), .ZN(n27144) );
  AOI22_X1 U30603 ( .A1(n29239), .A2(\xmem_data[54][1] ), .B1(n13481), .B2(
        \xmem_data[55][1] ), .ZN(n27143) );
  NAND4_X1 U30604 ( .A1(n27146), .A2(n27145), .A3(n27144), .A4(n27143), .ZN(
        n27147) );
  NOR2_X1 U30605 ( .A1(n27150), .A2(n27149), .ZN(n27152) );
  INV_X1 U30606 ( .A(n28361), .ZN(n27151) );
  AOI21_X1 U30607 ( .B1(n27153), .B2(n27152), .A(n27151), .ZN(n27154) );
  NOR2_X1 U30608 ( .A1(n27155), .A2(n27154), .ZN(n27212) );
  AOI22_X1 U30609 ( .A1(n28309), .A2(\xmem_data[78][1] ), .B1(n24639), .B2(
        \xmem_data[79][1] ), .ZN(n27166) );
  AOI22_X1 U30610 ( .A1(n30557), .A2(\xmem_data[88][1] ), .B1(n28291), .B2(
        \xmem_data[89][1] ), .ZN(n27160) );
  AOI22_X1 U30611 ( .A1(n3301), .A2(\xmem_data[90][1] ), .B1(n29245), .B2(
        \xmem_data[91][1] ), .ZN(n27159) );
  AOI22_X1 U30612 ( .A1(n28293), .A2(\xmem_data[92][1] ), .B1(n28292), .B2(
        \xmem_data[93][1] ), .ZN(n27158) );
  AND2_X1 U30613 ( .A1(n30498), .A2(\xmem_data[95][1] ), .ZN(n27156) );
  AOI21_X1 U30614 ( .B1(n30754), .B2(\xmem_data[94][1] ), .A(n27156), .ZN(
        n27157) );
  NAND4_X1 U30615 ( .A1(n27160), .A2(n27159), .A3(n27158), .A4(n27157), .ZN(
        n27164) );
  AOI22_X1 U30616 ( .A1(n22758), .A2(\xmem_data[72][1] ), .B1(n24633), .B2(
        \xmem_data[73][1] ), .ZN(n27162) );
  AOI22_X1 U30617 ( .A1(n30885), .A2(\xmem_data[76][1] ), .B1(n20982), .B2(
        \xmem_data[77][1] ), .ZN(n27161) );
  NAND2_X1 U30618 ( .A1(n27162), .A2(n27161), .ZN(n27163) );
  NOR2_X1 U30619 ( .A1(n27164), .A2(n27163), .ZN(n27165) );
  NAND2_X1 U30620 ( .A1(n27166), .A2(n27165), .ZN(n27172) );
  AOI22_X1 U30621 ( .A1(n21061), .A2(\xmem_data[64][1] ), .B1(n28317), .B2(
        \xmem_data[65][1] ), .ZN(n27170) );
  AOI22_X1 U30622 ( .A1(n3245), .A2(\xmem_data[66][1] ), .B1(n25442), .B2(
        \xmem_data[67][1] ), .ZN(n27169) );
  AOI22_X1 U30623 ( .A1(n28318), .A2(\xmem_data[68][1] ), .B1(n3218), .B2(
        \xmem_data[69][1] ), .ZN(n27168) );
  AOI22_X1 U30624 ( .A1(n28733), .A2(\xmem_data[70][1] ), .B1(n28319), .B2(
        \xmem_data[71][1] ), .ZN(n27167) );
  NAND4_X1 U30625 ( .A1(n27170), .A2(n27169), .A3(n27168), .A4(n27167), .ZN(
        n27171) );
  AOI22_X1 U30626 ( .A1(n28298), .A2(\xmem_data[80][1] ), .B1(n20584), .B2(
        \xmem_data[81][1] ), .ZN(n27176) );
  AOI22_X1 U30627 ( .A1(n28752), .A2(\xmem_data[82][1] ), .B1(n28299), .B2(
        \xmem_data[83][1] ), .ZN(n27175) );
  AOI22_X1 U30628 ( .A1(n20800), .A2(\xmem_data[84][1] ), .B1(n29048), .B2(
        \xmem_data[85][1] ), .ZN(n27174) );
  AOI22_X1 U30629 ( .A1(n28302), .A2(\xmem_data[86][1] ), .B1(n28301), .B2(
        \xmem_data[87][1] ), .ZN(n27173) );
  NAND4_X1 U30630 ( .A1(n27176), .A2(n27175), .A3(n27174), .A4(n27173), .ZN(
        n27179) );
  AOI22_X1 U30631 ( .A1(n28308), .A2(\xmem_data[74][1] ), .B1(n28307), .B2(
        \xmem_data[75][1] ), .ZN(n27177) );
  INV_X1 U30632 ( .A(n27177), .ZN(n27178) );
  NOR2_X1 U30633 ( .A1(n27179), .A2(n27178), .ZN(n27181) );
  INV_X1 U30634 ( .A(n28324), .ZN(n27180) );
  AOI21_X1 U30635 ( .B1(n27182), .B2(n27181), .A(n27180), .ZN(n27210) );
  AOI22_X1 U30636 ( .A1(n30698), .A2(\xmem_data[10][1] ), .B1(n28007), .B2(
        \xmem_data[11][1] ), .ZN(n27208) );
  AOI22_X1 U30637 ( .A1(n30663), .A2(\xmem_data[14][1] ), .B1(n28375), .B2(
        \xmem_data[15][1] ), .ZN(n27193) );
  AOI22_X1 U30638 ( .A1(n28374), .A2(\xmem_data[12][1] ), .B1(n3357), .B2(
        \xmem_data[13][1] ), .ZN(n27184) );
  AOI22_X1 U30639 ( .A1(n30883), .A2(\xmem_data[8][1] ), .B1(n28372), .B2(
        \xmem_data[9][1] ), .ZN(n27183) );
  NAND2_X1 U30640 ( .A1(n27184), .A2(n27183), .ZN(n27191) );
  AOI22_X1 U30641 ( .A1(n30674), .A2(\xmem_data[30][1] ), .B1(n21059), .B2(
        \xmem_data[31][1] ), .ZN(n27185) );
  INV_X1 U30642 ( .A(n27185), .ZN(n27190) );
  AOI22_X1 U30643 ( .A1(n28385), .A2(\xmem_data[24][1] ), .B1(n25716), .B2(
        \xmem_data[25][1] ), .ZN(n27188) );
  AOI22_X1 U30644 ( .A1(n30497), .A2(\xmem_data[28][1] ), .B1(n25723), .B2(
        \xmem_data[29][1] ), .ZN(n27187) );
  AOI22_X1 U30645 ( .A1(n30645), .A2(\xmem_data[26][1] ), .B1(n27975), .B2(
        \xmem_data[27][1] ), .ZN(n27186) );
  NOR3_X1 U30646 ( .A1(n27191), .A2(n27190), .A3(n27189), .ZN(n27192) );
  NAND2_X1 U30647 ( .A1(n27193), .A2(n27192), .ZN(n27205) );
  AOI22_X1 U30648 ( .A1(n30862), .A2(\xmem_data[0][1] ), .B1(n28366), .B2(
        \xmem_data[1][1] ), .ZN(n27197) );
  AOI22_X1 U30649 ( .A1(n3306), .A2(\xmem_data[2][1] ), .B1(n14875), .B2(
        \xmem_data[3][1] ), .ZN(n27196) );
  AOI22_X1 U30650 ( .A1(n28364), .A2(\xmem_data[4][1] ), .B1(n3222), .B2(
        \xmem_data[5][1] ), .ZN(n27195) );
  AOI22_X1 U30651 ( .A1(n28367), .A2(\xmem_data[6][1] ), .B1(n25562), .B2(
        \xmem_data[7][1] ), .ZN(n27194) );
  NAND4_X1 U30652 ( .A1(n27197), .A2(n27196), .A3(n27195), .A4(n27194), .ZN(
        n27203) );
  AOI22_X1 U30653 ( .A1(n17041), .A2(\xmem_data[16][1] ), .B1(n14898), .B2(
        \xmem_data[17][1] ), .ZN(n27201) );
  AOI22_X1 U30654 ( .A1(n3465), .A2(\xmem_data[18][1] ), .B1(n22677), .B2(
        \xmem_data[19][1] ), .ZN(n27200) );
  AOI22_X1 U30655 ( .A1(n24133), .A2(\xmem_data[20][1] ), .B1(n28492), .B2(
        \xmem_data[21][1] ), .ZN(n27199) );
  AOI22_X1 U30656 ( .A1(n29439), .A2(\xmem_data[22][1] ), .B1(n28380), .B2(
        \xmem_data[23][1] ), .ZN(n27198) );
  NAND4_X1 U30657 ( .A1(n27201), .A2(n27200), .A3(n27199), .A4(n27198), .ZN(
        n27202) );
  INV_X1 U30658 ( .A(n28395), .ZN(n27206) );
  AOI21_X1 U30659 ( .B1(n27208), .B2(n27207), .A(n27206), .ZN(n27209) );
  NOR2_X1 U30660 ( .A1(n27210), .A2(n27209), .ZN(n27211) );
  XNOR2_X1 U30661 ( .A(n32940), .B(\fmem_data[18][5] ), .ZN(n31165) );
  AOI22_X1 U30662 ( .A1(n28318), .A2(\xmem_data[100][2] ), .B1(n3221), .B2(
        \xmem_data[101][2] ), .ZN(n27216) );
  AOI22_X1 U30663 ( .A1(n3245), .A2(\xmem_data[98][2] ), .B1(n24439), .B2(
        \xmem_data[99][2] ), .ZN(n27215) );
  AOI22_X1 U30664 ( .A1(n25408), .A2(\xmem_data[96][2] ), .B1(n28317), .B2(
        \xmem_data[97][2] ), .ZN(n27214) );
  AOI22_X1 U30665 ( .A1(n25448), .A2(\xmem_data[102][2] ), .B1(n28319), .B2(
        \xmem_data[103][2] ), .ZN(n27213) );
  NAND4_X1 U30666 ( .A1(n27216), .A2(n27215), .A3(n27214), .A4(n27213), .ZN(
        n27233) );
  AOI22_X1 U30667 ( .A1(n28493), .A2(\xmem_data[120][2] ), .B1(n28291), .B2(
        \xmem_data[121][2] ), .ZN(n27220) );
  AOI22_X1 U30668 ( .A1(n3271), .A2(\xmem_data[122][2] ), .B1(n28098), .B2(
        \xmem_data[123][2] ), .ZN(n27219) );
  AOI22_X1 U30669 ( .A1(n28293), .A2(\xmem_data[124][2] ), .B1(n28292), .B2(
        \xmem_data[125][2] ), .ZN(n27218) );
  AOI22_X1 U30670 ( .A1(n28772), .A2(\xmem_data[126][2] ), .B1(n20579), .B2(
        \xmem_data[127][2] ), .ZN(n27217) );
  NAND4_X1 U30671 ( .A1(n27220), .A2(n27219), .A3(n27218), .A4(n27217), .ZN(
        n27231) );
  AOI22_X1 U30672 ( .A1(n28298), .A2(\xmem_data[112][2] ), .B1(n27536), .B2(
        \xmem_data[113][2] ), .ZN(n27224) );
  AOI22_X1 U30673 ( .A1(n30303), .A2(\xmem_data[114][2] ), .B1(n28299), .B2(
        \xmem_data[115][2] ), .ZN(n27223) );
  AOI22_X1 U30674 ( .A1(n21007), .A2(\xmem_data[116][2] ), .B1(n25398), .B2(
        \xmem_data[117][2] ), .ZN(n27222) );
  AOI22_X1 U30675 ( .A1(n28302), .A2(\xmem_data[118][2] ), .B1(n28301), .B2(
        \xmem_data[119][2] ), .ZN(n27221) );
  NAND4_X1 U30676 ( .A1(n27224), .A2(n27223), .A3(n27222), .A4(n27221), .ZN(
        n27230) );
  AOI22_X1 U30677 ( .A1(n23812), .A2(\xmem_data[104][2] ), .B1(n28372), .B2(
        \xmem_data[105][2] ), .ZN(n27228) );
  AOI22_X1 U30678 ( .A1(n28308), .A2(\xmem_data[106][2] ), .B1(n28307), .B2(
        \xmem_data[107][2] ), .ZN(n27227) );
  AOI22_X1 U30679 ( .A1(n25422), .A2(\xmem_data[108][2] ), .B1(n28373), .B2(
        \xmem_data[109][2] ), .ZN(n27226) );
  AOI22_X1 U30680 ( .A1(n28309), .A2(\xmem_data[110][2] ), .B1(n25423), .B2(
        \xmem_data[111][2] ), .ZN(n27225) );
  NAND4_X1 U30681 ( .A1(n27228), .A2(n27227), .A3(n27226), .A4(n27225), .ZN(
        n27229) );
  OR3_X1 U30682 ( .A1(n27231), .A2(n27230), .A3(n27229), .ZN(n27232) );
  OAI21_X1 U30683 ( .B1(n27233), .B2(n27232), .A(n28288), .ZN(n27303) );
  AOI22_X1 U30684 ( .A1(n28354), .A2(\xmem_data[32][2] ), .B1(n27499), .B2(
        \xmem_data[33][2] ), .ZN(n27237) );
  AOI22_X1 U30685 ( .A1(n3424), .A2(\xmem_data[34][2] ), .B1(n28501), .B2(
        \xmem_data[35][2] ), .ZN(n27236) );
  AOI22_X1 U30686 ( .A1(n28355), .A2(\xmem_data[36][2] ), .B1(n3220), .B2(
        \xmem_data[37][2] ), .ZN(n27235) );
  AOI22_X1 U30687 ( .A1(n29065), .A2(\xmem_data[38][2] ), .B1(n28356), .B2(
        \xmem_data[39][2] ), .ZN(n27234) );
  NAND4_X1 U30688 ( .A1(n27237), .A2(n27236), .A3(n27235), .A4(n27234), .ZN(
        n27254) );
  AOI22_X1 U30689 ( .A1(n24647), .A2(\xmem_data[56][2] ), .B1(n21009), .B2(
        \xmem_data[57][2] ), .ZN(n27241) );
  AOI22_X1 U30690 ( .A1(n3271), .A2(\xmem_data[58][2] ), .B1(n20507), .B2(
        \xmem_data[59][2] ), .ZN(n27240) );
  AOI22_X1 U30691 ( .A1(n3179), .A2(\xmem_data[60][2] ), .B1(n28328), .B2(
        \xmem_data[61][2] ), .ZN(n27239) );
  AOI22_X1 U30692 ( .A1(n30901), .A2(\xmem_data[62][2] ), .B1(n28329), .B2(
        \xmem_data[63][2] ), .ZN(n27238) );
  NAND4_X1 U30693 ( .A1(n27241), .A2(n27240), .A3(n27239), .A4(n27238), .ZN(
        n27252) );
  AOI22_X1 U30694 ( .A1(n28334), .A2(\xmem_data[48][2] ), .B1(n30541), .B2(
        \xmem_data[49][2] ), .ZN(n27245) );
  AOI22_X1 U30695 ( .A1(n28336), .A2(\xmem_data[50][2] ), .B1(n28335), .B2(
        \xmem_data[51][2] ), .ZN(n27244) );
  AOI22_X1 U30696 ( .A1(n28337), .A2(\xmem_data[52][2] ), .B1(n25398), .B2(
        \xmem_data[53][2] ), .ZN(n27243) );
  AOI22_X1 U30697 ( .A1(n21050), .A2(\xmem_data[54][2] ), .B1(n30871), .B2(
        \xmem_data[55][2] ), .ZN(n27242) );
  NAND4_X1 U30698 ( .A1(n27245), .A2(n27244), .A3(n27243), .A4(n27242), .ZN(
        n27251) );
  AOI22_X1 U30699 ( .A1(n30883), .A2(\xmem_data[40][2] ), .B1(n28342), .B2(
        \xmem_data[41][2] ), .ZN(n27249) );
  AOI22_X1 U30700 ( .A1(n28344), .A2(\xmem_data[42][2] ), .B1(n27547), .B2(
        \xmem_data[43][2] ), .ZN(n27248) );
  AOI22_X1 U30701 ( .A1(n25422), .A2(\xmem_data[44][2] ), .B1(n14996), .B2(
        \xmem_data[45][2] ), .ZN(n27247) );
  AOI22_X1 U30702 ( .A1(n28346), .A2(\xmem_data[46][2] ), .B1(n28345), .B2(
        \xmem_data[47][2] ), .ZN(n27246) );
  NAND4_X1 U30703 ( .A1(n27249), .A2(n27248), .A3(n27247), .A4(n27246), .ZN(
        n27250) );
  OR3_X1 U30704 ( .A1(n27252), .A2(n27251), .A3(n27250), .ZN(n27253) );
  OAI21_X1 U30705 ( .B1(n27254), .B2(n27253), .A(n28361), .ZN(n27302) );
  AOI22_X1 U30706 ( .A1(n28076), .A2(\xmem_data[0][2] ), .B1(n28366), .B2(
        \xmem_data[1][2] ), .ZN(n27258) );
  AOI22_X1 U30707 ( .A1(n3306), .A2(\xmem_data[2][2] ), .B1(n28501), .B2(
        \xmem_data[3][2] ), .ZN(n27257) );
  AOI22_X1 U30708 ( .A1(n28364), .A2(\xmem_data[4][2] ), .B1(n3218), .B2(
        \xmem_data[5][2] ), .ZN(n27256) );
  AOI22_X1 U30709 ( .A1(n28367), .A2(\xmem_data[6][2] ), .B1(n28508), .B2(
        \xmem_data[7][2] ), .ZN(n27255) );
  NAND4_X1 U30710 ( .A1(n27258), .A2(n27257), .A3(n27256), .A4(n27255), .ZN(
        n27275) );
  AOI22_X1 U30711 ( .A1(n24697), .A2(\xmem_data[8][2] ), .B1(n28372), .B2(
        \xmem_data[9][2] ), .ZN(n27262) );
  AOI22_X1 U30712 ( .A1(n29231), .A2(\xmem_data[10][2] ), .B1(n28343), .B2(
        \xmem_data[11][2] ), .ZN(n27261) );
  AOI22_X1 U30713 ( .A1(n28374), .A2(\xmem_data[12][2] ), .B1(n3358), .B2(
        \xmem_data[13][2] ), .ZN(n27260) );
  AOI22_X1 U30714 ( .A1(n28309), .A2(\xmem_data[14][2] ), .B1(n28375), .B2(
        \xmem_data[15][2] ), .ZN(n27259) );
  NAND4_X1 U30715 ( .A1(n27262), .A2(n27261), .A3(n27260), .A4(n27259), .ZN(
        n27274) );
  AOI22_X1 U30716 ( .A1(n28980), .A2(\xmem_data[16][2] ), .B1(n23715), .B2(
        \xmem_data[17][2] ), .ZN(n27266) );
  AOI22_X1 U30717 ( .A1(n28336), .A2(\xmem_data[18][2] ), .B1(n3212), .B2(
        \xmem_data[19][2] ), .ZN(n27265) );
  AOI22_X1 U30718 ( .A1(n25573), .A2(\xmem_data[20][2] ), .B1(n30544), .B2(
        \xmem_data[21][2] ), .ZN(n27264) );
  AOI22_X1 U30719 ( .A1(n21008), .A2(\xmem_data[22][2] ), .B1(n28380), .B2(
        \xmem_data[23][2] ), .ZN(n27263) );
  NAND4_X1 U30720 ( .A1(n27266), .A2(n27265), .A3(n27264), .A4(n27263), .ZN(
        n27273) );
  AOI22_X1 U30721 ( .A1(n28385), .A2(\xmem_data[24][2] ), .B1(n30598), .B2(
        \xmem_data[25][2] ), .ZN(n27271) );
  AOI22_X1 U30722 ( .A1(n28202), .A2(\xmem_data[26][2] ), .B1(n23723), .B2(
        \xmem_data[27][2] ), .ZN(n27270) );
  AOI22_X1 U30723 ( .A1(n3209), .A2(\xmem_data[28][2] ), .B1(n25527), .B2(
        \xmem_data[29][2] ), .ZN(n27269) );
  AND2_X1 U30724 ( .A1(n13487), .A2(\xmem_data[31][2] ), .ZN(n27267) );
  AOI21_X1 U30725 ( .B1(n23753), .B2(\xmem_data[30][2] ), .A(n27267), .ZN(
        n27268) );
  NAND4_X1 U30726 ( .A1(n27271), .A2(n27270), .A3(n27269), .A4(n27268), .ZN(
        n27272) );
  OR4_X1 U30727 ( .A1(n27275), .A2(n27274), .A3(n27273), .A4(n27272), .ZN(
        n27276) );
  NAND2_X1 U30728 ( .A1(n27276), .A2(n28395), .ZN(n27301) );
  AND2_X1 U30729 ( .A1(n3221), .A2(\xmem_data[69][2] ), .ZN(n27277) );
  AOI21_X1 U30730 ( .B1(n28318), .B2(\xmem_data[68][2] ), .A(n27277), .ZN(
        n27282) );
  AOI22_X1 U30731 ( .A1(n3245), .A2(\xmem_data[66][2] ), .B1(n23731), .B2(
        \xmem_data[67][2] ), .ZN(n27281) );
  AND2_X1 U30732 ( .A1(n27436), .A2(\xmem_data[64][2] ), .ZN(n27278) );
  AOI21_X1 U30733 ( .B1(n28317), .B2(\xmem_data[65][2] ), .A(n27278), .ZN(
        n27280) );
  AOI22_X1 U30734 ( .A1(n17033), .A2(\xmem_data[70][2] ), .B1(n28319), .B2(
        \xmem_data[71][2] ), .ZN(n27279) );
  NAND4_X1 U30735 ( .A1(n27282), .A2(n27281), .A3(n27280), .A4(n27279), .ZN(
        n27299) );
  AOI22_X1 U30736 ( .A1(n3178), .A2(\xmem_data[88][2] ), .B1(n28291), .B2(
        \xmem_data[89][2] ), .ZN(n27286) );
  AOI22_X1 U30737 ( .A1(n3307), .A2(\xmem_data[90][2] ), .B1(n24622), .B2(
        \xmem_data[91][2] ), .ZN(n27285) );
  AOI22_X1 U30738 ( .A1(n28293), .A2(\xmem_data[92][2] ), .B1(n28292), .B2(
        \xmem_data[93][2] ), .ZN(n27284) );
  AOI22_X1 U30739 ( .A1(n28467), .A2(\xmem_data[94][2] ), .B1(n20579), .B2(
        \xmem_data[95][2] ), .ZN(n27283) );
  NAND4_X1 U30740 ( .A1(n27286), .A2(n27285), .A3(n27284), .A4(n27283), .ZN(
        n27297) );
  AOI22_X1 U30741 ( .A1(n28298), .A2(\xmem_data[80][2] ), .B1(n22741), .B2(
        \xmem_data[81][2] ), .ZN(n27290) );
  AOI22_X1 U30742 ( .A1(n30303), .A2(\xmem_data[82][2] ), .B1(n28299), .B2(
        \xmem_data[83][2] ), .ZN(n27289) );
  AOI22_X1 U30743 ( .A1(n24509), .A2(\xmem_data[84][2] ), .B1(n25398), .B2(
        \xmem_data[85][2] ), .ZN(n27288) );
  AOI22_X1 U30744 ( .A1(n28302), .A2(\xmem_data[86][2] ), .B1(n28301), .B2(
        \xmem_data[87][2] ), .ZN(n27287) );
  NAND4_X1 U30745 ( .A1(n27290), .A2(n27289), .A3(n27288), .A4(n27287), .ZN(
        n27296) );
  AOI22_X1 U30746 ( .A1(n24141), .A2(\xmem_data[72][2] ), .B1(n3255), .B2(
        \xmem_data[73][2] ), .ZN(n27294) );
  AOI22_X1 U30747 ( .A1(n28308), .A2(\xmem_data[74][2] ), .B1(n28307), .B2(
        \xmem_data[75][2] ), .ZN(n27293) );
  AOI22_X1 U30748 ( .A1(n30607), .A2(\xmem_data[76][2] ), .B1(n30854), .B2(
        \xmem_data[77][2] ), .ZN(n27292) );
  AOI22_X1 U30749 ( .A1(n28309), .A2(\xmem_data[78][2] ), .B1(n20958), .B2(
        \xmem_data[79][2] ), .ZN(n27291) );
  NAND4_X1 U30750 ( .A1(n27294), .A2(n27293), .A3(n27292), .A4(n27291), .ZN(
        n27295) );
  OR3_X1 U30751 ( .A1(n27297), .A2(n27296), .A3(n27295), .ZN(n27298) );
  OAI21_X1 U30752 ( .B1(n27299), .B2(n27298), .A(n28324), .ZN(n27300) );
  XNOR2_X1 U30753 ( .A(n32596), .B(\fmem_data[18][5] ), .ZN(n27326) );
  OAI21_X1 U30754 ( .B1(n27309), .B2(n27310), .A(n27311), .ZN(n27307) );
  NAND2_X1 U30755 ( .A1(n27309), .A2(n27310), .ZN(n27306) );
  NAND2_X1 U30756 ( .A1(n27307), .A2(n27306), .ZN(n31772) );
  XNOR2_X1 U30757 ( .A(n27308), .B(n31772), .ZN(n35439) );
  XNOR2_X1 U30758 ( .A(n27310), .B(n27309), .ZN(n27312) );
  XNOR2_X1 U30759 ( .A(n27312), .B(n27311), .ZN(n31425) );
  FA_X1 U30760 ( .A(n27315), .B(n27314), .CI(n27313), .CO(n35215), .S(n31424)
         );
  XNOR2_X1 U30761 ( .A(n27317), .B(n27316), .ZN(n27319) );
  XNOR2_X1 U30762 ( .A(n27319), .B(n27318), .ZN(n34288) );
  FA_X1 U30763 ( .A(n27322), .B(n27321), .CI(n27320), .CO(n30136), .S(n30151)
         );
  XNOR2_X1 U30764 ( .A(n32440), .B(\fmem_data[7][5] ), .ZN(n32107) );
  XOR2_X1 U30765 ( .A(\fmem_data[7][4] ), .B(\fmem_data[7][5] ), .Z(n27323) );
  XNOR2_X1 U30766 ( .A(n32174), .B(\fmem_data[7][5] ), .ZN(n34232) );
  XNOR2_X1 U30767 ( .A(n35108), .B(\fmem_data[18][1] ), .ZN(n33265) );
  XNOR2_X1 U30768 ( .A(n31672), .B(\fmem_data[18][1] ), .ZN(n32146) );
  OAI22_X1 U30769 ( .A1(n33265), .A2(n3580), .B1(n32146), .B2(n36104), .ZN(
        n30798) );
  OAI22_X1 U30770 ( .A1(n27327), .A2(n35006), .B1(n27326), .B2(n35007), .ZN(
        n30796) );
  NAND2_X1 U30771 ( .A1(n27329), .A2(n27328), .ZN(n32444) );
  XNOR2_X1 U30772 ( .A(n32444), .B(\fmem_data[27][5] ), .ZN(n32308) );
  XNOR2_X1 U30773 ( .A(n3278), .B(\fmem_data[27][5] ), .ZN(n33167) );
  OAI22_X1 U30774 ( .A1(n32308), .A2(n34904), .B1(n33167), .B2(n34903), .ZN(
        n30801) );
  OAI22_X1 U30775 ( .A1(n32154), .A2(n34918), .B1(n27333), .B2(n34919), .ZN(
        n29691) );
  AOI22_X1 U30776 ( .A1(n25382), .A2(\xmem_data[24][0] ), .B1(n3464), .B2(
        \xmem_data[25][0] ), .ZN(n27337) );
  AOI22_X1 U30777 ( .A1(n29162), .A2(\xmem_data[26][0] ), .B1(n29317), .B2(
        \xmem_data[27][0] ), .ZN(n27336) );
  AOI22_X1 U30778 ( .A1(n31270), .A2(\xmem_data[28][0] ), .B1(n17044), .B2(
        \xmem_data[29][0] ), .ZN(n27335) );
  AOI22_X1 U30779 ( .A1(n30871), .A2(\xmem_data[30][0] ), .B1(n3178), .B2(
        \xmem_data[31][0] ), .ZN(n27334) );
  AOI22_X1 U30780 ( .A1(n30552), .A2(\xmem_data[22][0] ), .B1(n29023), .B2(
        \xmem_data[23][0] ), .ZN(n27345) );
  NAND2_X1 U30781 ( .A1(n25708), .A2(\xmem_data[21][0] ), .ZN(n27339) );
  NAND2_X1 U30782 ( .A1(n29157), .A2(\xmem_data[17][0] ), .ZN(n27338) );
  NAND2_X1 U30783 ( .A1(n27341), .A2(n27340), .ZN(n27342) );
  NOR2_X1 U30784 ( .A1(n27342), .A2(n3908), .ZN(n27344) );
  AOI22_X1 U30785 ( .A1(n25492), .A2(\xmem_data[18][0] ), .B1(n24638), .B2(
        \xmem_data[19][0] ), .ZN(n27343) );
  NAND4_X1 U30786 ( .A1(n3844), .A2(n27345), .A3(n27344), .A4(n27343), .ZN(
        n27359) );
  NAND2_X1 U30787 ( .A1(n29254), .A2(\xmem_data[11][0] ), .ZN(n27351) );
  AOI22_X1 U30788 ( .A1(n29118), .A2(\xmem_data[8][0] ), .B1(n3348), .B2(
        \xmem_data[9][0] ), .ZN(n27350) );
  AOI22_X1 U30789 ( .A1(n3218), .A2(\xmem_data[12][0] ), .B1(n25612), .B2(
        \xmem_data[13][0] ), .ZN(n27347) );
  AOI22_X1 U30790 ( .A1(n20992), .A2(\xmem_data[14][0] ), .B1(n14990), .B2(
        \xmem_data[15][0] ), .ZN(n27346) );
  NAND2_X1 U30791 ( .A1(n27347), .A2(n27346), .ZN(n27348) );
  NAND3_X1 U30792 ( .A1(n27351), .A2(n27350), .A3(n27349), .ZN(n27357) );
  AOI22_X1 U30793 ( .A1(n25581), .A2(\xmem_data[0][0] ), .B1(n25401), .B2(
        \xmem_data[1][0] ), .ZN(n27355) );
  AOI22_X1 U30794 ( .A1(n29126), .A2(\xmem_data[2][0] ), .B1(n29151), .B2(
        \xmem_data[3][0] ), .ZN(n27354) );
  AOI22_X1 U30795 ( .A1(n29136), .A2(\xmem_data[4][0] ), .B1(n25407), .B2(
        \xmem_data[5][0] ), .ZN(n27353) );
  AOI22_X1 U30796 ( .A1(n29125), .A2(\xmem_data[6][0] ), .B1(n29124), .B2(
        \xmem_data[7][0] ), .ZN(n27352) );
  NAND4_X1 U30797 ( .A1(n27355), .A2(n27354), .A3(n27353), .A4(n27352), .ZN(
        n27356) );
  OR2_X1 U30798 ( .A1(n27357), .A2(n27356), .ZN(n27358) );
  OAI21_X1 U30799 ( .B1(n27359), .B2(n27358), .A(n29143), .ZN(n27432) );
  AOI22_X1 U30800 ( .A1(n24132), .A2(\xmem_data[118][0] ), .B1(n28298), .B2(
        \xmem_data[119][0] ), .ZN(n27363) );
  AOI22_X1 U30801 ( .A1(n29180), .A2(\xmem_data[116][0] ), .B1(n29179), .B2(
        \xmem_data[117][0] ), .ZN(n27362) );
  AOI22_X1 U30802 ( .A1(n28307), .A2(\xmem_data[114][0] ), .B1(n30551), .B2(
        \xmem_data[115][0] ), .ZN(n27361) );
  AOI22_X1 U30803 ( .A1(n29181), .A2(\xmem_data[112][0] ), .B1(n27396), .B2(
        \xmem_data[113][0] ), .ZN(n27360) );
  AOI22_X1 U30804 ( .A1(n30598), .A2(\xmem_data[96][0] ), .B1(n3301), .B2(
        \xmem_data[97][0] ), .ZN(n27364) );
  INV_X1 U30805 ( .A(n27364), .ZN(n27369) );
  AOI22_X1 U30806 ( .A1(n17050), .A2(\xmem_data[102][0] ), .B1(n25630), .B2(
        \xmem_data[103][0] ), .ZN(n27367) );
  AOI22_X1 U30807 ( .A1(n27365), .A2(\xmem_data[98][0] ), .B1(n3172), .B2(
        \xmem_data[99][0] ), .ZN(n27366) );
  NAND2_X1 U30808 ( .A1(n27367), .A2(n27366), .ZN(n27368) );
  NOR2_X1 U30809 ( .A1(n27369), .A2(n27368), .ZN(n27375) );
  AOI22_X1 U30810 ( .A1(n27526), .A2(\xmem_data[100][0] ), .B1(n30754), .B2(
        \xmem_data[101][0] ), .ZN(n27374) );
  AOI22_X1 U30811 ( .A1(n20544), .A2(\xmem_data[120][0] ), .B1(n25461), .B2(
        \xmem_data[121][0] ), .ZN(n27373) );
  AOI22_X1 U30812 ( .A1(n29188), .A2(\xmem_data[122][0] ), .B1(n17020), .B2(
        \xmem_data[123][0] ), .ZN(n27372) );
  AOI22_X1 U30813 ( .A1(n24645), .A2(\xmem_data[124][0] ), .B1(n28302), .B2(
        \xmem_data[125][0] ), .ZN(n27371) );
  AOI22_X1 U30814 ( .A1(n29190), .A2(\xmem_data[126][0] ), .B1(n3206), .B2(
        \xmem_data[127][0] ), .ZN(n27370) );
  NAND4_X1 U30815 ( .A1(n3837), .A2(n27375), .A3(n27374), .A4(n3506), .ZN(
        n27381) );
  AOI22_X1 U30816 ( .A1(n31346), .A2(\xmem_data[104][0] ), .B1(n28039), .B2(
        \xmem_data[105][0] ), .ZN(n27379) );
  AOI22_X1 U30817 ( .A1(n29173), .A2(\xmem_data[106][0] ), .B1(n27902), .B2(
        \xmem_data[107][0] ), .ZN(n27378) );
  AOI22_X1 U30818 ( .A1(n3221), .A2(\xmem_data[108][0] ), .B1(n24632), .B2(
        \xmem_data[109][0] ), .ZN(n27377) );
  AOI22_X1 U30819 ( .A1(n20723), .A2(\xmem_data[110][0] ), .B1(n29174), .B2(
        \xmem_data[111][0] ), .ZN(n27376) );
  NAND4_X1 U30820 ( .A1(n27379), .A2(n27378), .A3(n27377), .A4(n27376), .ZN(
        n27380) );
  OAI21_X1 U30821 ( .B1(n27381), .B2(n27380), .A(n29171), .ZN(n27431) );
  AOI22_X1 U30822 ( .A1(n30495), .A2(\xmem_data[64][0] ), .B1(n24623), .B2(
        \xmem_data[65][0] ), .ZN(n27386) );
  AOI22_X1 U30823 ( .A1(n28495), .A2(\xmem_data[66][0] ), .B1(n24685), .B2(
        \xmem_data[67][0] ), .ZN(n27385) );
  AND2_X1 U30824 ( .A1(n25527), .A2(\xmem_data[68][0] ), .ZN(n27382) );
  AOI21_X1 U30825 ( .B1(n25628), .B2(\xmem_data[69][0] ), .A(n27382), .ZN(
        n27384) );
  AOI22_X1 U30826 ( .A1(n20769), .A2(\xmem_data[70][0] ), .B1(n20710), .B2(
        \xmem_data[71][0] ), .ZN(n27383) );
  NAND4_X1 U30827 ( .A1(n27386), .A2(n27385), .A3(n27384), .A4(n27383), .ZN(
        n27404) );
  AND2_X1 U30828 ( .A1(n29173), .A2(\xmem_data[74][0] ), .ZN(n27387) );
  AOI21_X1 U30829 ( .B1(n20576), .B2(\xmem_data[75][0] ), .A(n27387), .ZN(
        n27391) );
  AOI22_X1 U30830 ( .A1(n31262), .A2(\xmem_data[72][0] ), .B1(n3245), .B2(
        \xmem_data[73][0] ), .ZN(n27390) );
  AOI22_X1 U30831 ( .A1(n3217), .A2(\xmem_data[76][0] ), .B1(n24533), .B2(
        \xmem_data[77][0] ), .ZN(n27389) );
  AOI22_X1 U30832 ( .A1(n31367), .A2(\xmem_data[78][0] ), .B1(n29174), .B2(
        \xmem_data[79][0] ), .ZN(n27388) );
  NAND4_X1 U30833 ( .A1(n27391), .A2(n27390), .A3(n27389), .A4(n27388), .ZN(
        n27403) );
  AOI22_X1 U30834 ( .A1(n30541), .A2(\xmem_data[88][0] ), .B1(n25607), .B2(
        \xmem_data[89][0] ), .ZN(n27395) );
  AOI22_X1 U30835 ( .A1(n29162), .A2(\xmem_data[90][0] ), .B1(n24133), .B2(
        \xmem_data[91][0] ), .ZN(n27394) );
  AOI22_X1 U30836 ( .A1(n29048), .A2(\xmem_data[92][0] ), .B1(n24115), .B2(
        \xmem_data[93][0] ), .ZN(n27393) );
  AOI22_X1 U30837 ( .A1(n29190), .A2(\xmem_data[94][0] ), .B1(n3205), .B2(
        \xmem_data[95][0] ), .ZN(n27392) );
  NAND4_X1 U30838 ( .A1(n27395), .A2(n27394), .A3(n27393), .A4(n27392), .ZN(
        n27402) );
  AOI22_X1 U30839 ( .A1(n29180), .A2(\xmem_data[84][0] ), .B1(n29179), .B2(
        \xmem_data[85][0] ), .ZN(n27400) );
  AOI22_X1 U30840 ( .A1(n15011), .A2(\xmem_data[82][0] ), .B1(n23813), .B2(
        \xmem_data[83][0] ), .ZN(n27399) );
  AOI22_X1 U30841 ( .A1(n29181), .A2(\xmem_data[80][0] ), .B1(n27396), .B2(
        \xmem_data[81][0] ), .ZN(n27398) );
  AOI22_X1 U30842 ( .A1(n14998), .A2(\xmem_data[86][0] ), .B1(n25710), .B2(
        \xmem_data[87][0] ), .ZN(n27397) );
  NAND4_X1 U30843 ( .A1(n27400), .A2(n27399), .A3(n27398), .A4(n27397), .ZN(
        n27401) );
  OR4_X1 U30844 ( .A1(n27404), .A2(n27403), .A3(n27402), .A4(n27401), .ZN(
        n27405) );
  NAND2_X1 U30845 ( .A1(n27405), .A2(n29201), .ZN(n27430) );
  NAND2_X1 U30846 ( .A1(n29151), .A2(\xmem_data[35][0] ), .ZN(n27407) );
  NAND2_X1 U30847 ( .A1(n29126), .A2(\xmem_data[34][0] ), .ZN(n27406) );
  NAND2_X1 U30848 ( .A1(n27407), .A2(n27406), .ZN(n27408) );
  AOI21_X1 U30849 ( .B1(n27568), .B2(\xmem_data[37][0] ), .A(n27408), .ZN(
        n27411) );
  AOI22_X1 U30850 ( .A1(n29089), .A2(\xmem_data[32][0] ), .B1(n24571), .B2(
        \xmem_data[33][0] ), .ZN(n27410) );
  AOI22_X1 U30851 ( .A1(n27567), .A2(\xmem_data[38][0] ), .B1(n25441), .B2(
        \xmem_data[39][0] ), .ZN(n27409) );
  NAND4_X1 U30852 ( .A1(n27411), .A2(n27410), .A3(n27409), .A4(n3975), .ZN(
        n27422) );
  AOI22_X1 U30853 ( .A1(n28375), .A2(\xmem_data[54][0] ), .B1(n29109), .B2(
        \xmem_data[55][0] ), .ZN(n27415) );
  AOI22_X1 U30854 ( .A1(n29103), .A2(\xmem_data[50][0] ), .B1(n27447), .B2(
        \xmem_data[51][0] ), .ZN(n27414) );
  AOI22_X1 U30855 ( .A1(n3358), .A2(\xmem_data[52][0] ), .B1(n20545), .B2(
        \xmem_data[53][0] ), .ZN(n27413) );
  AOI22_X1 U30856 ( .A1(n29104), .A2(\xmem_data[48][0] ), .B1(n29157), .B2(
        \xmem_data[49][0] ), .ZN(n27412) );
  NAND4_X1 U30857 ( .A1(n27415), .A2(n27414), .A3(n27413), .A4(n27412), .ZN(
        n27421) );
  AOI22_X1 U30858 ( .A1(n27516), .A2(\xmem_data[58][0] ), .B1(n20585), .B2(
        \xmem_data[59][0] ), .ZN(n27419) );
  AOI22_X1 U30859 ( .A1(n27536), .A2(\xmem_data[56][0] ), .B1(n20776), .B2(
        \xmem_data[57][0] ), .ZN(n27418) );
  AOI22_X1 U30860 ( .A1(n31270), .A2(\xmem_data[60][0] ), .B1(n29047), .B2(
        \xmem_data[61][0] ), .ZN(n27417) );
  AOI22_X1 U30861 ( .A1(n24190), .A2(\xmem_data[63][0] ), .B1(
        \xmem_data[62][0] ), .B2(n29101), .ZN(n27416) );
  NAND4_X1 U30862 ( .A1(n27419), .A2(n27418), .A3(n27417), .A4(n27416), .ZN(
        n27420) );
  AOI22_X1 U30863 ( .A1(n25357), .A2(\xmem_data[40][0] ), .B1(n25443), .B2(
        \xmem_data[41][0] ), .ZN(n27426) );
  AOI22_X1 U30864 ( .A1(n24172), .A2(\xmem_data[42][0] ), .B1(n27502), .B2(
        \xmem_data[43][0] ), .ZN(n27425) );
  AOI22_X1 U30865 ( .A1(n3221), .A2(\xmem_data[44][0] ), .B1(n29422), .B2(
        \xmem_data[45][0] ), .ZN(n27424) );
  AOI22_X1 U30866 ( .A1(n29095), .A2(\xmem_data[46][0] ), .B1(n17010), .B2(
        \xmem_data[47][0] ), .ZN(n27423) );
  NAND4_X1 U30867 ( .A1(n27426), .A2(n27425), .A3(n27424), .A4(n27423), .ZN(
        n27427) );
  OAI21_X1 U30868 ( .B1(n27428), .B2(n27427), .A(n29145), .ZN(n27429) );
  XNOR2_X1 U30869 ( .A(n35021), .B(\fmem_data[9][1] ), .ZN(n32226) );
  XNOR2_X1 U30870 ( .A(n35338), .B(\fmem_data[9][1] ), .ZN(n33197) );
  OAI22_X1 U30871 ( .A1(n32226), .A2(n34476), .B1(n3579), .B2(n33197), .ZN(
        n30491) );
  XNOR2_X1 U30872 ( .A(n32014), .B(\fmem_data[2][1] ), .ZN(n30982) );
  OAI22_X1 U30873 ( .A1(n33271), .A2(n3578), .B1(n30982), .B2(n34343), .ZN(
        n30490) );
  INV_X1 U30874 ( .A(n27434), .ZN(n29689) );
  XNOR2_X1 U30875 ( .A(n35340), .B(\fmem_data[20][1] ), .ZN(n33196) );
  AOI22_X1 U30876 ( .A1(n23730), .A2(\xmem_data[96][6] ), .B1(n27435), .B2(
        \xmem_data[97][6] ), .ZN(n27443) );
  AOI22_X1 U30877 ( .A1(n27436), .A2(\xmem_data[98][6] ), .B1(n28075), .B2(
        \xmem_data[99][6] ), .ZN(n27442) );
  AOI22_X1 U30878 ( .A1(n3306), .A2(\xmem_data[100][6] ), .B1(n27437), .B2(
        \xmem_data[101][6] ), .ZN(n27441) );
  AND2_X1 U30879 ( .A1(n3220), .A2(\xmem_data[103][6] ), .ZN(n27438) );
  AOI21_X1 U30880 ( .B1(n27439), .B2(\xmem_data[102][6] ), .A(n27438), .ZN(
        n27440) );
  NAND4_X1 U30881 ( .A1(n27443), .A2(n27442), .A3(n27441), .A4(n27440), .ZN(
        n27471) );
  AOI22_X1 U30882 ( .A1(n27445), .A2(\xmem_data[104][6] ), .B1(n27444), .B2(
        \xmem_data[105][6] ), .ZN(n27451) );
  AOI22_X1 U30883 ( .A1(n29257), .A2(\xmem_data[106][6] ), .B1(n28509), .B2(
        \xmem_data[107][6] ), .ZN(n27450) );
  AOI22_X1 U30884 ( .A1(n30295), .A2(\xmem_data[108][6] ), .B1(n27446), .B2(
        \xmem_data[109][6] ), .ZN(n27449) );
  AOI22_X1 U30885 ( .A1(n27447), .A2(\xmem_data[110][6] ), .B1(n20982), .B2(
        \xmem_data[111][6] ), .ZN(n27448) );
  NAND4_X1 U30886 ( .A1(n27451), .A2(n27450), .A3(n27449), .A4(n27448), .ZN(
        n27470) );
  AOI22_X1 U30887 ( .A1(n27453), .A2(\xmem_data[112][6] ), .B1(n27452), .B2(
        \xmem_data[113][6] ), .ZN(n27459) );
  AOI22_X1 U30888 ( .A1(n28298), .A2(\xmem_data[114][6] ), .B1(n30541), .B2(
        \xmem_data[115][6] ), .ZN(n27458) );
  AOI22_X1 U30889 ( .A1(n23795), .A2(\xmem_data[116][6] ), .B1(n27454), .B2(
        \xmem_data[117][6] ), .ZN(n27457) );
  AOI22_X1 U30890 ( .A1(n24509), .A2(\xmem_data[118][6] ), .B1(n28492), .B2(
        \xmem_data[119][6] ), .ZN(n27456) );
  NAND4_X1 U30891 ( .A1(n27459), .A2(n27458), .A3(n27457), .A4(n27456), .ZN(
        n27469) );
  AOI22_X1 U30892 ( .A1(n25678), .A2(\xmem_data[120][6] ), .B1(n27460), .B2(
        \xmem_data[121][6] ), .ZN(n27467) );
  AOI22_X1 U30893 ( .A1(n27462), .A2(\xmem_data[122][6] ), .B1(n27461), .B2(
        \xmem_data[123][6] ), .ZN(n27466) );
  AOI22_X1 U30894 ( .A1(n25401), .A2(\xmem_data[124][6] ), .B1(n24570), .B2(
        \xmem_data[125][6] ), .ZN(n27465) );
  AOI22_X1 U30895 ( .A1(n25526), .A2(\xmem_data[126][6] ), .B1(n27463), .B2(
        \xmem_data[127][6] ), .ZN(n27464) );
  NAND4_X1 U30896 ( .A1(n27467), .A2(n27466), .A3(n27465), .A4(n27464), .ZN(
        n27468) );
  OR4_X1 U30897 ( .A1(n27471), .A2(n27470), .A3(n27469), .A4(n27468), .ZN(
        n27497) );
  AOI22_X1 U30898 ( .A1(n27498), .A2(\xmem_data[64][6] ), .B1(n24468), .B2(
        \xmem_data[65][6] ), .ZN(n27476) );
  AOI22_X1 U30899 ( .A1(n27500), .A2(\xmem_data[66][6] ), .B1(n27499), .B2(
        \xmem_data[67][6] ), .ZN(n27475) );
  AOI22_X1 U30900 ( .A1(n27813), .A2(\xmem_data[68][6] ), .B1(n27501), .B2(
        \xmem_data[69][6] ), .ZN(n27474) );
  AND2_X1 U30901 ( .A1(n3217), .A2(\xmem_data[71][6] ), .ZN(n27472) );
  AOI21_X1 U30902 ( .B1(n27502), .B2(\xmem_data[70][6] ), .A(n27472), .ZN(
        n27473) );
  NAND4_X1 U30903 ( .A1(n27476), .A2(n27475), .A3(n27474), .A4(n27473), .ZN(
        n27493) );
  AOI22_X1 U30904 ( .A1(n30872), .A2(\xmem_data[88][6] ), .B1(n27523), .B2(
        \xmem_data[89][6] ), .ZN(n27480) );
  AOI22_X1 U30905 ( .A1(n27524), .A2(\xmem_data[90][6] ), .B1(n24117), .B2(
        \xmem_data[91][6] ), .ZN(n27479) );
  AOI22_X1 U30906 ( .A1(n28202), .A2(\xmem_data[92][6] ), .B1(n27525), .B2(
        \xmem_data[93][6] ), .ZN(n27478) );
  AOI22_X1 U30907 ( .A1(n3209), .A2(\xmem_data[94][6] ), .B1(n27526), .B2(
        \xmem_data[95][6] ), .ZN(n27477) );
  NAND4_X1 U30908 ( .A1(n27480), .A2(n27479), .A3(n27478), .A4(n27477), .ZN(
        n27491) );
  AOI22_X1 U30909 ( .A1(n27514), .A2(\xmem_data[80][6] ), .B1(n27513), .B2(
        \xmem_data[81][6] ), .ZN(n27484) );
  AOI22_X1 U30910 ( .A1(n27515), .A2(\xmem_data[82][6] ), .B1(n22703), .B2(
        \xmem_data[83][6] ), .ZN(n27483) );
  AOI22_X1 U30911 ( .A1(n29396), .A2(\xmem_data[84][6] ), .B1(n27516), .B2(
        \xmem_data[85][6] ), .ZN(n27482) );
  AOI22_X1 U30912 ( .A1(n24133), .A2(\xmem_data[86][6] ), .B1(n27518), .B2(
        \xmem_data[87][6] ), .ZN(n27481) );
  NAND4_X1 U30913 ( .A1(n27484), .A2(n27483), .A3(n27482), .A4(n27481), .ZN(
        n27490) );
  AOI22_X1 U30914 ( .A1(n24533), .A2(\xmem_data[72][6] ), .B1(n27507), .B2(
        \xmem_data[73][6] ), .ZN(n27488) );
  AOI22_X1 U30915 ( .A1(n24697), .A2(\xmem_data[74][6] ), .B1(n13444), .B2(
        \xmem_data[75][6] ), .ZN(n27487) );
  AOI22_X1 U30916 ( .A1(n3282), .A2(\xmem_data[76][6] ), .B1(n15011), .B2(
        \xmem_data[77][6] ), .ZN(n27486) );
  AOI22_X1 U30917 ( .A1(n27508), .A2(\xmem_data[78][6] ), .B1(n25456), .B2(
        \xmem_data[79][6] ), .ZN(n27485) );
  NAND4_X1 U30918 ( .A1(n27488), .A2(n27487), .A3(n27486), .A4(n27485), .ZN(
        n27489) );
  OR3_X1 U30919 ( .A1(n27491), .A2(n27490), .A3(n27489), .ZN(n27492) );
  OR2_X1 U30920 ( .A1(n27493), .A2(n27492), .ZN(n27495) );
  AOI22_X1 U30921 ( .A1(n27497), .A2(n27496), .B1(n27495), .B2(n27494), .ZN(
        n27580) );
  AOI22_X1 U30922 ( .A1(n27498), .A2(\xmem_data[32][6] ), .B1(n25388), .B2(
        \xmem_data[33][6] ), .ZN(n27506) );
  AOI22_X1 U30923 ( .A1(n27500), .A2(\xmem_data[34][6] ), .B1(n27499), .B2(
        \xmem_data[35][6] ), .ZN(n27505) );
  AOI22_X1 U30924 ( .A1(n3449), .A2(\xmem_data[36][6] ), .B1(n27501), .B2(
        \xmem_data[37][6] ), .ZN(n27504) );
  AOI22_X1 U30925 ( .A1(n27502), .A2(\xmem_data[38][6] ), .B1(n3220), .B2(
        \xmem_data[39][6] ), .ZN(n27503) );
  NAND4_X1 U30926 ( .A1(n27506), .A2(n27505), .A3(n27504), .A4(n27503), .ZN(
        n27534) );
  AOI22_X1 U30927 ( .A1(n29256), .A2(\xmem_data[40][6] ), .B1(n27507), .B2(
        \xmem_data[41][6] ), .ZN(n27512) );
  AOI22_X1 U30928 ( .A1(n20807), .A2(\xmem_data[42][6] ), .B1(n13444), .B2(
        \xmem_data[43][6] ), .ZN(n27511) );
  AOI22_X1 U30929 ( .A1(n3140), .A2(\xmem_data[44][6] ), .B1(n31252), .B2(
        \xmem_data[45][6] ), .ZN(n27510) );
  AOI22_X1 U30930 ( .A1(n27508), .A2(\xmem_data[46][6] ), .B1(n3357), .B2(
        \xmem_data[47][6] ), .ZN(n27509) );
  NAND4_X1 U30931 ( .A1(n27512), .A2(n27511), .A3(n27510), .A4(n27509), .ZN(
        n27533) );
  AOI22_X1 U30932 ( .A1(n27514), .A2(\xmem_data[48][6] ), .B1(n27513), .B2(
        \xmem_data[49][6] ), .ZN(n27522) );
  AOI22_X1 U30933 ( .A1(n27515), .A2(\xmem_data[50][6] ), .B1(n28517), .B2(
        \xmem_data[51][6] ), .ZN(n27521) );
  AOI22_X1 U30934 ( .A1(n25461), .A2(\xmem_data[52][6] ), .B1(n27516), .B2(
        \xmem_data[53][6] ), .ZN(n27520) );
  AOI22_X1 U30935 ( .A1(n29317), .A2(\xmem_data[54][6] ), .B1(n27518), .B2(
        \xmem_data[55][6] ), .ZN(n27519) );
  NAND4_X1 U30936 ( .A1(n27522), .A2(n27521), .A3(n27520), .A4(n27519), .ZN(
        n27532) );
  AOI22_X1 U30937 ( .A1(n29047), .A2(\xmem_data[56][6] ), .B1(n27523), .B2(
        \xmem_data[57][6] ), .ZN(n27530) );
  AOI22_X1 U30938 ( .A1(n27524), .A2(\xmem_data[58][6] ), .B1(n30955), .B2(
        \xmem_data[59][6] ), .ZN(n27529) );
  AOI22_X1 U30939 ( .A1(n29297), .A2(\xmem_data[60][6] ), .B1(n27525), .B2(
        \xmem_data[61][6] ), .ZN(n27528) );
  AOI22_X1 U30940 ( .A1(n22719), .A2(\xmem_data[62][6] ), .B1(n27526), .B2(
        \xmem_data[63][6] ), .ZN(n27527) );
  NAND4_X1 U30941 ( .A1(n27530), .A2(n27529), .A3(n27528), .A4(n27527), .ZN(
        n27531) );
  OR4_X1 U30942 ( .A1(n27534), .A2(n27533), .A3(n27532), .A4(n27531), .ZN(
        n27578) );
  AOI22_X1 U30943 ( .A1(n20545), .A2(\xmem_data[16][6] ), .B1(n27535), .B2(
        \xmem_data[17][6] ), .ZN(n27541) );
  AOI22_X1 U30944 ( .A1(n20541), .A2(\xmem_data[18][6] ), .B1(n27536), .B2(
        \xmem_data[19][6] ), .ZN(n27540) );
  AOI22_X1 U30945 ( .A1(n25519), .A2(\xmem_data[20][6] ), .B1(n27516), .B2(
        \xmem_data[21][6] ), .ZN(n27539) );
  AOI22_X1 U30946 ( .A1(n20585), .A2(\xmem_data[22][6] ), .B1(n14970), .B2(
        \xmem_data[23][6] ), .ZN(n27538) );
  NAND4_X1 U30947 ( .A1(n27541), .A2(n27540), .A3(n27539), .A4(n27538), .ZN(
        n27549) );
  AOI22_X1 U30948 ( .A1(n22682), .A2(\xmem_data[24][6] ), .B1(n13452), .B2(
        \xmem_data[25][6] ), .ZN(n27546) );
  AOI22_X1 U30949 ( .A1(n14972), .A2(\xmem_data[26][6] ), .B1(n23778), .B2(
        \xmem_data[27][6] ), .ZN(n27545) );
  AOI22_X1 U30950 ( .A1(n29054), .A2(\xmem_data[28][6] ), .B1(n14975), .B2(
        \xmem_data[29][6] ), .ZN(n27544) );
  AOI22_X1 U30951 ( .A1(n27542), .A2(\xmem_data[30][6] ), .B1(n28979), .B2(
        \xmem_data[31][6] ), .ZN(n27543) );
  NAND4_X1 U30952 ( .A1(n27546), .A2(n27545), .A3(n27544), .A4(n27543), .ZN(
        n27548) );
  OR3_X1 U30953 ( .A1(n27549), .A2(n27548), .A3(n3977), .ZN(n27560) );
  AOI22_X1 U30954 ( .A1(n25449), .A2(\xmem_data[10][6] ), .B1(n27550), .B2(
        \xmem_data[11][6] ), .ZN(n27558) );
  AOI22_X1 U30955 ( .A1(n27551), .A2(\xmem_data[14][6] ), .B1(n14996), .B2(
        \xmem_data[15][6] ), .ZN(n27552) );
  INV_X1 U30956 ( .A(n27552), .ZN(n27556) );
  AND2_X1 U30957 ( .A1(n3375), .A2(\xmem_data[12][6] ), .ZN(n27555) );
  AOI22_X1 U30958 ( .A1(n29698), .A2(\xmem_data[8][6] ), .B1(n20500), .B2(
        \xmem_data[9][6] ), .ZN(n27553) );
  INV_X1 U30959 ( .A(n27553), .ZN(n27554) );
  NOR3_X1 U30960 ( .A1(n27556), .A2(n27555), .A3(n27554), .ZN(n27557) );
  NAND2_X1 U30961 ( .A1(n27558), .A2(n27557), .ZN(n27559) );
  NOR2_X1 U30962 ( .A1(n27560), .A2(n27559), .ZN(n27575) );
  AND2_X1 U30963 ( .A1(n3221), .A2(\xmem_data[7][6] ), .ZN(n27561) );
  AOI21_X1 U30964 ( .B1(n28470), .B2(\xmem_data[6][6] ), .A(n27561), .ZN(
        n27562) );
  INV_X1 U30965 ( .A(n27562), .ZN(n27572) );
  AOI22_X1 U30966 ( .A1(n27564), .A2(\xmem_data[2][6] ), .B1(n27563), .B2(
        \xmem_data[3][6] ), .ZN(n27566) );
  AOI22_X1 U30967 ( .A1(n3317), .A2(\xmem_data[4][6] ), .B1(n25360), .B2(
        \xmem_data[5][6] ), .ZN(n27565) );
  NAND2_X1 U30968 ( .A1(n27566), .A2(n27565), .ZN(n27571) );
  AOI22_X1 U30969 ( .A1(n27568), .A2(\xmem_data[0][6] ), .B1(n27567), .B2(
        \xmem_data[1][6] ), .ZN(n27569) );
  INV_X1 U30970 ( .A(n27569), .ZN(n27570) );
  NOR3_X1 U30971 ( .A1(n27572), .A2(n27571), .A3(n27570), .ZN(n27574) );
  AOI21_X1 U30972 ( .B1(n27575), .B2(n27574), .A(n27573), .ZN(n27576) );
  AOI21_X1 U30973 ( .B1(n27578), .B2(n27577), .A(n27576), .ZN(n27579) );
  XNOR2_X1 U30974 ( .A(n35178), .B(\fmem_data[20][1] ), .ZN(n33877) );
  OAI22_X1 U30975 ( .A1(n33196), .A2(n3647), .B1(n33877), .B2(n36227), .ZN(
        n28937) );
  XNOR2_X1 U30976 ( .A(n35324), .B(\fmem_data[4][1] ), .ZN(n33162) );
  XNOR2_X1 U30977 ( .A(n33055), .B(\fmem_data[4][1] ), .ZN(n31896) );
  OAI22_X1 U30978 ( .A1(n33162), .A2(n3569), .B1(n31896), .B2(n34598), .ZN(
        n28935) );
  XNOR2_X1 U30979 ( .A(n32025), .B(\fmem_data[12][3] ), .ZN(n32236) );
  AOI22_X1 U30980 ( .A1(n28680), .A2(\xmem_data[44][0] ), .B1(n30266), .B2(
        \xmem_data[45][0] ), .ZN(n27584) );
  AOI22_X1 U30981 ( .A1(n29630), .A2(\xmem_data[60][0] ), .B1(n30776), .B2(
        \xmem_data[61][0] ), .ZN(n27587) );
  AOI22_X1 U30982 ( .A1(n3162), .A2(\xmem_data[40][0] ), .B1(n3186), .B2(
        \xmem_data[41][0] ), .ZN(n27586) );
  AOI22_X1 U30983 ( .A1(n3174), .A2(\xmem_data[36][0] ), .B1(n29768), .B2(
        \xmem_data[37][0] ), .ZN(n27585) );
  NAND3_X1 U30984 ( .A1(n27587), .A2(n27586), .A3(n27585), .ZN(n27588) );
  NOR2_X1 U30985 ( .A1(n27589), .A2(n27588), .ZN(n27612) );
  AOI22_X1 U30986 ( .A1(n29641), .A2(\xmem_data[46][0] ), .B1(n29246), .B2(
        \xmem_data[47][0] ), .ZN(n27590) );
  INV_X1 U30987 ( .A(n27590), .ZN(n27596) );
  AOI22_X1 U30988 ( .A1(n29616), .A2(\xmem_data[48][0] ), .B1(n29579), .B2(
        \xmem_data[49][0] ), .ZN(n27594) );
  AOI22_X1 U30989 ( .A1(n29617), .A2(\xmem_data[50][0] ), .B1(n21060), .B2(
        \xmem_data[51][0] ), .ZN(n27593) );
  AOI22_X1 U30990 ( .A1(n29619), .A2(\xmem_data[52][0] ), .B1(n29618), .B2(
        \xmem_data[53][0] ), .ZN(n27592) );
  AOI22_X1 U30991 ( .A1(n29621), .A2(\xmem_data[54][0] ), .B1(n3142), .B2(
        \xmem_data[55][0] ), .ZN(n27591) );
  NAND4_X1 U30992 ( .A1(n27594), .A2(n27593), .A3(n27592), .A4(n27591), .ZN(
        n27595) );
  NOR2_X1 U30993 ( .A1(n27596), .A2(n27595), .ZN(n27611) );
  AOI22_X1 U30994 ( .A1(n29667), .A2(\xmem_data[62][0] ), .B1(n30698), .B2(
        \xmem_data[63][0] ), .ZN(n27599) );
  AOI22_X1 U30995 ( .A1(n29649), .A2(\xmem_data[38][0] ), .B1(n30948), .B2(
        \xmem_data[39][0] ), .ZN(n27598) );
  AOI22_X1 U30996 ( .A1(n29603), .A2(\xmem_data[34][0] ), .B1(n28089), .B2(
        \xmem_data[35][0] ), .ZN(n27597) );
  NAND3_X1 U30997 ( .A1(n27599), .A2(n27598), .A3(n27597), .ZN(n27602) );
  AOI22_X1 U30998 ( .A1(n28755), .A2(\xmem_data[42][0] ), .B1(n29439), .B2(
        \xmem_data[43][0] ), .ZN(n27600) );
  INV_X1 U30999 ( .A(n27600), .ZN(n27601) );
  NOR2_X1 U31000 ( .A1(n27602), .A2(n27601), .ZN(n27610) );
  NAND2_X1 U31001 ( .A1(n28665), .A2(\xmem_data[33][0] ), .ZN(n27604) );
  NAND2_X1 U31002 ( .A1(n29481), .A2(\xmem_data[32][0] ), .ZN(n27603) );
  NAND2_X1 U31003 ( .A1(n27604), .A2(n27603), .ZN(n27608) );
  AOI22_X1 U31004 ( .A1(n29628), .A2(\xmem_data[58][0] ), .B1(n29627), .B2(
        \xmem_data[59][0] ), .ZN(n27606) );
  AOI22_X1 U31005 ( .A1(n28136), .A2(\xmem_data[56][0] ), .B1(n29672), .B2(
        \xmem_data[57][0] ), .ZN(n27605) );
  NAND2_X1 U31006 ( .A1(n27606), .A2(n27605), .ZN(n27607) );
  NOR2_X1 U31007 ( .A1(n27608), .A2(n27607), .ZN(n27609) );
  NAND4_X1 U31008 ( .A1(n27612), .A2(n27611), .A3(n27610), .A4(n27609), .ZN(
        n27613) );
  NAND2_X1 U31009 ( .A1(n27613), .A2(n29683), .ZN(n27697) );
  AOI22_X1 U31010 ( .A1(n30070), .A2(\xmem_data[106][0] ), .B1(n29639), .B2(
        \xmem_data[107][0] ), .ZN(n27633) );
  NAND2_X1 U31011 ( .A1(n27761), .A2(\xmem_data[97][0] ), .ZN(n27615) );
  NAND2_X1 U31012 ( .A1(n30191), .A2(\xmem_data[96][0] ), .ZN(n27614) );
  NAND2_X1 U31013 ( .A1(n27615), .A2(n27614), .ZN(n27625) );
  AOI22_X1 U31014 ( .A1(n29593), .A2(\xmem_data[102][0] ), .B1(n3120), .B2(
        \xmem_data[103][0] ), .ZN(n27618) );
  AOI22_X1 U31015 ( .A1(n29574), .A2(\xmem_data[110][0] ), .B1(n29573), .B2(
        \xmem_data[111][0] ), .ZN(n27617) );
  AOI22_X1 U31016 ( .A1(n3239), .A2(\xmem_data[98][0] ), .B1(n29591), .B2(
        \xmem_data[99][0] ), .ZN(n27616) );
  NAND3_X1 U31017 ( .A1(n27618), .A2(n27617), .A3(n27616), .ZN(n27624) );
  AOI22_X1 U31018 ( .A1(n29580), .A2(\xmem_data[112][0] ), .B1(n29615), .B2(
        \xmem_data[113][0] ), .ZN(n27622) );
  AOI22_X1 U31019 ( .A1(n29581), .A2(\xmem_data[114][0] ), .B1(n29657), .B2(
        \xmem_data[115][0] ), .ZN(n27621) );
  AOI22_X1 U31020 ( .A1(n29583), .A2(\xmem_data[116][0] ), .B1(n29582), .B2(
        \xmem_data[117][0] ), .ZN(n27620) );
  AOI22_X1 U31021 ( .A1(n29584), .A2(\xmem_data[118][0] ), .B1(n3144), .B2(
        \xmem_data[119][0] ), .ZN(n27619) );
  NAND4_X1 U31022 ( .A1(n27622), .A2(n27621), .A3(n27620), .A4(n27619), .ZN(
        n27623) );
  NOR3_X1 U31023 ( .A1(n27625), .A2(n27624), .A3(n27623), .ZN(n27632) );
  AOI22_X1 U31024 ( .A1(n27754), .A2(\xmem_data[100][0] ), .B1(n29768), .B2(
        \xmem_data[101][0] ), .ZN(n27626) );
  AOI22_X1 U31025 ( .A1(n3162), .A2(\xmem_data[104][0] ), .B1(n3182), .B2(
        \xmem_data[105][0] ), .ZN(n27627) );
  INV_X1 U31026 ( .A(n27627), .ZN(n27630) );
  AOI22_X1 U31027 ( .A1(n29363), .A2(\xmem_data[108][0] ), .B1(n30266), .B2(
        \xmem_data[109][0] ), .ZN(n27628) );
  INV_X1 U31028 ( .A(n27628), .ZN(n27629) );
  NOR2_X1 U31029 ( .A1(n27630), .A2(n27629), .ZN(n27631) );
  NAND4_X1 U31030 ( .A1(n27633), .A2(n27632), .A3(n27626), .A4(n27631), .ZN(
        n27639) );
  AOI22_X1 U31031 ( .A1(n29421), .A2(\xmem_data[120][0] ), .B1(n26616), .B2(
        \xmem_data[121][0] ), .ZN(n27637) );
  AOI22_X1 U31032 ( .A1(n28138), .A2(\xmem_data[122][0] ), .B1(n29565), .B2(
        \xmem_data[123][0] ), .ZN(n27636) );
  AOI22_X1 U31033 ( .A1(n29566), .A2(\xmem_data[124][0] ), .B1(n28208), .B2(
        \xmem_data[125][0] ), .ZN(n27635) );
  AOI22_X1 U31034 ( .A1(n29568), .A2(\xmem_data[126][0] ), .B1(n3345), .B2(
        \xmem_data[127][0] ), .ZN(n27634) );
  NAND4_X1 U31035 ( .A1(n27637), .A2(n27636), .A3(n27635), .A4(n27634), .ZN(
        n27638) );
  AOI22_X1 U31036 ( .A1(n3165), .A2(\xmem_data[8][0] ), .B1(n3184), .B2(
        \xmem_data[9][0] ), .ZN(n27640) );
  AOI22_X1 U31037 ( .A1(n29649), .A2(\xmem_data[6][0] ), .B1(n20776), .B2(
        \xmem_data[7][0] ), .ZN(n27643) );
  AOI22_X1 U31038 ( .A1(n29641), .A2(\xmem_data[14][0] ), .B1(n29054), .B2(
        \xmem_data[15][0] ), .ZN(n27642) );
  AOI22_X1 U31039 ( .A1(n28689), .A2(\xmem_data[10][0] ), .B1(n17021), .B2(
        \xmem_data[11][0] ), .ZN(n27641) );
  NAND3_X1 U31040 ( .A1(n27643), .A2(n27642), .A3(n27641), .ZN(n27644) );
  NOR2_X1 U31041 ( .A1(n27645), .A2(n27644), .ZN(n27664) );
  AND2_X1 U31042 ( .A1(n28751), .A2(\xmem_data[4][0] ), .ZN(n27648) );
  AOI22_X1 U31043 ( .A1(n3239), .A2(\xmem_data[2][0] ), .B1(n28233), .B2(
        \xmem_data[3][0] ), .ZN(n27646) );
  INV_X1 U31044 ( .A(n27646), .ZN(n27647) );
  AOI22_X1 U31045 ( .A1(\xmem_data[22][0] ), .A2(n29662), .B1(n29617), .B2(
        \xmem_data[18][0] ), .ZN(n27650) );
  AOI22_X1 U31046 ( .A1(\xmem_data[21][0] ), .A2(n29659), .B1(n29616), .B2(
        \xmem_data[16][0] ), .ZN(n27649) );
  NOR2_X1 U31047 ( .A1(n3973), .A2(n27651), .ZN(n27663) );
  AOI22_X1 U31048 ( .A1(n30248), .A2(\xmem_data[0][0] ), .B1(n3369), .B2(
        \xmem_data[1][0] ), .ZN(n27652) );
  AOI22_X1 U31049 ( .A1(n29488), .A2(\xmem_data[12][0] ), .B1(n30266), .B2(
        \xmem_data[13][0] ), .ZN(n27653) );
  INV_X1 U31050 ( .A(n27653), .ZN(n27661) );
  NAND2_X1 U31051 ( .A1(n29657), .A2(\xmem_data[19][0] ), .ZN(n27655) );
  NAND2_X1 U31052 ( .A1(n29661), .A2(\xmem_data[23][0] ), .ZN(n27654) );
  NAND2_X1 U31053 ( .A1(n27655), .A2(n27654), .ZN(n27656) );
  AOI21_X1 U31054 ( .B1(n29615), .B2(\xmem_data[17][0] ), .A(n27656), .ZN(
        n27659) );
  NAND2_X1 U31055 ( .A1(n29660), .A2(\xmem_data[20][0] ), .ZN(n27658) );
  NAND2_X1 U31056 ( .A1(n26884), .A2(\xmem_data[5][0] ), .ZN(n27657) );
  NAND3_X1 U31057 ( .A1(n27659), .A2(n27658), .A3(n27657), .ZN(n27660) );
  NOR2_X1 U31058 ( .A1(n27661), .A2(n27660), .ZN(n27662) );
  NAND4_X1 U31059 ( .A1(n27664), .A2(n27663), .A3(n27652), .A4(n27662), .ZN(
        n27670) );
  AOI22_X1 U31060 ( .A1(n27710), .A2(\xmem_data[24][0] ), .B1(n28766), .B2(
        \xmem_data[25][0] ), .ZN(n27668) );
  AOI22_X1 U31061 ( .A1(n30279), .A2(\xmem_data[26][0] ), .B1(n31368), .B2(
        \xmem_data[27][0] ), .ZN(n27667) );
  AOI22_X1 U31062 ( .A1(n29630), .A2(\xmem_data[28][0] ), .B1(n28667), .B2(
        \xmem_data[29][0] ), .ZN(n27666) );
  AOI22_X1 U31063 ( .A1(n29667), .A2(\xmem_data[30][0] ), .B1(n3345), .B2(
        \xmem_data[31][0] ), .ZN(n27665) );
  NAND4_X1 U31064 ( .A1(n27668), .A2(n27667), .A3(n27666), .A4(n27665), .ZN(
        n27669) );
  OAI21_X1 U31065 ( .B1(n27670), .B2(n27669), .A(n29681), .ZN(n27695) );
  AOI22_X1 U31066 ( .A1(n29647), .A2(\xmem_data[64][0] ), .B1(n28665), .B2(
        \xmem_data[65][0] ), .ZN(n27681) );
  AOI22_X1 U31067 ( .A1(n27754), .A2(\xmem_data[68][0] ), .B1(n29739), .B2(
        \xmem_data[69][0] ), .ZN(n27680) );
  AOI22_X1 U31068 ( .A1(n29656), .A2(\xmem_data[80][0] ), .B1(n29579), .B2(
        \xmem_data[81][0] ), .ZN(n27674) );
  AOI22_X1 U31069 ( .A1(n29658), .A2(\xmem_data[82][0] ), .B1(n27498), .B2(
        \xmem_data[83][0] ), .ZN(n27673) );
  AOI22_X1 U31070 ( .A1(n29583), .A2(\xmem_data[84][0] ), .B1(n29582), .B2(
        \xmem_data[85][0] ), .ZN(n27672) );
  AOI22_X1 U31071 ( .A1(n29584), .A2(\xmem_data[86][0] ), .B1(n3449), .B2(
        \xmem_data[87][0] ), .ZN(n27671) );
  NAND4_X1 U31072 ( .A1(n27674), .A2(n27673), .A3(n27672), .A4(n27671), .ZN(
        n27678) );
  AOI22_X1 U31073 ( .A1(n29593), .A2(\xmem_data[70][0] ), .B1(n24213), .B2(
        \xmem_data[71][0] ), .ZN(n27676) );
  AOI22_X1 U31074 ( .A1(n3239), .A2(\xmem_data[66][0] ), .B1(n29591), .B2(
        \xmem_data[67][0] ), .ZN(n27675) );
  NAND2_X1 U31075 ( .A1(n27676), .A2(n27675), .ZN(n27677) );
  NOR2_X1 U31076 ( .A1(n27678), .A2(n27677), .ZN(n27679) );
  NAND3_X1 U31077 ( .A1(n27681), .A2(n27680), .A3(n27679), .ZN(n27687) );
  AOI22_X1 U31078 ( .A1(n3168), .A2(\xmem_data[72][0] ), .B1(n3186), .B2(
        \xmem_data[73][0] ), .ZN(n27685) );
  AOI22_X1 U31079 ( .A1(n28755), .A2(\xmem_data[74][0] ), .B1(n24115), .B2(
        \xmem_data[75][0] ), .ZN(n27684) );
  AOI22_X1 U31080 ( .A1(n27713), .A2(\xmem_data[76][0] ), .B1(n30644), .B2(
        \xmem_data[77][0] ), .ZN(n27683) );
  AOI22_X1 U31081 ( .A1(n29574), .A2(\xmem_data[78][0] ), .B1(n29573), .B2(
        \xmem_data[79][0] ), .ZN(n27682) );
  NAND4_X1 U31082 ( .A1(n27685), .A2(n27684), .A3(n27683), .A4(n27682), .ZN(
        n27686) );
  AOI22_X1 U31083 ( .A1(n29433), .A2(\xmem_data[88][0] ), .B1(n30100), .B2(
        \xmem_data[89][0] ), .ZN(n27691) );
  AOI22_X1 U31084 ( .A1(n28207), .A2(\xmem_data[90][0] ), .B1(n29565), .B2(
        \xmem_data[91][0] ), .ZN(n27690) );
  AOI22_X1 U31085 ( .A1(n29674), .A2(\xmem_data[92][0] ), .B1(n3170), .B2(
        \xmem_data[93][0] ), .ZN(n27689) );
  AOI22_X1 U31086 ( .A1(n29568), .A2(\xmem_data[94][0] ), .B1(n3345), .B2(
        \xmem_data[95][0] ), .ZN(n27688) );
  NAND4_X1 U31087 ( .A1(n27691), .A2(n27690), .A3(n27689), .A4(n27688), .ZN(
        n27692) );
  INV_X1 U31088 ( .A(n35619), .ZN(n27698) );
  XNOR2_X1 U31089 ( .A(n31673), .B(\fmem_data[10][1] ), .ZN(n32583) );
  XNOR2_X1 U31090 ( .A(n31674), .B(\fmem_data[10][1] ), .ZN(n32729) );
  OAI22_X1 U31091 ( .A1(n32583), .A2(n36114), .B1(n32729), .B2(n3561), .ZN(
        n31142) );
  AOI22_X1 U31092 ( .A1(n27701), .A2(\xmem_data[48][0] ), .B1(n3198), .B2(
        \xmem_data[49][0] ), .ZN(n27707) );
  AOI22_X1 U31093 ( .A1(n27702), .A2(\xmem_data[50][0] ), .B1(n3140), .B2(
        \xmem_data[51][0] ), .ZN(n27706) );
  AOI22_X1 U31094 ( .A1(n29801), .A2(\xmem_data[52][0] ), .B1(n28238), .B2(
        \xmem_data[53][0] ), .ZN(n27705) );
  AOI22_X1 U31095 ( .A1(n29709), .A2(\xmem_data[54][0] ), .B1(n27763), .B2(
        \xmem_data[55][0] ), .ZN(n27704) );
  NAND4_X1 U31096 ( .A1(n27707), .A2(n27706), .A3(n27705), .A4(n27704), .ZN(
        n27739) );
  AND2_X1 U31097 ( .A1(n27708), .A2(\xmem_data[47][0] ), .ZN(n27709) );
  AOI21_X1 U31098 ( .B1(n29423), .B2(\xmem_data[46][0] ), .A(n27709), .ZN(
        n27712) );
  NAND2_X1 U31099 ( .A1(n27710), .A2(\xmem_data[44][0] ), .ZN(n27711) );
  AND2_X1 U31100 ( .A1(n27712), .A2(n27711), .ZN(n27736) );
  AOI22_X1 U31101 ( .A1(n29722), .A2(\xmem_data[32][0] ), .B1(n30266), .B2(
        \xmem_data[33][0] ), .ZN(n27722) );
  AOI22_X1 U31102 ( .A1(n27714), .A2(\xmem_data[34][0] ), .B1(n21056), .B2(
        \xmem_data[35][0] ), .ZN(n27721) );
  AOI22_X1 U31103 ( .A1(n27716), .A2(\xmem_data[36][0] ), .B1(n27715), .B2(
        \xmem_data[37][0] ), .ZN(n27720) );
  AOI22_X1 U31104 ( .A1(n27718), .A2(\xmem_data[38][0] ), .B1(n27717), .B2(
        \xmem_data[39][0] ), .ZN(n27719) );
  AOI22_X1 U31105 ( .A1(n28765), .A2(\xmem_data[40][0] ), .B1(n27723), .B2(
        \xmem_data[41][0] ), .ZN(n27726) );
  AOI22_X1 U31106 ( .A1(n27742), .A2(\xmem_data[42][0] ), .B1(n3149), .B2(
        \xmem_data[43][0] ), .ZN(n27725) );
  NAND2_X1 U31107 ( .A1(n27726), .A2(n27725), .ZN(n27727) );
  AOI22_X1 U31108 ( .A1(n29714), .A2(\xmem_data[56][0] ), .B1(n30301), .B2(
        \xmem_data[57][0] ), .ZN(n27734) );
  AOI22_X1 U31109 ( .A1(n27729), .A2(\xmem_data[58][0] ), .B1(n27455), .B2(
        \xmem_data[59][0] ), .ZN(n27733) );
  AOI22_X1 U31110 ( .A1(n3166), .A2(\xmem_data[60][0] ), .B1(n3187), .B2(
        \xmem_data[61][0] ), .ZN(n27732) );
  AND2_X1 U31111 ( .A1(n27825), .A2(\xmem_data[63][0] ), .ZN(n27730) );
  AOI21_X1 U31112 ( .B1(n29810), .B2(\xmem_data[62][0] ), .A(n27730), .ZN(
        n27731) );
  NAND4_X1 U31113 ( .A1(n27736), .A2(n3809), .A3(n27735), .A4(n3512), .ZN(
        n27738) );
  OAI21_X1 U31114 ( .B1(n27739), .B2(n27738), .A(n27737), .ZN(n27845) );
  NAND2_X1 U31115 ( .A1(n29790), .A2(\xmem_data[14][0] ), .ZN(n27752) );
  NAND2_X1 U31116 ( .A1(n29788), .A2(\xmem_data[12][0] ), .ZN(n27751) );
  AOI22_X1 U31117 ( .A1(n27742), .A2(\xmem_data[10][0] ), .B1(n3142), .B2(
        \xmem_data[11][0] ), .ZN(n27750) );
  AOI22_X1 U31118 ( .A1(n29419), .A2(\xmem_data[8][0] ), .B1(n27743), .B2(
        \xmem_data[9][0] ), .ZN(n27744) );
  INV_X1 U31119 ( .A(n27744), .ZN(n27748) );
  NAND2_X1 U31120 ( .A1(n26510), .A2(\xmem_data[13][0] ), .ZN(n27746) );
  NAND2_X1 U31121 ( .A1(n29565), .A2(\xmem_data[15][0] ), .ZN(n27745) );
  NAND2_X1 U31122 ( .A1(n27746), .A2(n27745), .ZN(n27747) );
  NOR2_X1 U31123 ( .A1(n27748), .A2(n27747), .ZN(n27749) );
  AOI22_X1 U31124 ( .A1(n30635), .A2(\xmem_data[24][0] ), .B1(n29768), .B2(
        \xmem_data[25][0] ), .ZN(n27760) );
  AOI22_X1 U31125 ( .A1(n27756), .A2(\xmem_data[26][0] ), .B1(n30303), .B2(
        \xmem_data[27][0] ), .ZN(n27759) );
  AOI22_X1 U31126 ( .A1(n3164), .A2(\xmem_data[28][0] ), .B1(n3189), .B2(
        \xmem_data[29][0] ), .ZN(n27758) );
  AOI22_X1 U31127 ( .A1(n30062), .A2(\xmem_data[30][0] ), .B1(n30617), .B2(
        \xmem_data[31][0] ), .ZN(n27757) );
  NAND4_X1 U31128 ( .A1(n27760), .A2(n27759), .A3(n27758), .A4(n27757), .ZN(
        n27769) );
  NAND2_X1 U31129 ( .A1(n30190), .A2(\xmem_data[21][0] ), .ZN(n27767) );
  AOI22_X1 U31130 ( .A1(n3223), .A2(\xmem_data[18][0] ), .B1(n3140), .B2(
        \xmem_data[19][0] ), .ZN(n27766) );
  AOI22_X1 U31131 ( .A1(n29500), .A2(\xmem_data[22][0] ), .B1(n27763), .B2(
        \xmem_data[23][0] ), .ZN(n27765) );
  NAND2_X1 U31132 ( .A1(n29647), .A2(\xmem_data[20][0] ), .ZN(n27764) );
  NAND4_X1 U31133 ( .A1(n27767), .A2(n27766), .A3(n27765), .A4(n27764), .ZN(
        n27768) );
  NOR2_X1 U31134 ( .A1(n27769), .A2(n27768), .ZN(n27777) );
  AOI22_X1 U31135 ( .A1(n27771), .A2(\xmem_data[16][0] ), .B1(n29495), .B2(
        \xmem_data[17][0] ), .ZN(n27776) );
  AOI22_X1 U31136 ( .A1(n30717), .A2(\xmem_data[0][0] ), .B1(n30765), .B2(
        \xmem_data[1][0] ), .ZN(n27775) );
  AOI22_X1 U31137 ( .A1(n7446), .A2(\xmem_data[2][0] ), .B1(n3151), .B2(
        \xmem_data[3][0] ), .ZN(n27774) );
  AOI22_X1 U31138 ( .A1(n29724), .A2(\xmem_data[4][0] ), .B1(n28696), .B2(
        \xmem_data[5][0] ), .ZN(n27773) );
  AOI22_X1 U31139 ( .A1(n29489), .A2(\xmem_data[6][0] ), .B1(n14982), .B2(
        \xmem_data[7][0] ), .ZN(n27772) );
  NAND4_X1 U31140 ( .A1(n3875), .A2(n27777), .A3(n27776), .A4(n3523), .ZN(
        n27779) );
  NAND2_X1 U31141 ( .A1(n27779), .A2(n27778), .ZN(n27844) );
  AOI22_X1 U31142 ( .A1(n27811), .A2(\xmem_data[120][0] ), .B1(n30249), .B2(
        \xmem_data[121][0] ), .ZN(n27785) );
  AOI22_X1 U31143 ( .A1(n3168), .A2(\xmem_data[124][0] ), .B1(n3183), .B2(
        \xmem_data[125][0] ), .ZN(n27784) );
  AOI22_X1 U31144 ( .A1(n3223), .A2(\xmem_data[114][0] ), .B1(n3146), .B2(
        \xmem_data[115][0] ), .ZN(n27782) );
  AOI22_X1 U31145 ( .A1(n27819), .A2(\xmem_data[122][0] ), .B1(n30892), .B2(
        \xmem_data[123][0] ), .ZN(n27781) );
  AOI22_X1 U31146 ( .A1(n29500), .A2(\xmem_data[118][0] ), .B1(n31353), .B2(
        \xmem_data[119][0] ), .ZN(n27780) );
  NAND3_X1 U31147 ( .A1(n27785), .A2(n27784), .A3(n27783), .ZN(n27788) );
  AOI22_X1 U31148 ( .A1(n23901), .A2(\xmem_data[126][0] ), .B1(n28781), .B2(
        \xmem_data[127][0] ), .ZN(n27786) );
  INV_X1 U31149 ( .A(n27786), .ZN(n27787) );
  NOR2_X1 U31150 ( .A1(n27788), .A2(n27787), .ZN(n27796) );
  AOI22_X1 U31151 ( .A1(n29488), .A2(\xmem_data[96][0] ), .B1(n29640), .B2(
        \xmem_data[97][0] ), .ZN(n27792) );
  AOI22_X1 U31152 ( .A1(n27804), .A2(\xmem_data[98][0] ), .B1(n28226), .B2(
        \xmem_data[99][0] ), .ZN(n27791) );
  AOI22_X1 U31153 ( .A1(n28725), .A2(\xmem_data[100][0] ), .B1(n27805), .B2(
        \xmem_data[101][0] ), .ZN(n27790) );
  AOI22_X1 U31154 ( .A1(n27806), .A2(\xmem_data[102][0] ), .B1(n27852), .B2(
        \xmem_data[103][0] ), .ZN(n27789) );
  AOI22_X1 U31155 ( .A1(n27834), .A2(\xmem_data[112][0] ), .B1(n3170), .B2(
        \xmem_data[113][0] ), .ZN(n27794) );
  AOI22_X1 U31156 ( .A1(\xmem_data[117][0] ), .A2(n28665), .B1(n3249), .B2(
        \xmem_data[116][0] ), .ZN(n27793) );
  AND2_X1 U31157 ( .A1(n27794), .A2(n27793), .ZN(n27795) );
  NAND3_X1 U31158 ( .A1(n27796), .A2(n3797), .A3(n27795), .ZN(n27803) );
  AOI22_X1 U31159 ( .A1(n7451), .A2(\xmem_data[104][0] ), .B1(n27812), .B2(
        \xmem_data[105][0] ), .ZN(n27800) );
  AOI22_X1 U31160 ( .A1(n27814), .A2(\xmem_data[106][0] ), .B1(n27813), .B2(
        \xmem_data[107][0] ), .ZN(n27799) );
  AOI22_X1 U31161 ( .A1(n27741), .A2(\xmem_data[108][0] ), .B1(n30775), .B2(
        \xmem_data[109][0] ), .ZN(n27798) );
  AOI22_X1 U31162 ( .A1(n3392), .A2(\xmem_data[110][0] ), .B1(n27831), .B2(
        \xmem_data[111][0] ), .ZN(n27797) );
  NAND4_X1 U31163 ( .A1(n27800), .A2(n27799), .A3(n27798), .A4(n27797), .ZN(
        n27802) );
  OAI21_X1 U31164 ( .B1(n27803), .B2(n27802), .A(n27801), .ZN(n27843) );
  AOI22_X1 U31165 ( .A1(n30198), .A2(\xmem_data[64][0] ), .B1(n29721), .B2(
        \xmem_data[65][0] ), .ZN(n27810) );
  AOI22_X1 U31166 ( .A1(n27804), .A2(\xmem_data[66][0] ), .B1(n31315), .B2(
        \xmem_data[67][0] ), .ZN(n27809) );
  AOI22_X1 U31167 ( .A1(n29819), .A2(\xmem_data[68][0] ), .B1(n27805), .B2(
        \xmem_data[69][0] ), .ZN(n27808) );
  AOI22_X1 U31168 ( .A1(n27806), .A2(\xmem_data[70][0] ), .B1(n20577), .B2(
        \xmem_data[71][0] ), .ZN(n27807) );
  AOI22_X1 U31169 ( .A1(n27754), .A2(\xmem_data[88][0] ), .B1(n30090), .B2(
        \xmem_data[89][0] ), .ZN(n27830) );
  AOI22_X1 U31170 ( .A1(n7451), .A2(\xmem_data[72][0] ), .B1(n27812), .B2(
        \xmem_data[73][0] ), .ZN(n27816) );
  AOI22_X1 U31171 ( .A1(n27814), .A2(\xmem_data[74][0] ), .B1(n27813), .B2(
        \xmem_data[75][0] ), .ZN(n27815) );
  NAND2_X1 U31172 ( .A1(n27816), .A2(n27815), .ZN(n27824) );
  AOI22_X1 U31173 ( .A1(n3223), .A2(\xmem_data[82][0] ), .B1(n3146), .B2(
        \xmem_data[83][0] ), .ZN(n27822) );
  AOI22_X1 U31174 ( .A1(n27819), .A2(\xmem_data[90][0] ), .B1(n21005), .B2(
        \xmem_data[91][0] ), .ZN(n27821) );
  AOI22_X1 U31175 ( .A1(n29500), .A2(\xmem_data[86][0] ), .B1(n20587), .B2(
        \xmem_data[87][0] ), .ZN(n27820) );
  AOI22_X1 U31176 ( .A1(n3167), .A2(\xmem_data[92][0] ), .B1(n3185), .B2(
        \xmem_data[93][0] ), .ZN(n27827) );
  AOI22_X1 U31177 ( .A1(n30715), .A2(\xmem_data[94][0] ), .B1(n27825), .B2(
        \xmem_data[95][0] ), .ZN(n27826) );
  NAND4_X1 U31178 ( .A1(n3839), .A2(n27830), .A3(n27829), .A4(n27828), .ZN(
        n27841) );
  AOI22_X1 U31179 ( .A1(n29628), .A2(\xmem_data[78][0] ), .B1(n27831), .B2(
        \xmem_data[79][0] ), .ZN(n27838) );
  AOI22_X1 U31180 ( .A1(n28734), .A2(\xmem_data[76][0] ), .B1(n27832), .B2(
        \xmem_data[77][0] ), .ZN(n27837) );
  AOI22_X1 U31181 ( .A1(n27834), .A2(\xmem_data[80][0] ), .B1(n27833), .B2(
        \xmem_data[81][0] ), .ZN(n27836) );
  AOI22_X1 U31182 ( .A1(n29705), .A2(\xmem_data[84][0] ), .B1(n3117), .B2(
        \xmem_data[85][0] ), .ZN(n27835) );
  NAND4_X1 U31183 ( .A1(n27838), .A2(n27837), .A3(n27836), .A4(n27835), .ZN(
        n27840) );
  OAI21_X1 U31184 ( .B1(n27841), .B2(n27840), .A(n27839), .ZN(n27842) );
  NAND4_X2 U31185 ( .A1(n27845), .A2(n27844), .A3(n27843), .A4(n27842), .ZN(
        n36316) );
  INV_X1 U31186 ( .A(n35642), .ZN(n27846) );
  AND2_X1 U31187 ( .A1(n36316), .A2(n27846), .ZN(n31141) );
  AOI22_X1 U31188 ( .A1(n28354), .A2(\xmem_data[28][1] ), .B1(n28317), .B2(
        \xmem_data[29][1] ), .ZN(n27854) );
  AND2_X1 U31189 ( .A1(n30900), .A2(\xmem_data[27][1] ), .ZN(n27851) );
  AOI22_X1 U31190 ( .A1(n27847), .A2(\xmem_data[24][1] ), .B1(n11008), .B2(
        \xmem_data[25][1] ), .ZN(n27849) );
  AOI22_X1 U31191 ( .A1(n3382), .A2(\xmem_data[30][1] ), .B1(n28501), .B2(
        \xmem_data[31][1] ), .ZN(n27848) );
  NAND2_X1 U31192 ( .A1(n27848), .A2(n27849), .ZN(n27850) );
  AOI211_X1 U31193 ( .C1(\xmem_data[26][1] ), .C2(n27852), .A(n27851), .B(
        n27850), .ZN(n27853) );
  NAND2_X1 U31194 ( .A1(n27853), .A2(n27854), .ZN(n27862) );
  AOI22_X1 U31195 ( .A1(n30949), .A2(\xmem_data[16][1] ), .B1(n28427), .B2(
        \xmem_data[17][1] ), .ZN(n27860) );
  AOI22_X1 U31196 ( .A1(n27855), .A2(\xmem_data[18][1] ), .B1(n29280), .B2(
        \xmem_data[19][1] ), .ZN(n27859) );
  AOI22_X1 U31197 ( .A1(n29240), .A2(\xmem_data[20][1] ), .B1(n21051), .B2(
        \xmem_data[21][1] ), .ZN(n27858) );
  AOI22_X1 U31198 ( .A1(n30269), .A2(\xmem_data[22][1] ), .B1(n27365), .B2(
        \xmem_data[23][1] ), .ZN(n27857) );
  NAND4_X1 U31199 ( .A1(n27860), .A2(n27859), .A3(n27858), .A4(n27857), .ZN(
        n27861) );
  AOI22_X1 U31200 ( .A1(n31276), .A2(\xmem_data[8][1] ), .B1(n27863), .B2(
        \xmem_data[9][1] ), .ZN(n27868) );
  AOI22_X1 U31201 ( .A1(n30744), .A2(\xmem_data[10][1] ), .B1(n24448), .B2(
        \xmem_data[11][1] ), .ZN(n27867) );
  AOI22_X1 U31202 ( .A1(n16986), .A2(\xmem_data[12][1] ), .B1(n30541), .B2(
        \xmem_data[13][1] ), .ZN(n27866) );
  AOI22_X1 U31203 ( .A1(n16988), .A2(\xmem_data[14][1] ), .B1(n27864), .B2(
        \xmem_data[15][1] ), .ZN(n27865) );
  NAND4_X1 U31204 ( .A1(n27868), .A2(n27867), .A3(n27866), .A4(n27865), .ZN(
        n27876) );
  AOI22_X1 U31205 ( .A1(n24694), .A2(\xmem_data[0][1] ), .B1(n3219), .B2(
        \xmem_data[1][1] ), .ZN(n27873) );
  AOI22_X1 U31206 ( .A1(n3322), .A2(\xmem_data[4][1] ), .B1(n30550), .B2(
        \xmem_data[5][1] ), .ZN(n27871) );
  AOI22_X1 U31207 ( .A1(n28367), .A2(\xmem_data[2][1] ), .B1(n27869), .B2(
        \xmem_data[3][1] ), .ZN(n27870) );
  NAND2_X1 U31208 ( .A1(n27873), .A2(n27872), .ZN(n27875) );
  AND2_X1 U31209 ( .A1(n3375), .A2(\xmem_data[6][1] ), .ZN(n27874) );
  AOI21_X1 U31210 ( .B1(n27879), .B2(n39020), .A(n27877), .ZN(n27881) );
  INV_X1 U31211 ( .A(n29103), .ZN(n27878) );
  NAND2_X1 U31212 ( .A1(n27879), .A2(n27878), .ZN(n27880) );
  NAND2_X1 U31213 ( .A1(n27881), .A2(n27880), .ZN(n27972) );
  AOI22_X1 U31214 ( .A1(n27902), .A2(\xmem_data[96][1] ), .B1(n3222), .B2(
        \xmem_data[97][1] ), .ZN(n27885) );
  AOI22_X1 U31215 ( .A1(n31368), .A2(\xmem_data[98][1] ), .B1(n25491), .B2(
        \xmem_data[99][1] ), .ZN(n27884) );
  AOI22_X1 U31216 ( .A1(n27904), .A2(\xmem_data[100][1] ), .B1(n27903), .B2(
        \xmem_data[101][1] ), .ZN(n27883) );
  AOI22_X1 U31217 ( .A1(n27905), .A2(\xmem_data[102][1] ), .B1(n28307), .B2(
        \xmem_data[103][1] ), .ZN(n27882) );
  NAND4_X1 U31218 ( .A1(n27885), .A2(n27884), .A3(n27883), .A4(n27882), .ZN(
        n27901) );
  AOI22_X1 U31219 ( .A1(n27910), .A2(\xmem_data[104][1] ), .B1(n3358), .B2(
        \xmem_data[105][1] ), .ZN(n27889) );
  AOI22_X1 U31220 ( .A1(n27911), .A2(\xmem_data[106][1] ), .B1(n24212), .B2(
        \xmem_data[107][1] ), .ZN(n27888) );
  AOI22_X1 U31221 ( .A1(n3176), .A2(\xmem_data[108][1] ), .B1(n27912), .B2(
        \xmem_data[109][1] ), .ZN(n27887) );
  AOI22_X1 U31222 ( .A1(n31328), .A2(\xmem_data[110][1] ), .B1(n29279), .B2(
        \xmem_data[111][1] ), .ZN(n27886) );
  NAND4_X1 U31223 ( .A1(n27889), .A2(n27888), .A3(n27887), .A4(n27886), .ZN(
        n27900) );
  AOI22_X1 U31224 ( .A1(n27919), .A2(\xmem_data[112][1] ), .B1(n27918), .B2(
        \xmem_data[113][1] ), .ZN(n27893) );
  AOI22_X1 U31225 ( .A1(n20815), .A2(\xmem_data[114][1] ), .B1(n27920), .B2(
        \xmem_data[115][1] ), .ZN(n27892) );
  AOI22_X1 U31226 ( .A1(n3177), .A2(\xmem_data[116][1] ), .B1(n25581), .B2(
        \xmem_data[117][1] ), .ZN(n27891) );
  AOI22_X1 U31227 ( .A1(n3308), .A2(\xmem_data[118][1] ), .B1(n28098), .B2(
        \xmem_data[119][1] ), .ZN(n27890) );
  NAND4_X1 U31228 ( .A1(n27893), .A2(n27892), .A3(n27891), .A4(n27890), .ZN(
        n27899) );
  AOI22_X1 U31229 ( .A1(n21058), .A2(\xmem_data[120][1] ), .B1(n25527), .B2(
        \xmem_data[121][1] ), .ZN(n27897) );
  AOI22_X1 U31230 ( .A1(n20826), .A2(\xmem_data[122][1] ), .B1(n20707), .B2(
        \xmem_data[123][1] ), .ZN(n27896) );
  AOI22_X1 U31231 ( .A1(n27925), .A2(\xmem_data[124][1] ), .B1(n27499), .B2(
        \xmem_data[125][1] ), .ZN(n27895) );
  AOI22_X1 U31232 ( .A1(n16980), .A2(\xmem_data[126][1] ), .B1(n31347), .B2(
        \xmem_data[127][1] ), .ZN(n27894) );
  NAND4_X1 U31233 ( .A1(n27897), .A2(n27896), .A3(n27895), .A4(n27894), .ZN(
        n27898) );
  OR4_X1 U31234 ( .A1(n27901), .A2(n27900), .A3(n27899), .A4(n27898), .ZN(
        n27936) );
  AOI22_X1 U31235 ( .A1(n27902), .A2(\xmem_data[64][1] ), .B1(n3219), .B2(
        \xmem_data[65][1] ), .ZN(n27909) );
  AOI22_X1 U31236 ( .A1(n25448), .A2(\xmem_data[66][1] ), .B1(n25562), .B2(
        \xmem_data[67][1] ), .ZN(n27908) );
  AOI22_X1 U31237 ( .A1(n27904), .A2(\xmem_data[68][1] ), .B1(n27903), .B2(
        \xmem_data[69][1] ), .ZN(n27907) );
  AOI22_X1 U31238 ( .A1(n27905), .A2(\xmem_data[70][1] ), .B1(n28045), .B2(
        \xmem_data[71][1] ), .ZN(n27906) );
  NAND4_X1 U31239 ( .A1(n27909), .A2(n27908), .A3(n27907), .A4(n27906), .ZN(
        n27933) );
  AOI22_X1 U31240 ( .A1(n27910), .A2(\xmem_data[72][1] ), .B1(n25481), .B2(
        \xmem_data[73][1] ), .ZN(n27917) );
  AOI22_X1 U31241 ( .A1(n27911), .A2(\xmem_data[74][1] ), .B1(n24212), .B2(
        \xmem_data[75][1] ), .ZN(n27916) );
  AOI22_X1 U31242 ( .A1(n3176), .A2(\xmem_data[76][1] ), .B1(n27912), .B2(
        \xmem_data[77][1] ), .ZN(n27915) );
  AOI22_X1 U31243 ( .A1(n28516), .A2(\xmem_data[78][1] ), .B1(n27864), .B2(
        \xmem_data[79][1] ), .ZN(n27914) );
  NAND4_X1 U31244 ( .A1(n27917), .A2(n27916), .A3(n27915), .A4(n27914), .ZN(
        n27932) );
  AOI22_X1 U31245 ( .A1(n27919), .A2(\xmem_data[80][1] ), .B1(n27918), .B2(
        \xmem_data[81][1] ), .ZN(n27924) );
  AOI22_X1 U31246 ( .A1(n25400), .A2(\xmem_data[82][1] ), .B1(n27920), .B2(
        \xmem_data[83][1] ), .ZN(n27923) );
  AOI22_X1 U31247 ( .A1(n24647), .A2(\xmem_data[84][1] ), .B1(n28429), .B2(
        \xmem_data[85][1] ), .ZN(n27922) );
  AOI22_X1 U31248 ( .A1(n29816), .A2(\xmem_data[86][1] ), .B1(n28495), .B2(
        \xmem_data[87][1] ), .ZN(n27921) );
  NAND4_X1 U31249 ( .A1(n27924), .A2(n27923), .A3(n27922), .A4(n27921), .ZN(
        n27931) );
  AOI22_X1 U31250 ( .A1(n30497), .A2(\xmem_data[88][1] ), .B1(n25359), .B2(
        \xmem_data[89][1] ), .ZN(n27929) );
  AOI22_X1 U31251 ( .A1(n24687), .A2(\xmem_data[90][1] ), .B1(n27567), .B2(
        \xmem_data[91][1] ), .ZN(n27928) );
  AOI22_X1 U31252 ( .A1(n27925), .A2(\xmem_data[92][1] ), .B1(n30861), .B2(
        \xmem_data[93][1] ), .ZN(n27927) );
  AOI22_X1 U31253 ( .A1(n28039), .A2(\xmem_data[94][1] ), .B1(n27437), .B2(
        \xmem_data[95][1] ), .ZN(n27926) );
  NAND4_X1 U31254 ( .A1(n27929), .A2(n27928), .A3(n27927), .A4(n27926), .ZN(
        n27930) );
  OR4_X1 U31255 ( .A1(n27933), .A2(n27932), .A3(n27931), .A4(n27930), .ZN(
        n27934) );
  AOI22_X1 U31256 ( .A1(n27937), .A2(n27936), .B1(n27935), .B2(n27934), .ZN(
        n27971) );
  AOI22_X1 U31257 ( .A1(n25354), .A2(\xmem_data[32][1] ), .B1(n3221), .B2(
        \xmem_data[33][1] ), .ZN(n27942) );
  AOI22_X1 U31258 ( .A1(n22708), .A2(\xmem_data[34][1] ), .B1(n25491), .B2(
        \xmem_data[35][1] ), .ZN(n27941) );
  AOI22_X1 U31259 ( .A1(n27938), .A2(\xmem_data[36][1] ), .B1(n3256), .B2(
        \xmem_data[37][1] ), .ZN(n27940) );
  AOI22_X1 U31260 ( .A1(n16973), .A2(\xmem_data[38][1] ), .B1(n27446), .B2(
        \xmem_data[39][1] ), .ZN(n27939) );
  NAND4_X1 U31261 ( .A1(n27942), .A2(n27941), .A3(n27940), .A4(n27939), .ZN(
        n27967) );
  AOI22_X1 U31262 ( .A1(n25422), .A2(\xmem_data[40][1] ), .B1(n20546), .B2(
        \xmem_data[41][1] ), .ZN(n27949) );
  AOI22_X1 U31263 ( .A1(n27944), .A2(\xmem_data[42][1] ), .B1(n24212), .B2(
        \xmem_data[43][1] ), .ZN(n27948) );
  AOI22_X1 U31264 ( .A1(n30891), .A2(\xmem_data[44][1] ), .B1(n25572), .B2(
        \xmem_data[45][1] ), .ZN(n27947) );
  AOI22_X1 U31265 ( .A1(n29437), .A2(\xmem_data[46][1] ), .B1(n23716), .B2(
        \xmem_data[47][1] ), .ZN(n27946) );
  NAND4_X1 U31266 ( .A1(n27949), .A2(n27948), .A3(n27947), .A4(n27946), .ZN(
        n27966) );
  AOI22_X1 U31267 ( .A1(n28337), .A2(\xmem_data[48][1] ), .B1(n25398), .B2(
        \xmem_data[49][1] ), .ZN(n27956) );
  AOI22_X1 U31268 ( .A1(n28994), .A2(\xmem_data[50][1] ), .B1(n27950), .B2(
        \xmem_data[51][1] ), .ZN(n27955) );
  AOI22_X1 U31269 ( .A1(n27952), .A2(\xmem_data[52][1] ), .B1(n27951), .B2(
        \xmem_data[53][1] ), .ZN(n27954) );
  AOI22_X1 U31270 ( .A1(n20732), .A2(\xmem_data[54][1] ), .B1(n24167), .B2(
        \xmem_data[55][1] ), .ZN(n27953) );
  NAND4_X1 U31271 ( .A1(n27956), .A2(n27955), .A3(n27954), .A4(n27953), .ZN(
        n27965) );
  AOI22_X1 U31272 ( .A1(n3179), .A2(\xmem_data[56][1] ), .B1(n28500), .B2(
        \xmem_data[57][1] ), .ZN(n27963) );
  AOI22_X1 U31273 ( .A1(n31345), .A2(\xmem_data[58][1] ), .B1(n27957), .B2(
        \xmem_data[59][1] ), .ZN(n27962) );
  AOI22_X1 U31274 ( .A1(n27959), .A2(\xmem_data[60][1] ), .B1(n27958), .B2(
        \xmem_data[61][1] ), .ZN(n27961) );
  AOI22_X1 U31275 ( .A1(n25725), .A2(\xmem_data[62][1] ), .B1(n23731), .B2(
        \xmem_data[63][1] ), .ZN(n27960) );
  NAND4_X1 U31276 ( .A1(n27963), .A2(n27962), .A3(n27961), .A4(n27960), .ZN(
        n27964) );
  OR4_X1 U31277 ( .A1(n27967), .A2(n27966), .A3(n27965), .A4(n27964), .ZN(
        n27969) );
  NAND2_X1 U31278 ( .A1(n27969), .A2(n27968), .ZN(n27970) );
  XNOR2_X1 U31279 ( .A(n32165), .B(\fmem_data[2][5] ), .ZN(n34036) );
  XNOR2_X1 U31280 ( .A(n32787), .B(\fmem_data[2][5] ), .ZN(n32286) );
  OAI22_X1 U31281 ( .A1(n34036), .A2(n35019), .B1(n32286), .B2(n35018), .ZN(
        n30430) );
  XNOR2_X1 U31282 ( .A(n35106), .B(\fmem_data[26][1] ), .ZN(n32752) );
  XNOR2_X1 U31283 ( .A(n31670), .B(\fmem_data[26][1] ), .ZN(n32164) );
  AOI22_X1 U31284 ( .A1(n24708), .A2(\xmem_data[24][1] ), .B1(n28492), .B2(
        \xmem_data[25][1] ), .ZN(n27980) );
  AOI22_X1 U31285 ( .A1(n29639), .A2(\xmem_data[26][1] ), .B1(n24116), .B2(
        \xmem_data[27][1] ), .ZN(n27979) );
  AOI22_X1 U31286 ( .A1(n27974), .A2(\xmem_data[28][1] ), .B1(n28462), .B2(
        \xmem_data[29][1] ), .ZN(n27978) );
  AOI22_X1 U31287 ( .A1(n3330), .A2(\xmem_data[30][1] ), .B1(n27975), .B2(
        \xmem_data[31][1] ), .ZN(n27977) );
  NAND4_X1 U31288 ( .A1(n27980), .A2(n27979), .A3(n27978), .A4(n27977), .ZN(
        n27987) );
  AOI22_X1 U31289 ( .A1(n24685), .A2(\xmem_data[0][1] ), .B1(n27981), .B2(
        \xmem_data[1][1] ), .ZN(n27985) );
  AOI22_X1 U31290 ( .A1(n30674), .A2(\xmem_data[2][1] ), .B1(n31261), .B2(
        \xmem_data[3][1] ), .ZN(n27984) );
  AOI22_X1 U31291 ( .A1(n28354), .A2(\xmem_data[4][1] ), .B1(n28075), .B2(
        \xmem_data[5][1] ), .ZN(n27983) );
  AOI22_X1 U31292 ( .A1(n3228), .A2(\xmem_data[6][1] ), .B1(n27437), .B2(
        \xmem_data[7][1] ), .ZN(n27982) );
  NAND4_X1 U31293 ( .A1(n27985), .A2(n27984), .A3(n27983), .A4(n27982), .ZN(
        n27986) );
  OR2_X1 U31294 ( .A1(n27987), .A2(n27986), .ZN(n28004) );
  AOI22_X1 U31295 ( .A1(n20809), .A2(\xmem_data[16][1] ), .B1(n27988), .B2(
        \xmem_data[17][1] ), .ZN(n27993) );
  AOI22_X1 U31296 ( .A1(n29451), .A2(\xmem_data[18][1] ), .B1(n28416), .B2(
        \xmem_data[19][1] ), .ZN(n27992) );
  AOI22_X1 U31297 ( .A1(n3176), .A2(\xmem_data[20][1] ), .B1(n22703), .B2(
        \xmem_data[21][1] ), .ZN(n27991) );
  AOI22_X1 U31298 ( .A1(n29605), .A2(\xmem_data[22][1] ), .B1(n27989), .B2(
        \xmem_data[23][1] ), .ZN(n27990) );
  AOI22_X1 U31299 ( .A1(n25490), .A2(\xmem_data[12][1] ), .B1(n27994), .B2(
        \xmem_data[13][1] ), .ZN(n27996) );
  NAND2_X1 U31300 ( .A1(n28344), .A2(\xmem_data[14][1] ), .ZN(n27995) );
  NAND2_X1 U31301 ( .A1(n27996), .A2(n27995), .ZN(n28001) );
  AOI22_X1 U31302 ( .A1(n28355), .A2(\xmem_data[8][1] ), .B1(n3221), .B2(
        \xmem_data[9][1] ), .ZN(n27997) );
  INV_X1 U31303 ( .A(n27997), .ZN(n28000) );
  AOI22_X1 U31304 ( .A1(n29422), .A2(\xmem_data[10][1] ), .B1(n25562), .B2(
        \xmem_data[11][1] ), .ZN(n27998) );
  INV_X1 U31305 ( .A(n27998), .ZN(n27999) );
  NOR3_X1 U31306 ( .A1(n28001), .A2(n28000), .A3(n27999), .ZN(n28002) );
  NAND2_X1 U31307 ( .A1(n3817), .A2(n28002), .ZN(n28003) );
  NOR2_X1 U31308 ( .A1(n28004), .A2(n28003), .ZN(n28005) );
  NOR2_X1 U31309 ( .A1(n28005), .A2(n24043), .ZN(n28009) );
  NOR2_X1 U31310 ( .A1(n24043), .A2(n39016), .ZN(n28006) );
  AND2_X1 U31311 ( .A1(n23771), .A2(n28006), .ZN(n28008) );
  NOR2_X1 U31312 ( .A1(n28009), .A2(n28008), .ZN(n34589) );
  AOI22_X1 U31313 ( .A1(n24572), .A2(\xmem_data[64][1] ), .B1(n27526), .B2(
        \xmem_data[65][1] ), .ZN(n28013) );
  AOI22_X1 U31314 ( .A1(n28036), .A2(\xmem_data[66][1] ), .B1(n28035), .B2(
        \xmem_data[67][1] ), .ZN(n28012) );
  AOI22_X1 U31315 ( .A1(n28038), .A2(\xmem_data[68][1] ), .B1(n28037), .B2(
        \xmem_data[69][1] ), .ZN(n28011) );
  AOI22_X1 U31316 ( .A1(n28039), .A2(\xmem_data[70][1] ), .B1(n24439), .B2(
        \xmem_data[71][1] ), .ZN(n28010) );
  NAND4_X1 U31317 ( .A1(n28013), .A2(n28012), .A3(n28011), .A4(n28010), .ZN(
        n28032) );
  AOI22_X1 U31318 ( .A1(n28044), .A2(\xmem_data[72][1] ), .B1(n3222), .B2(
        \xmem_data[73][1] ), .ZN(n28020) );
  AOI22_X1 U31319 ( .A1(n29288), .A2(\xmem_data[74][1] ), .B1(n30534), .B2(
        \xmem_data[75][1] ), .ZN(n28015) );
  AOI22_X1 U31320 ( .A1(n14991), .A2(\xmem_data[78][1] ), .B1(n14928), .B2(
        \xmem_data[79][1] ), .ZN(n28014) );
  NAND2_X1 U31321 ( .A1(n28015), .A2(n28014), .ZN(n28018) );
  AOI22_X1 U31322 ( .A1(n24141), .A2(\xmem_data[76][1] ), .B1(n13444), .B2(
        \xmem_data[77][1] ), .ZN(n28016) );
  INV_X1 U31323 ( .A(n28016), .ZN(n28017) );
  NOR2_X1 U31324 ( .A1(n28018), .A2(n28017), .ZN(n28019) );
  NAND2_X1 U31325 ( .A1(n28020), .A2(n28019), .ZN(n28031) );
  AOI22_X1 U31326 ( .A1(n28050), .A2(\xmem_data[80][1] ), .B1(n27943), .B2(
        \xmem_data[81][1] ), .ZN(n28024) );
  AOI22_X1 U31327 ( .A1(n28051), .A2(\xmem_data[82][1] ), .B1(n24132), .B2(
        \xmem_data[83][1] ), .ZN(n28023) );
  AOI22_X1 U31328 ( .A1(n28298), .A2(\xmem_data[84][1] ), .B1(n28052), .B2(
        \xmem_data[85][1] ), .ZN(n28022) );
  AOI22_X1 U31329 ( .A1(n31354), .A2(\xmem_data[86][1] ), .B1(n28993), .B2(
        \xmem_data[87][1] ), .ZN(n28021) );
  NAND4_X1 U31330 ( .A1(n28024), .A2(n28023), .A3(n28022), .A4(n28021), .ZN(
        n28030) );
  AOI22_X1 U31331 ( .A1(n28059), .A2(\xmem_data[88][1] ), .B1(n28058), .B2(
        \xmem_data[89][1] ), .ZN(n28028) );
  AOI22_X1 U31332 ( .A1(n28302), .A2(\xmem_data[90][1] ), .B1(n29318), .B2(
        \xmem_data[91][1] ), .ZN(n28027) );
  AOI22_X1 U31333 ( .A1(n28061), .A2(\xmem_data[92][1] ), .B1(n28060), .B2(
        \xmem_data[93][1] ), .ZN(n28026) );
  AOI22_X1 U31334 ( .A1(n23780), .A2(\xmem_data[94][1] ), .B1(n28062), .B2(
        \xmem_data[95][1] ), .ZN(n28025) );
  NAND4_X1 U31335 ( .A1(n28028), .A2(n28027), .A3(n28026), .A4(n28025), .ZN(
        n28029) );
  OR4_X1 U31336 ( .A1(n28032), .A2(n28031), .A3(n28030), .A4(n28029), .ZN(
        n28034) );
  NAND2_X1 U31337 ( .A1(n28034), .A2(n28033), .ZN(n28074) );
  AOI22_X1 U31338 ( .A1(n20782), .A2(\xmem_data[96][1] ), .B1(n29136), .B2(
        \xmem_data[97][1] ), .ZN(n28043) );
  AOI22_X1 U31339 ( .A1(n28036), .A2(\xmem_data[98][1] ), .B1(n28035), .B2(
        \xmem_data[99][1] ), .ZN(n28042) );
  AOI22_X1 U31340 ( .A1(n28038), .A2(\xmem_data[100][1] ), .B1(n28037), .B2(
        \xmem_data[101][1] ), .ZN(n28041) );
  AOI22_X1 U31341 ( .A1(n28039), .A2(\xmem_data[102][1] ), .B1(n29286), .B2(
        \xmem_data[103][1] ), .ZN(n28040) );
  NAND4_X1 U31342 ( .A1(n28043), .A2(n28042), .A3(n28041), .A4(n28040), .ZN(
        n28070) );
  AOI22_X1 U31343 ( .A1(n28044), .A2(\xmem_data[104][1] ), .B1(n3221), .B2(
        \xmem_data[105][1] ), .ZN(n28049) );
  AOI22_X1 U31344 ( .A1(n17033), .A2(\xmem_data[106][1] ), .B1(n29028), .B2(
        \xmem_data[107][1] ), .ZN(n28048) );
  AOI22_X1 U31345 ( .A1(n24697), .A2(\xmem_data[108][1] ), .B1(n17061), .B2(
        \xmem_data[109][1] ), .ZN(n28047) );
  AOI22_X1 U31346 ( .A1(n20808), .A2(\xmem_data[110][1] ), .B1(n25450), .B2(
        \xmem_data[111][1] ), .ZN(n28046) );
  NAND4_X1 U31347 ( .A1(n28049), .A2(n28048), .A3(n28047), .A4(n28046), .ZN(
        n28069) );
  AOI22_X1 U31348 ( .A1(n28050), .A2(\xmem_data[112][1] ), .B1(n3358), .B2(
        \xmem_data[113][1] ), .ZN(n28057) );
  AOI22_X1 U31349 ( .A1(n28051), .A2(\xmem_data[114][1] ), .B1(n28416), .B2(
        \xmem_data[115][1] ), .ZN(n28056) );
  AOI22_X1 U31350 ( .A1(n30891), .A2(\xmem_data[116][1] ), .B1(n28052), .B2(
        \xmem_data[117][1] ), .ZN(n28055) );
  AOI22_X1 U31351 ( .A1(n27517), .A2(\xmem_data[118][1] ), .B1(n30615), .B2(
        \xmem_data[119][1] ), .ZN(n28054) );
  NAND4_X1 U31352 ( .A1(n28057), .A2(n28056), .A3(n28055), .A4(n28054), .ZN(
        n28068) );
  AOI22_X1 U31353 ( .A1(n28059), .A2(\xmem_data[120][1] ), .B1(n28058), .B2(
        \xmem_data[121][1] ), .ZN(n28066) );
  AOI22_X1 U31354 ( .A1(n20942), .A2(\xmem_data[122][1] ), .B1(n23801), .B2(
        \xmem_data[123][1] ), .ZN(n28065) );
  AOI22_X1 U31355 ( .A1(n28061), .A2(\xmem_data[124][1] ), .B1(n28060), .B2(
        \xmem_data[125][1] ), .ZN(n28064) );
  AOI22_X1 U31356 ( .A1(n24571), .A2(\xmem_data[126][1] ), .B1(n28062), .B2(
        \xmem_data[127][1] ), .ZN(n28063) );
  NAND4_X1 U31357 ( .A1(n28066), .A2(n28065), .A3(n28064), .A4(n28063), .ZN(
        n28067) );
  OR4_X1 U31358 ( .A1(n28070), .A2(n28069), .A3(n28068), .A4(n28067), .ZN(
        n28072) );
  NAND2_X1 U31359 ( .A1(n28072), .A2(n28071), .ZN(n28073) );
  NAND2_X1 U31360 ( .A1(n28074), .A2(n28073), .ZN(n28109) );
  AOI22_X1 U31361 ( .A1(n24467), .A2(\xmem_data[32][1] ), .B1(n20488), .B2(
        \xmem_data[33][1] ), .ZN(n28081) );
  AOI22_X1 U31362 ( .A1(n30901), .A2(\xmem_data[34][1] ), .B1(n27435), .B2(
        \xmem_data[35][1] ), .ZN(n28080) );
  AOI22_X1 U31363 ( .A1(n28076), .A2(\xmem_data[36][1] ), .B1(n28075), .B2(
        \xmem_data[37][1] ), .ZN(n28079) );
  AOI22_X1 U31364 ( .A1(n3434), .A2(\xmem_data[38][1] ), .B1(n3247), .B2(
        \xmem_data[39][1] ), .ZN(n28078) );
  NAND4_X1 U31365 ( .A1(n28081), .A2(n28080), .A3(n28079), .A4(n28078), .ZN(
        n28106) );
  AOI22_X1 U31366 ( .A1(n28082), .A2(\xmem_data[40][1] ), .B1(n3221), .B2(
        \xmem_data[41][1] ), .ZN(n28088) );
  AOI22_X1 U31367 ( .A1(n22708), .A2(\xmem_data[42][1] ), .B1(n25509), .B2(
        \xmem_data[43][1] ), .ZN(n28087) );
  AOI22_X1 U31368 ( .A1(n28083), .A2(\xmem_data[44][1] ), .B1(n27550), .B2(
        \xmem_data[45][1] ), .ZN(n28086) );
  AOI22_X1 U31369 ( .A1(n28084), .A2(\xmem_data[46][1] ), .B1(n25514), .B2(
        \xmem_data[47][1] ), .ZN(n28085) );
  NAND4_X1 U31370 ( .A1(n28088), .A2(n28087), .A3(n28086), .A4(n28085), .ZN(
        n28105) );
  AOI22_X1 U31371 ( .A1(n27551), .A2(\xmem_data[48][1] ), .B1(n13475), .B2(
        \xmem_data[49][1] ), .ZN(n28095) );
  AOI22_X1 U31372 ( .A1(n28089), .A2(\xmem_data[50][1] ), .B1(n24448), .B2(
        \xmem_data[51][1] ), .ZN(n28094) );
  AOI22_X1 U31373 ( .A1(n30514), .A2(\xmem_data[52][1] ), .B1(n28090), .B2(
        \xmem_data[53][1] ), .ZN(n28093) );
  AOI22_X1 U31374 ( .A1(n29807), .A2(\xmem_data[54][1] ), .B1(n24457), .B2(
        \xmem_data[55][1] ), .ZN(n28092) );
  NAND4_X1 U31375 ( .A1(n28095), .A2(n28094), .A3(n28093), .A4(n28092), .ZN(
        n28104) );
  AOI22_X1 U31376 ( .A1(n28096), .A2(\xmem_data[56][1] ), .B1(n31329), .B2(
        \xmem_data[57][1] ), .ZN(n28102) );
  AOI22_X1 U31377 ( .A1(n24710), .A2(\xmem_data[58][1] ), .B1(n28097), .B2(
        \xmem_data[59][1] ), .ZN(n28101) );
  AOI22_X1 U31378 ( .A1(n24511), .A2(\xmem_data[60][1] ), .B1(n23778), .B2(
        \xmem_data[61][1] ), .ZN(n28100) );
  AOI22_X1 U31379 ( .A1(n3301), .A2(\xmem_data[62][1] ), .B1(n28098), .B2(
        \xmem_data[63][1] ), .ZN(n28099) );
  NAND4_X1 U31380 ( .A1(n28102), .A2(n28101), .A3(n28100), .A4(n28099), .ZN(
        n28103) );
  OR4_X1 U31381 ( .A1(n28106), .A2(n28105), .A3(n28104), .A4(n28103), .ZN(
        n28108) );
  NAND2_X1 U31382 ( .A1(n34589), .A2(n34588), .ZN(n31946) );
  XNOR2_X1 U31383 ( .A(n31946), .B(\fmem_data[22][5] ), .ZN(n32080) );
  XNOR2_X1 U31384 ( .A(n32124), .B(\fmem_data[22][5] ), .ZN(n33962) );
  OAI22_X1 U31385 ( .A1(n32080), .A2(n33961), .B1(n33962), .B2(n33963), .ZN(
        n31214) );
  AOI22_X1 U31386 ( .A1(n30076), .A2(\xmem_data[100][0] ), .B1(n30765), .B2(
        \xmem_data[101][0] ), .ZN(n28124) );
  AOI22_X1 U31387 ( .A1(n29769), .A2(\xmem_data[124][0] ), .B1(n30193), .B2(
        \xmem_data[125][0] ), .ZN(n28123) );
  AOI22_X1 U31388 ( .A1(n3161), .A2(\xmem_data[96][0] ), .B1(n3190), .B2(
        \xmem_data[97][0] ), .ZN(n28122) );
  AOI22_X1 U31389 ( .A1(n28240), .A2(\xmem_data[104][0] ), .B1(n28239), .B2(
        \xmem_data[105][0] ), .ZN(n28115) );
  AOI22_X1 U31390 ( .A1(n28242), .A2(\xmem_data[106][0] ), .B1(n28241), .B2(
        \xmem_data[107][0] ), .ZN(n28114) );
  AOI22_X1 U31391 ( .A1(n28244), .A2(\xmem_data[108][0] ), .B1(n28243), .B2(
        \xmem_data[109][0] ), .ZN(n28113) );
  AOI22_X1 U31392 ( .A1(n28111), .A2(\xmem_data[110][0] ), .B1(n28245), .B2(
        \xmem_data[111][0] ), .ZN(n28112) );
  NAND4_X1 U31393 ( .A1(n28115), .A2(n28114), .A3(n28113), .A4(n28112), .ZN(
        n28120) );
  AOI22_X1 U31394 ( .A1(n3233), .A2(\xmem_data[102][0] ), .B1(n28226), .B2(
        \xmem_data[103][0] ), .ZN(n28118) );
  AOI22_X1 U31395 ( .A1(n3241), .A2(\xmem_data[122][0] ), .B1(n28233), .B2(
        \xmem_data[123][0] ), .ZN(n28117) );
  AOI22_X1 U31396 ( .A1(n3240), .A2(\xmem_data[126][0] ), .B1(n28231), .B2(
        \xmem_data[127][0] ), .ZN(n28116) );
  NAND3_X1 U31397 ( .A1(n28118), .A2(n28117), .A3(n28116), .ZN(n28119) );
  NOR2_X1 U31398 ( .A1(n28120), .A2(n28119), .ZN(n28121) );
  NAND4_X1 U31399 ( .A1(n28124), .A2(n28123), .A3(n28122), .A4(n28121), .ZN(
        n28128) );
  AOI22_X1 U31400 ( .A1(n29801), .A2(\xmem_data[120][0] ), .B1(n28145), .B2(
        \xmem_data[121][0] ), .ZN(n28126) );
  AOI22_X1 U31401 ( .A1(n30684), .A2(\xmem_data[98][0] ), .B1(n28232), .B2(
        \xmem_data[99][0] ), .ZN(n28125) );
  NAND2_X1 U31402 ( .A1(n28126), .A2(n28125), .ZN(n28127) );
  OR2_X1 U31403 ( .A1(n28128), .A2(n28127), .ZN(n28135) );
  AOI22_X1 U31404 ( .A1(n27710), .A2(\xmem_data[112][0] ), .B1(n30775), .B2(
        \xmem_data[113][0] ), .ZN(n28132) );
  AOI22_X1 U31405 ( .A1(n27740), .A2(\xmem_data[114][0] ), .B1(n28218), .B2(
        \xmem_data[115][0] ), .ZN(n28131) );
  AOI22_X1 U31406 ( .A1(n28219), .A2(\xmem_data[116][0] ), .B1(n29495), .B2(
        \xmem_data[117][0] ), .ZN(n28130) );
  AOI22_X1 U31407 ( .A1(n28220), .A2(\xmem_data[118][0] ), .B1(n30698), .B2(
        \xmem_data[119][0] ), .ZN(n28129) );
  NAND4_X1 U31408 ( .A1(n28132), .A2(n28131), .A3(n28130), .A4(n28129), .ZN(
        n28134) );
  AOI22_X1 U31409 ( .A1(n29421), .A2(\xmem_data[48][0] ), .B1(n28766), .B2(
        \xmem_data[49][0] ), .ZN(n28144) );
  AOI22_X1 U31410 ( .A1(n27740), .A2(\xmem_data[50][0] ), .B1(n28137), .B2(
        \xmem_data[51][0] ), .ZN(n28143) );
  AOI22_X1 U31411 ( .A1(n28139), .A2(\xmem_data[52][0] ), .B1(n29761), .B2(
        \xmem_data[53][0] ), .ZN(n28142) );
  AOI22_X1 U31412 ( .A1(n28140), .A2(\xmem_data[54][0] ), .B1(n24702), .B2(
        \xmem_data[55][0] ), .ZN(n28141) );
  NAND4_X1 U31413 ( .A1(n28144), .A2(n28143), .A3(n28142), .A4(n28141), .ZN(
        n28179) );
  AOI22_X1 U31414 ( .A1(n29590), .A2(\xmem_data[56][0] ), .B1(n29589), .B2(
        \xmem_data[57][0] ), .ZN(n28149) );
  AOI22_X1 U31415 ( .A1(n29476), .A2(\xmem_data[34][0] ), .B1(n28147), .B2(
        \xmem_data[35][0] ), .ZN(n28148) );
  AOI22_X1 U31416 ( .A1(n3162), .A2(\xmem_data[32][0] ), .B1(n3187), .B2(
        \xmem_data[33][0] ), .ZN(n28150) );
  INV_X1 U31417 ( .A(n28150), .ZN(n28172) );
  AOI22_X1 U31418 ( .A1(n28151), .A2(\xmem_data[38][0] ), .B1(n29246), .B2(
        \xmem_data[39][0] ), .ZN(n28158) );
  AOI22_X1 U31419 ( .A1(n28153), .A2(\xmem_data[58][0] ), .B1(n28152), .B2(
        \xmem_data[59][0] ), .ZN(n28157) );
  AOI22_X1 U31420 ( .A1(n28155), .A2(\xmem_data[62][0] ), .B1(n28154), .B2(
        \xmem_data[63][0] ), .ZN(n28156) );
  NAND3_X1 U31421 ( .A1(n28158), .A2(n28157), .A3(n28156), .ZN(n28171) );
  AOI22_X1 U31422 ( .A1(n28160), .A2(\xmem_data[40][0] ), .B1(n28159), .B2(
        \xmem_data[41][0] ), .ZN(n28169) );
  AOI22_X1 U31423 ( .A1(n28161), .A2(\xmem_data[42][0] ), .B1(n23730), .B2(
        \xmem_data[43][0] ), .ZN(n28168) );
  AOI22_X1 U31424 ( .A1(n28163), .A2(\xmem_data[44][0] ), .B1(n28162), .B2(
        \xmem_data[45][0] ), .ZN(n28167) );
  AOI22_X1 U31425 ( .A1(n28165), .A2(\xmem_data[46][0] ), .B1(n28164), .B2(
        \xmem_data[47][0] ), .ZN(n28166) );
  NAND4_X1 U31426 ( .A1(n28169), .A2(n28168), .A3(n28167), .A4(n28166), .ZN(
        n28170) );
  NOR3_X1 U31427 ( .A1(n28172), .A2(n28171), .A3(n28170), .ZN(n28176) );
  AOI22_X1 U31428 ( .A1(n29547), .A2(\xmem_data[36][0] ), .B1(n30765), .B2(
        \xmem_data[37][0] ), .ZN(n28175) );
  AOI22_X1 U31429 ( .A1(n27754), .A2(\xmem_data[60][0] ), .B1(n28684), .B2(
        \xmem_data[61][0] ), .ZN(n28174) );
  NAND4_X1 U31430 ( .A1(n3942), .A2(n28176), .A3(n28175), .A4(n28174), .ZN(
        n28178) );
  OAI21_X1 U31431 ( .B1(n28179), .B2(n28178), .A(n28177), .ZN(n28263) );
  AOI22_X1 U31432 ( .A1(n29481), .A2(\xmem_data[24][0] ), .B1(n3368), .B2(
        \xmem_data[25][0] ), .ZN(n28184) );
  AOI22_X1 U31433 ( .A1(n3241), .A2(\xmem_data[26][0] ), .B1(n30663), .B2(
        \xmem_data[27][0] ), .ZN(n28183) );
  AOI22_X1 U31434 ( .A1(n30635), .A2(\xmem_data[28][0] ), .B1(n27753), .B2(
        \xmem_data[29][0] ), .ZN(n28182) );
  AOI22_X1 U31435 ( .A1(n3240), .A2(\xmem_data[30][0] ), .B1(n28091), .B2(
        \xmem_data[31][0] ), .ZN(n28181) );
  NAND2_X1 U31436 ( .A1(n30685), .A2(\xmem_data[5][0] ), .ZN(n28187) );
  NAND2_X1 U31437 ( .A1(n3182), .A2(\xmem_data[1][0] ), .ZN(n28186) );
  NAND2_X1 U31438 ( .A1(n3166), .A2(\xmem_data[0][0] ), .ZN(n28185) );
  NAND3_X1 U31439 ( .A1(n28187), .A2(n28186), .A3(n28185), .ZN(n28189) );
  AND2_X1 U31440 ( .A1(n29610), .A2(\xmem_data[2][0] ), .ZN(n28188) );
  AOI22_X1 U31441 ( .A1(n28191), .A2(\xmem_data[8][0] ), .B1(n28190), .B2(
        \xmem_data[9][0] ), .ZN(n28200) );
  AOI22_X1 U31442 ( .A1(n28193), .A2(\xmem_data[10][0] ), .B1(n28192), .B2(
        \xmem_data[11][0] ), .ZN(n28199) );
  AOI22_X1 U31443 ( .A1(n28195), .A2(\xmem_data[12][0] ), .B1(n28194), .B2(
        \xmem_data[13][0] ), .ZN(n28198) );
  AOI22_X1 U31444 ( .A1(n28196), .A2(\xmem_data[14][0] ), .B1(n3351), .B2(
        \xmem_data[15][0] ), .ZN(n28197) );
  AND2_X1 U31445 ( .A1(n28147), .A2(\xmem_data[3][0] ), .ZN(n28201) );
  AOI21_X1 U31446 ( .B1(n27713), .B2(\xmem_data[4][0] ), .A(n28201), .ZN(
        n28204) );
  AOI22_X1 U31447 ( .A1(n3233), .A2(\xmem_data[6][0] ), .B1(n28202), .B2(
        \xmem_data[7][0] ), .ZN(n28203) );
  NAND3_X1 U31448 ( .A1(n3824), .A2(n28205), .A3(n3551), .ZN(n28217) );
  AOI22_X1 U31449 ( .A1(n28734), .A2(\xmem_data[16][0] ), .B1(n30775), .B2(
        \xmem_data[17][0] ), .ZN(n28214) );
  AOI22_X1 U31450 ( .A1(n30215), .A2(\xmem_data[18][0] ), .B1(n30292), .B2(
        \xmem_data[19][0] ), .ZN(n28213) );
  AOI22_X1 U31451 ( .A1(n28209), .A2(\xmem_data[20][0] ), .B1(n29556), .B2(
        \xmem_data[21][0] ), .ZN(n28212) );
  AOI22_X1 U31452 ( .A1(n28210), .A2(\xmem_data[22][0] ), .B1(n3132), .B2(
        \xmem_data[23][0] ), .ZN(n28211) );
  NAND4_X1 U31453 ( .A1(n28214), .A2(n28213), .A3(n28212), .A4(n28211), .ZN(
        n28216) );
  AOI22_X1 U31454 ( .A1(n29421), .A2(\xmem_data[80][0] ), .B1(n30654), .B2(
        \xmem_data[81][0] ), .ZN(n28224) );
  AOI22_X1 U31455 ( .A1(n30279), .A2(\xmem_data[82][0] ), .B1(n28218), .B2(
        \xmem_data[83][0] ), .ZN(n28223) );
  AOI22_X1 U31456 ( .A1(n28219), .A2(\xmem_data[84][0] ), .B1(n3198), .B2(
        \xmem_data[85][0] ), .ZN(n28222) );
  AOI22_X1 U31457 ( .A1(n28220), .A2(\xmem_data[86][0] ), .B1(n20962), .B2(
        \xmem_data[87][0] ), .ZN(n28221) );
  NAND4_X1 U31458 ( .A1(n28224), .A2(n28223), .A3(n28222), .A4(n28221), .ZN(
        n28260) );
  AOI22_X1 U31459 ( .A1(\xmem_data[88][0] ), .A2(n27703), .B1(n30764), .B2(
        \xmem_data[66][0] ), .ZN(n28257) );
  AOI22_X1 U31460 ( .A1(n28685), .A2(\xmem_data[92][0] ), .B1(n28778), .B2(
        \xmem_data[93][0] ), .ZN(n28225) );
  INV_X1 U31461 ( .A(n28225), .ZN(n28230) );
  AOI22_X1 U31462 ( .A1(n30076), .A2(\xmem_data[68][0] ), .B1(n30644), .B2(
        \xmem_data[69][0] ), .ZN(n28228) );
  AOI22_X1 U31463 ( .A1(n3233), .A2(\xmem_data[70][0] ), .B1(n28226), .B2(
        \xmem_data[71][0] ), .ZN(n28227) );
  NAND2_X1 U31464 ( .A1(n28228), .A2(n28227), .ZN(n28229) );
  NOR2_X1 U31465 ( .A1(n28230), .A2(n28229), .ZN(n28256) );
  AOI22_X1 U31466 ( .A1(n3240), .A2(\xmem_data[94][0] ), .B1(n28231), .B2(
        \xmem_data[95][0] ), .ZN(n28236) );
  NAND2_X1 U31467 ( .A1(n28232), .A2(\xmem_data[67][0] ), .ZN(n28235) );
  AOI22_X1 U31468 ( .A1(n3241), .A2(\xmem_data[90][0] ), .B1(n28233), .B2(
        \xmem_data[91][0] ), .ZN(n28234) );
  NAND3_X1 U31469 ( .A1(n28236), .A2(n28235), .A3(n28234), .ZN(n28237) );
  AOI21_X1 U31470 ( .B1(n27761), .B2(\xmem_data[89][0] ), .A(n28237), .ZN(
        n28255) );
  AOI22_X1 U31471 ( .A1(n28240), .A2(\xmem_data[72][0] ), .B1(n28239), .B2(
        \xmem_data[73][0] ), .ZN(n28250) );
  AOI22_X1 U31472 ( .A1(n28242), .A2(\xmem_data[74][0] ), .B1(n28241), .B2(
        \xmem_data[75][0] ), .ZN(n28249) );
  AOI22_X1 U31473 ( .A1(n28244), .A2(\xmem_data[76][0] ), .B1(n28243), .B2(
        \xmem_data[77][0] ), .ZN(n28248) );
  AOI22_X1 U31474 ( .A1(n28246), .A2(\xmem_data[78][0] ), .B1(n28245), .B2(
        \xmem_data[79][0] ), .ZN(n28247) );
  NAND4_X1 U31475 ( .A1(n28250), .A2(n28249), .A3(n28248), .A4(n28247), .ZN(
        n28253) );
  AOI22_X1 U31476 ( .A1(n3165), .A2(\xmem_data[64][0] ), .B1(n3190), .B2(
        \xmem_data[65][0] ), .ZN(n28251) );
  INV_X1 U31477 ( .A(n28251), .ZN(n28252) );
  NOR2_X1 U31478 ( .A1(n28253), .A2(n28252), .ZN(n28254) );
  NAND4_X1 U31479 ( .A1(n28257), .A2(n28256), .A3(n28255), .A4(n28254), .ZN(
        n28259) );
  OAI21_X1 U31480 ( .B1(n28260), .B2(n28259), .A(n28258), .ZN(n28261) );
  XNOR2_X1 U31481 ( .A(n31940), .B(\fmem_data[23][3] ), .ZN(n32257) );
  OAI22_X1 U31482 ( .A1(n32257), .A2(n34410), .B1(n28266), .B2(n34412), .ZN(
        n28931) );
  OR2_X1 U31483 ( .A1(n34624), .A2(n3659), .ZN(n28267) );
  OAI22_X1 U31484 ( .A1(n28267), .A2(n35761), .B1(n35760), .B2(n3659), .ZN(
        n29847) );
  AOI22_X1 U31485 ( .A1(n28061), .A2(\xmem_data[120][0] ), .B1(n28291), .B2(
        \xmem_data[121][0] ), .ZN(n28272) );
  AOI22_X1 U31486 ( .A1(n29573), .A2(\xmem_data[122][0] ), .B1(n28062), .B2(
        \xmem_data[123][0] ), .ZN(n28271) );
  AOI22_X1 U31487 ( .A1(n28293), .A2(\xmem_data[124][0] ), .B1(n28292), .B2(
        \xmem_data[125][0] ), .ZN(n28270) );
  AND2_X1 U31488 ( .A1(n30601), .A2(\xmem_data[127][0] ), .ZN(n28268) );
  AOI21_X1 U31489 ( .B1(n29657), .B2(\xmem_data[126][0] ), .A(n28268), .ZN(
        n28269) );
  NAND4_X1 U31490 ( .A1(n28272), .A2(n28271), .A3(n28270), .A4(n28269), .ZN(
        n28283) );
  AOI22_X1 U31491 ( .A1(n28298), .A2(\xmem_data[112][0] ), .B1(n29309), .B2(
        \xmem_data[113][0] ), .ZN(n28276) );
  AOI22_X1 U31492 ( .A1(n31354), .A2(\xmem_data[114][0] ), .B1(n28299), .B2(
        \xmem_data[115][0] ), .ZN(n28275) );
  AOI22_X1 U31493 ( .A1(n29317), .A2(\xmem_data[116][0] ), .B1(n31355), .B2(
        \xmem_data[117][0] ), .ZN(n28274) );
  AOI22_X1 U31494 ( .A1(n28302), .A2(\xmem_data[118][0] ), .B1(n28301), .B2(
        \xmem_data[119][0] ), .ZN(n28273) );
  NAND4_X1 U31495 ( .A1(n28276), .A2(n28275), .A3(n28274), .A4(n28273), .ZN(
        n28282) );
  AOI22_X1 U31496 ( .A1(n24534), .A2(\xmem_data[104][0] ), .B1(n30550), .B2(
        \xmem_data[105][0] ), .ZN(n28280) );
  AOI22_X1 U31497 ( .A1(n28308), .A2(\xmem_data[106][0] ), .B1(n28307), .B2(
        \xmem_data[107][0] ), .ZN(n28279) );
  AOI22_X1 U31498 ( .A1(n27447), .A2(\xmem_data[108][0] ), .B1(n14996), .B2(
        \xmem_data[109][0] ), .ZN(n28278) );
  AOI22_X1 U31499 ( .A1(n28309), .A2(\xmem_data[110][0] ), .B1(n20958), .B2(
        \xmem_data[111][0] ), .ZN(n28277) );
  NAND4_X1 U31500 ( .A1(n28280), .A2(n28279), .A3(n28278), .A4(n28277), .ZN(
        n28281) );
  AOI22_X1 U31501 ( .A1(n30909), .A2(\xmem_data[96][0] ), .B1(n28317), .B2(
        \xmem_data[97][0] ), .ZN(n28287) );
  AOI22_X1 U31502 ( .A1(n3424), .A2(\xmem_data[98][0] ), .B1(n25687), .B2(
        \xmem_data[99][0] ), .ZN(n28286) );
  AOI22_X1 U31503 ( .A1(n28318), .A2(\xmem_data[100][0] ), .B1(n3220), .B2(
        \xmem_data[101][0] ), .ZN(n28285) );
  AOI22_X1 U31504 ( .A1(n27445), .A2(\xmem_data[102][0] ), .B1(n28319), .B2(
        \xmem_data[103][0] ), .ZN(n28284) );
  NAND4_X1 U31505 ( .A1(n28287), .A2(n28286), .A3(n28285), .A4(n28284), .ZN(
        n28289) );
  AOI22_X1 U31506 ( .A1(n28428), .A2(\xmem_data[88][0] ), .B1(n28291), .B2(
        \xmem_data[89][0] ), .ZN(n28297) );
  AOI22_X1 U31507 ( .A1(n24623), .A2(\xmem_data[90][0] ), .B1(n24622), .B2(
        \xmem_data[91][0] ), .ZN(n28296) );
  AOI22_X1 U31508 ( .A1(n28293), .A2(\xmem_data[92][0] ), .B1(n28292), .B2(
        \xmem_data[93][0] ), .ZN(n28295) );
  AOI22_X1 U31509 ( .A1(n20985), .A2(\xmem_data[94][0] ), .B1(n29125), .B2(
        \xmem_data[95][0] ), .ZN(n28294) );
  NAND4_X1 U31510 ( .A1(n28297), .A2(n28296), .A3(n28295), .A4(n28294), .ZN(
        n28316) );
  AOI22_X1 U31511 ( .A1(n28298), .A2(\xmem_data[80][0] ), .B1(n22703), .B2(
        \xmem_data[81][0] ), .ZN(n28306) );
  AOI22_X1 U31512 ( .A1(n29396), .A2(\xmem_data[82][0] ), .B1(n28299), .B2(
        \xmem_data[83][0] ), .ZN(n28305) );
  AOI22_X1 U31513 ( .A1(n25573), .A2(\xmem_data[84][0] ), .B1(n25398), .B2(
        \xmem_data[85][0] ), .ZN(n28304) );
  AOI22_X1 U31514 ( .A1(n28302), .A2(\xmem_data[86][0] ), .B1(n28301), .B2(
        \xmem_data[87][0] ), .ZN(n28303) );
  NAND4_X1 U31515 ( .A1(n28306), .A2(n28305), .A3(n28304), .A4(n28303), .ZN(
        n28315) );
  AOI22_X1 U31516 ( .A1(n20725), .A2(\xmem_data[72][0] ), .B1(n25616), .B2(
        \xmem_data[73][0] ), .ZN(n28313) );
  AOI22_X1 U31517 ( .A1(n28308), .A2(\xmem_data[74][0] ), .B1(n28307), .B2(
        \xmem_data[75][0] ), .ZN(n28312) );
  AOI22_X1 U31518 ( .A1(n25422), .A2(\xmem_data[76][0] ), .B1(n14996), .B2(
        \xmem_data[77][0] ), .ZN(n28311) );
  AOI22_X1 U31519 ( .A1(n28309), .A2(\xmem_data[78][0] ), .B1(n24555), .B2(
        \xmem_data[79][0] ), .ZN(n28310) );
  NAND4_X1 U31520 ( .A1(n28313), .A2(n28312), .A3(n28311), .A4(n28310), .ZN(
        n28314) );
  AOI22_X1 U31521 ( .A1(n20827), .A2(\xmem_data[64][0] ), .B1(n28317), .B2(
        \xmem_data[65][0] ), .ZN(n28323) );
  AOI22_X1 U31522 ( .A1(n3424), .A2(\xmem_data[66][0] ), .B1(n31347), .B2(
        \xmem_data[67][0] ), .ZN(n28322) );
  AOI22_X1 U31523 ( .A1(n28318), .A2(\xmem_data[68][0] ), .B1(n3221), .B2(
        \xmem_data[69][0] ), .ZN(n28321) );
  AOI22_X1 U31524 ( .A1(n28137), .A2(\xmem_data[70][0] ), .B1(n28319), .B2(
        \xmem_data[71][0] ), .ZN(n28320) );
  NAND4_X1 U31525 ( .A1(n28323), .A2(n28322), .A3(n28321), .A4(n28320), .ZN(
        n28325) );
  AOI22_X1 U31526 ( .A1(n27524), .A2(\xmem_data[56][0] ), .B1(n25581), .B2(
        \xmem_data[57][0] ), .ZN(n28333) );
  AOI22_X1 U31527 ( .A1(n31315), .A2(\xmem_data[58][0] ), .B1(n14975), .B2(
        \xmem_data[59][0] ), .ZN(n28332) );
  AOI22_X1 U31528 ( .A1(n3179), .A2(\xmem_data[60][0] ), .B1(n28328), .B2(
        \xmem_data[61][0] ), .ZN(n28331) );
  AOI22_X1 U31529 ( .A1(n30674), .A2(\xmem_data[62][0] ), .B1(n28329), .B2(
        \xmem_data[63][0] ), .ZN(n28330) );
  NAND4_X1 U31530 ( .A1(n28333), .A2(n28332), .A3(n28331), .A4(n28330), .ZN(
        n28353) );
  AOI22_X1 U31531 ( .A1(n28334), .A2(\xmem_data[48][0] ), .B1(n24160), .B2(
        \xmem_data[49][0] ), .ZN(n28341) );
  AOI22_X1 U31532 ( .A1(n28336), .A2(\xmem_data[50][0] ), .B1(n28335), .B2(
        \xmem_data[51][0] ), .ZN(n28340) );
  AOI22_X1 U31533 ( .A1(n28337), .A2(\xmem_data[52][0] ), .B1(n29048), .B2(
        \xmem_data[53][0] ), .ZN(n28339) );
  AOI22_X1 U31534 ( .A1(n27855), .A2(\xmem_data[54][0] ), .B1(n24646), .B2(
        \xmem_data[55][0] ), .ZN(n28338) );
  NAND4_X1 U31535 ( .A1(n28341), .A2(n28340), .A3(n28339), .A4(n28338), .ZN(
        n28352) );
  AOI22_X1 U31536 ( .A1(n25490), .A2(\xmem_data[40][0] ), .B1(n28342), .B2(
        \xmem_data[41][0] ), .ZN(n28350) );
  AOI22_X1 U31537 ( .A1(n28344), .A2(\xmem_data[42][0] ), .B1(n28007), .B2(
        \xmem_data[43][0] ), .ZN(n28349) );
  AOI22_X1 U31538 ( .A1(n25422), .A2(\xmem_data[44][0] ), .B1(n27988), .B2(
        \xmem_data[45][0] ), .ZN(n28348) );
  AOI22_X1 U31539 ( .A1(n28346), .A2(\xmem_data[46][0] ), .B1(n28345), .B2(
        \xmem_data[47][0] ), .ZN(n28347) );
  NAND4_X1 U31540 ( .A1(n28350), .A2(n28349), .A3(n28348), .A4(n28347), .ZN(
        n28351) );
  AOI22_X1 U31541 ( .A1(n28354), .A2(\xmem_data[32][0] ), .B1(n25561), .B2(
        \xmem_data[33][0] ), .ZN(n28360) );
  AOI22_X1 U31542 ( .A1(n24693), .A2(\xmem_data[34][0] ), .B1(n14875), .B2(
        \xmem_data[35][0] ), .ZN(n28359) );
  AOI22_X1 U31543 ( .A1(n28355), .A2(\xmem_data[36][0] ), .B1(n3222), .B2(
        \xmem_data[37][0] ), .ZN(n28358) );
  AOI22_X1 U31544 ( .A1(n25414), .A2(\xmem_data[38][0] ), .B1(n28356), .B2(
        \xmem_data[39][0] ), .ZN(n28357) );
  NAND4_X1 U31545 ( .A1(n28360), .A2(n28359), .A3(n28358), .A4(n28357), .ZN(
        n28362) );
  AOI22_X1 U31546 ( .A1(n28364), .A2(\xmem_data[4][0] ), .B1(n3219), .B2(
        \xmem_data[5][0] ), .ZN(n28371) );
  AOI22_X1 U31547 ( .A1(n3305), .A2(\xmem_data[2][0] ), .B1(n25360), .B2(
        \xmem_data[3][0] ), .ZN(n28370) );
  AOI22_X1 U31548 ( .A1(n25630), .A2(\xmem_data[0][0] ), .B1(n28366), .B2(
        \xmem_data[1][0] ), .ZN(n28369) );
  AOI22_X1 U31549 ( .A1(n28367), .A2(\xmem_data[6][0] ), .B1(n22667), .B2(
        \xmem_data[7][0] ), .ZN(n28368) );
  NAND4_X1 U31550 ( .A1(n28371), .A2(n28370), .A3(n28369), .A4(n28368), .ZN(
        n28394) );
  AOI22_X1 U31551 ( .A1(n29289), .A2(\xmem_data[8][0] ), .B1(n28372), .B2(
        \xmem_data[9][0] ), .ZN(n28379) );
  AOI22_X1 U31552 ( .A1(n16973), .A2(\xmem_data[10][0] ), .B1(n24657), .B2(
        \xmem_data[11][0] ), .ZN(n28378) );
  AOI22_X1 U31553 ( .A1(n28374), .A2(\xmem_data[12][0] ), .B1(n3357), .B2(
        \xmem_data[13][0] ), .ZN(n28377) );
  AOI22_X1 U31554 ( .A1(n17064), .A2(\xmem_data[14][0] ), .B1(n28375), .B2(
        \xmem_data[15][0] ), .ZN(n28376) );
  NAND4_X1 U31555 ( .A1(n28379), .A2(n28378), .A3(n28377), .A4(n28376), .ZN(
        n28393) );
  AOI22_X1 U31556 ( .A1(n28053), .A2(\xmem_data[18][0] ), .B1(n13188), .B2(
        \xmem_data[19][0] ), .ZN(n28384) );
  AOI22_X1 U31557 ( .A1(n24131), .A2(\xmem_data[16][0] ), .B1(n22703), .B2(
        \xmem_data[17][0] ), .ZN(n28383) );
  AOI22_X1 U31558 ( .A1(n13149), .A2(\xmem_data[20][0] ), .B1(n20505), .B2(
        \xmem_data[21][0] ), .ZN(n28382) );
  AOI22_X1 U31559 ( .A1(n22682), .A2(\xmem_data[22][0] ), .B1(n28380), .B2(
        \xmem_data[23][0] ), .ZN(n28381) );
  NAND4_X1 U31560 ( .A1(n28384), .A2(n28383), .A3(n28382), .A4(n28381), .ZN(
        n28392) );
  AOI22_X1 U31561 ( .A1(n28385), .A2(\xmem_data[24][0] ), .B1(n20816), .B2(
        \xmem_data[25][0] ), .ZN(n28390) );
  AOI22_X1 U31562 ( .A1(n29054), .A2(\xmem_data[26][0] ), .B1(n14975), .B2(
        \xmem_data[27][0] ), .ZN(n28389) );
  AOI22_X1 U31563 ( .A1(n27542), .A2(\xmem_data[28][0] ), .B1(n28979), .B2(
        \xmem_data[29][0] ), .ZN(n28388) );
  AND2_X1 U31564 ( .A1(n10456), .A2(\xmem_data[31][0] ), .ZN(n28386) );
  AOI21_X1 U31565 ( .B1(n14982), .B2(\xmem_data[30][0] ), .A(n28386), .ZN(
        n28387) );
  NAND4_X1 U31566 ( .A1(n28390), .A2(n28389), .A3(n28388), .A4(n28387), .ZN(
        n28391) );
  OR4_X1 U31567 ( .A1(n28394), .A2(n28393), .A3(n28392), .A4(n28391), .ZN(
        n28396) );
  NAND2_X1 U31568 ( .A1(n28396), .A2(n28395), .ZN(n28397) );
  NAND4_X4 U31569 ( .A1(n28400), .A2(n28399), .A3(n28398), .A4(n28397), .ZN(
        n36105) );
  XNOR2_X1 U31570 ( .A(n3366), .B(\fmem_data[3][3] ), .ZN(n32195) );
  OAI21_X1 U31571 ( .B1(n31208), .B2(n31210), .A(n31209), .ZN(n28405) );
  NAND2_X1 U31572 ( .A1(n31208), .A2(n31210), .ZN(n28404) );
  NAND2_X1 U31573 ( .A1(n28405), .A2(n28404), .ZN(n30149) );
  FA_X1 U31574 ( .A(n28408), .B(n28407), .CI(n28406), .CO(n34166), .S(n33626)
         );
  XNOR2_X1 U31575 ( .A(n30451), .B(\fmem_data[6][1] ), .ZN(n34018) );
  XNOR2_X1 U31576 ( .A(n33556), .B(\fmem_data[16][5] ), .ZN(n32565) );
  AOI22_X1 U31577 ( .A1(n27981), .A2(\xmem_data[8][0] ), .B1(n20952), .B2(
        \xmem_data[9][0] ), .ZN(n28413) );
  AOI22_X1 U31578 ( .A1(n24524), .A2(\xmem_data[10][0] ), .B1(n30862), .B2(
        \xmem_data[11][0] ), .ZN(n28412) );
  AOI22_X1 U31579 ( .A1(n25629), .A2(\xmem_data[12][0] ), .B1(n28677), .B2(
        \xmem_data[13][0] ), .ZN(n28411) );
  AOI22_X1 U31580 ( .A1(n3247), .A2(\xmem_data[14][0] ), .B1(n28082), .B2(
        \xmem_data[15][0] ), .ZN(n28410) );
  AOI22_X1 U31581 ( .A1(n28007), .A2(\xmem_data[22][0] ), .B1(n25422), .B2(
        \xmem_data[23][0] ), .ZN(n28414) );
  INV_X1 U31582 ( .A(n28414), .ZN(n28426) );
  AOI22_X1 U31583 ( .A1(n28415), .A2(\xmem_data[24][0] ), .B1(n27911), .B2(
        \xmem_data[25][0] ), .ZN(n28420) );
  AOI22_X1 U31584 ( .A1(n28416), .A2(\xmem_data[26][0] ), .B1(n30514), .B2(
        \xmem_data[27][0] ), .ZN(n28419) );
  AOI22_X1 U31585 ( .A1(n25382), .A2(\xmem_data[28][0] ), .B1(n3465), .B2(
        \xmem_data[29][0] ), .ZN(n28418) );
  AOI22_X1 U31586 ( .A1(n13188), .A2(\xmem_data[30][0] ), .B1(n24509), .B2(
        \xmem_data[31][0] ), .ZN(n28417) );
  NAND4_X1 U31587 ( .A1(n28420), .A2(n28419), .A3(n28418), .A4(n28417), .ZN(
        n28425) );
  AOI22_X1 U31588 ( .A1(n23811), .A2(\xmem_data[20][0] ), .B1(n29706), .B2(
        \xmem_data[21][0] ), .ZN(n28423) );
  AOI22_X1 U31589 ( .A1(n25562), .A2(\xmem_data[18][0] ), .B1(n27904), .B2(
        \xmem_data[19][0] ), .ZN(n28422) );
  AOI22_X1 U31590 ( .A1(n3222), .A2(\xmem_data[16][0] ), .B1(n29789), .B2(
        \xmem_data[17][0] ), .ZN(n28421) );
  NAND3_X1 U31591 ( .A1(n28423), .A2(n28422), .A3(n28421), .ZN(n28424) );
  OR3_X1 U31592 ( .A1(n28426), .A2(n28425), .A3(n28424), .ZN(n28435) );
  AOI22_X1 U31593 ( .A1(n28427), .A2(\xmem_data[0][0] ), .B1(n29439), .B2(
        \xmem_data[1][0] ), .ZN(n28433) );
  AOI22_X1 U31594 ( .A1(n23776), .A2(\xmem_data[2][0] ), .B1(n28428), .B2(
        \xmem_data[3][0] ), .ZN(n28432) );
  AOI22_X1 U31595 ( .A1(n21009), .A2(\xmem_data[4][0] ), .B1(n29816), .B2(
        \xmem_data[5][0] ), .ZN(n28431) );
  AOI22_X1 U31596 ( .A1(n31362), .A2(\xmem_data[6][0] ), .B1(n14976), .B2(
        \xmem_data[7][0] ), .ZN(n28430) );
  NAND4_X1 U31597 ( .A1(n28433), .A2(n28432), .A3(n28431), .A4(n28430), .ZN(
        n28434) );
  NOR2_X1 U31598 ( .A1(n28435), .A2(n28434), .ZN(n28436) );
  AOI21_X1 U31599 ( .B1(n3749), .B2(n28436), .A(n15043), .ZN(n28437) );
  AOI22_X1 U31600 ( .A1(n28492), .A2(\xmem_data[96][0] ), .B1(n29239), .B2(
        \xmem_data[97][0] ), .ZN(n28441) );
  AOI22_X1 U31601 ( .A1(n29238), .A2(\xmem_data[98][0] ), .B1(n28493), .B2(
        \xmem_data[99][0] ), .ZN(n28440) );
  AOI22_X1 U31602 ( .A1(n28494), .A2(\xmem_data[100][0] ), .B1(n3271), .B2(
        \xmem_data[101][0] ), .ZN(n28439) );
  AOI22_X1 U31603 ( .A1(n28495), .A2(\xmem_data[102][0] ), .B1(n24685), .B2(
        \xmem_data[103][0] ), .ZN(n28438) );
  NAND4_X1 U31604 ( .A1(n28441), .A2(n28440), .A3(n28439), .A4(n28438), .ZN(
        n28457) );
  AOI22_X1 U31605 ( .A1(n28500), .A2(\xmem_data[104][0] ), .B1(n27717), .B2(
        \xmem_data[105][0] ), .ZN(n28445) );
  AOI22_X1 U31606 ( .A1(n25388), .A2(\xmem_data[106][0] ), .B1(n20710), .B2(
        \xmem_data[107][0] ), .ZN(n28444) );
  AOI22_X1 U31607 ( .A1(n22752), .A2(\xmem_data[108][0] ), .B1(n3352), .B2(
        \xmem_data[109][0] ), .ZN(n28443) );
  AOI22_X1 U31608 ( .A1(n28501), .A2(\xmem_data[110][0] ), .B1(n28503), .B2(
        \xmem_data[111][0] ), .ZN(n28442) );
  NAND4_X1 U31609 ( .A1(n28445), .A2(n28444), .A3(n28443), .A4(n28442), .ZN(
        n28456) );
  AOI22_X1 U31610 ( .A1(n3220), .A2(\xmem_data[112][0] ), .B1(n24696), .B2(
        \xmem_data[113][0] ), .ZN(n28449) );
  AOI22_X1 U31611 ( .A1(n28508), .A2(\xmem_data[114][0] ), .B1(n3322), .B2(
        \xmem_data[115][0] ), .ZN(n28448) );
  AOI22_X1 U31612 ( .A1(n28509), .A2(\xmem_data[116][0] ), .B1(n30698), .B2(
        \xmem_data[117][0] ), .ZN(n28447) );
  AOI22_X1 U31613 ( .A1(n28343), .A2(\xmem_data[118][0] ), .B1(n28374), .B2(
        \xmem_data[119][0] ), .ZN(n28446) );
  NAND4_X1 U31614 ( .A1(n28449), .A2(n28448), .A3(n28447), .A4(n28446), .ZN(
        n28455) );
  AOI22_X1 U31615 ( .A1(n3358), .A2(\xmem_data[120][0] ), .B1(n20716), .B2(
        \xmem_data[121][0] ), .ZN(n28453) );
  AOI22_X1 U31616 ( .A1(n28515), .A2(\xmem_data[122][0] ), .B1(n17041), .B2(
        \xmem_data[123][0] ), .ZN(n28452) );
  AOI22_X1 U31617 ( .A1(n28517), .A2(\xmem_data[124][0] ), .B1(n27818), .B2(
        \xmem_data[125][0] ), .ZN(n28451) );
  AOI22_X1 U31618 ( .A1(n28299), .A2(\xmem_data[126][0] ), .B1(n24509), .B2(
        \xmem_data[127][0] ), .ZN(n28450) );
  NAND4_X1 U31619 ( .A1(n28453), .A2(n28452), .A3(n28451), .A4(n28450), .ZN(
        n28454) );
  OR4_X1 U31620 ( .A1(n28457), .A2(n28456), .A3(n28455), .A4(n28454), .ZN(
        n28459) );
  AOI22_X1 U31621 ( .A1(n24645), .A2(\xmem_data[32][0] ), .B1(n28302), .B2(
        \xmem_data[33][0] ), .ZN(n28466) );
  AOI22_X1 U31622 ( .A1(n29238), .A2(\xmem_data[34][0] ), .B1(n3326), .B2(
        \xmem_data[35][0] ), .ZN(n28465) );
  AOI22_X1 U31623 ( .A1(n28462), .A2(\xmem_data[36][0] ), .B1(n28461), .B2(
        \xmem_data[37][0] ), .ZN(n28464) );
  AOI22_X1 U31624 ( .A1(n24521), .A2(\xmem_data[38][0] ), .B1(n24685), .B2(
        \xmem_data[39][0] ), .ZN(n28463) );
  NAND4_X1 U31625 ( .A1(n28466), .A2(n28465), .A3(n28464), .A4(n28463), .ZN(
        n28489) );
  AOI22_X1 U31626 ( .A1(n28468), .A2(\xmem_data[40][0] ), .B1(n28467), .B2(
        \xmem_data[41][0] ), .ZN(n28474) );
  AOI22_X1 U31627 ( .A1(n25528), .A2(\xmem_data[42][0] ), .B1(n30588), .B2(
        \xmem_data[43][0] ), .ZN(n28473) );
  AOI22_X1 U31628 ( .A1(n24573), .A2(\xmem_data[44][0] ), .B1(n28718), .B2(
        \xmem_data[45][0] ), .ZN(n28472) );
  AND2_X1 U31629 ( .A1(n25360), .A2(\xmem_data[46][0] ), .ZN(n28469) );
  AOI21_X1 U31630 ( .B1(n28470), .B2(\xmem_data[47][0] ), .A(n28469), .ZN(
        n28471) );
  NAND4_X1 U31631 ( .A1(n28474), .A2(n28473), .A3(n28472), .A4(n28471), .ZN(
        n28488) );
  AOI22_X1 U31632 ( .A1(n3220), .A2(\xmem_data[48][0] ), .B1(n29422), .B2(
        \xmem_data[49][0] ), .ZN(n28480) );
  AOI22_X1 U31633 ( .A1(n28476), .A2(\xmem_data[50][0] ), .B1(n28475), .B2(
        \xmem_data[51][0] ), .ZN(n28479) );
  AOI22_X1 U31634 ( .A1(n20559), .A2(\xmem_data[52][0] ), .B1(n3132), .B2(
        \xmem_data[53][0] ), .ZN(n28478) );
  AOI22_X1 U31635 ( .A1(n25514), .A2(\xmem_data[54][0] ), .B1(n27551), .B2(
        \xmem_data[55][0] ), .ZN(n28477) );
  NAND4_X1 U31636 ( .A1(n28480), .A2(n28479), .A3(n28478), .A4(n28477), .ZN(
        n28487) );
  AOI22_X1 U31637 ( .A1(n28481), .A2(\xmem_data[56][0] ), .B1(n28152), .B2(
        \xmem_data[57][0] ), .ZN(n28485) );
  AOI22_X1 U31638 ( .A1(n14998), .A2(\xmem_data[58][0] ), .B1(n28298), .B2(
        \xmem_data[59][0] ), .ZN(n28484) );
  AOI22_X1 U31639 ( .A1(n29009), .A2(\xmem_data[60][0] ), .B1(n29237), .B2(
        \xmem_data[61][0] ), .ZN(n28483) );
  AOI22_X1 U31640 ( .A1(n27516), .A2(\xmem_data[62][0] ), .B1(n23717), .B2(
        \xmem_data[63][0] ), .ZN(n28482) );
  NAND4_X1 U31641 ( .A1(n28485), .A2(n28484), .A3(n28483), .A4(n28482), .ZN(
        n28486) );
  OR4_X1 U31642 ( .A1(n28489), .A2(n28488), .A3(n28487), .A4(n28486), .ZN(
        n28491) );
  AOI22_X1 U31643 ( .A1(n28492), .A2(\xmem_data[64][0] ), .B1(n23722), .B2(
        \xmem_data[65][0] ), .ZN(n28499) );
  AOI22_X1 U31644 ( .A1(n24460), .A2(\xmem_data[66][0] ), .B1(n28493), .B2(
        \xmem_data[67][0] ), .ZN(n28498) );
  AOI22_X1 U31645 ( .A1(n28494), .A2(\xmem_data[68][0] ), .B1(n17004), .B2(
        \xmem_data[69][0] ), .ZN(n28497) );
  AOI22_X1 U31646 ( .A1(n28495), .A2(\xmem_data[70][0] ), .B1(n24606), .B2(
        \xmem_data[71][0] ), .ZN(n28496) );
  NAND4_X1 U31647 ( .A1(n28499), .A2(n28498), .A3(n28497), .A4(n28496), .ZN(
        n28525) );
  AOI22_X1 U31648 ( .A1(n28500), .A2(\xmem_data[72][0] ), .B1(n29383), .B2(
        \xmem_data[73][0] ), .ZN(n28507) );
  AOI22_X1 U31649 ( .A1(n24468), .A2(\xmem_data[74][0] ), .B1(n28076), .B2(
        \xmem_data[75][0] ), .ZN(n28506) );
  AOI22_X1 U31650 ( .A1(n29328), .A2(\xmem_data[76][0] ), .B1(n3412), .B2(
        \xmem_data[77][0] ), .ZN(n28505) );
  AND2_X1 U31651 ( .A1(n28501), .A2(\xmem_data[78][0] ), .ZN(n28502) );
  AOI21_X1 U31652 ( .B1(n28503), .B2(\xmem_data[79][0] ), .A(n28502), .ZN(
        n28504) );
  NAND4_X1 U31653 ( .A1(n28507), .A2(n28506), .A3(n28505), .A4(n28504), .ZN(
        n28524) );
  AOI22_X1 U31654 ( .A1(n3218), .A2(\xmem_data[80][0] ), .B1(n27445), .B2(
        \xmem_data[81][0] ), .ZN(n28514) );
  AOI22_X1 U31655 ( .A1(n28508), .A2(\xmem_data[82][0] ), .B1(n3342), .B2(
        \xmem_data[83][0] ), .ZN(n28513) );
  AOI22_X1 U31656 ( .A1(n28509), .A2(\xmem_data[84][0] ), .B1(n30295), .B2(
        \xmem_data[85][0] ), .ZN(n28512) );
  AOI22_X1 U31657 ( .A1(n27547), .A2(\xmem_data[86][0] ), .B1(n28374), .B2(
        \xmem_data[87][0] ), .ZN(n28511) );
  NAND4_X1 U31658 ( .A1(n28514), .A2(n28513), .A3(n28512), .A4(n28511), .ZN(
        n28523) );
  AOI22_X1 U31659 ( .A1(n3358), .A2(\xmem_data[88][0] ), .B1(n29591), .B2(
        \xmem_data[89][0] ), .ZN(n28521) );
  AOI22_X1 U31660 ( .A1(n28515), .A2(\xmem_data[90][0] ), .B1(n29310), .B2(
        \xmem_data[91][0] ), .ZN(n28520) );
  AOI22_X1 U31661 ( .A1(n28517), .A2(\xmem_data[92][0] ), .B1(n29237), .B2(
        \xmem_data[93][0] ), .ZN(n28519) );
  AOI22_X1 U31662 ( .A1(n24134), .A2(\xmem_data[94][0] ), .B1(n24509), .B2(
        \xmem_data[95][0] ), .ZN(n28518) );
  NAND4_X1 U31663 ( .A1(n28521), .A2(n28520), .A3(n28519), .A4(n28518), .ZN(
        n28522) );
  OR4_X1 U31664 ( .A1(n28525), .A2(n28524), .A3(n28523), .A4(n28522), .ZN(
        n28527) );
  NAND2_X1 U31665 ( .A1(n28527), .A2(n28526), .ZN(n28528) );
  INV_X1 U31666 ( .A(n35083), .ZN(n28532) );
  XNOR2_X1 U31667 ( .A(n28534), .B(n28533), .ZN(n31509) );
  XNOR2_X1 U31668 ( .A(n33555), .B(\fmem_data[21][3] ), .ZN(n32067) );
  XNOR2_X1 U31669 ( .A(n32057), .B(\fmem_data[21][3] ), .ZN(n34200) );
  XNOR2_X1 U31670 ( .A(n28538), .B(n28537), .ZN(n31465) );
  XNOR2_X1 U31671 ( .A(n30846), .B(\fmem_data[13][1] ), .ZN(n32056) );
  XNOR2_X1 U31672 ( .A(n28539), .B(\fmem_data[13][1] ), .ZN(n32240) );
  XNOR2_X1 U31673 ( .A(n31897), .B(\fmem_data[28][1] ), .ZN(n32071) );
  XNOR2_X1 U31674 ( .A(n31219), .B(\fmem_data[26][3] ), .ZN(n32144) );
  AOI22_X1 U31675 ( .A1(n30514), .A2(\xmem_data[56][2] ), .B1(n30513), .B2(
        \xmem_data[57][2] ), .ZN(n28546) );
  AOI22_X1 U31676 ( .A1(n28154), .A2(\xmem_data[58][2] ), .B1(n3208), .B2(
        \xmem_data[59][2] ), .ZN(n28545) );
  AOI22_X1 U31677 ( .A1(n24593), .A2(\xmem_data[60][2] ), .B1(n21006), .B2(
        \xmem_data[61][2] ), .ZN(n28544) );
  AOI22_X1 U31678 ( .A1(n25678), .A2(\xmem_data[62][2] ), .B1(n30515), .B2(
        \xmem_data[63][2] ), .ZN(n28543) );
  NAND4_X1 U31679 ( .A1(n28546), .A2(n28545), .A3(n28544), .A4(n28543), .ZN(
        n28549) );
  AOI22_X1 U31680 ( .A1(n24688), .A2(\xmem_data[40][2] ), .B1(n30908), .B2(
        \xmem_data[41][2] ), .ZN(n28547) );
  INV_X1 U31681 ( .A(n28547), .ZN(n28548) );
  NOR2_X1 U31682 ( .A1(n28549), .A2(n28548), .ZN(n28554) );
  AOI22_X1 U31683 ( .A1(n24647), .A2(\xmem_data[32][2] ), .B1(n30495), .B2(
        \xmem_data[33][2] ), .ZN(n28553) );
  AOI22_X1 U31684 ( .A1(n14974), .A2(\xmem_data[34][2] ), .B1(n20949), .B2(
        \xmem_data[35][2] ), .ZN(n28552) );
  AOI22_X1 U31685 ( .A1(n30497), .A2(\xmem_data[36][2] ), .B1(n30496), .B2(
        \xmem_data[37][2] ), .ZN(n28551) );
  AOI22_X1 U31686 ( .A1(n24687), .A2(\xmem_data[38][2] ), .B1(n30498), .B2(
        \xmem_data[39][2] ), .ZN(n28550) );
  NAND2_X1 U31687 ( .A1(n28554), .A2(n3747), .ZN(n28566) );
  AOI22_X1 U31688 ( .A1(n20725), .A2(\xmem_data[48][2] ), .B1(n3256), .B2(
        \xmem_data[49][2] ), .ZN(n28558) );
  AOI22_X1 U31689 ( .A1(n22668), .A2(\xmem_data[50][2] ), .B1(n29103), .B2(
        \xmem_data[51][2] ), .ZN(n28557) );
  AOI22_X1 U31690 ( .A1(n24638), .A2(\xmem_data[52][2] ), .B1(n22701), .B2(
        \xmem_data[53][2] ), .ZN(n28556) );
  AOI22_X1 U31691 ( .A1(n30508), .A2(\xmem_data[54][2] ), .B1(n24212), .B2(
        \xmem_data[55][2] ), .ZN(n28555) );
  NAND4_X1 U31692 ( .A1(n28558), .A2(n28557), .A3(n28556), .A4(n28555), .ZN(
        n28562) );
  AOI22_X1 U31693 ( .A1(n25612), .A2(\xmem_data[46][2] ), .B1(n29095), .B2(
        \xmem_data[47][2] ), .ZN(n28560) );
  AOI22_X1 U31694 ( .A1(n28039), .A2(\xmem_data[42][2] ), .B1(n29286), .B2(
        \xmem_data[43][2] ), .ZN(n28559) );
  NAND2_X1 U31695 ( .A1(n28560), .A2(n28559), .ZN(n28561) );
  NOR2_X1 U31696 ( .A1(n28562), .A2(n28561), .ZN(n28564) );
  AOI22_X1 U31697 ( .A1(n30503), .A2(\xmem_data[44][2] ), .B1(n3217), .B2(
        \xmem_data[45][2] ), .ZN(n28563) );
  NAND2_X1 U31698 ( .A1(n28564), .A2(n28563), .ZN(n28565) );
  OAI21_X1 U31699 ( .B1(n28566), .B2(n28565), .A(n30565), .ZN(n28635) );
  AND2_X1 U31700 ( .A1(n3218), .A2(\xmem_data[77][2] ), .ZN(n28567) );
  AOI21_X1 U31701 ( .B1(n30592), .B2(\xmem_data[76][2] ), .A(n28567), .ZN(
        n28571) );
  AOI22_X1 U31702 ( .A1(n3229), .A2(\xmem_data[74][2] ), .B1(n30589), .B2(
        \xmem_data[75][2] ), .ZN(n28570) );
  AOI22_X1 U31703 ( .A1(n30588), .A2(\xmem_data[72][2] ), .B1(n20578), .B2(
        \xmem_data[73][2] ), .ZN(n28569) );
  AOI22_X1 U31704 ( .A1(n30593), .A2(\xmem_data[78][2] ), .B1(n20558), .B2(
        \xmem_data[79][2] ), .ZN(n28568) );
  NAND4_X1 U31705 ( .A1(n28571), .A2(n28570), .A3(n28569), .A4(n28568), .ZN(
        n28587) );
  AOI22_X1 U31706 ( .A1(n30849), .A2(\xmem_data[64][2] ), .B1(n25716), .B2(
        \xmem_data[65][2] ), .ZN(n28575) );
  AOI22_X1 U31707 ( .A1(n30600), .A2(\xmem_data[66][2] ), .B1(n30599), .B2(
        \xmem_data[67][2] ), .ZN(n28574) );
  AOI22_X1 U31708 ( .A1(n20782), .A2(\xmem_data[68][2] ), .B1(n31256), .B2(
        \xmem_data[69][2] ), .ZN(n28573) );
  AOI22_X1 U31709 ( .A1(n25628), .A2(\xmem_data[70][2] ), .B1(n30601), .B2(
        \xmem_data[71][2] ), .ZN(n28572) );
  NAND4_X1 U31710 ( .A1(n28575), .A2(n28574), .A3(n28573), .A4(n28572), .ZN(
        n28586) );
  AOI22_X1 U31711 ( .A1(n30606), .A2(\xmem_data[80][2] ), .B1(n3255), .B2(
        \xmem_data[81][2] ), .ZN(n28579) );
  AOI22_X1 U31712 ( .A1(n29231), .A2(\xmem_data[82][2] ), .B1(n28045), .B2(
        \xmem_data[83][2] ), .ZN(n28578) );
  AOI22_X1 U31713 ( .A1(n30607), .A2(\xmem_data[84][2] ), .B1(n27863), .B2(
        \xmem_data[85][2] ), .ZN(n28577) );
  AOI22_X1 U31714 ( .A1(n30608), .A2(\xmem_data[86][2] ), .B1(n22675), .B2(
        \xmem_data[87][2] ), .ZN(n28576) );
  NAND4_X1 U31715 ( .A1(n28579), .A2(n28578), .A3(n28577), .A4(n28576), .ZN(
        n28585) );
  AOI22_X1 U31716 ( .A1(n30614), .A2(\xmem_data[88][2] ), .B1(n30613), .B2(
        \xmem_data[89][2] ), .ZN(n28583) );
  AOI22_X1 U31717 ( .A1(n3157), .A2(\xmem_data[90][2] ), .B1(n30615), .B2(
        \xmem_data[91][2] ), .ZN(n28582) );
  AOI22_X1 U31718 ( .A1(n24547), .A2(\xmem_data[92][2] ), .B1(n20505), .B2(
        \xmem_data[93][2] ), .ZN(n28581) );
  AOI22_X1 U31719 ( .A1(n30617), .A2(\xmem_data[94][2] ), .B1(n30616), .B2(
        \xmem_data[95][2] ), .ZN(n28580) );
  NAND4_X1 U31720 ( .A1(n28583), .A2(n28582), .A3(n28581), .A4(n28580), .ZN(
        n28584) );
  OR4_X1 U31721 ( .A1(n28587), .A2(n28586), .A3(n28585), .A4(n28584), .ZN(
        n28588) );
  NAND2_X1 U31722 ( .A1(n28588), .A2(n30628), .ZN(n28634) );
  AOI22_X1 U31723 ( .A1(n28038), .A2(\xmem_data[8][2] ), .B1(n28317), .B2(
        \xmem_data[9][2] ), .ZN(n28592) );
  AOI22_X1 U31724 ( .A1(n3412), .A2(\xmem_data[10][2] ), .B1(n28501), .B2(
        \xmem_data[11][2] ), .ZN(n28591) );
  AOI22_X1 U31725 ( .A1(n20991), .A2(\xmem_data[12][2] ), .B1(n3221), .B2(
        \xmem_data[13][2] ), .ZN(n28590) );
  AOI22_X1 U31726 ( .A1(n28733), .A2(\xmem_data[14][2] ), .B1(n30534), .B2(
        \xmem_data[15][2] ), .ZN(n28589) );
  NAND4_X1 U31727 ( .A1(n28592), .A2(n28591), .A3(n28590), .A4(n28589), .ZN(
        n28608) );
  AOI22_X1 U31728 ( .A1(n30557), .A2(\xmem_data[0][2] ), .B1(n28291), .B2(
        \xmem_data[1][2] ), .ZN(n28596) );
  AOI22_X1 U31729 ( .A1(n3307), .A2(\xmem_data[2][2] ), .B1(n24223), .B2(
        \xmem_data[3][2] ), .ZN(n28595) );
  AOI22_X1 U31730 ( .A1(n3171), .A2(\xmem_data[4][2] ), .B1(n20488), .B2(
        \xmem_data[5][2] ), .ZN(n28594) );
  AOI22_X1 U31731 ( .A1(n20826), .A2(\xmem_data[6][2] ), .B1(n30524), .B2(
        \xmem_data[7][2] ), .ZN(n28593) );
  NAND4_X1 U31732 ( .A1(n28596), .A2(n28595), .A3(n28594), .A4(n28593), .ZN(
        n28607) );
  AOI22_X1 U31733 ( .A1(n3322), .A2(\xmem_data[16][2] ), .B1(n30550), .B2(
        \xmem_data[17][2] ), .ZN(n28600) );
  AOI22_X1 U31734 ( .A1(n25451), .A2(\xmem_data[18][2] ), .B1(n13474), .B2(
        \xmem_data[19][2] ), .ZN(n28599) );
  AOI22_X1 U31735 ( .A1(n30551), .A2(\xmem_data[20][2] ), .B1(n27863), .B2(
        \xmem_data[21][2] ), .ZN(n28598) );
  AOI22_X1 U31736 ( .A1(n30508), .A2(\xmem_data[22][2] ), .B1(n30552), .B2(
        \xmem_data[23][2] ), .ZN(n28597) );
  NAND4_X1 U31737 ( .A1(n28600), .A2(n28599), .A3(n28598), .A4(n28597), .ZN(
        n28606) );
  AOI22_X1 U31738 ( .A1(n28298), .A2(\xmem_data[24][2] ), .B1(n30541), .B2(
        \xmem_data[25][2] ), .ZN(n28604) );
  AOI22_X1 U31739 ( .A1(n27755), .A2(\xmem_data[26][2] ), .B1(n30542), .B2(
        \xmem_data[27][2] ), .ZN(n28603) );
  AOI22_X1 U31740 ( .A1(n24708), .A2(\xmem_data[28][2] ), .B1(n30544), .B2(
        \xmem_data[29][2] ), .ZN(n28602) );
  AOI22_X1 U31741 ( .A1(n17044), .A2(\xmem_data[30][2] ), .B1(n30545), .B2(
        \xmem_data[31][2] ), .ZN(n28601) );
  NAND4_X1 U31742 ( .A1(n28604), .A2(n28603), .A3(n28602), .A4(n28601), .ZN(
        n28605) );
  OR4_X1 U31743 ( .A1(n28608), .A2(n28607), .A3(n28606), .A4(n28605), .ZN(
        n28609) );
  NAND2_X1 U31744 ( .A1(n28609), .A2(n30563), .ZN(n28633) );
  AOI22_X1 U31745 ( .A1(n30592), .A2(\xmem_data[108][2] ), .B1(n3222), .B2(
        \xmem_data[109][2] ), .ZN(n28613) );
  AOI22_X1 U31746 ( .A1(n3348), .A2(\xmem_data[106][2] ), .B1(n30589), .B2(
        \xmem_data[107][2] ), .ZN(n28612) );
  AOI22_X1 U31747 ( .A1(n30588), .A2(\xmem_data[104][2] ), .B1(n30571), .B2(
        \xmem_data[105][2] ), .ZN(n28611) );
  AOI22_X1 U31748 ( .A1(n30593), .A2(\xmem_data[110][2] ), .B1(n20992), .B2(
        \xmem_data[111][2] ), .ZN(n28610) );
  NAND4_X1 U31749 ( .A1(n28613), .A2(n28612), .A3(n28611), .A4(n28610), .ZN(
        n28631) );
  AOI22_X1 U31750 ( .A1(n24647), .A2(\xmem_data[96][2] ), .B1(n25581), .B2(
        \xmem_data[97][2] ), .ZN(n28617) );
  AOI22_X1 U31751 ( .A1(n30600), .A2(\xmem_data[98][2] ), .B1(n30599), .B2(
        \xmem_data[99][2] ), .ZN(n28616) );
  AOI22_X1 U31752 ( .A1(n22719), .A2(\xmem_data[100][2] ), .B1(n25359), .B2(
        \xmem_data[101][2] ), .ZN(n28615) );
  AOI22_X1 U31753 ( .A1(n21060), .A2(\xmem_data[102][2] ), .B1(n30601), .B2(
        \xmem_data[103][2] ), .ZN(n28614) );
  NAND4_X1 U31754 ( .A1(n28617), .A2(n28616), .A3(n28615), .A4(n28614), .ZN(
        n28629) );
  AOI22_X1 U31755 ( .A1(n20718), .A2(\xmem_data[122][2] ), .B1(n30615), .B2(
        \xmem_data[123][2] ), .ZN(n28621) );
  AOI22_X1 U31756 ( .A1(n30614), .A2(\xmem_data[120][2] ), .B1(n30613), .B2(
        \xmem_data[121][2] ), .ZN(n28620) );
  AOI22_X1 U31757 ( .A1(n30617), .A2(\xmem_data[126][2] ), .B1(n30616), .B2(
        \xmem_data[127][2] ), .ZN(n28619) );
  AOI22_X1 U31758 ( .A1(n20585), .A2(\xmem_data[124][2] ), .B1(n20505), .B2(
        \xmem_data[125][2] ), .ZN(n28618) );
  NAND4_X1 U31759 ( .A1(n28621), .A2(n28620), .A3(n28619), .A4(n28618), .ZN(
        n28627) );
  AOI22_X1 U31760 ( .A1(n30606), .A2(\xmem_data[112][2] ), .B1(n30882), .B2(
        \xmem_data[113][2] ), .ZN(n28625) );
  AOI22_X1 U31761 ( .A1(n3282), .A2(\xmem_data[114][2] ), .B1(n31252), .B2(
        \xmem_data[115][2] ), .ZN(n28624) );
  AOI22_X1 U31762 ( .A1(n30607), .A2(\xmem_data[116][2] ), .B1(n13475), .B2(
        \xmem_data[117][2] ), .ZN(n28623) );
  AOI22_X1 U31763 ( .A1(n30608), .A2(\xmem_data[118][2] ), .B1(n27513), .B2(
        \xmem_data[119][2] ), .ZN(n28622) );
  NAND4_X1 U31764 ( .A1(n28625), .A2(n28624), .A3(n28623), .A4(n28622), .ZN(
        n28626) );
  OR2_X1 U31765 ( .A1(n28627), .A2(n28626), .ZN(n28628) );
  OR2_X1 U31766 ( .A1(n28629), .A2(n28628), .ZN(n28630) );
  OAI21_X1 U31767 ( .B1(n28631), .B2(n28630), .A(n30626), .ZN(n28632) );
  XNOR2_X1 U31768 ( .A(n32554), .B(\fmem_data[26][3] ), .ZN(n31399) );
  OAI22_X1 U31769 ( .A1(n32144), .A2(n32780), .B1(n31399), .B2(n32779), .ZN(
        n33986) );
  XNOR2_X1 U31770 ( .A(n33750), .B(\fmem_data[17][3] ), .ZN(n32069) );
  XNOR2_X1 U31771 ( .A(n31512), .B(\fmem_data[17][3] ), .ZN(n32133) );
  OAI22_X1 U31772 ( .A1(n32069), .A2(n33249), .B1(n33250), .B2(n32133), .ZN(
        n33687) );
  AOI22_X1 U31773 ( .A1(n30076), .A2(\xmem_data[80][0] ), .B1(n29487), .B2(
        \xmem_data[81][0] ), .ZN(n28637) );
  AOI22_X1 U31774 ( .A1(n3249), .A2(\xmem_data[68][0] ), .B1(n27761), .B2(
        \xmem_data[69][0] ), .ZN(n28636) );
  AOI22_X1 U31775 ( .A1(n27710), .A2(\xmem_data[92][0] ), .B1(n30106), .B2(
        \xmem_data[93][0] ), .ZN(n28650) );
  AOI22_X1 U31776 ( .A1(n28725), .A2(\xmem_data[84][0] ), .B1(n28724), .B2(
        \xmem_data[85][0] ), .ZN(n28638) );
  INV_X1 U31777 ( .A(n28638), .ZN(n28647) );
  AOI22_X1 U31778 ( .A1(n28727), .A2(\xmem_data[86][0] ), .B1(n20826), .B2(
        \xmem_data[87][0] ), .ZN(n28640) );
  AOI22_X1 U31779 ( .A1(n29786), .A2(\xmem_data[88][0] ), .B1(n3124), .B2(
        \xmem_data[89][0] ), .ZN(n28639) );
  NAND2_X1 U31780 ( .A1(n28640), .A2(n28639), .ZN(n28646) );
  AOI22_X1 U31781 ( .A1(n28719), .A2(\xmem_data[90][0] ), .B1(n28718), .B2(
        \xmem_data[91][0] ), .ZN(n28644) );
  AOI22_X1 U31782 ( .A1(n28720), .A2(\xmem_data[82][0] ), .B1(n3151), .B2(
        \xmem_data[83][0] ), .ZN(n28643) );
  AOI22_X1 U31783 ( .A1(n28744), .A2(\xmem_data[70][0] ), .B1(n28743), .B2(
        \xmem_data[71][0] ), .ZN(n28642) );
  AOI22_X1 U31784 ( .A1(n3244), .A2(\xmem_data[66][0] ), .B1(n3126), .B2(
        \xmem_data[67][0] ), .ZN(n28641) );
  NAND4_X1 U31785 ( .A1(n28644), .A2(n28643), .A3(n28642), .A4(n28641), .ZN(
        n28645) );
  NOR3_X1 U31786 ( .A1(n28647), .A2(n28646), .A3(n28645), .ZN(n28649) );
  AOI22_X1 U31787 ( .A1(n28138), .A2(\xmem_data[94][0] ), .B1(n28733), .B2(
        \xmem_data[95][0] ), .ZN(n28648) );
  NAND4_X1 U31788 ( .A1(n28651), .A2(n28650), .A3(n28649), .A4(n28648), .ZN(
        n28664) );
  AOI22_X1 U31789 ( .A1(n28740), .A2(\xmem_data[64][0] ), .B1(n29761), .B2(
        \xmem_data[65][0] ), .ZN(n28652) );
  AOI22_X1 U31790 ( .A1(n30764), .A2(\xmem_data[78][0] ), .B1(n28687), .B2(
        \xmem_data[79][0] ), .ZN(n28653) );
  INV_X1 U31791 ( .A(n28653), .ZN(n28660) );
  AOI22_X1 U31792 ( .A1(n28753), .A2(\xmem_data[74][0] ), .B1(n30666), .B2(
        \xmem_data[75][0] ), .ZN(n28655) );
  AOI22_X1 U31793 ( .A1(n29604), .A2(\xmem_data[72][0] ), .B1(n29648), .B2(
        \xmem_data[73][0] ), .ZN(n28654) );
  NAND2_X1 U31794 ( .A1(n28655), .A2(n28654), .ZN(n28659) );
  NAND2_X1 U31795 ( .A1(n3188), .A2(\xmem_data[77][0] ), .ZN(n28657) );
  NAND2_X1 U31796 ( .A1(n3165), .A2(\xmem_data[76][0] ), .ZN(n28656) );
  NAND2_X1 U31797 ( .A1(n28657), .A2(n28656), .ZN(n28658) );
  NOR3_X1 U31798 ( .A1(n28660), .A2(n28659), .A3(n28658), .ZN(n28661) );
  NAND2_X1 U31799 ( .A1(n28652), .A2(n28661), .ZN(n28663) );
  OAI21_X1 U31800 ( .B1(n28664), .B2(n28663), .A(n28662), .ZN(n28799) );
  AOI22_X1 U31801 ( .A1(n28739), .A2(\xmem_data[36][0] ), .B1(n28145), .B2(
        \xmem_data[37][0] ), .ZN(n28666) );
  INV_X1 U31802 ( .A(n28666), .ZN(n28676) );
  NAND2_X1 U31803 ( .A1(n3197), .A2(\xmem_data[33][0] ), .ZN(n28669) );
  NAND2_X1 U31804 ( .A1(n27771), .A2(\xmem_data[32][0] ), .ZN(n28668) );
  NAND2_X1 U31805 ( .A1(n28669), .A2(n28668), .ZN(n28675) );
  AOI22_X1 U31806 ( .A1(n28670), .A2(\xmem_data[34][0] ), .B1(n29350), .B2(
        \xmem_data[35][0] ), .ZN(n28673) );
  AOI22_X1 U31807 ( .A1(n28744), .A2(\xmem_data[38][0] ), .B1(n28671), .B2(
        \xmem_data[39][0] ), .ZN(n28672) );
  NAND2_X1 U31808 ( .A1(n28673), .A2(n28672), .ZN(n28674) );
  NOR3_X1 U31809 ( .A1(n28676), .A2(n28675), .A3(n28674), .ZN(n28712) );
  AOI22_X1 U31810 ( .A1(n3227), .A2(\xmem_data[58][0] ), .B1(n28677), .B2(
        \xmem_data[59][0] ), .ZN(n28678) );
  INV_X1 U31811 ( .A(n28678), .ZN(n28679) );
  AOI21_X1 U31812 ( .B1(\xmem_data[48][0] ), .B2(n27713), .A(n28679), .ZN(
        n28683) );
  AOI22_X1 U31813 ( .A1(n28681), .A2(\xmem_data[54][0] ), .B1(n23730), .B2(
        \xmem_data[55][0] ), .ZN(n28682) );
  AOI22_X1 U31814 ( .A1(n3167), .A2(\xmem_data[44][0] ), .B1(n3191), .B2(
        \xmem_data[45][0] ), .ZN(n28693) );
  AOI22_X1 U31815 ( .A1(n27811), .A2(\xmem_data[40][0] ), .B1(n30301), .B2(
        \xmem_data[41][0] ), .ZN(n28692) );
  AOI22_X1 U31816 ( .A1(n28686), .A2(\xmem_data[42][0] ), .B1(n27945), .B2(
        \xmem_data[43][0] ), .ZN(n28691) );
  AND2_X1 U31817 ( .A1(n28687), .A2(\xmem_data[47][0] ), .ZN(n28688) );
  AOI21_X1 U31818 ( .B1(n28689), .B2(\xmem_data[46][0] ), .A(n28688), .ZN(
        n28690) );
  NAND4_X1 U31819 ( .A1(n28693), .A2(n28692), .A3(n28691), .A4(n28690), .ZN(
        n28694) );
  NOR2_X1 U31820 ( .A1(n28695), .A2(n28694), .ZN(n28711) );
  AOI22_X1 U31821 ( .A1(n29724), .A2(\xmem_data[52][0] ), .B1(n28696), .B2(
        \xmem_data[53][0] ), .ZN(n28699) );
  AOI22_X1 U31822 ( .A1(n28765), .A2(\xmem_data[56][0] ), .B1(n29497), .B2(
        \xmem_data[57][0] ), .ZN(n28698) );
  NAND2_X1 U31823 ( .A1(n29626), .A2(\xmem_data[60][0] ), .ZN(n28697) );
  NAND2_X1 U31824 ( .A1(n29640), .A2(\xmem_data[49][0] ), .ZN(n28706) );
  AOI22_X1 U31825 ( .A1(n28702), .A2(\xmem_data[50][0] ), .B1(n28701), .B2(
        \xmem_data[51][0] ), .ZN(n28705) );
  NAND2_X1 U31826 ( .A1(n29672), .A2(\xmem_data[61][0] ), .ZN(n28704) );
  NAND2_X1 U31827 ( .A1(n29627), .A2(\xmem_data[63][0] ), .ZN(n28703) );
  NAND4_X1 U31828 ( .A1(n28706), .A2(n28705), .A3(n28704), .A4(n28703), .ZN(
        n28707) );
  NOR2_X1 U31829 ( .A1(n28708), .A2(n28707), .ZN(n28709) );
  NAND4_X1 U31830 ( .A1(n28712), .A2(n28711), .A3(n28710), .A4(n28709), .ZN(
        n28714) );
  NAND2_X1 U31831 ( .A1(n28714), .A2(n28713), .ZN(n28798) );
  NAND2_X1 U31832 ( .A1(n30765), .A2(\xmem_data[113][0] ), .ZN(n28716) );
  NAND2_X1 U31833 ( .A1(n30717), .A2(\xmem_data[112][0] ), .ZN(n28715) );
  NAND2_X1 U31834 ( .A1(n28716), .A2(n28715), .ZN(n28732) );
  AOI22_X1 U31835 ( .A1(n28765), .A2(\xmem_data[120][0] ), .B1(n3124), .B2(
        \xmem_data[121][0] ), .ZN(n28723) );
  AOI22_X1 U31836 ( .A1(n28719), .A2(\xmem_data[122][0] ), .B1(n28718), .B2(
        \xmem_data[123][0] ), .ZN(n28722) );
  AOI22_X1 U31837 ( .A1(n28720), .A2(\xmem_data[114][0] ), .B1(n3337), .B2(
        \xmem_data[115][0] ), .ZN(n28721) );
  AOI22_X1 U31838 ( .A1(n28725), .A2(\xmem_data[116][0] ), .B1(n28724), .B2(
        \xmem_data[117][0] ), .ZN(n28729) );
  AND2_X1 U31839 ( .A1(n28467), .A2(\xmem_data[119][0] ), .ZN(n28726) );
  AOI21_X1 U31840 ( .B1(n28727), .B2(\xmem_data[118][0] ), .A(n28726), .ZN(
        n28728) );
  NAND2_X1 U31841 ( .A1(n28729), .A2(n28728), .ZN(n28730) );
  NOR3_X1 U31842 ( .A1(n28732), .A2(n28731), .A3(n28730), .ZN(n28737) );
  AOI22_X1 U31843 ( .A1(n29423), .A2(\xmem_data[126][0] ), .B1(n28733), .B2(
        \xmem_data[127][0] ), .ZN(n28736) );
  AOI22_X1 U31844 ( .A1(n29421), .A2(\xmem_data[124][0] ), .B1(n26616), .B2(
        \xmem_data[125][0] ), .ZN(n28735) );
  AOI22_X1 U31845 ( .A1(n3249), .A2(\xmem_data[100][0] ), .B1(n29646), .B2(
        \xmem_data[101][0] ), .ZN(n28750) );
  AOI22_X1 U31846 ( .A1(n28740), .A2(\xmem_data[96][0] ), .B1(n29556), .B2(
        \xmem_data[97][0] ), .ZN(n28749) );
  AOI22_X1 U31847 ( .A1(n3244), .A2(\xmem_data[98][0] ), .B1(n3126), .B2(
        \xmem_data[99][0] ), .ZN(n28742) );
  AOI22_X1 U31848 ( .A1(n28744), .A2(\xmem_data[102][0] ), .B1(n28743), .B2(
        \xmem_data[103][0] ), .ZN(n28745) );
  NOR2_X1 U31849 ( .A1(n28747), .A2(n28746), .ZN(n28748) );
  NAND3_X1 U31850 ( .A1(n28750), .A2(n28749), .A3(n28748), .ZN(n28761) );
  AOI22_X1 U31851 ( .A1(n27811), .A2(\xmem_data[104][0] ), .B1(n26884), .B2(
        \xmem_data[105][0] ), .ZN(n28759) );
  AOI22_X1 U31852 ( .A1(n28753), .A2(\xmem_data[106][0] ), .B1(n3466), .B2(
        \xmem_data[107][0] ), .ZN(n28758) );
  AOI22_X1 U31853 ( .A1(n3163), .A2(\xmem_data[108][0] ), .B1(n3188), .B2(
        \xmem_data[109][0] ), .ZN(n28757) );
  AOI22_X1 U31854 ( .A1(n28755), .A2(\xmem_data[110][0] ), .B1(n28754), .B2(
        \xmem_data[111][0] ), .ZN(n28756) );
  NAND4_X1 U31855 ( .A1(n28759), .A2(n28758), .A3(n28757), .A4(n28756), .ZN(
        n28760) );
  OR2_X1 U31856 ( .A1(n28761), .A2(n28760), .ZN(n28763) );
  AOI22_X1 U31857 ( .A1(n28765), .A2(\xmem_data[24][0] ), .B1(n27743), .B2(
        \xmem_data[25][0] ), .ZN(n28770) );
  AOI22_X1 U31858 ( .A1(n3227), .A2(\xmem_data[26][0] ), .B1(n3144), .B2(
        \xmem_data[27][0] ), .ZN(n28769) );
  AOI22_X1 U31859 ( .A1(n27710), .A2(\xmem_data[28][0] ), .B1(n28766), .B2(
        \xmem_data[29][0] ), .ZN(n28768) );
  AOI22_X1 U31860 ( .A1(n29790), .A2(\xmem_data[30][0] ), .B1(n30278), .B2(
        \xmem_data[31][0] ), .ZN(n28767) );
  AOI22_X1 U31861 ( .A1(n29815), .A2(\xmem_data[16][0] ), .B1(n30266), .B2(
        \xmem_data[17][0] ), .ZN(n28771) );
  INV_X1 U31862 ( .A(n28771), .ZN(n28777) );
  AOI22_X1 U31863 ( .A1(n29819), .A2(\xmem_data[20][0] ), .B1(n27805), .B2(
        \xmem_data[21][0] ), .ZN(n28775) );
  AOI22_X1 U31864 ( .A1(n29464), .A2(\xmem_data[22][0] ), .B1(n28772), .B2(
        \xmem_data[23][0] ), .ZN(n28774) );
  AOI22_X1 U31865 ( .A1(n28702), .A2(\xmem_data[18][0] ), .B1(n28701), .B2(
        \xmem_data[19][0] ), .ZN(n28773) );
  NOR2_X1 U31866 ( .A1(n28777), .A2(n28776), .ZN(n28793) );
  AOI22_X1 U31867 ( .A1(n30302), .A2(\xmem_data[8][0] ), .B1(n29592), .B2(
        \xmem_data[9][0] ), .ZN(n28785) );
  AOI22_X1 U31868 ( .A1(n28780), .A2(\xmem_data[10][0] ), .B1(n30948), .B2(
        \xmem_data[11][0] ), .ZN(n28784) );
  AOI22_X1 U31869 ( .A1(n3166), .A2(\xmem_data[12][0] ), .B1(n3187), .B2(
        \xmem_data[13][0] ), .ZN(n28783) );
  AOI22_X1 U31870 ( .A1(n30062), .A2(\xmem_data[14][0] ), .B1(n28781), .B2(
        \xmem_data[15][0] ), .ZN(n28782) );
  AOI22_X1 U31871 ( .A1(n28787), .A2(\xmem_data[0][0] ), .B1(n30776), .B2(
        \xmem_data[1][0] ), .ZN(n28792) );
  AOI22_X1 U31872 ( .A1(n3244), .A2(\xmem_data[2][0] ), .B1(n30295), .B2(
        \xmem_data[3][0] ), .ZN(n28791) );
  AOI22_X1 U31873 ( .A1(n28180), .A2(\xmem_data[4][0] ), .B1(n28665), .B2(
        \xmem_data[5][0] ), .ZN(n28790) );
  AOI22_X1 U31874 ( .A1(n28788), .A2(\xmem_data[6][0] ), .B1(n27514), .B2(
        \xmem_data[7][0] ), .ZN(n28789) );
  NAND4_X1 U31875 ( .A1(n3857), .A2(n28793), .A3(n3156), .A4(n3515), .ZN(
        n28795) );
  NAND2_X1 U31876 ( .A1(n28795), .A2(n28794), .ZN(n28796) );
  NAND4_X2 U31877 ( .A1(n28799), .A2(n28798), .A3(n28797), .A4(n28796), .ZN(
        n36313) );
  INV_X1 U31878 ( .A(n34932), .ZN(n28800) );
  AND2_X1 U31879 ( .A1(n36313), .A2(n28800), .ZN(n33686) );
  AOI22_X1 U31880 ( .A1(n30849), .A2(\xmem_data[16][1] ), .B1(n21009), .B2(
        \xmem_data[17][1] ), .ZN(n28804) );
  AOI22_X1 U31881 ( .A1(n31315), .A2(\xmem_data[18][1] ), .B1(n14975), .B2(
        \xmem_data[19][1] ), .ZN(n28803) );
  AOI22_X1 U31882 ( .A1(n20734), .A2(\xmem_data[20][1] ), .B1(n27981), .B2(
        \xmem_data[21][1] ), .ZN(n28802) );
  AOI22_X1 U31883 ( .A1(n30674), .A2(\xmem_data[22][1] ), .B1(n22727), .B2(
        \xmem_data[23][1] ), .ZN(n28801) );
  NAND4_X1 U31884 ( .A1(n28804), .A2(n28803), .A3(n28802), .A4(n28801), .ZN(
        n28813) );
  AOI22_X1 U31885 ( .A1(n24157), .A2(\xmem_data[6][1] ), .B1(n24212), .B2(
        \xmem_data[7][1] ), .ZN(n28811) );
  AOI22_X1 U31886 ( .A1(n3342), .A2(\xmem_data[0][1] ), .B1(n30550), .B2(
        \xmem_data[1][1] ), .ZN(n28805) );
  INV_X1 U31887 ( .A(n28805), .ZN(n28809) );
  AOI22_X1 U31888 ( .A1(n23813), .A2(\xmem_data[4][1] ), .B1(n30854), .B2(
        \xmem_data[5][1] ), .ZN(n28807) );
  NAND2_X1 U31889 ( .A1(n25377), .A2(\xmem_data[2][1] ), .ZN(n28806) );
  NAND2_X1 U31890 ( .A1(n28807), .A2(n28806), .ZN(n28808) );
  NOR2_X1 U31891 ( .A1(n28809), .A2(n28808), .ZN(n28810) );
  NAND2_X1 U31892 ( .A1(n28811), .A2(n28810), .ZN(n28812) );
  OR2_X1 U31893 ( .A1(n28813), .A2(n28812), .ZN(n28825) );
  AOI22_X1 U31894 ( .A1(n27502), .A2(\xmem_data[28][1] ), .B1(n3222), .B2(
        \xmem_data[29][1] ), .ZN(n28817) );
  AOI22_X1 U31895 ( .A1(n30864), .A2(\xmem_data[26][1] ), .B1(n30863), .B2(
        \xmem_data[27][1] ), .ZN(n28816) );
  AOI22_X1 U31896 ( .A1(n30862), .A2(\xmem_data[24][1] ), .B1(n30861), .B2(
        \xmem_data[25][1] ), .ZN(n28815) );
  AOI22_X1 U31897 ( .A1(n22708), .A2(\xmem_data[30][1] ), .B1(n22710), .B2(
        \xmem_data[31][1] ), .ZN(n28814) );
  NAND4_X1 U31898 ( .A1(n28817), .A2(n28816), .A3(n28815), .A4(n28814), .ZN(
        n28823) );
  AOI22_X1 U31899 ( .A1(n25459), .A2(\xmem_data[8][1] ), .B1(n29309), .B2(
        \xmem_data[9][1] ), .ZN(n28821) );
  AOI22_X1 U31900 ( .A1(n30948), .A2(\xmem_data[10][1] ), .B1(n24457), .B2(
        \xmem_data[11][1] ), .ZN(n28820) );
  AOI22_X1 U31901 ( .A1(n24547), .A2(\xmem_data[12][1] ), .B1(n24219), .B2(
        \xmem_data[13][1] ), .ZN(n28819) );
  AOI22_X1 U31902 ( .A1(n30872), .A2(\xmem_data[14][1] ), .B1(n30871), .B2(
        \xmem_data[15][1] ), .ZN(n28818) );
  NAND4_X1 U31903 ( .A1(n28821), .A2(n28820), .A3(n28819), .A4(n28818), .ZN(
        n28822) );
  OR2_X1 U31904 ( .A1(n28823), .A2(n28822), .ZN(n28824) );
  NOR2_X1 U31905 ( .A1(n28825), .A2(n28824), .ZN(n28826) );
  AOI22_X1 U31906 ( .A1(n30606), .A2(\xmem_data[96][1] ), .B1(n22759), .B2(
        \xmem_data[97][1] ), .ZN(n28830) );
  AOI22_X1 U31907 ( .A1(n3128), .A2(\xmem_data[98][1] ), .B1(n28007), .B2(
        \xmem_data[99][1] ), .ZN(n28829) );
  AOI22_X1 U31908 ( .A1(n27551), .A2(\xmem_data[100][1] ), .B1(n27988), .B2(
        \xmem_data[101][1] ), .ZN(n28828) );
  AOI22_X1 U31909 ( .A1(n30943), .A2(\xmem_data[102][1] ), .B1(n13168), .B2(
        \xmem_data[103][1] ), .ZN(n28827) );
  NAND4_X1 U31910 ( .A1(n28830), .A2(n28829), .A3(n28828), .A4(n28827), .ZN(
        n28846) );
  AOI22_X1 U31911 ( .A1(n30514), .A2(\xmem_data[104][1] ), .B1(n22741), .B2(
        \xmem_data[105][1] ), .ZN(n28834) );
  AOI22_X1 U31912 ( .A1(n29237), .A2(\xmem_data[106][1] ), .B1(n24134), .B2(
        \xmem_data[107][1] ), .ZN(n28833) );
  AOI22_X1 U31913 ( .A1(n30949), .A2(\xmem_data[108][1] ), .B1(n28427), .B2(
        \xmem_data[109][1] ), .ZN(n28832) );
  AOI22_X1 U31914 ( .A1(n30950), .A2(\xmem_data[110][1] ), .B1(n25435), .B2(
        \xmem_data[111][1] ), .ZN(n28831) );
  NAND4_X1 U31915 ( .A1(n28834), .A2(n28833), .A3(n28832), .A4(n28831), .ZN(
        n28845) );
  AOI22_X1 U31916 ( .A1(n30956), .A2(\xmem_data[112][1] ), .B1(n30955), .B2(
        \xmem_data[113][1] ), .ZN(n28838) );
  AOI22_X1 U31917 ( .A1(n3337), .A2(\xmem_data[114][1] ), .B1(n28495), .B2(
        \xmem_data[115][1] ), .ZN(n28837) );
  AOI22_X1 U31918 ( .A1(n25582), .A2(\xmem_data[116][1] ), .B1(n31256), .B2(
        \xmem_data[117][1] ), .ZN(n28836) );
  AOI22_X1 U31919 ( .A1(n23730), .A2(\xmem_data[118][1] ), .B1(n24686), .B2(
        \xmem_data[119][1] ), .ZN(n28835) );
  NAND4_X1 U31920 ( .A1(n28838), .A2(n28837), .A3(n28836), .A4(n28835), .ZN(
        n28844) );
  AOI22_X1 U31921 ( .A1(n17030), .A2(\xmem_data[120][1] ), .B1(n25357), .B2(
        \xmem_data[121][1] ), .ZN(n28842) );
  AOI22_X1 U31922 ( .A1(n3332), .A2(\xmem_data[122][1] ), .B1(n20568), .B2(
        \xmem_data[123][1] ), .ZN(n28841) );
  AOI22_X1 U31923 ( .A1(n30962), .A2(\xmem_data[124][1] ), .B1(n3217), .B2(
        \xmem_data[125][1] ), .ZN(n28840) );
  AOI22_X1 U31924 ( .A1(n30964), .A2(\xmem_data[126][1] ), .B1(n30963), .B2(
        \xmem_data[127][1] ), .ZN(n28839) );
  NAND4_X1 U31925 ( .A1(n28842), .A2(n28841), .A3(n28840), .A4(n28839), .ZN(
        n28843) );
  OR4_X1 U31926 ( .A1(n28846), .A2(n28845), .A3(n28844), .A4(n28843), .ZN(
        n28868) );
  AOI22_X1 U31927 ( .A1(n29174), .A2(\xmem_data[64][1] ), .B1(n27994), .B2(
        \xmem_data[65][1] ), .ZN(n28850) );
  AOI22_X1 U31928 ( .A1(n3129), .A2(\xmem_data[66][1] ), .B1(n28045), .B2(
        \xmem_data[67][1] ), .ZN(n28849) );
  AOI22_X1 U31929 ( .A1(n27551), .A2(\xmem_data[68][1] ), .B1(n27988), .B2(
        \xmem_data[69][1] ), .ZN(n28848) );
  AOI22_X1 U31930 ( .A1(n30943), .A2(\xmem_data[70][1] ), .B1(n13168), .B2(
        \xmem_data[71][1] ), .ZN(n28847) );
  NAND4_X1 U31931 ( .A1(n28850), .A2(n28849), .A3(n28848), .A4(n28847), .ZN(
        n28866) );
  AOI22_X1 U31932 ( .A1(n3176), .A2(\xmem_data[72][1] ), .B1(n30513), .B2(
        \xmem_data[73][1] ), .ZN(n28854) );
  AOI22_X1 U31933 ( .A1(n3466), .A2(\xmem_data[74][1] ), .B1(n24457), .B2(
        \xmem_data[75][1] ), .ZN(n28853) );
  AOI22_X1 U31934 ( .A1(n30949), .A2(\xmem_data[76][1] ), .B1(n25715), .B2(
        \xmem_data[77][1] ), .ZN(n28852) );
  AOI22_X1 U31935 ( .A1(n30950), .A2(\xmem_data[78][1] ), .B1(n28380), .B2(
        \xmem_data[79][1] ), .ZN(n28851) );
  NAND4_X1 U31936 ( .A1(n28854), .A2(n28853), .A3(n28852), .A4(n28851), .ZN(
        n28865) );
  AOI22_X1 U31937 ( .A1(n30956), .A2(\xmem_data[80][1] ), .B1(n30955), .B2(
        \xmem_data[81][1] ), .ZN(n28858) );
  AOI22_X1 U31938 ( .A1(n30686), .A2(\xmem_data[82][1] ), .B1(n24622), .B2(
        \xmem_data[83][1] ), .ZN(n28857) );
  AOI22_X1 U31939 ( .A1(n27847), .A2(\xmem_data[84][1] ), .B1(n27981), .B2(
        \xmem_data[85][1] ), .ZN(n28856) );
  AOI22_X1 U31940 ( .A1(n21060), .A2(\xmem_data[86][1] ), .B1(n24524), .B2(
        \xmem_data[87][1] ), .ZN(n28855) );
  NAND4_X1 U31941 ( .A1(n28858), .A2(n28857), .A3(n28856), .A4(n28855), .ZN(
        n28864) );
  AOI22_X1 U31942 ( .A1(n30962), .A2(\xmem_data[92][1] ), .B1(n3220), .B2(
        \xmem_data[93][1] ), .ZN(n28862) );
  AOI22_X1 U31943 ( .A1(n3332), .A2(\xmem_data[90][1] ), .B1(n20711), .B2(
        \xmem_data[91][1] ), .ZN(n28861) );
  AOI22_X1 U31944 ( .A1(n24526), .A2(\xmem_data[88][1] ), .B1(n31346), .B2(
        \xmem_data[89][1] ), .ZN(n28860) );
  AOI22_X1 U31945 ( .A1(n30964), .A2(\xmem_data[94][1] ), .B1(n30963), .B2(
        \xmem_data[95][1] ), .ZN(n28859) );
  NAND4_X1 U31946 ( .A1(n28862), .A2(n28861), .A3(n28860), .A4(n28859), .ZN(
        n28863) );
  OR4_X1 U31947 ( .A1(n28866), .A2(n28865), .A3(n28864), .A4(n28863), .ZN(
        n28867) );
  AOI22_X1 U31948 ( .A1(n30976), .A2(n28868), .B1(n30974), .B2(n28867), .ZN(
        n28892) );
  AOI22_X1 U31949 ( .A1(n30883), .A2(\xmem_data[32][1] ), .B1(n30882), .B2(
        \xmem_data[33][1] ), .ZN(n28872) );
  AOI22_X1 U31950 ( .A1(n3375), .A2(\xmem_data[34][1] ), .B1(n25514), .B2(
        \xmem_data[35][1] ), .ZN(n28871) );
  AOI22_X1 U31951 ( .A1(n30885), .A2(\xmem_data[36][1] ), .B1(n30884), .B2(
        \xmem_data[37][1] ), .ZN(n28870) );
  AOI22_X1 U31952 ( .A1(n30886), .A2(\xmem_data[38][1] ), .B1(n22702), .B2(
        \xmem_data[39][1] ), .ZN(n28869) );
  NAND4_X1 U31953 ( .A1(n28872), .A2(n28871), .A3(n28870), .A4(n28869), .ZN(
        n28888) );
  AOI22_X1 U31954 ( .A1(n30891), .A2(\xmem_data[40][1] ), .B1(n14898), .B2(
        \xmem_data[41][1] ), .ZN(n28876) );
  AOI22_X1 U31955 ( .A1(n23795), .A2(\xmem_data[42][1] ), .B1(n28335), .B2(
        \xmem_data[43][1] ), .ZN(n28875) );
  AOI22_X1 U31956 ( .A1(n23764), .A2(\xmem_data[44][1] ), .B1(n16989), .B2(
        \xmem_data[45][1] ), .ZN(n28874) );
  AOI22_X1 U31957 ( .A1(n30893), .A2(\xmem_data[46][1] ), .B1(n25399), .B2(
        \xmem_data[47][1] ), .ZN(n28873) );
  NAND4_X1 U31958 ( .A1(n28876), .A2(n28875), .A3(n28874), .A4(n28873), .ZN(
        n28887) );
  AOI22_X1 U31959 ( .A1(n24220), .A2(\xmem_data[48][1] ), .B1(n30898), .B2(
        \xmem_data[49][1] ), .ZN(n28880) );
  AOI22_X1 U31960 ( .A1(n3302), .A2(\xmem_data[50][1] ), .B1(n28495), .B2(
        \xmem_data[51][1] ), .ZN(n28879) );
  AOI22_X1 U31961 ( .A1(n20552), .A2(\xmem_data[52][1] ), .B1(n11008), .B2(
        \xmem_data[53][1] ), .ZN(n28878) );
  AOI22_X1 U31962 ( .A1(n30901), .A2(\xmem_data[54][1] ), .B1(n30900), .B2(
        \xmem_data[55][1] ), .ZN(n28877) );
  NAND4_X1 U31963 ( .A1(n28880), .A2(n28879), .A3(n28878), .A4(n28877), .ZN(
        n28886) );
  AOI22_X1 U31964 ( .A1(n30909), .A2(\xmem_data[56][1] ), .B1(n30908), .B2(
        \xmem_data[57][1] ), .ZN(n28884) );
  AOI22_X1 U31965 ( .A1(n3351), .A2(\xmem_data[58][1] ), .B1(n27437), .B2(
        \xmem_data[59][1] ), .ZN(n28883) );
  AOI22_X1 U31966 ( .A1(n30906), .A2(\xmem_data[60][1] ), .B1(n3218), .B2(
        \xmem_data[61][1] ), .ZN(n28882) );
  AOI22_X1 U31967 ( .A1(n28733), .A2(\xmem_data[62][1] ), .B1(n24207), .B2(
        \xmem_data[63][1] ), .ZN(n28881) );
  NAND4_X1 U31968 ( .A1(n28884), .A2(n28883), .A3(n28882), .A4(n28881), .ZN(
        n28885) );
  OR4_X1 U31969 ( .A1(n28888), .A2(n28887), .A3(n28886), .A4(n28885), .ZN(
        n28890) );
  NOR2_X1 U31970 ( .A1(n30879), .A2(n39029), .ZN(n28889) );
  AOI21_X1 U31971 ( .B1(n28890), .B2(n30918), .A(n3894), .ZN(n28891) );
  XNOR2_X1 U31972 ( .A(n31452), .B(\fmem_data[10][3] ), .ZN(n32571) );
  OAI22_X1 U31973 ( .A1(n33590), .A2(n33690), .B1(n32571), .B2(n34736), .ZN(
        n33685) );
  OAI21_X1 U31974 ( .B1(n31466), .B2(n31465), .A(n31467), .ZN(n28894) );
  NAND2_X1 U31975 ( .A1(n31466), .A2(n31465), .ZN(n28893) );
  NAND2_X1 U31976 ( .A1(n28894), .A2(n28893), .ZN(n33625) );
  FA_X1 U31977 ( .A(n28897), .B(n28896), .CI(n28895), .CO(n28917), .S(n33659)
         );
  FA_X1 U31978 ( .A(n28900), .B(n28899), .CI(n28898), .CO(n33628), .S(n33658)
         );
  FA_X1 U31979 ( .A(n28903), .B(n28902), .CI(n28901), .CO(n28922), .S(n33657)
         );
  FA_X1 U31980 ( .A(n28909), .B(n28908), .CI(n3729), .CO(n24842), .S(n30130)
         );
  FA_X1 U31981 ( .A(n28912), .B(n28911), .CI(n28910), .CO(n24841), .S(n30129)
         );
  FA_X1 U31982 ( .A(n28913), .B(n28914), .CI(n28915), .CO(n34169), .S(n33623)
         );
  XNOR2_X1 U31983 ( .A(n28917), .B(n28916), .ZN(n28919) );
  XNOR2_X1 U31984 ( .A(n28921), .B(n28920), .ZN(n28923) );
  XNOR2_X1 U31985 ( .A(n28923), .B(n28922), .ZN(n33621) );
  OAI21_X1 U31986 ( .B1(n31626), .B2(n31624), .A(n31625), .ZN(n28924) );
  NAND2_X1 U31987 ( .A1(n28925), .A2(n28924), .ZN(n34286) );
  FA_X1 U31988 ( .A(n28928), .B(n28927), .CI(n28926), .CO(n31846), .S(n31414)
         );
  FA_X1 U31989 ( .A(n28931), .B(n28930), .CI(n28929), .CO(n30141), .S(n31209)
         );
  FA_X1 U31990 ( .A(n28934), .B(n28933), .CI(n28932), .CO(n30154), .S(n30142)
         );
  XNOR2_X1 U31991 ( .A(n30141), .B(n30142), .ZN(n28939) );
  XNOR2_X1 U31992 ( .A(n31250), .B(\fmem_data[1][3] ), .ZN(n32177) );
  XNOR2_X1 U31993 ( .A(n31892), .B(\fmem_data[1][3] ), .ZN(n33189) );
  FA_X1 U31994 ( .A(n28937), .B(n28936), .CI(n28935), .CO(n28941), .S(n31129)
         );
  XNOR2_X1 U31995 ( .A(n32438), .B(\fmem_data[31][5] ), .ZN(n32190) );
  OAI22_X1 U31996 ( .A1(n32190), .A2(n34945), .B1(n28938), .B2(n34944), .ZN(
        n28940) );
  XNOR2_X1 U31997 ( .A(n28939), .B(n30143), .ZN(n31133) );
  FA_X1 U31998 ( .A(n28942), .B(n28941), .CI(n28940), .CO(n30143), .S(n31406)
         );
  AOI22_X1 U31999 ( .A1(n13474), .A2(\xmem_data[98][3] ), .B1(n20961), .B2(
        \xmem_data[99][3] ), .ZN(n28971) );
  AOI22_X1 U32000 ( .A1(n29009), .A2(\xmem_data[104][3] ), .B1(n29008), .B2(
        \xmem_data[105][3] ), .ZN(n28946) );
  AOI22_X1 U32001 ( .A1(n3213), .A2(\xmem_data[106][3] ), .B1(n29010), .B2(
        \xmem_data[107][3] ), .ZN(n28945) );
  AOI22_X1 U32002 ( .A1(n28427), .A2(\xmem_data[108][3] ), .B1(n29012), .B2(
        \xmem_data[109][3] ), .ZN(n28944) );
  AOI22_X1 U32003 ( .A1(n23776), .A2(\xmem_data[110][3] ), .B1(n24548), .B2(
        \xmem_data[111][3] ), .ZN(n28943) );
  NAND4_X1 U32004 ( .A1(n28946), .A2(n28945), .A3(n28944), .A4(n28943), .ZN(
        n28967) );
  AOI22_X1 U32005 ( .A1(n27988), .A2(\xmem_data[100][3] ), .B1(n27911), .B2(
        \xmem_data[101][3] ), .ZN(n28965) );
  AOI22_X1 U32006 ( .A1(n28947), .A2(\xmem_data[120][3] ), .B1(n3142), .B2(
        \xmem_data[121][3] ), .ZN(n28951) );
  AOI22_X1 U32007 ( .A1(n25360), .A2(\xmem_data[122][3] ), .B1(n29064), .B2(
        \xmem_data[123][3] ), .ZN(n28950) );
  AOI22_X1 U32008 ( .A1(n3220), .A2(\xmem_data[124][3] ), .B1(n29026), .B2(
        \xmem_data[125][3] ), .ZN(n28949) );
  AOI22_X1 U32009 ( .A1(n29028), .A2(\xmem_data[126][3] ), .B1(n29027), .B2(
        \xmem_data[127][3] ), .ZN(n28948) );
  NAND4_X1 U32010 ( .A1(n28951), .A2(n28950), .A3(n28949), .A4(n28948), .ZN(
        n28963) );
  AOI22_X1 U32011 ( .A1(n31275), .A2(\xmem_data[96][3] ), .B1(n28952), .B2(
        \xmem_data[97][3] ), .ZN(n28954) );
  AOI22_X1 U32012 ( .A1(n24639), .A2(\xmem_data[102][3] ), .B1(n28980), .B2(
        \xmem_data[103][3] ), .ZN(n28953) );
  NAND2_X1 U32013 ( .A1(n28954), .A2(n28953), .ZN(n28961) );
  AOI22_X1 U32014 ( .A1(n28327), .A2(\xmem_data[112][3] ), .B1(n28955), .B2(
        \xmem_data[113][3] ), .ZN(n28959) );
  AOI22_X1 U32015 ( .A1(n24622), .A2(\xmem_data[114][3] ), .B1(n24572), .B2(
        \xmem_data[115][3] ), .ZN(n28958) );
  AOI22_X1 U32016 ( .A1(n29017), .A2(\xmem_data[116][3] ), .B1(n29725), .B2(
        \xmem_data[117][3] ), .ZN(n28957) );
  AOI22_X1 U32017 ( .A1(n25440), .A2(\xmem_data[118][3] ), .B1(n25358), .B2(
        \xmem_data[119][3] ), .ZN(n28956) );
  NAND4_X1 U32018 ( .A1(n28959), .A2(n28958), .A3(n28957), .A4(n28956), .ZN(
        n28960) );
  OR2_X1 U32019 ( .A1(n28961), .A2(n28960), .ZN(n28962) );
  NOR2_X1 U32020 ( .A1(n28963), .A2(n28962), .ZN(n28964) );
  NAND2_X1 U32021 ( .A1(n28965), .A2(n28964), .ZN(n28966) );
  NOR2_X1 U32022 ( .A1(n28967), .A2(n28966), .ZN(n28970) );
  INV_X1 U32023 ( .A(n28968), .ZN(n28969) );
  AOI21_X1 U32024 ( .B1(n28971), .B2(n28970), .A(n28969), .ZN(n29007) );
  AOI22_X1 U32025 ( .A1(n25514), .A2(\xmem_data[2][3] ), .B1(n28972), .B2(
        \xmem_data[3][3] ), .ZN(n29005) );
  AOI22_X1 U32026 ( .A1(n28974), .A2(\xmem_data[24][3] ), .B1(n3144), .B2(
        \xmem_data[25][3] ), .ZN(n28978) );
  AOI22_X1 U32027 ( .A1(n31347), .A2(\xmem_data[26][3] ), .B1(n29064), .B2(
        \xmem_data[27][3] ), .ZN(n28977) );
  AOI22_X1 U32028 ( .A1(n3222), .A2(\xmem_data[28][3] ), .B1(n29789), .B2(
        \xmem_data[29][3] ), .ZN(n28976) );
  AOI22_X1 U32029 ( .A1(n29028), .A2(\xmem_data[30][3] ), .B1(n30883), .B2(
        \xmem_data[31][3] ), .ZN(n28975) );
  NAND4_X1 U32030 ( .A1(n28978), .A2(n28977), .A3(n28976), .A4(n28975), .ZN(
        n28992) );
  AOI22_X1 U32031 ( .A1(n28979), .A2(\xmem_data[20][3] ), .B1(n29820), .B2(
        \xmem_data[21][3] ), .ZN(n28990) );
  AOI22_X1 U32032 ( .A1(n31275), .A2(\xmem_data[0][3] ), .B1(n25417), .B2(
        \xmem_data[1][3] ), .ZN(n28982) );
  AOI22_X1 U32033 ( .A1(n25423), .A2(\xmem_data[6][3] ), .B1(n24131), .B2(
        \xmem_data[7][3] ), .ZN(n28981) );
  NAND2_X1 U32034 ( .A1(n28982), .A2(n28981), .ZN(n28988) );
  AOI22_X1 U32035 ( .A1(n21051), .A2(\xmem_data[16][3] ), .B1(n3328), .B2(
        \xmem_data[17][3] ), .ZN(n28986) );
  AOI22_X1 U32036 ( .A1(n24686), .A2(\xmem_data[22][3] ), .B1(n20986), .B2(
        \xmem_data[23][3] ), .ZN(n28985) );
  AOI22_X1 U32037 ( .A1(n28983), .A2(\xmem_data[18][3] ), .B1(n3172), .B2(
        \xmem_data[19][3] ), .ZN(n28984) );
  NAND3_X1 U32038 ( .A1(n28986), .A2(n28985), .A3(n28984), .ZN(n28987) );
  AOI22_X1 U32039 ( .A1(n23793), .A2(\xmem_data[8][3] ), .B1(n27517), .B2(
        \xmem_data[9][3] ), .ZN(n28998) );
  AOI22_X1 U32040 ( .A1(n28993), .A2(\xmem_data[10][3] ), .B1(n20585), .B2(
        \xmem_data[11][3] ), .ZN(n28997) );
  AOI22_X1 U32041 ( .A1(n24707), .A2(\xmem_data[12][3] ), .B1(n28994), .B2(
        \xmem_data[13][3] ), .ZN(n28996) );
  AOI22_X1 U32042 ( .A1(n31254), .A2(\xmem_data[14][3] ), .B1(n24220), .B2(
        \xmem_data[15][3] ), .ZN(n28995) );
  NAND4_X1 U32043 ( .A1(n28998), .A2(n28997), .A3(n28996), .A4(n28995), .ZN(
        n29001) );
  AOI22_X1 U32044 ( .A1(n27863), .A2(\xmem_data[4][3] ), .B1(n30663), .B2(
        \xmem_data[5][3] ), .ZN(n28999) );
  INV_X1 U32045 ( .A(n28999), .ZN(n29000) );
  NOR3_X1 U32046 ( .A1(n3951), .A2(n29001), .A3(n29000), .ZN(n29004) );
  INV_X1 U32047 ( .A(n29002), .ZN(n29003) );
  AOI21_X1 U32048 ( .B1(n29005), .B2(n29004), .A(n29003), .ZN(n29006) );
  NOR2_X1 U32049 ( .A1(n29007), .A2(n29006), .ZN(n29085) );
  AOI22_X1 U32050 ( .A1(n28045), .A2(\xmem_data[66][3] ), .B1(n27508), .B2(
        \xmem_data[67][3] ), .ZN(n29044) );
  AOI22_X1 U32051 ( .A1(n29009), .A2(\xmem_data[72][3] ), .B1(n29008), .B2(
        \xmem_data[73][3] ), .ZN(n29016) );
  AOI22_X1 U32052 ( .A1(n3213), .A2(\xmem_data[74][3] ), .B1(n29010), .B2(
        \xmem_data[75][3] ), .ZN(n29015) );
  AOI22_X1 U32053 ( .A1(n28492), .A2(\xmem_data[76][3] ), .B1(n29012), .B2(
        \xmem_data[77][3] ), .ZN(n29014) );
  AOI22_X1 U32054 ( .A1(n29238), .A2(\xmem_data[78][3] ), .B1(n27974), .B2(
        \xmem_data[79][3] ), .ZN(n29013) );
  NAND4_X1 U32055 ( .A1(n29016), .A2(n29015), .A3(n29014), .A4(n29013), .ZN(
        n29040) );
  AOI22_X1 U32056 ( .A1(n3357), .A2(\xmem_data[68][3] ), .B1(n29308), .B2(
        \xmem_data[69][3] ), .ZN(n29038) );
  AOI22_X1 U32057 ( .A1(n25364), .A2(\xmem_data[80][3] ), .B1(n29246), .B2(
        \xmem_data[81][3] ), .ZN(n29022) );
  AOI22_X1 U32058 ( .A1(n24521), .A2(\xmem_data[82][3] ), .B1(n3172), .B2(
        \xmem_data[83][3] ), .ZN(n29021) );
  AND2_X1 U32059 ( .A1(n29017), .A2(\xmem_data[84][3] ), .ZN(n29018) );
  AOI21_X1 U32060 ( .B1(n21060), .B2(\xmem_data[85][3] ), .A(n29018), .ZN(
        n29020) );
  AOI22_X1 U32061 ( .A1(n21059), .A2(\xmem_data[86][3] ), .B1(n30862), .B2(
        \xmem_data[87][3] ), .ZN(n29019) );
  NAND4_X1 U32062 ( .A1(n29022), .A2(n29021), .A3(n29020), .A4(n29019), .ZN(
        n29036) );
  AOI22_X1 U32063 ( .A1(n28509), .A2(\xmem_data[64][3] ), .B1(n29350), .B2(
        \xmem_data[65][3] ), .ZN(n29025) );
  AOI22_X1 U32064 ( .A1(n27513), .A2(\xmem_data[70][3] ), .B1(n28980), .B2(
        \xmem_data[71][3] ), .ZN(n29024) );
  NAND2_X1 U32065 ( .A1(n29025), .A2(n29024), .ZN(n29034) );
  AOI22_X1 U32066 ( .A1(n31347), .A2(\xmem_data[90][3] ), .B1(n29064), .B2(
        \xmem_data[91][3] ), .ZN(n29032) );
  AOI22_X1 U32067 ( .A1(n3203), .A2(\xmem_data[88][3] ), .B1(n3413), .B2(
        \xmem_data[89][3] ), .ZN(n29031) );
  AOI22_X1 U32068 ( .A1(n3217), .A2(\xmem_data[92][3] ), .B1(n29026), .B2(
        \xmem_data[93][3] ), .ZN(n29030) );
  AOI22_X1 U32069 ( .A1(n29028), .A2(\xmem_data[94][3] ), .B1(n29027), .B2(
        \xmem_data[95][3] ), .ZN(n29029) );
  NAND4_X1 U32070 ( .A1(n29032), .A2(n29031), .A3(n29030), .A4(n29029), .ZN(
        n29033) );
  NAND2_X1 U32071 ( .A1(n29038), .A2(n29037), .ZN(n29039) );
  NOR2_X1 U32072 ( .A1(n29040), .A2(n29039), .ZN(n29043) );
  INV_X1 U32073 ( .A(n29041), .ZN(n29042) );
  AOI21_X1 U32074 ( .B1(n29044), .B2(n29043), .A(n29042), .ZN(n29083) );
  AOI22_X1 U32075 ( .A1(n29045), .A2(\xmem_data[34][3] ), .B1(n30885), .B2(
        \xmem_data[35][3] ), .ZN(n29081) );
  AOI22_X1 U32076 ( .A1(n29046), .A2(\xmem_data[40][3] ), .B1(n30892), .B2(
        \xmem_data[41][3] ), .ZN(n29053) );
  AOI22_X1 U32077 ( .A1(n29162), .A2(\xmem_data[42][3] ), .B1(n20585), .B2(
        \xmem_data[43][3] ), .ZN(n29052) );
  AOI22_X1 U32078 ( .A1(n29048), .A2(\xmem_data[44][3] ), .B1(n29047), .B2(
        \xmem_data[45][3] ), .ZN(n29051) );
  AOI22_X1 U32079 ( .A1(n29049), .A2(\xmem_data[46][3] ), .B1(n28428), .B2(
        \xmem_data[47][3] ), .ZN(n29050) );
  NAND4_X1 U32080 ( .A1(n29053), .A2(n29052), .A3(n29051), .A4(n29050), .ZN(
        n29077) );
  AOI22_X1 U32081 ( .A1(n29307), .A2(\xmem_data[36][3] ), .B1(n30083), .B2(
        \xmem_data[37][3] ), .ZN(n29075) );
  AOI22_X1 U32082 ( .A1(n29055), .A2(\xmem_data[48][3] ), .B1(n29054), .B2(
        \xmem_data[49][3] ), .ZN(n29061) );
  AOI22_X1 U32083 ( .A1(n27525), .A2(\xmem_data[50][3] ), .B1(n3179), .B2(
        \xmem_data[51][3] ), .ZN(n29060) );
  AND2_X1 U32084 ( .A1(n28500), .A2(\xmem_data[52][3] ), .ZN(n29056) );
  AOI21_X1 U32085 ( .B1(n28772), .B2(\xmem_data[53][3] ), .A(n29056), .ZN(
        n29059) );
  AOI22_X1 U32086 ( .A1(n29248), .A2(\xmem_data[54][3] ), .B1(n29057), .B2(
        \xmem_data[55][3] ), .ZN(n29058) );
  NAND4_X1 U32087 ( .A1(n29061), .A2(n29060), .A3(n29059), .A4(n29058), .ZN(
        n29073) );
  AOI22_X1 U32088 ( .A1(n3256), .A2(\xmem_data[32][3] ), .B1(n3375), .B2(
        \xmem_data[33][3] ), .ZN(n29063) );
  AOI22_X1 U32089 ( .A1(n13168), .A2(\xmem_data[38][3] ), .B1(n28298), .B2(
        \xmem_data[39][3] ), .ZN(n29062) );
  NAND2_X1 U32090 ( .A1(n29063), .A2(n29062), .ZN(n29071) );
  AOI22_X1 U32091 ( .A1(n22753), .A2(\xmem_data[58][3] ), .B1(n29064), .B2(
        \xmem_data[59][3] ), .ZN(n29069) );
  AOI22_X1 U32092 ( .A1(n29118), .A2(\xmem_data[56][3] ), .B1(n3412), .B2(
        \xmem_data[57][3] ), .ZN(n29068) );
  AOI22_X1 U32093 ( .A1(n3220), .A2(\xmem_data[60][3] ), .B1(n29065), .B2(
        \xmem_data[61][3] ), .ZN(n29067) );
  AOI22_X1 U32094 ( .A1(n20723), .A2(\xmem_data[62][3] ), .B1(n24438), .B2(
        \xmem_data[63][3] ), .ZN(n29066) );
  NAND4_X1 U32095 ( .A1(n29069), .A2(n29068), .A3(n29067), .A4(n29066), .ZN(
        n29070) );
  NAND2_X1 U32096 ( .A1(n29075), .A2(n29074), .ZN(n29076) );
  NOR2_X1 U32097 ( .A1(n29077), .A2(n29076), .ZN(n29080) );
  INV_X1 U32098 ( .A(n29078), .ZN(n29079) );
  AOI21_X1 U32099 ( .B1(n29081), .B2(n29080), .A(n29079), .ZN(n29082) );
  NOR2_X1 U32100 ( .A1(n29083), .A2(n29082), .ZN(n29084) );
  XNOR2_X1 U32101 ( .A(n32616), .B(\fmem_data[9][5] ), .ZN(n32139) );
  OAI22_X1 U32102 ( .A1(n32139), .A2(n35040), .B1(n30360), .B2(n35041), .ZN(
        n30367) );
  XNOR2_X1 U32103 ( .A(n3371), .B(\fmem_data[18][3] ), .ZN(n30393) );
  XNOR2_X1 U32104 ( .A(n3442), .B(\fmem_data[18][3] ), .ZN(n32284) );
  OAI22_X1 U32105 ( .A1(n30393), .A2(n33681), .B1(n32284), .B2(n33679), .ZN(
        n30845) );
  XNOR2_X1 U32106 ( .A(n36110), .B(\fmem_data[25][7] ), .ZN(n29207) );
  AND2_X1 U32107 ( .A1(n29086), .A2(\xmem_data[36][1] ), .ZN(n29087) );
  AOI21_X1 U32108 ( .B1(n29298), .B2(\xmem_data[37][1] ), .A(n29087), .ZN(
        n29088) );
  INV_X1 U32109 ( .A(n29088), .ZN(n29094) );
  AOI22_X1 U32110 ( .A1(n29089), .A2(\xmem_data[32][1] ), .B1(n29297), .B2(
        \xmem_data[33][1] ), .ZN(n29092) );
  AOI22_X1 U32111 ( .A1(n28035), .A2(\xmem_data[38][1] ), .B1(n24688), .B2(
        \xmem_data[39][1] ), .ZN(n29091) );
  AOI22_X1 U32112 ( .A1(n29126), .A2(\xmem_data[34][1] ), .B1(n3179), .B2(
        \xmem_data[35][1] ), .ZN(n29090) );
  NOR2_X1 U32113 ( .A1(n29094), .A2(n29093), .ZN(n29117) );
  AOI22_X1 U32114 ( .A1(n20711), .A2(\xmem_data[42][1] ), .B1(n20518), .B2(
        \xmem_data[43][1] ), .ZN(n29099) );
  AOI22_X1 U32115 ( .A1(n22729), .A2(\xmem_data[40][1] ), .B1(n3306), .B2(
        \xmem_data[41][1] ), .ZN(n29098) );
  AOI22_X1 U32116 ( .A1(n3217), .A2(\xmem_data[44][1] ), .B1(n28137), .B2(
        \xmem_data[45][1] ), .ZN(n29097) );
  AOI22_X1 U32117 ( .A1(n29095), .A2(\xmem_data[46][1] ), .B1(n25694), .B2(
        \xmem_data[47][1] ), .ZN(n29096) );
  AOI22_X1 U32118 ( .A1(n29101), .A2(\xmem_data[62][1] ), .B1(n28460), .B2(
        \xmem_data[63][1] ), .ZN(n29102) );
  INV_X1 U32119 ( .A(n29102), .ZN(n29115) );
  AOI22_X1 U32120 ( .A1(n30854), .A2(\xmem_data[52][1] ), .B1(n20587), .B2(
        \xmem_data[53][1] ), .ZN(n29108) );
  AOI22_X1 U32121 ( .A1(n29103), .A2(\xmem_data[50][1] ), .B1(n27447), .B2(
        \xmem_data[51][1] ), .ZN(n29107) );
  AOI22_X1 U32122 ( .A1(n29104), .A2(\xmem_data[48][1] ), .B1(n29157), .B2(
        \xmem_data[49][1] ), .ZN(n29106) );
  AOI22_X1 U32123 ( .A1(n29009), .A2(\xmem_data[56][1] ), .B1(n3464), .B2(
        \xmem_data[57][1] ), .ZN(n29105) );
  NAND4_X1 U32124 ( .A1(n29108), .A2(n29107), .A3(n29106), .A4(n29105), .ZN(
        n29114) );
  AOI22_X1 U32125 ( .A1(n28416), .A2(\xmem_data[54][1] ), .B1(n29109), .B2(
        \xmem_data[55][1] ), .ZN(n29112) );
  AOI22_X1 U32126 ( .A1(n28058), .A2(\xmem_data[60][1] ), .B1(n29319), .B2(
        \xmem_data[61][1] ), .ZN(n29111) );
  AOI22_X1 U32127 ( .A1(n29162), .A2(\xmem_data[58][1] ), .B1(n21007), .B2(
        \xmem_data[59][1] ), .ZN(n29110) );
  NOR3_X1 U32128 ( .A1(n29115), .A2(n29114), .A3(n29113), .ZN(n29116) );
  NAND3_X1 U32129 ( .A1(n29117), .A2(n3808), .A3(n29116), .ZN(n29146) );
  AOI22_X1 U32130 ( .A1(n29118), .A2(\xmem_data[8][1] ), .B1(n28973), .B2(
        \xmem_data[9][1] ), .ZN(n29122) );
  AOI22_X1 U32131 ( .A1(n27437), .A2(\xmem_data[10][1] ), .B1(n24631), .B2(
        \xmem_data[11][1] ), .ZN(n29121) );
  AOI22_X1 U32132 ( .A1(n3222), .A2(\xmem_data[12][1] ), .B1(n28733), .B2(
        \xmem_data[13][1] ), .ZN(n29120) );
  AOI22_X1 U32133 ( .A1(n25562), .A2(\xmem_data[14][1] ), .B1(n27904), .B2(
        \xmem_data[15][1] ), .ZN(n29119) );
  AOI22_X1 U32134 ( .A1(n25576), .A2(\xmem_data[30][1] ), .B1(n24190), .B2(
        \xmem_data[31][1] ), .ZN(n29123) );
  INV_X1 U32135 ( .A(n29123), .ZN(n29135) );
  AOI22_X1 U32136 ( .A1(n20544), .A2(\xmem_data[24][1] ), .B1(n3464), .B2(
        \xmem_data[25][1] ), .ZN(n29129) );
  AOI22_X1 U32137 ( .A1(n29125), .A2(\xmem_data[6][1] ), .B1(n29124), .B2(
        \xmem_data[7][1] ), .ZN(n29128) );
  AOI22_X1 U32138 ( .A1(n29126), .A2(\xmem_data[2][1] ), .B1(n3172), .B2(
        \xmem_data[3][1] ), .ZN(n29127) );
  AOI22_X1 U32139 ( .A1(n29089), .A2(\xmem_data[0][1] ), .B1(n30600), .B2(
        \xmem_data[1][1] ), .ZN(n29132) );
  AOI22_X1 U32140 ( .A1(n30544), .A2(\xmem_data[28][1] ), .B1(n24115), .B2(
        \xmem_data[29][1] ), .ZN(n29131) );
  AOI22_X1 U32141 ( .A1(n22742), .A2(\xmem_data[26][1] ), .B1(n25635), .B2(
        \xmem_data[27][1] ), .ZN(n29130) );
  NOR3_X1 U32142 ( .A1(n29135), .A2(n29134), .A3(n29133), .ZN(n29142) );
  AOI22_X1 U32143 ( .A1(n29136), .A2(\xmem_data[4][1] ), .B1(n29725), .B2(
        \xmem_data[5][1] ), .ZN(n29141) );
  AOI22_X1 U32144 ( .A1(n20993), .A2(\xmem_data[16][1] ), .B1(n3375), .B2(
        \xmem_data[17][1] ), .ZN(n29140) );
  AOI22_X1 U32145 ( .A1(n27547), .A2(\xmem_data[18][1] ), .B1(n27447), .B2(
        \xmem_data[19][1] ), .ZN(n29139) );
  AOI22_X1 U32146 ( .A1(n25481), .A2(\xmem_data[20][1] ), .B1(n30886), .B2(
        \xmem_data[21][1] ), .ZN(n29138) );
  AOI22_X1 U32147 ( .A1(n17012), .A2(\xmem_data[22][1] ), .B1(n16986), .B2(
        \xmem_data[23][1] ), .ZN(n29137) );
  NAND4_X1 U32148 ( .A1(n3868), .A2(n29142), .A3(n29141), .A4(n3516), .ZN(
        n29144) );
  AOI22_X1 U32149 ( .A1(n29146), .A2(n29145), .B1(n29144), .B2(n29143), .ZN(
        n29206) );
  AOI22_X1 U32150 ( .A1(n29173), .A2(\xmem_data[106][1] ), .B1(n29064), .B2(
        \xmem_data[107][1] ), .ZN(n29150) );
  AOI22_X1 U32151 ( .A1(n28037), .A2(\xmem_data[104][1] ), .B1(n16980), .B2(
        \xmem_data[105][1] ), .ZN(n29149) );
  AOI22_X1 U32152 ( .A1(n3222), .A2(\xmem_data[108][1] ), .B1(n27445), .B2(
        \xmem_data[109][1] ), .ZN(n29148) );
  AOI22_X1 U32153 ( .A1(n23769), .A2(\xmem_data[110][1] ), .B1(n29174), .B2(
        \xmem_data[111][1] ), .ZN(n29147) );
  AND4_X1 U32154 ( .A1(n29150), .A2(n29149), .A3(n29148), .A4(n29147), .ZN(
        n29170) );
  AOI22_X1 U32155 ( .A1(n28462), .A2(\xmem_data[96][1] ), .B1(n30686), .B2(
        \xmem_data[97][1] ), .ZN(n29156) );
  AOI22_X1 U32156 ( .A1(n24622), .A2(\xmem_data[98][1] ), .B1(n29151), .B2(
        \xmem_data[99][1] ), .ZN(n29155) );
  AND2_X1 U32157 ( .A1(n11008), .A2(\xmem_data[100][1] ), .ZN(n29152) );
  AOI21_X1 U32158 ( .B1(n20567), .B2(\xmem_data[101][1] ), .A(n29152), .ZN(
        n29154) );
  AOI22_X1 U32159 ( .A1(n30498), .A2(\xmem_data[102][1] ), .B1(n30588), .B2(
        \xmem_data[103][1] ), .ZN(n29153) );
  AND4_X1 U32160 ( .A1(n29156), .A2(n29155), .A3(n29154), .A4(n29153), .ZN(
        n29169) );
  AOI22_X1 U32161 ( .A1(n29181), .A2(\xmem_data[112][1] ), .B1(n29157), .B2(
        \xmem_data[113][1] ), .ZN(n29161) );
  AOI22_X1 U32162 ( .A1(n29103), .A2(\xmem_data[114][1] ), .B1(n30551), .B2(
        \xmem_data[115][1] ), .ZN(n29160) );
  AOI22_X1 U32163 ( .A1(n29180), .A2(\xmem_data[116][1] ), .B1(n29179), .B2(
        \xmem_data[117][1] ), .ZN(n29159) );
  AOI22_X1 U32164 ( .A1(n25423), .A2(\xmem_data[118][1] ), .B1(n28980), .B2(
        \xmem_data[119][1] ), .ZN(n29158) );
  AND4_X1 U32165 ( .A1(n29161), .A2(n29160), .A3(n29159), .A4(n29158), .ZN(
        n29168) );
  AOI22_X1 U32166 ( .A1(n14898), .A2(\xmem_data[120][1] ), .B1(n3464), .B2(
        \xmem_data[121][1] ), .ZN(n29166) );
  AOI22_X1 U32167 ( .A1(n29162), .A2(\xmem_data[122][1] ), .B1(n28059), .B2(
        \xmem_data[123][1] ), .ZN(n29165) );
  AOI22_X1 U32168 ( .A1(n30544), .A2(\xmem_data[124][1] ), .B1(n17044), .B2(
        \xmem_data[125][1] ), .ZN(n29164) );
  AOI22_X1 U32169 ( .A1(n29190), .A2(\xmem_data[126][1] ), .B1(n3206), .B2(
        \xmem_data[127][1] ), .ZN(n29163) );
  AND4_X1 U32170 ( .A1(n29166), .A2(n29165), .A3(n29164), .A4(n29163), .ZN(
        n29167) );
  NAND4_X1 U32171 ( .A1(n29170), .A2(n29169), .A3(n29168), .A4(n29167), .ZN(
        n29172) );
  AOI22_X1 U32172 ( .A1(n24470), .A2(\xmem_data[72][1] ), .B1(n3306), .B2(
        \xmem_data[73][1] ), .ZN(n29178) );
  AOI22_X1 U32173 ( .A1(n29173), .A2(\xmem_data[74][1] ), .B1(n28503), .B2(
        \xmem_data[75][1] ), .ZN(n29177) );
  AOI22_X1 U32174 ( .A1(n3222), .A2(\xmem_data[76][1] ), .B1(n29789), .B2(
        \xmem_data[77][1] ), .ZN(n29176) );
  AOI22_X1 U32175 ( .A1(n22710), .A2(\xmem_data[78][1] ), .B1(n29174), .B2(
        \xmem_data[79][1] ), .ZN(n29175) );
  AND4_X1 U32176 ( .A1(n29178), .A2(n29177), .A3(n29176), .A4(n29175), .ZN(
        n29186) );
  AOI22_X1 U32177 ( .A1(n29180), .A2(\xmem_data[84][1] ), .B1(n29179), .B2(
        \xmem_data[85][1] ), .ZN(n29185) );
  AOI22_X1 U32178 ( .A1(n29181), .A2(\xmem_data[80][1] ), .B1(n30710), .B2(
        \xmem_data[81][1] ), .ZN(n29182) );
  AOI22_X1 U32179 ( .A1(n22740), .A2(\xmem_data[86][1] ), .B1(n3176), .B2(
        \xmem_data[87][1] ), .ZN(n29183) );
  NAND3_X1 U32180 ( .A1(n29186), .A2(n29185), .A3(n29184), .ZN(n29203) );
  AOI22_X1 U32181 ( .A1(n28090), .A2(\xmem_data[88][1] ), .B1(n29187), .B2(
        \xmem_data[89][1] ), .ZN(n29194) );
  AOI22_X1 U32182 ( .A1(n29188), .A2(\xmem_data[90][1] ), .B1(n20800), .B2(
        \xmem_data[91][1] ), .ZN(n29193) );
  AOI22_X1 U32183 ( .A1(n28058), .A2(\xmem_data[92][1] ), .B1(n30950), .B2(
        \xmem_data[93][1] ), .ZN(n29192) );
  AOI22_X1 U32184 ( .A1(n29190), .A2(\xmem_data[94][1] ), .B1(n3205), .B2(
        \xmem_data[95][1] ), .ZN(n29191) );
  AOI22_X1 U32185 ( .A1(n21009), .A2(\xmem_data[64][1] ), .B1(n3269), .B2(
        \xmem_data[65][1] ), .ZN(n29197) );
  AOI22_X1 U32186 ( .A1(n31261), .A2(\xmem_data[70][1] ), .B1(n24607), .B2(
        \xmem_data[71][1] ), .ZN(n29196) );
  AOI22_X1 U32187 ( .A1(n27975), .A2(\xmem_data[66][1] ), .B1(n22684), .B2(
        \xmem_data[67][1] ), .ZN(n29195) );
  NAND3_X1 U32188 ( .A1(n29197), .A2(n29196), .A3(n29195), .ZN(n29198) );
  NOR2_X1 U32189 ( .A1(n3920), .A2(n29198), .ZN(n29200) );
  AOI22_X1 U32190 ( .A1(n28292), .A2(\xmem_data[68][1] ), .B1(n30674), .B2(
        \xmem_data[69][1] ), .ZN(n29199) );
  OAI21_X1 U32191 ( .B1(n29203), .B2(n29202), .A(n29201), .ZN(n29204) );
  XNOR2_X1 U32192 ( .A(n32078), .B(\fmem_data[25][7] ), .ZN(n30395) );
  OAI22_X1 U32193 ( .A1(n29207), .A2(n35744), .B1(n30395), .B2(n35745), .ZN(
        n30844) );
  OAI22_X1 U32194 ( .A1(n29209), .A2(n33057), .B1(n33059), .B2(n29208), .ZN(
        n30843) );
  XNOR2_X1 U32195 ( .A(n31386), .B(\fmem_data[31][3] ), .ZN(n32111) );
  OAI22_X1 U32196 ( .A1(n32111), .A2(n34468), .B1(n29210), .B2(n34470), .ZN(
        n30365) );
  AOI22_X1 U32197 ( .A1(n29231), .A2(\xmem_data[96][2] ), .B1(n29103), .B2(
        \xmem_data[97][2] ), .ZN(n29214) );
  AOI22_X1 U32198 ( .A1(n25422), .A2(\xmem_data[98][2] ), .B1(n3358), .B2(
        \xmem_data[99][2] ), .ZN(n29213) );
  AOI22_X1 U32199 ( .A1(n28346), .A2(\xmem_data[100][2] ), .B1(n29232), .B2(
        \xmem_data[101][2] ), .ZN(n29212) );
  AOI22_X1 U32200 ( .A1(n28980), .A2(\xmem_data[102][2] ), .B1(n23715), .B2(
        \xmem_data[103][2] ), .ZN(n29211) );
  NAND4_X1 U32201 ( .A1(n29214), .A2(n29213), .A3(n29212), .A4(n29211), .ZN(
        n29230) );
  AOI22_X1 U32202 ( .A1(n20776), .A2(\xmem_data[104][2] ), .B1(n3213), .B2(
        \xmem_data[105][2] ), .ZN(n29218) );
  AOI22_X1 U32203 ( .A1(n13149), .A2(\xmem_data[106][2] ), .B1(n28058), .B2(
        \xmem_data[107][2] ), .ZN(n29217) );
  AOI22_X1 U32204 ( .A1(n29239), .A2(\xmem_data[108][2] ), .B1(n29238), .B2(
        \xmem_data[109][2] ), .ZN(n29216) );
  AOI22_X1 U32205 ( .A1(n29240), .A2(\xmem_data[110][2] ), .B1(n28429), .B2(
        \xmem_data[111][2] ), .ZN(n29215) );
  NAND4_X1 U32206 ( .A1(n29218), .A2(n29217), .A3(n29216), .A4(n29215), .ZN(
        n29229) );
  AOI22_X1 U32207 ( .A1(n29246), .A2(\xmem_data[112][2] ), .B1(n29245), .B2(
        \xmem_data[113][2] ), .ZN(n29222) );
  AOI22_X1 U32208 ( .A1(n20782), .A2(\xmem_data[114][2] ), .B1(n29247), .B2(
        \xmem_data[115][2] ), .ZN(n29221) );
  AOI22_X1 U32209 ( .A1(n28467), .A2(\xmem_data[116][2] ), .B1(n29248), .B2(
        \xmem_data[117][2] ), .ZN(n29220) );
  AOI22_X1 U32210 ( .A1(n24526), .A2(\xmem_data[118][2] ), .B1(n30861), .B2(
        \xmem_data[119][2] ), .ZN(n29219) );
  NAND4_X1 U32211 ( .A1(n29222), .A2(n29221), .A3(n29220), .A4(n29219), .ZN(
        n29228) );
  AOI22_X1 U32212 ( .A1(n28677), .A2(\xmem_data[120][2] ), .B1(n29253), .B2(
        \xmem_data[121][2] ), .ZN(n29226) );
  AOI22_X1 U32213 ( .A1(n29254), .A2(\xmem_data[122][2] ), .B1(n3222), .B2(
        \xmem_data[123][2] ), .ZN(n29225) );
  AOI22_X1 U32214 ( .A1(n29256), .A2(\xmem_data[124][2] ), .B1(n29255), .B2(
        \xmem_data[125][2] ), .ZN(n29224) );
  AOI22_X1 U32215 ( .A1(n29257), .A2(\xmem_data[126][2] ), .B1(n27994), .B2(
        \xmem_data[127][2] ), .ZN(n29223) );
  NAND4_X1 U32216 ( .A1(n29226), .A2(n29225), .A3(n29224), .A4(n29223), .ZN(
        n29227) );
  OR4_X1 U32217 ( .A1(n29230), .A2(n29229), .A3(n29228), .A4(n29227), .ZN(
        n29268) );
  AOI22_X1 U32218 ( .A1(n29231), .A2(\xmem_data[64][2] ), .B1(n23771), .B2(
        \xmem_data[65][2] ), .ZN(n29236) );
  AOI22_X1 U32219 ( .A1(n27508), .A2(\xmem_data[66][2] ), .B1(n14996), .B2(
        \xmem_data[67][2] ), .ZN(n29235) );
  AOI22_X1 U32220 ( .A1(n27514), .A2(\xmem_data[68][2] ), .B1(n29232), .B2(
        \xmem_data[69][2] ), .ZN(n29234) );
  AOI22_X1 U32221 ( .A1(n20959), .A2(\xmem_data[70][2] ), .B1(n25606), .B2(
        \xmem_data[71][2] ), .ZN(n29233) );
  NAND4_X1 U32222 ( .A1(n29236), .A2(n29235), .A3(n29234), .A4(n29233), .ZN(
        n29265) );
  AOI22_X1 U32223 ( .A1(n28516), .A2(\xmem_data[72][2] ), .B1(n23716), .B2(
        \xmem_data[73][2] ), .ZN(n29244) );
  AOI22_X1 U32224 ( .A1(n13149), .A2(\xmem_data[74][2] ), .B1(n23796), .B2(
        \xmem_data[75][2] ), .ZN(n29243) );
  AOI22_X1 U32225 ( .A1(n29239), .A2(\xmem_data[76][2] ), .B1(n29238), .B2(
        \xmem_data[77][2] ), .ZN(n29242) );
  AOI22_X1 U32226 ( .A1(n29240), .A2(\xmem_data[78][2] ), .B1(n30955), .B2(
        \xmem_data[79][2] ), .ZN(n29241) );
  NAND4_X1 U32227 ( .A1(n29244), .A2(n29243), .A3(n29242), .A4(n29241), .ZN(
        n29264) );
  AOI22_X1 U32228 ( .A1(n29246), .A2(\xmem_data[80][2] ), .B1(n29245), .B2(
        \xmem_data[81][2] ), .ZN(n29252) );
  AOI22_X1 U32229 ( .A1(n29325), .A2(\xmem_data[82][2] ), .B1(n29247), .B2(
        \xmem_data[83][2] ), .ZN(n29251) );
  AOI22_X1 U32230 ( .A1(n20708), .A2(\xmem_data[84][2] ), .B1(n29248), .B2(
        \xmem_data[85][2] ), .ZN(n29250) );
  AOI22_X1 U32231 ( .A1(n25441), .A2(\xmem_data[86][2] ), .B1(n12471), .B2(
        \xmem_data[87][2] ), .ZN(n29249) );
  NAND4_X1 U32232 ( .A1(n29252), .A2(n29251), .A3(n29250), .A4(n29249), .ZN(
        n29263) );
  AOI22_X1 U32233 ( .A1(n25624), .A2(\xmem_data[88][2] ), .B1(n29253), .B2(
        \xmem_data[89][2] ), .ZN(n29261) );
  AOI22_X1 U32234 ( .A1(n29254), .A2(\xmem_data[90][2] ), .B1(n3220), .B2(
        \xmem_data[91][2] ), .ZN(n29260) );
  AOI22_X1 U32235 ( .A1(n29256), .A2(\xmem_data[92][2] ), .B1(n29255), .B2(
        \xmem_data[93][2] ), .ZN(n29259) );
  AOI22_X1 U32236 ( .A1(n29257), .A2(\xmem_data[94][2] ), .B1(n25486), .B2(
        \xmem_data[95][2] ), .ZN(n29258) );
  NAND4_X1 U32237 ( .A1(n29261), .A2(n29260), .A3(n29259), .A4(n29258), .ZN(
        n29262) );
  OR4_X1 U32238 ( .A1(n29265), .A2(n29264), .A3(n29263), .A4(n29262), .ZN(
        n29266) );
  AOI22_X1 U32239 ( .A1(n29269), .A2(n29268), .B1(n29267), .B2(n29266), .ZN(
        n29346) );
  AOI22_X1 U32240 ( .A1(n31327), .A2(\xmem_data[4][2] ), .B1(n27535), .B2(
        \xmem_data[5][2] ), .ZN(n29270) );
  INV_X1 U32241 ( .A(n29270), .ZN(n29278) );
  AOI22_X1 U32242 ( .A1(n29272), .A2(\xmem_data[6][2] ), .B1(n29271), .B2(
        \xmem_data[7][2] ), .ZN(n29273) );
  INV_X1 U32243 ( .A(n29273), .ZN(n29277) );
  AOI22_X1 U32244 ( .A1(n25422), .A2(\xmem_data[2][2] ), .B1(n3358), .B2(
        \xmem_data[3][2] ), .ZN(n29275) );
  NAND2_X1 U32245 ( .A1(n17063), .A2(\xmem_data[0][2] ), .ZN(n29274) );
  NAND2_X1 U32246 ( .A1(n29275), .A2(n29274), .ZN(n29276) );
  OR3_X1 U32247 ( .A1(n29278), .A2(n29277), .A3(n29276), .ZN(n29296) );
  AOI22_X1 U32248 ( .A1(n3158), .A2(\xmem_data[8][2] ), .B1(n29279), .B2(
        \xmem_data[9][2] ), .ZN(n29285) );
  AOI22_X1 U32249 ( .A1(n28096), .A2(\xmem_data[10][2] ), .B1(n31329), .B2(
        \xmem_data[11][2] ), .ZN(n29284) );
  AOI22_X1 U32250 ( .A1(n22717), .A2(\xmem_data[12][2] ), .B1(n29280), .B2(
        \xmem_data[13][2] ), .ZN(n29283) );
  AOI22_X1 U32251 ( .A1(n24615), .A2(\xmem_data[14][2] ), .B1(n3372), .B2(
        \xmem_data[15][2] ), .ZN(n29282) );
  NAND4_X1 U32252 ( .A1(n29285), .A2(n29284), .A3(n29283), .A4(n29282), .ZN(
        n29295) );
  AOI22_X1 U32253 ( .A1(n3335), .A2(\xmem_data[24][2] ), .B1(n29286), .B2(
        \xmem_data[25][2] ), .ZN(n29293) );
  AND2_X1 U32254 ( .A1(n3217), .A2(\xmem_data[27][2] ), .ZN(n29287) );
  AOI21_X1 U32255 ( .B1(n28082), .B2(\xmem_data[26][2] ), .A(n29287), .ZN(
        n29292) );
  AOI22_X1 U32256 ( .A1(n29288), .A2(\xmem_data[28][2] ), .B1(n23739), .B2(
        \xmem_data[29][2] ), .ZN(n29291) );
  AOI22_X1 U32257 ( .A1(n29289), .A2(\xmem_data[30][2] ), .B1(n24564), .B2(
        \xmem_data[31][2] ), .ZN(n29290) );
  NAND4_X1 U32258 ( .A1(n29293), .A2(n29292), .A3(n29291), .A4(n29290), .ZN(
        n29294) );
  OR3_X1 U32259 ( .A1(n29296), .A2(n29295), .A3(n29294), .ZN(n29304) );
  AOI22_X1 U32260 ( .A1(n29297), .A2(\xmem_data[16][2] ), .B1(n20507), .B2(
        \xmem_data[17][2] ), .ZN(n29302) );
  AOI22_X1 U32261 ( .A1(n24467), .A2(\xmem_data[18][2] ), .B1(n17049), .B2(
        \xmem_data[19][2] ), .ZN(n29301) );
  AOI22_X1 U32262 ( .A1(n29298), .A2(\xmem_data[20][2] ), .B1(n24524), .B2(
        \xmem_data[21][2] ), .ZN(n29300) );
  AOI22_X1 U32263 ( .A1(n17030), .A2(\xmem_data[22][2] ), .B1(n22729), .B2(
        \xmem_data[23][2] ), .ZN(n29299) );
  NAND4_X1 U32264 ( .A1(n29302), .A2(n29301), .A3(n29300), .A4(n29299), .ZN(
        n29303) );
  NOR2_X1 U32265 ( .A1(n29304), .A2(n29303), .ZN(n29305) );
  AOI22_X1 U32266 ( .A1(n28952), .A2(\xmem_data[32][2] ), .B1(n25450), .B2(
        \xmem_data[33][2] ), .ZN(n29314) );
  AOI22_X1 U32267 ( .A1(n28050), .A2(\xmem_data[34][2] ), .B1(n29307), .B2(
        \xmem_data[35][2] ), .ZN(n29313) );
  AOI22_X1 U32268 ( .A1(n29308), .A2(\xmem_data[36][2] ), .B1(n25605), .B2(
        \xmem_data[37][2] ), .ZN(n29312) );
  AOI22_X1 U32269 ( .A1(n29310), .A2(\xmem_data[38][2] ), .B1(n29309), .B2(
        \xmem_data[39][2] ), .ZN(n29311) );
  NAND4_X1 U32270 ( .A1(n29314), .A2(n29313), .A3(n29312), .A4(n29311), .ZN(
        n29340) );
  AOI22_X1 U32271 ( .A1(n30303), .A2(\xmem_data[40][2] ), .B1(n29011), .B2(
        \xmem_data[41][2] ), .ZN(n29323) );
  AOI22_X1 U32272 ( .A1(n29317), .A2(\xmem_data[42][2] ), .B1(n29316), .B2(
        \xmem_data[43][2] ), .ZN(n29322) );
  AOI22_X1 U32273 ( .A1(n29319), .A2(\xmem_data[44][2] ), .B1(n29318), .B2(
        \xmem_data[45][2] ), .ZN(n29321) );
  AOI22_X1 U32274 ( .A1(n21010), .A2(\xmem_data[46][2] ), .B1(n28429), .B2(
        \xmem_data[47][2] ), .ZN(n29320) );
  NAND4_X1 U32275 ( .A1(n29323), .A2(n29322), .A3(n29321), .A4(n29320), .ZN(
        n29339) );
  AOI22_X1 U32276 ( .A1(n29324), .A2(\xmem_data[48][2] ), .B1(n14975), .B2(
        \xmem_data[49][2] ), .ZN(n29332) );
  AOI22_X1 U32277 ( .A1(n29325), .A2(\xmem_data[50][2] ), .B1(n23781), .B2(
        \xmem_data[51][2] ), .ZN(n29331) );
  AOI22_X1 U32278 ( .A1(n29327), .A2(\xmem_data[52][2] ), .B1(n29326), .B2(
        \xmem_data[53][2] ), .ZN(n29330) );
  AOI22_X1 U32279 ( .A1(n27564), .A2(\xmem_data[54][2] ), .B1(n29328), .B2(
        \xmem_data[55][2] ), .ZN(n29329) );
  NAND4_X1 U32280 ( .A1(n29332), .A2(n29331), .A3(n29330), .A4(n29329), .ZN(
        n29338) );
  AOI22_X1 U32281 ( .A1(n3384), .A2(\xmem_data[56][2] ), .B1(n31347), .B2(
        \xmem_data[57][2] ), .ZN(n29336) );
  AOI22_X1 U32282 ( .A1(n25354), .A2(\xmem_data[58][2] ), .B1(n3218), .B2(
        \xmem_data[59][2] ), .ZN(n29335) );
  AOI22_X1 U32283 ( .A1(n17033), .A2(\xmem_data[60][2] ), .B1(n30963), .B2(
        \xmem_data[61][2] ), .ZN(n29334) );
  AOI22_X1 U32284 ( .A1(n22709), .A2(\xmem_data[62][2] ), .B1(n24140), .B2(
        \xmem_data[63][2] ), .ZN(n29333) );
  NAND4_X1 U32285 ( .A1(n29336), .A2(n29335), .A3(n29334), .A4(n29333), .ZN(
        n29337) );
  OR4_X1 U32286 ( .A1(n29340), .A2(n29339), .A3(n29338), .A4(n29337), .ZN(
        n29344) );
  NOR2_X1 U32287 ( .A1(n29341), .A2(n39036), .ZN(n29342) );
  AOI21_X1 U32288 ( .B1(n29344), .B2(n29343), .A(n3902), .ZN(n29345) );
  XNOR2_X1 U32289 ( .A(n32899), .B(\fmem_data[8][5] ), .ZN(n30818) );
  OAI22_X1 U32290 ( .A1(n32130), .A2(n35004), .B1(n30818), .B2(n35003), .ZN(
        n31389) );
  NAND2_X1 U32291 ( .A1(n29646), .A2(\xmem_data[93][0] ), .ZN(n29349) );
  NAND2_X1 U32292 ( .A1(n27703), .A2(\xmem_data[92][0] ), .ZN(n29348) );
  NAND2_X1 U32293 ( .A1(n29349), .A2(n29348), .ZN(n29354) );
  AOI22_X1 U32294 ( .A1(n29402), .A2(\xmem_data[90][0] ), .B1(n29350), .B2(
        \xmem_data[91][0] ), .ZN(n29352) );
  AOI22_X1 U32295 ( .A1(n29404), .A2(\xmem_data[94][0] ), .B1(n29403), .B2(
        \xmem_data[95][0] ), .ZN(n29351) );
  NAND2_X1 U32296 ( .A1(n29352), .A2(n29351), .ZN(n29353) );
  NOR2_X1 U32297 ( .A1(n29354), .A2(n29353), .ZN(n29371) );
  AOI22_X1 U32298 ( .A1(n29400), .A2(\xmem_data[88][0] ), .B1(n30293), .B2(
        \xmem_data[89][0] ), .ZN(n29370) );
  AOI22_X1 U32299 ( .A1(n3165), .A2(\xmem_data[68][0] ), .B1(n3182), .B2(
        \xmem_data[69][0] ), .ZN(n29355) );
  INV_X1 U32300 ( .A(n29355), .ZN(n29362) );
  AOI22_X1 U32301 ( .A1(n30635), .A2(\xmem_data[64][0] ), .B1(n29648), .B2(
        \xmem_data[65][0] ), .ZN(n29357) );
  AOI22_X1 U32302 ( .A1(n29397), .A2(\xmem_data[66][0] ), .B1(n27517), .B2(
        \xmem_data[67][0] ), .ZN(n29356) );
  NAND2_X1 U32303 ( .A1(n29357), .A2(n29356), .ZN(n29361) );
  NAND2_X1 U32304 ( .A1(n30075), .A2(\xmem_data[70][0] ), .ZN(n29359) );
  NAND2_X1 U32305 ( .A1(n29410), .A2(\xmem_data[71][0] ), .ZN(n29358) );
  NAND2_X1 U32306 ( .A1(n29359), .A2(n29358), .ZN(n29360) );
  NOR3_X1 U32307 ( .A1(n29362), .A2(n29361), .A3(n29360), .ZN(n29369) );
  AOI22_X1 U32308 ( .A1(n29363), .A2(\xmem_data[72][0] ), .B1(n30765), .B2(
        \xmem_data[73][0] ), .ZN(n29367) );
  AOI22_X1 U32309 ( .A1(n29380), .A2(\xmem_data[74][0] ), .B1(n29379), .B2(
        \xmem_data[75][0] ), .ZN(n29366) );
  AOI22_X1 U32310 ( .A1(n29382), .A2(\xmem_data[76][0] ), .B1(n29381), .B2(
        \xmem_data[77][0] ), .ZN(n29365) );
  AOI22_X1 U32311 ( .A1(n29384), .A2(\xmem_data[78][0] ), .B1(n29383), .B2(
        \xmem_data[79][0] ), .ZN(n29364) );
  NAND4_X1 U32312 ( .A1(n29371), .A2(n29370), .A3(n29369), .A4(n29368), .ZN(
        n29378) );
  AOI22_X1 U32313 ( .A1(n29419), .A2(\xmem_data[80][0] ), .B1(n29418), .B2(
        \xmem_data[81][0] ), .ZN(n29375) );
  AOI22_X1 U32314 ( .A1(n29420), .A2(\xmem_data[82][0] ), .B1(n28718), .B2(
        \xmem_data[83][0] ), .ZN(n29374) );
  AOI22_X1 U32315 ( .A1(n29433), .A2(\xmem_data[84][0] ), .B1(n27013), .B2(
        \xmem_data[85][0] ), .ZN(n29373) );
  AOI22_X1 U32316 ( .A1(n3392), .A2(\xmem_data[86][0] ), .B1(n29422), .B2(
        \xmem_data[87][0] ), .ZN(n29372) );
  NAND4_X1 U32317 ( .A1(n29375), .A2(n29374), .A3(n29373), .A4(n29372), .ZN(
        n29377) );
  OAI21_X1 U32318 ( .B1(n29378), .B2(n29377), .A(n29376), .ZN(n29516) );
  AOI22_X1 U32319 ( .A1(n29363), .A2(\xmem_data[104][0] ), .B1(n29487), .B2(
        \xmem_data[105][0] ), .ZN(n29388) );
  AOI22_X1 U32320 ( .A1(n29380), .A2(\xmem_data[106][0] ), .B1(n29379), .B2(
        \xmem_data[107][0] ), .ZN(n29387) );
  AOI22_X1 U32321 ( .A1(n29382), .A2(\xmem_data[108][0] ), .B1(n29381), .B2(
        \xmem_data[109][0] ), .ZN(n29386) );
  AOI22_X1 U32322 ( .A1(n29384), .A2(\xmem_data[110][0] ), .B1(n29383), .B2(
        \xmem_data[111][0] ), .ZN(n29385) );
  NAND4_X1 U32323 ( .A1(n29388), .A2(n29387), .A3(n29386), .A4(n29385), .ZN(
        n29394) );
  NAND2_X1 U32324 ( .A1(n29482), .A2(\xmem_data[125][0] ), .ZN(n29392) );
  NAND2_X1 U32325 ( .A1(n28180), .A2(\xmem_data[124][0] ), .ZN(n29391) );
  NAND2_X1 U32326 ( .A1(n29392), .A2(n29391), .ZN(n29393) );
  NOR2_X1 U32327 ( .A1(n29394), .A2(n29393), .ZN(n29417) );
  AOI22_X1 U32328 ( .A1(n29395), .A2(\xmem_data[96][0] ), .B1(n28778), .B2(
        \xmem_data[97][0] ), .ZN(n29399) );
  AOI22_X1 U32329 ( .A1(n29397), .A2(\xmem_data[98][0] ), .B1(n23795), .B2(
        \xmem_data[99][0] ), .ZN(n29398) );
  NAND2_X1 U32330 ( .A1(n29399), .A2(n29398), .ZN(n29409) );
  AOI22_X1 U32331 ( .A1(n29400), .A2(\xmem_data[120][0] ), .B1(n3170), .B2(
        \xmem_data[121][0] ), .ZN(n29407) );
  AOI22_X1 U32332 ( .A1(n29402), .A2(\xmem_data[122][0] ), .B1(n3135), .B2(
        \xmem_data[123][0] ), .ZN(n29406) );
  AOI22_X1 U32333 ( .A1(n29404), .A2(\xmem_data[126][0] ), .B1(n29403), .B2(
        \xmem_data[127][0] ), .ZN(n29405) );
  NAND2_X1 U32334 ( .A1(n29407), .A2(n4009), .ZN(n29408) );
  NOR2_X1 U32335 ( .A1(n29409), .A2(n29408), .ZN(n29416) );
  AOI22_X1 U32336 ( .A1(n30075), .A2(\xmem_data[102][0] ), .B1(n29410), .B2(
        \xmem_data[103][0] ), .ZN(n29411) );
  INV_X1 U32337 ( .A(n29411), .ZN(n29414) );
  AOI22_X1 U32338 ( .A1(n3163), .A2(\xmem_data[100][0] ), .B1(n3185), .B2(
        \xmem_data[101][0] ), .ZN(n29412) );
  INV_X1 U32339 ( .A(n29412), .ZN(n29413) );
  NOR2_X1 U32340 ( .A1(n29414), .A2(n29413), .ZN(n29415) );
  NAND3_X1 U32341 ( .A1(n29417), .A2(n29416), .A3(n29415), .ZN(n29430) );
  AOI22_X1 U32342 ( .A1(n29419), .A2(\xmem_data[112][0] ), .B1(n29418), .B2(
        \xmem_data[113][0] ), .ZN(n29427) );
  AOI22_X1 U32343 ( .A1(n29420), .A2(\xmem_data[114][0] ), .B1(n22728), .B2(
        \xmem_data[115][0] ), .ZN(n29426) );
  AOI22_X1 U32344 ( .A1(n30223), .A2(\xmem_data[116][0] ), .B1(n30775), .B2(
        \xmem_data[117][0] ), .ZN(n29425) );
  AOI22_X1 U32345 ( .A1(n28138), .A2(\xmem_data[118][0] ), .B1(n29422), .B2(
        \xmem_data[119][0] ), .ZN(n29424) );
  NAND4_X1 U32346 ( .A1(n29427), .A2(n29426), .A3(n29425), .A4(n29424), .ZN(
        n29429) );
  OAI21_X1 U32347 ( .B1(n29430), .B2(n29429), .A(n29428), .ZN(n29515) );
  AOI22_X1 U32348 ( .A1(n29423), .A2(\xmem_data[54][0] ), .B1(n29431), .B2(
        \xmem_data[55][0] ), .ZN(n29435) );
  AOI22_X1 U32349 ( .A1(n30223), .A2(\xmem_data[52][0] ), .B1(n30290), .B2(
        \xmem_data[53][0] ), .ZN(n29434) );
  AOI22_X1 U32350 ( .A1(n3163), .A2(\xmem_data[36][0] ), .B1(n3187), .B2(
        \xmem_data[37][0] ), .ZN(n29444) );
  AOI22_X1 U32351 ( .A1(n29604), .A2(\xmem_data[32][0] ), .B1(n29648), .B2(
        \xmem_data[33][0] ), .ZN(n29443) );
  AOI22_X1 U32352 ( .A1(n29438), .A2(\xmem_data[34][0] ), .B1(n30892), .B2(
        \xmem_data[35][0] ), .ZN(n29442) );
  AND2_X1 U32353 ( .A1(n29439), .A2(\xmem_data[39][0] ), .ZN(n29440) );
  AOI21_X1 U32354 ( .B1(n30070), .B2(\xmem_data[38][0] ), .A(n29440), .ZN(
        n29441) );
  NAND2_X1 U32355 ( .A1(n29445), .A2(n3757), .ZN(n29473) );
  AOI22_X1 U32356 ( .A1(n28787), .A2(\xmem_data[56][0] ), .B1(n29495), .B2(
        \xmem_data[57][0] ), .ZN(n29459) );
  AOI22_X1 U32357 ( .A1(n30743), .A2(\xmem_data[60][0] ), .B1(n29389), .B2(
        \xmem_data[61][0] ), .ZN(n29458) );
  AOI22_X1 U32358 ( .A1(n29447), .A2(\xmem_data[48][0] ), .B1(n29497), .B2(
        \xmem_data[49][0] ), .ZN(n29448) );
  AOI22_X1 U32359 ( .A1(n29449), .A2(\xmem_data[50][0] ), .B1(n23754), .B2(
        \xmem_data[51][0] ), .ZN(n29454) );
  AOI22_X1 U32360 ( .A1(n29450), .A2(\xmem_data[58][0] ), .B1(n3375), .B2(
        \xmem_data[59][0] ), .ZN(n29453) );
  AOI22_X1 U32361 ( .A1(n7282), .A2(\xmem_data[62][0] ), .B1(n29451), .B2(
        \xmem_data[63][0] ), .ZN(n29452) );
  NAND3_X1 U32362 ( .A1(n29454), .A2(n29453), .A3(n29452), .ZN(n29455) );
  NOR2_X1 U32363 ( .A1(n29456), .A2(n29455), .ZN(n29457) );
  NAND3_X1 U32364 ( .A1(n29459), .A2(n29458), .A3(n29457), .ZN(n29470) );
  AOI22_X1 U32365 ( .A1(n30766), .A2(\xmem_data[40][0] ), .B1(n30685), .B2(
        \xmem_data[41][0] ), .ZN(n29468) );
  AOI22_X1 U32366 ( .A1(n29461), .A2(\xmem_data[42][0] ), .B1(n3151), .B2(
        \xmem_data[43][0] ), .ZN(n29467) );
  AOI22_X1 U32367 ( .A1(n29463), .A2(\xmem_data[44][0] ), .B1(n29462), .B2(
        \xmem_data[45][0] ), .ZN(n29466) );
  AOI22_X1 U32368 ( .A1(n29464), .A2(\xmem_data[46][0] ), .B1(n31345), .B2(
        \xmem_data[47][0] ), .ZN(n29465) );
  NAND4_X1 U32369 ( .A1(n29468), .A2(n29467), .A3(n29466), .A4(n29465), .ZN(
        n29469) );
  AOI22_X1 U32370 ( .A1(n29436), .A2(\xmem_data[0][0] ), .B1(n29739), .B2(
        \xmem_data[1][0] ), .ZN(n29480) );
  AOI22_X1 U32371 ( .A1(n29475), .A2(\xmem_data[2][0] ), .B1(n29807), .B2(
        \xmem_data[3][0] ), .ZN(n29479) );
  AOI22_X1 U32372 ( .A1(n3164), .A2(\xmem_data[4][0] ), .B1(n3185), .B2(
        \xmem_data[5][0] ), .ZN(n29478) );
  AOI22_X1 U32373 ( .A1(n29476), .A2(\xmem_data[6][0] ), .B1(n28232), .B2(
        \xmem_data[7][0] ), .ZN(n29477) );
  NAND4_X1 U32374 ( .A1(n29480), .A2(n29479), .A3(n29478), .A4(n29477), .ZN(
        n29486) );
  AOI22_X1 U32375 ( .A1(n29347), .A2(\xmem_data[29][0] ), .B1(n29647), .B2(
        \xmem_data[28][0] ), .ZN(n29484) );
  AOI22_X1 U32376 ( .A1(n30291), .A2(\xmem_data[20][0] ), .B1(n29831), .B2(
        \xmem_data[21][0] ), .ZN(n29483) );
  NAND2_X1 U32377 ( .A1(n29484), .A2(n29483), .ZN(n29485) );
  NOR2_X1 U32378 ( .A1(n29486), .A2(n29485), .ZN(n29510) );
  AOI22_X1 U32379 ( .A1(n30076), .A2(\xmem_data[8][0] ), .B1(n30266), .B2(
        \xmem_data[9][0] ), .ZN(n29493) );
  AOI22_X1 U32380 ( .A1(n7270), .A2(\xmem_data[10][0] ), .B1(n30311), .B2(
        \xmem_data[11][0] ), .ZN(n29492) );
  AOI22_X1 U32381 ( .A1(n29463), .A2(\xmem_data[12][0] ), .B1(n29818), .B2(
        \xmem_data[13][0] ), .ZN(n29491) );
  AOI22_X1 U32382 ( .A1(n29489), .A2(\xmem_data[14][0] ), .B1(n30754), .B2(
        \xmem_data[15][0] ), .ZN(n29490) );
  AOI22_X1 U32383 ( .A1(n29699), .A2(\xmem_data[22][0] ), .B1(n29494), .B2(
        \xmem_data[23][0] ), .ZN(n29509) );
  AOI22_X1 U32384 ( .A1(n29674), .A2(\xmem_data[24][0] ), .B1(n29495), .B2(
        \xmem_data[25][0] ), .ZN(n29496) );
  INV_X1 U32385 ( .A(n29496), .ZN(n29507) );
  AOI22_X1 U32386 ( .A1(n28717), .A2(\xmem_data[16][0] ), .B1(n29497), .B2(
        \xmem_data[17][0] ), .ZN(n29498) );
  INV_X1 U32387 ( .A(n29498), .ZN(n29506) );
  AOI22_X1 U32388 ( .A1(n29499), .A2(\xmem_data[18][0] ), .B1(n3153), .B2(
        \xmem_data[19][0] ), .ZN(n29504) );
  AOI22_X1 U32389 ( .A1(n29500), .A2(\xmem_data[30][0] ), .B1(n23762), .B2(
        \xmem_data[31][0] ), .ZN(n29503) );
  AOI22_X1 U32390 ( .A1(n29501), .A2(\xmem_data[26][0] ), .B1(n3375), .B2(
        \xmem_data[27][0] ), .ZN(n29502) );
  NOR3_X1 U32391 ( .A1(n29507), .A2(n29506), .A3(n29505), .ZN(n29508) );
  NAND4_X1 U32392 ( .A1(n29510), .A2(n3780), .A3(n29509), .A4(n29508), .ZN(
        n29512) );
  NAND2_X1 U32393 ( .A1(n29512), .A2(n29511), .ZN(n29513) );
  INV_X1 U32394 ( .A(n35638), .ZN(n29517) );
  XNOR2_X1 U32395 ( .A(n35326), .B(\fmem_data[25][1] ), .ZN(n33178) );
  XNOR2_X1 U32396 ( .A(n34982), .B(\fmem_data[25][1] ), .ZN(n32147) );
  OAI22_X1 U32397 ( .A1(n33178), .A2(n3483), .B1(n32147), .B2(n34440), .ZN(
        n29686) );
  XNOR2_X1 U32398 ( .A(n31996), .B(\fmem_data[8][1] ), .ZN(n29519) );
  XNOR2_X1 U32399 ( .A(n35328), .B(\fmem_data[8][1] ), .ZN(n33263) );
  OAI22_X1 U32400 ( .A1(n29519), .A2(n34625), .B1(n33263), .B2(n3574), .ZN(
        n29685) );
  XNOR2_X1 U32401 ( .A(n31957), .B(\fmem_data[6][3] ), .ZN(n32118) );
  XNOR2_X1 U32402 ( .A(n31958), .B(\fmem_data[6][3] ), .ZN(n31880) );
  OAI22_X1 U32403 ( .A1(n32118), .A2(n33598), .B1(n31880), .B2(n33596), .ZN(
        n31229) );
  XNOR2_X1 U32404 ( .A(n31668), .B(\fmem_data[13][1] ), .ZN(n32241) );
  OAI22_X1 U32405 ( .A1(n32241), .A2(n34742), .B1(n33927), .B2(n3571), .ZN(
        n31227) );
  XNOR2_X1 U32406 ( .A(n29521), .B(n29520), .ZN(n29523) );
  XNOR2_X1 U32407 ( .A(n29523), .B(n29522), .ZN(n31409) );
  FA_X1 U32408 ( .A(n29526), .B(n29525), .CI(n29524), .CO(n27321), .S(n31408)
         );
  FA_X1 U32409 ( .A(n29529), .B(n29528), .CI(n29527), .CO(n29522), .S(n31236)
         );
  FA_X1 U32410 ( .A(n29532), .B(n29531), .CI(n29530), .CO(n28906), .S(n31235)
         );
  FA_X1 U32411 ( .A(n29535), .B(n29534), .CI(n29533), .CO(n28910), .S(n31234)
         );
  NAND2_X1 U32412 ( .A1(n31414), .A2(n31413), .ZN(n30133) );
  FA_X1 U32413 ( .A(n29538), .B(n29537), .CI(n29536), .CO(n30139), .S(n30337)
         );
  FA_X1 U32414 ( .A(n29541), .B(n29540), .CI(n29539), .CO(n26035), .S(n30338)
         );
  XNOR2_X1 U32415 ( .A(n33027), .B(\fmem_data[7][3] ), .ZN(n32175) );
  OAI22_X1 U32416 ( .A1(n32175), .A2(n34503), .B1(n29542), .B2(n34505), .ZN(
        n29694) );
  AOI22_X1 U32417 ( .A1(n29647), .A2(\xmem_data[64][1] ), .B1(n28238), .B2(
        \xmem_data[65][1] ), .ZN(n29546) );
  AOI22_X1 U32418 ( .A1(n3239), .A2(\xmem_data[66][1] ), .B1(n29591), .B2(
        \xmem_data[67][1] ), .ZN(n29545) );
  AOI22_X1 U32419 ( .A1(n3173), .A2(\xmem_data[68][1] ), .B1(n28110), .B2(
        \xmem_data[69][1] ), .ZN(n29544) );
  AOI22_X1 U32420 ( .A1(n29593), .A2(\xmem_data[70][1] ), .B1(n29315), .B2(
        \xmem_data[71][1] ), .ZN(n29543) );
  NAND4_X1 U32421 ( .A1(n29546), .A2(n29545), .A3(n29544), .A4(n29543), .ZN(
        n29564) );
  AOI22_X1 U32422 ( .A1(n3160), .A2(\xmem_data[72][1] ), .B1(n3189), .B2(
        \xmem_data[73][1] ), .ZN(n29551) );
  AOI22_X1 U32423 ( .A1(n23901), .A2(\xmem_data[74][1] ), .B1(n29047), .B2(
        \xmem_data[75][1] ), .ZN(n29550) );
  AOI22_X1 U32424 ( .A1(n28173), .A2(\xmem_data[76][1] ), .B1(n30644), .B2(
        \xmem_data[77][1] ), .ZN(n29549) );
  AOI22_X1 U32425 ( .A1(n29574), .A2(\xmem_data[78][1] ), .B1(n29573), .B2(
        \xmem_data[79][1] ), .ZN(n29548) );
  NAND4_X1 U32426 ( .A1(n29551), .A2(n29550), .A3(n29549), .A4(n29548), .ZN(
        n29563) );
  AOI22_X1 U32427 ( .A1(n29656), .A2(\xmem_data[80][1] ), .B1(n29615), .B2(
        \xmem_data[81][1] ), .ZN(n29555) );
  AOI22_X1 U32428 ( .A1(n29658), .A2(\xmem_data[82][1] ), .B1(n14982), .B2(
        \xmem_data[83][1] ), .ZN(n29554) );
  AOI22_X1 U32429 ( .A1(n29583), .A2(\xmem_data[84][1] ), .B1(n29582), .B2(
        \xmem_data[85][1] ), .ZN(n29553) );
  AOI22_X1 U32430 ( .A1(n29584), .A2(\xmem_data[86][1] ), .B1(n25624), .B2(
        \xmem_data[87][1] ), .ZN(n29552) );
  NAND4_X1 U32431 ( .A1(n29555), .A2(n29554), .A3(n29553), .A4(n29552), .ZN(
        n29562) );
  AOI22_X1 U32432 ( .A1(n28207), .A2(\xmem_data[90][1] ), .B1(n29565), .B2(
        \xmem_data[91][1] ), .ZN(n29560) );
  AOI22_X1 U32433 ( .A1(n29674), .A2(\xmem_data[92][1] ), .B1(n29708), .B2(
        \xmem_data[93][1] ), .ZN(n29559) );
  AOI22_X1 U32434 ( .A1(n29626), .A2(\xmem_data[88][1] ), .B1(n30654), .B2(
        \xmem_data[89][1] ), .ZN(n29558) );
  AOI22_X1 U32435 ( .A1(n29568), .A2(\xmem_data[94][1] ), .B1(n3345), .B2(
        \xmem_data[95][1] ), .ZN(n29557) );
  NAND4_X1 U32436 ( .A1(n29560), .A2(n29559), .A3(n29558), .A4(n29557), .ZN(
        n29561) );
  AOI22_X1 U32437 ( .A1(n27710), .A2(\xmem_data[120][1] ), .B1(n29831), .B2(
        \xmem_data[121][1] ), .ZN(n29572) );
  AOI22_X1 U32438 ( .A1(n29628), .A2(\xmem_data[122][1] ), .B1(n29565), .B2(
        \xmem_data[123][1] ), .ZN(n29571) );
  AOI22_X1 U32439 ( .A1(n29566), .A2(\xmem_data[124][1] ), .B1(n29556), .B2(
        \xmem_data[125][1] ), .ZN(n29570) );
  AOI22_X1 U32440 ( .A1(n29568), .A2(\xmem_data[126][1] ), .B1(n3345), .B2(
        \xmem_data[127][1] ), .ZN(n29569) );
  AOI22_X1 U32441 ( .A1(n3166), .A2(\xmem_data[104][1] ), .B1(n3187), .B2(
        \xmem_data[105][1] ), .ZN(n29578) );
  AOI22_X1 U32442 ( .A1(n30764), .A2(\xmem_data[106][1] ), .B1(n29639), .B2(
        \xmem_data[107][1] ), .ZN(n29577) );
  AOI22_X1 U32443 ( .A1(n29547), .A2(\xmem_data[108][1] ), .B1(n29640), .B2(
        \xmem_data[109][1] ), .ZN(n29576) );
  AOI22_X1 U32444 ( .A1(n29574), .A2(\xmem_data[110][1] ), .B1(n29573), .B2(
        \xmem_data[111][1] ), .ZN(n29575) );
  AOI22_X1 U32445 ( .A1(n29580), .A2(\xmem_data[112][1] ), .B1(n29615), .B2(
        \xmem_data[113][1] ), .ZN(n29588) );
  AOI22_X1 U32446 ( .A1(n29581), .A2(\xmem_data[114][1] ), .B1(n17051), .B2(
        \xmem_data[115][1] ), .ZN(n29587) );
  AOI22_X1 U32447 ( .A1(n29583), .A2(\xmem_data[116][1] ), .B1(n29582), .B2(
        \xmem_data[117][1] ), .ZN(n29586) );
  AOI22_X1 U32448 ( .A1(n29584), .A2(\xmem_data[118][1] ), .B1(n22728), .B2(
        \xmem_data[119][1] ), .ZN(n29585) );
  AOI22_X1 U32449 ( .A1(n30743), .A2(\xmem_data[96][1] ), .B1(n29347), .B2(
        \xmem_data[97][1] ), .ZN(n29597) );
  AOI22_X1 U32450 ( .A1(n3239), .A2(\xmem_data[98][1] ), .B1(n29591), .B2(
        \xmem_data[99][1] ), .ZN(n29596) );
  AOI22_X1 U32451 ( .A1(n29604), .A2(\xmem_data[100][1] ), .B1(n28778), .B2(
        \xmem_data[101][1] ), .ZN(n29595) );
  AOI22_X1 U32452 ( .A1(n29593), .A2(\xmem_data[102][1] ), .B1(n27945), .B2(
        \xmem_data[103][1] ), .ZN(n29594) );
  AOI22_X2 U32453 ( .A1(n29601), .A2(n29600), .B1(n29599), .B2(n29598), .ZN(
        n33454) );
  AOI22_X1 U32454 ( .A1(n30191), .A2(\xmem_data[32][1] ), .B1(n29347), .B2(
        \xmem_data[33][1] ), .ZN(n29609) );
  AOI22_X1 U32455 ( .A1(n29603), .A2(\xmem_data[34][1] ), .B1(n30508), .B2(
        \xmem_data[35][1] ), .ZN(n29608) );
  AOI22_X1 U32456 ( .A1(n30665), .A2(\xmem_data[36][1] ), .B1(n30634), .B2(
        \xmem_data[37][1] ), .ZN(n29607) );
  AOI22_X1 U32457 ( .A1(n29649), .A2(\xmem_data[38][1] ), .B1(n3158), .B2(
        \xmem_data[39][1] ), .ZN(n29606) );
  NAND4_X1 U32458 ( .A1(n29609), .A2(n29608), .A3(n29607), .A4(n29606), .ZN(
        n29638) );
  AOI22_X1 U32459 ( .A1(n3161), .A2(\xmem_data[40][1] ), .B1(n3184), .B2(
        \xmem_data[41][1] ), .ZN(n29614) );
  AOI22_X1 U32460 ( .A1(n29610), .A2(\xmem_data[42][1] ), .B1(n29239), .B2(
        \xmem_data[43][1] ), .ZN(n29613) );
  AOI22_X1 U32461 ( .A1(n30766), .A2(\xmem_data[44][1] ), .B1(n30644), .B2(
        \xmem_data[45][1] ), .ZN(n29612) );
  AOI22_X1 U32462 ( .A1(n29641), .A2(\xmem_data[46][1] ), .B1(n3300), .B2(
        \xmem_data[47][1] ), .ZN(n29611) );
  NAND4_X1 U32463 ( .A1(n29614), .A2(n29613), .A3(n29612), .A4(n29611), .ZN(
        n29637) );
  AOI22_X1 U32464 ( .A1(n29616), .A2(\xmem_data[48][1] ), .B1(n29579), .B2(
        \xmem_data[49][1] ), .ZN(n29625) );
  AOI22_X1 U32465 ( .A1(n29617), .A2(\xmem_data[50][1] ), .B1(n27498), .B2(
        \xmem_data[51][1] ), .ZN(n29624) );
  AOI22_X1 U32466 ( .A1(n29619), .A2(\xmem_data[52][1] ), .B1(n29618), .B2(
        \xmem_data[53][1] ), .ZN(n29623) );
  AOI22_X1 U32467 ( .A1(n29621), .A2(\xmem_data[54][1] ), .B1(n3142), .B2(
        \xmem_data[55][1] ), .ZN(n29622) );
  NAND4_X1 U32468 ( .A1(n29625), .A2(n29624), .A3(n29623), .A4(n29622), .ZN(
        n29636) );
  AOI22_X1 U32469 ( .A1(n29788), .A2(\xmem_data[56][1] ), .B1(n30182), .B2(
        \xmem_data[57][1] ), .ZN(n29634) );
  AOI22_X1 U32470 ( .A1(n30215), .A2(\xmem_data[58][1] ), .B1(n29627), .B2(
        \xmem_data[59][1] ), .ZN(n29633) );
  AOI22_X1 U32471 ( .A1(n29630), .A2(\xmem_data[60][1] ), .B1(n27833), .B2(
        \xmem_data[61][1] ), .ZN(n29632) );
  AOI22_X1 U32472 ( .A1(n29667), .A2(\xmem_data[62][1] ), .B1(n3137), .B2(
        \xmem_data[63][1] ), .ZN(n29631) );
  NAND4_X1 U32473 ( .A1(n29634), .A2(n29633), .A3(n29632), .A4(n29631), .ZN(
        n29635) );
  OR4_X2 U32474 ( .A1(n29638), .A2(n29637), .A3(n29636), .A4(n29635), .ZN(
        n29682) );
  AOI22_X1 U32475 ( .A1(n3162), .A2(\xmem_data[8][1] ), .B1(n3184), .B2(
        \xmem_data[9][1] ), .ZN(n29645) );
  AOI22_X1 U32476 ( .A1(n30764), .A2(\xmem_data[10][1] ), .B1(n29639), .B2(
        \xmem_data[11][1] ), .ZN(n29644) );
  AOI22_X1 U32477 ( .A1(n29363), .A2(\xmem_data[12][1] ), .B1(n30765), .B2(
        \xmem_data[13][1] ), .ZN(n29643) );
  AOI22_X1 U32478 ( .A1(n29641), .A2(\xmem_data[14][1] ), .B1(n3302), .B2(
        \xmem_data[15][1] ), .ZN(n29642) );
  AOI22_X1 U32479 ( .A1(n27703), .A2(\xmem_data[0][1] ), .B1(n30730), .B2(
        \xmem_data[1][1] ), .ZN(n29653) );
  AOI22_X1 U32480 ( .A1(n3239), .A2(\xmem_data[2][1] ), .B1(n30083), .B2(
        \xmem_data[3][1] ), .ZN(n29652) );
  AOI22_X1 U32481 ( .A1(n27754), .A2(\xmem_data[4][1] ), .B1(n29739), .B2(
        \xmem_data[5][1] ), .ZN(n29651) );
  AOI22_X1 U32482 ( .A1(n29649), .A2(\xmem_data[6][1] ), .B1(n20776), .B2(
        \xmem_data[7][1] ), .ZN(n29650) );
  AOI22_X1 U32483 ( .A1(n28700), .A2(\xmem_data[26][1] ), .B1(n30292), .B2(
        \xmem_data[27][1] ), .ZN(n29654) );
  INV_X1 U32484 ( .A(n29654), .ZN(n29671) );
  AOI22_X1 U32485 ( .A1(n29656), .A2(\xmem_data[16][1] ), .B1(n29579), .B2(
        \xmem_data[17][1] ), .ZN(n29666) );
  AOI22_X1 U32486 ( .A1(n29658), .A2(\xmem_data[18][1] ), .B1(n29657), .B2(
        \xmem_data[19][1] ), .ZN(n29665) );
  AOI22_X1 U32487 ( .A1(n29660), .A2(\xmem_data[20][1] ), .B1(n29659), .B2(
        \xmem_data[21][1] ), .ZN(n29664) );
  AOI22_X1 U32488 ( .A1(n29662), .A2(\xmem_data[22][1] ), .B1(n29661), .B2(
        \xmem_data[23][1] ), .ZN(n29663) );
  NAND4_X1 U32489 ( .A1(n29666), .A2(n29665), .A3(n29664), .A4(n29663), .ZN(
        n29670) );
  AOI22_X1 U32490 ( .A1(n29667), .A2(\xmem_data[30][1] ), .B1(n3138), .B2(
        \xmem_data[31][1] ), .ZN(n29668) );
  INV_X1 U32491 ( .A(n29668), .ZN(n29669) );
  NOR3_X1 U32492 ( .A1(n29671), .A2(n29670), .A3(n29669), .ZN(n29679) );
  AOI22_X1 U32493 ( .A1(n27710), .A2(\xmem_data[24][1] ), .B1(n29753), .B2(
        \xmem_data[25][1] ), .ZN(n29673) );
  INV_X1 U32494 ( .A(n29673), .ZN(n29677) );
  AOI22_X1 U32495 ( .A1(n29674), .A2(\xmem_data[28][1] ), .B1(n29761), .B2(
        \xmem_data[29][1] ), .ZN(n29675) );
  INV_X1 U32496 ( .A(n29675), .ZN(n29676) );
  NOR2_X1 U32497 ( .A1(n29677), .A2(n29676), .ZN(n29678) );
  NAND4_X1 U32498 ( .A1(n3858), .A2(n3536), .A3(n29679), .A4(n29678), .ZN(
        n29680) );
  AOI22_X1 U32499 ( .A1(n29683), .A2(n29682), .B1(n29681), .B2(n29680), .ZN(
        n33455) );
  NAND2_X1 U32500 ( .A1(n33454), .A2(n33455), .ZN(n32603) );
  XNOR2_X1 U32501 ( .A(n32603), .B(\fmem_data[7][7] ), .ZN(n32193) );
  OAI22_X1 U32502 ( .A1(n32193), .A2(n35618), .B1(n29684), .B2(n35619), .ZN(
        n29693) );
  FA_X1 U32503 ( .A(n29687), .B(n29686), .CI(n29685), .CO(n29692), .S(n31185)
         );
  XNOR2_X1 U32504 ( .A(n29688), .B(n30339), .ZN(n31241) );
  FA_X1 U32505 ( .A(n29691), .B(n29690), .CI(n29689), .CO(n30146), .S(n31207)
         );
  FA_X1 U32506 ( .A(n29694), .B(n29693), .CI(n29692), .CO(n30339), .S(n31206)
         );
  XNOR2_X1 U32507 ( .A(n31658), .B(\fmem_data[30][1] ), .ZN(n32574) );
  XNOR2_X1 U32508 ( .A(n31659), .B(\fmem_data[30][1] ), .ZN(n33977) );
  OAI22_X1 U32509 ( .A1(n32574), .A2(n34788), .B1(n3560), .B2(n33977), .ZN(
        n31136) );
  AOI22_X1 U32510 ( .A1(n28717), .A2(\xmem_data[0][0] ), .B1(n29695), .B2(
        \xmem_data[1][0] ), .ZN(n29703) );
  AOI22_X1 U32511 ( .A1(n29696), .A2(\xmem_data[2][0] ), .B1(n3144), .B2(
        \xmem_data[3][0] ), .ZN(n29702) );
  AOI22_X1 U32512 ( .A1(n28136), .A2(\xmem_data[4][0] ), .B1(n26510), .B2(
        \xmem_data[5][0] ), .ZN(n29701) );
  AOI22_X1 U32513 ( .A1(n29790), .A2(\xmem_data[6][0] ), .B1(n29698), .B2(
        \xmem_data[7][0] ), .ZN(n29700) );
  AND4_X1 U32514 ( .A1(n29703), .A2(n29702), .A3(n29701), .A4(n29700), .ZN(
        n29732) );
  AOI22_X1 U32515 ( .A1(n29446), .A2(\xmem_data[12][0] ), .B1(n28738), .B2(
        \xmem_data[13][0] ), .ZN(n29713) );
  AOI22_X1 U32516 ( .A1(n29707), .A2(\xmem_data[10][0] ), .B1(n29706), .B2(
        \xmem_data[11][0] ), .ZN(n29712) );
  AOI22_X1 U32517 ( .A1(n29674), .A2(\xmem_data[8][0] ), .B1(n28786), .B2(
        \xmem_data[9][0] ), .ZN(n29711) );
  AOI22_X1 U32518 ( .A1(n29709), .A2(\xmem_data[14][0] ), .B1(n24640), .B2(
        \xmem_data[15][0] ), .ZN(n29710) );
  AOI22_X1 U32519 ( .A1(n3162), .A2(\xmem_data[20][0] ), .B1(n3187), .B2(
        \xmem_data[21][0] ), .ZN(n29720) );
  AOI22_X1 U32520 ( .A1(n29740), .A2(\xmem_data[18][0] ), .B1(n30892), .B2(
        \xmem_data[19][0] ), .ZN(n29719) );
  AOI22_X1 U32521 ( .A1(n27811), .A2(\xmem_data[16][0] ), .B1(n30090), .B2(
        \xmem_data[17][0] ), .ZN(n29718) );
  AND2_X1 U32522 ( .A1(n28754), .A2(\xmem_data[23][0] ), .ZN(n29715) );
  AOI21_X1 U32523 ( .B1(n29716), .B2(\xmem_data[22][0] ), .A(n29715), .ZN(
        n29717) );
  AOI22_X1 U32524 ( .A1(n28680), .A2(\xmem_data[24][0] ), .B1(n30644), .B2(
        \xmem_data[25][0] ), .ZN(n29730) );
  AOI22_X1 U32525 ( .A1(n3226), .A2(\xmem_data[26][0] ), .B1(n3307), .B2(
        \xmem_data[27][0] ), .ZN(n29729) );
  AOI22_X1 U32526 ( .A1(n29724), .A2(\xmem_data[28][0] ), .B1(n29723), .B2(
        \xmem_data[29][0] ), .ZN(n29728) );
  AOI22_X1 U32527 ( .A1(n29726), .A2(\xmem_data[30][0] ), .B1(n29725), .B2(
        \xmem_data[31][0] ), .ZN(n29727) );
  NAND4_X1 U32528 ( .A1(n29732), .A2(n29731), .A3(n3513), .A4(n3769), .ZN(
        n29734) );
  NAND2_X1 U32529 ( .A1(n29734), .A2(n29733), .ZN(n29843) );
  AOI22_X1 U32530 ( .A1(n29799), .A2(\xmem_data[72][0] ), .B1(n3170), .B2(
        \xmem_data[73][0] ), .ZN(n29738) );
  AOI22_X1 U32531 ( .A1(n29800), .A2(\xmem_data[74][0] ), .B1(n29762), .B2(
        \xmem_data[75][0] ), .ZN(n29737) );
  AOI22_X1 U32532 ( .A1(n29705), .A2(\xmem_data[76][0] ), .B1(n28238), .B2(
        \xmem_data[77][0] ), .ZN(n29736) );
  AOI22_X1 U32533 ( .A1(n29802), .A2(\xmem_data[78][0] ), .B1(n20716), .B2(
        \xmem_data[79][0] ), .ZN(n29735) );
  NAND4_X1 U32534 ( .A1(n29738), .A2(n29737), .A3(n29736), .A4(n29735), .ZN(
        n29752) );
  AOI22_X1 U32535 ( .A1(n30635), .A2(\xmem_data[80][0] ), .B1(n29592), .B2(
        \xmem_data[81][0] ), .ZN(n29745) );
  AOI22_X1 U32536 ( .A1(n29740), .A2(\xmem_data[82][0] ), .B1(n29807), .B2(
        \xmem_data[83][0] ), .ZN(n29744) );
  AOI22_X1 U32537 ( .A1(n3165), .A2(\xmem_data[84][0] ), .B1(n3191), .B2(
        \xmem_data[85][0] ), .ZN(n29743) );
  AND2_X1 U32538 ( .A1(n29639), .A2(\xmem_data[87][0] ), .ZN(n29741) );
  AOI21_X1 U32539 ( .B1(n30715), .B2(\xmem_data[86][0] ), .A(n29741), .ZN(
        n29742) );
  NAND4_X1 U32540 ( .A1(n29745), .A2(n29744), .A3(n29743), .A4(n29742), .ZN(
        n29751) );
  AOI22_X1 U32541 ( .A1(n28680), .A2(\xmem_data[88][0] ), .B1(n30266), .B2(
        \xmem_data[89][0] ), .ZN(n29749) );
  AOI22_X1 U32542 ( .A1(n29817), .A2(\xmem_data[90][0] ), .B1(n3271), .B2(
        \xmem_data[91][0] ), .ZN(n29748) );
  AOI22_X1 U32543 ( .A1(n29777), .A2(\xmem_data[92][0] ), .B1(n29776), .B2(
        \xmem_data[93][0] ), .ZN(n29747) );
  AOI22_X1 U32544 ( .A1(n27806), .A2(\xmem_data[94][0] ), .B1(n14982), .B2(
        \xmem_data[95][0] ), .ZN(n29746) );
  NAND4_X1 U32545 ( .A1(n29749), .A2(n29748), .A3(n29747), .A4(n29746), .ZN(
        n29750) );
  AOI22_X1 U32546 ( .A1(n28765), .A2(\xmem_data[64][0] ), .B1(n29695), .B2(
        \xmem_data[65][0] ), .ZN(n29757) );
  AOI22_X1 U32547 ( .A1(n29830), .A2(\xmem_data[66][0] ), .B1(n21308), .B2(
        \xmem_data[67][0] ), .ZN(n29756) );
  AOI22_X1 U32548 ( .A1(n29788), .A2(\xmem_data[68][0] ), .B1(n29672), .B2(
        \xmem_data[69][0] ), .ZN(n29755) );
  AOI22_X1 U32549 ( .A1(n29790), .A2(\xmem_data[70][0] ), .B1(n29832), .B2(
        \xmem_data[71][0] ), .ZN(n29754) );
  NAND4_X1 U32550 ( .A1(n29757), .A2(n29756), .A3(n29755), .A4(n29754), .ZN(
        n29759) );
  AOI22_X1 U32551 ( .A1(n29400), .A2(\xmem_data[40][0] ), .B1(n27833), .B2(
        \xmem_data[41][0] ), .ZN(n29767) );
  AOI22_X1 U32552 ( .A1(n29707), .A2(\xmem_data[42][0] ), .B1(n29762), .B2(
        \xmem_data[43][0] ), .ZN(n29766) );
  AOI22_X1 U32553 ( .A1(n29390), .A2(\xmem_data[44][0] ), .B1(n29704), .B2(
        \xmem_data[45][0] ), .ZN(n29765) );
  AOI22_X1 U32554 ( .A1(n29763), .A2(\xmem_data[46][0] ), .B1(n23792), .B2(
        \xmem_data[47][0] ), .ZN(n29764) );
  NAND4_X1 U32555 ( .A1(n29767), .A2(n29766), .A3(n29765), .A4(n29764), .ZN(
        n29784) );
  AOI22_X1 U32556 ( .A1(n29604), .A2(\xmem_data[48][0] ), .B1(n30249), .B2(
        \xmem_data[49][0] ), .ZN(n29775) );
  AOI22_X1 U32557 ( .A1(n29771), .A2(\xmem_data[50][0] ), .B1(n25607), .B2(
        \xmem_data[51][0] ), .ZN(n29774) );
  AOI22_X1 U32558 ( .A1(n3164), .A2(\xmem_data[52][0] ), .B1(n3183), .B2(
        \xmem_data[53][0] ), .ZN(n29773) );
  AOI22_X1 U32559 ( .A1(n30062), .A2(\xmem_data[54][0] ), .B1(n20815), .B2(
        \xmem_data[55][0] ), .ZN(n29772) );
  NAND4_X1 U32560 ( .A1(n29775), .A2(n29774), .A3(n29773), .A4(n29772), .ZN(
        n29783) );
  AOI22_X1 U32561 ( .A1(n29815), .A2(\xmem_data[56][0] ), .B1(n30716), .B2(
        \xmem_data[57][0] ), .ZN(n29781) );
  AOI22_X1 U32562 ( .A1(n3226), .A2(\xmem_data[58][0] ), .B1(n3151), .B2(
        \xmem_data[59][0] ), .ZN(n29780) );
  AOI22_X1 U32563 ( .A1(n29777), .A2(\xmem_data[60][0] ), .B1(n29776), .B2(
        \xmem_data[61][0] ), .ZN(n29779) );
  AOI22_X1 U32564 ( .A1(n28681), .A2(\xmem_data[62][0] ), .B1(n17051), .B2(
        \xmem_data[63][0] ), .ZN(n29778) );
  NAND4_X1 U32565 ( .A1(n29781), .A2(n29780), .A3(n29779), .A4(n29778), .ZN(
        n29782) );
  AOI22_X1 U32566 ( .A1(n29786), .A2(\xmem_data[32][0] ), .B1(n29785), .B2(
        \xmem_data[33][0] ), .ZN(n29794) );
  AOI22_X1 U32567 ( .A1(n29787), .A2(\xmem_data[34][0] ), .B1(n20828), .B2(
        \xmem_data[35][0] ), .ZN(n29793) );
  AOI22_X1 U32568 ( .A1(n28136), .A2(\xmem_data[36][0] ), .B1(n30100), .B2(
        \xmem_data[37][0] ), .ZN(n29792) );
  AOI22_X1 U32569 ( .A1(n28138), .A2(\xmem_data[38][0] ), .B1(n29789), .B2(
        \xmem_data[39][0] ), .ZN(n29791) );
  NAND4_X1 U32570 ( .A1(n29794), .A2(n29793), .A3(n29792), .A4(n29791), .ZN(
        n29796) );
  AOI22_X1 U32571 ( .A1(n29799), .A2(\xmem_data[104][0] ), .B1(n29495), .B2(
        \xmem_data[105][0] ), .ZN(n29806) );
  AOI22_X1 U32572 ( .A1(n29800), .A2(\xmem_data[106][0] ), .B1(n3375), .B2(
        \xmem_data[107][0] ), .ZN(n29805) );
  AOI22_X1 U32573 ( .A1(n30191), .A2(\xmem_data[108][0] ), .B1(n29482), .B2(
        \xmem_data[109][0] ), .ZN(n29804) );
  AOI22_X1 U32574 ( .A1(n29802), .A2(\xmem_data[110][0] ), .B1(n24556), .B2(
        \xmem_data[111][0] ), .ZN(n29803) );
  NAND4_X1 U32575 ( .A1(n29806), .A2(n29805), .A3(n29804), .A4(n29803), .ZN(
        n29828) );
  AOI22_X1 U32576 ( .A1(n3167), .A2(\xmem_data[116][0] ), .B1(n3190), .B2(
        \xmem_data[117][0] ), .ZN(n29814) );
  AOI22_X1 U32577 ( .A1(n29808), .A2(\xmem_data[114][0] ), .B1(n29807), .B2(
        \xmem_data[115][0] ), .ZN(n29813) );
  AOI22_X1 U32578 ( .A1(n30250), .A2(\xmem_data[112][0] ), .B1(n29768), .B2(
        \xmem_data[113][0] ), .ZN(n29812) );
  AND2_X1 U32579 ( .A1(n30309), .A2(\xmem_data[119][0] ), .ZN(n29809) );
  AOI21_X1 U32580 ( .B1(n29810), .B2(\xmem_data[118][0] ), .A(n29809), .ZN(
        n29811) );
  NAND4_X1 U32581 ( .A1(n29814), .A2(n29813), .A3(n29812), .A4(n29811), .ZN(
        n29827) );
  AOI22_X1 U32582 ( .A1(n30717), .A2(\xmem_data[120][0] ), .B1(n30716), .B2(
        \xmem_data[121][0] ), .ZN(n29825) );
  AOI22_X1 U32583 ( .A1(n29817), .A2(\xmem_data[122][0] ), .B1(n29816), .B2(
        \xmem_data[123][0] ), .ZN(n29824) );
  AOI22_X1 U32584 ( .A1(n29819), .A2(\xmem_data[124][0] ), .B1(n29818), .B2(
        \xmem_data[125][0] ), .ZN(n29823) );
  AOI22_X1 U32585 ( .A1(n29821), .A2(\xmem_data[126][0] ), .B1(n29820), .B2(
        \xmem_data[127][0] ), .ZN(n29822) );
  NAND4_X1 U32586 ( .A1(n29825), .A2(n29824), .A3(n29823), .A4(n29822), .ZN(
        n29826) );
  AOI22_X1 U32587 ( .A1(n28765), .A2(\xmem_data[96][0] ), .B1(n29695), .B2(
        \xmem_data[97][0] ), .ZN(n29836) );
  AOI22_X1 U32588 ( .A1(n29830), .A2(\xmem_data[98][0] ), .B1(n27813), .B2(
        \xmem_data[99][0] ), .ZN(n29835) );
  AOI22_X1 U32589 ( .A1(n28734), .A2(\xmem_data[100][0] ), .B1(n29831), .B2(
        \xmem_data[101][0] ), .ZN(n29834) );
  AOI22_X1 U32590 ( .A1(n30279), .A2(\xmem_data[102][0] ), .B1(n29832), .B2(
        \xmem_data[103][0] ), .ZN(n29833) );
  NAND4_X1 U32591 ( .A1(n29836), .A2(n29835), .A3(n29834), .A4(n29833), .ZN(
        n29838) );
  INV_X1 U32592 ( .A(n35656), .ZN(n29844) );
  OAI22_X1 U32593 ( .A1(n32576), .A2(n33954), .B1(n33955), .B2(n33956), .ZN(
        n31134) );
  FA_X1 U32594 ( .A(n29847), .B(n29846), .CI(n29845), .CO(n28930), .S(n31144)
         );
  OR2_X1 U32595 ( .A1(n31143), .A2(n31144), .ZN(n30126) );
  XNOR2_X1 U32596 ( .A(n32023), .B(\fmem_data[11][3] ), .ZN(n32234) );
  XNOR2_X1 U32597 ( .A(n31247), .B(\fmem_data[11][3] ), .ZN(n32260) );
  AOI22_X1 U32598 ( .A1(n29849), .A2(\xmem_data[32][0] ), .B1(n29848), .B2(
        \xmem_data[33][0] ), .ZN(n29859) );
  AOI22_X1 U32599 ( .A1(n29851), .A2(\xmem_data[34][0] ), .B1(n29850), .B2(
        \xmem_data[35][0] ), .ZN(n29858) );
  AOI22_X1 U32600 ( .A1(n29853), .A2(\xmem_data[36][0] ), .B1(n29852), .B2(
        \xmem_data[37][0] ), .ZN(n29857) );
  AOI22_X1 U32601 ( .A1(n29855), .A2(\xmem_data[38][0] ), .B1(n29854), .B2(
        \xmem_data[39][0] ), .ZN(n29856) );
  NAND4_X1 U32602 ( .A1(n29859), .A2(n29858), .A3(n29857), .A4(n29856), .ZN(
        n29891) );
  AOI22_X1 U32603 ( .A1(n29860), .A2(\xmem_data[40][0] ), .B1(n29942), .B2(
        \xmem_data[41][0] ), .ZN(n29864) );
  AOI22_X1 U32604 ( .A1(n29943), .A2(\xmem_data[42][0] ), .B1(n3194), .B2(
        \xmem_data[43][0] ), .ZN(n29863) );
  AOI22_X1 U32605 ( .A1(n29945), .A2(\xmem_data[44][0] ), .B1(n29944), .B2(
        \xmem_data[45][0] ), .ZN(n29862) );
  AOI22_X1 U32606 ( .A1(n29947), .A2(\xmem_data[46][0] ), .B1(n29946), .B2(
        \xmem_data[47][0] ), .ZN(n29861) );
  NAND4_X1 U32607 ( .A1(n29864), .A2(n29863), .A3(n29862), .A4(n29861), .ZN(
        n29890) );
  AOI22_X1 U32608 ( .A1(n29866), .A2(\xmem_data[48][0] ), .B1(n29865), .B2(
        \xmem_data[49][0] ), .ZN(n29875) );
  AOI22_X1 U32609 ( .A1(n29868), .A2(\xmem_data[50][0] ), .B1(n29867), .B2(
        \xmem_data[51][0] ), .ZN(n29874) );
  AOI22_X1 U32610 ( .A1(n29870), .A2(\xmem_data[52][0] ), .B1(n29869), .B2(
        \xmem_data[53][0] ), .ZN(n29873) );
  AOI22_X1 U32611 ( .A1(n29871), .A2(\xmem_data[54][0] ), .B1(n29920), .B2(
        \xmem_data[55][0] ), .ZN(n29872) );
  NAND4_X1 U32612 ( .A1(n29875), .A2(n29874), .A3(n29873), .A4(n29872), .ZN(
        n29889) );
  AOI22_X1 U32613 ( .A1(n29877), .A2(\xmem_data[56][0] ), .B1(n29876), .B2(
        \xmem_data[57][0] ), .ZN(n29887) );
  AOI22_X1 U32614 ( .A1(n29879), .A2(\xmem_data[58][0] ), .B1(n29878), .B2(
        \xmem_data[59][0] ), .ZN(n29886) );
  AOI22_X1 U32615 ( .A1(n29881), .A2(\xmem_data[60][0] ), .B1(n29880), .B2(
        \xmem_data[61][0] ), .ZN(n29885) );
  AOI22_X1 U32616 ( .A1(n29883), .A2(\xmem_data[62][0] ), .B1(n29882), .B2(
        \xmem_data[63][0] ), .ZN(n29884) );
  NAND4_X1 U32617 ( .A1(n29887), .A2(n29886), .A3(n29885), .A4(n29884), .ZN(
        n29888) );
  OR4_X1 U32618 ( .A1(n29891), .A2(n29890), .A3(n29889), .A4(n29888), .ZN(
        n29936) );
  AOI22_X1 U32619 ( .A1(n29893), .A2(\xmem_data[0][0] ), .B1(n29892), .B2(
        \xmem_data[1][0] ), .ZN(n29903) );
  AOI22_X1 U32620 ( .A1(n29895), .A2(\xmem_data[2][0] ), .B1(n29894), .B2(
        \xmem_data[3][0] ), .ZN(n29902) );
  AOI22_X1 U32621 ( .A1(n29897), .A2(\xmem_data[4][0] ), .B1(n29896), .B2(
        \xmem_data[5][0] ), .ZN(n29901) );
  AOI22_X1 U32622 ( .A1(n29899), .A2(\xmem_data[6][0] ), .B1(n29898), .B2(
        \xmem_data[7][0] ), .ZN(n29900) );
  NAND4_X1 U32623 ( .A1(n29903), .A2(n29902), .A3(n29901), .A4(n29900), .ZN(
        n29933) );
  AOI22_X1 U32624 ( .A1(n29904), .A2(\xmem_data[8][0] ), .B1(n29976), .B2(
        \xmem_data[9][0] ), .ZN(n29913) );
  AOI22_X1 U32625 ( .A1(n29905), .A2(\xmem_data[10][0] ), .B1(n3194), .B2(
        \xmem_data[11][0] ), .ZN(n29912) );
  AOI22_X1 U32626 ( .A1(n29907), .A2(\xmem_data[12][0] ), .B1(n29906), .B2(
        \xmem_data[13][0] ), .ZN(n29911) );
  AOI22_X1 U32627 ( .A1(n29909), .A2(\xmem_data[14][0] ), .B1(n29908), .B2(
        \xmem_data[15][0] ), .ZN(n29910) );
  NAND4_X1 U32628 ( .A1(n29913), .A2(n29912), .A3(n29911), .A4(n29910), .ZN(
        n29932) );
  AOI22_X1 U32629 ( .A1(n29915), .A2(\xmem_data[16][0] ), .B1(n29914), .B2(
        \xmem_data[17][0] ), .ZN(n29925) );
  AOI22_X1 U32630 ( .A1(n29917), .A2(\xmem_data[18][0] ), .B1(n29916), .B2(
        \xmem_data[19][0] ), .ZN(n29924) );
  AOI22_X1 U32631 ( .A1(n29919), .A2(\xmem_data[20][0] ), .B1(n29918), .B2(
        \xmem_data[21][0] ), .ZN(n29923) );
  AOI22_X1 U32632 ( .A1(n29921), .A2(\xmem_data[22][0] ), .B1(n29920), .B2(
        \xmem_data[23][0] ), .ZN(n29922) );
  NAND4_X1 U32633 ( .A1(n29925), .A2(n29924), .A3(n29923), .A4(n29922), .ZN(
        n29931) );
  AOI22_X1 U32634 ( .A1(n3243), .A2(\xmem_data[24][0] ), .B1(n3242), .B2(
        \xmem_data[25][0] ), .ZN(n29929) );
  AOI22_X1 U32635 ( .A1(n3235), .A2(\xmem_data[26][0] ), .B1(n3238), .B2(
        \xmem_data[27][0] ), .ZN(n29928) );
  AOI22_X1 U32636 ( .A1(n3236), .A2(\xmem_data[28][0] ), .B1(n3225), .B2(
        \xmem_data[29][0] ), .ZN(n29927) );
  AOI22_X1 U32637 ( .A1(n3237), .A2(\xmem_data[30][0] ), .B1(n3234), .B2(
        \xmem_data[31][0] ), .ZN(n29926) );
  NAND4_X1 U32638 ( .A1(n29929), .A2(n29928), .A3(n29927), .A4(n29926), .ZN(
        n29930) );
  OR4_X1 U32639 ( .A1(n29933), .A2(n29932), .A3(n29931), .A4(n29930), .ZN(
        n29934) );
  AOI22_X1 U32640 ( .A1(n29937), .A2(n29936), .B1(n29935), .B2(n29934), .ZN(
        n30012) );
  AOI22_X1 U32641 ( .A1(n29966), .A2(\xmem_data[64][0] ), .B1(n29965), .B2(
        \xmem_data[65][0] ), .ZN(n29941) );
  AOI22_X1 U32642 ( .A1(n29968), .A2(\xmem_data[66][0] ), .B1(n29967), .B2(
        \xmem_data[67][0] ), .ZN(n29940) );
  AOI22_X1 U32643 ( .A1(n29969), .A2(\xmem_data[68][0] ), .B1(n29896), .B2(
        \xmem_data[69][0] ), .ZN(n29939) );
  AOI22_X1 U32644 ( .A1(n29971), .A2(\xmem_data[70][0] ), .B1(n29970), .B2(
        \xmem_data[71][0] ), .ZN(n29938) );
  NAND4_X1 U32645 ( .A1(n29941), .A2(n29940), .A3(n29939), .A4(n29938), .ZN(
        n29964) );
  AOI22_X1 U32646 ( .A1(n29977), .A2(\xmem_data[72][0] ), .B1(n29942), .B2(
        \xmem_data[73][0] ), .ZN(n29951) );
  AOI22_X1 U32647 ( .A1(n29943), .A2(\xmem_data[74][0] ), .B1(n3194), .B2(
        \xmem_data[75][0] ), .ZN(n29950) );
  AOI22_X1 U32648 ( .A1(n29945), .A2(\xmem_data[76][0] ), .B1(n29944), .B2(
        \xmem_data[77][0] ), .ZN(n29949) );
  AOI22_X1 U32649 ( .A1(n29947), .A2(\xmem_data[78][0] ), .B1(n29946), .B2(
        \xmem_data[79][0] ), .ZN(n29948) );
  NAND4_X1 U32650 ( .A1(n29951), .A2(n29950), .A3(n29949), .A4(n29948), .ZN(
        n29963) );
  AOI22_X1 U32651 ( .A1(n29988), .A2(\xmem_data[80][0] ), .B1(n29987), .B2(
        \xmem_data[81][0] ), .ZN(n29956) );
  AOI22_X1 U32652 ( .A1(n29990), .A2(\xmem_data[82][0] ), .B1(n29989), .B2(
        \xmem_data[83][0] ), .ZN(n29955) );
  AOI22_X1 U32653 ( .A1(n29992), .A2(\xmem_data[84][0] ), .B1(n29991), .B2(
        \xmem_data[85][0] ), .ZN(n29954) );
  AOI22_X1 U32654 ( .A1(n29994), .A2(\xmem_data[86][0] ), .B1(n29952), .B2(
        \xmem_data[87][0] ), .ZN(n29953) );
  NAND4_X1 U32655 ( .A1(n29956), .A2(n29955), .A3(n29954), .A4(n29953), .ZN(
        n29962) );
  AOI22_X1 U32656 ( .A1(n3243), .A2(\xmem_data[88][0] ), .B1(n3242), .B2(
        \xmem_data[89][0] ), .ZN(n29960) );
  AOI22_X1 U32657 ( .A1(n3235), .A2(\xmem_data[90][0] ), .B1(n3238), .B2(
        \xmem_data[91][0] ), .ZN(n29959) );
  AOI22_X1 U32658 ( .A1(n3236), .A2(\xmem_data[92][0] ), .B1(n3225), .B2(
        \xmem_data[93][0] ), .ZN(n29958) );
  AOI22_X1 U32659 ( .A1(n3237), .A2(\xmem_data[94][0] ), .B1(n3234), .B2(
        \xmem_data[95][0] ), .ZN(n29957) );
  NAND4_X1 U32660 ( .A1(n29960), .A2(n29959), .A3(n29958), .A4(n29957), .ZN(
        n29961) );
  OR4_X1 U32661 ( .A1(n29964), .A2(n29963), .A3(n29962), .A4(n29961), .ZN(
        n30010) );
  AOI22_X1 U32662 ( .A1(n29966), .A2(\xmem_data[96][0] ), .B1(n29965), .B2(
        \xmem_data[97][0] ), .ZN(n29975) );
  AOI22_X1 U32663 ( .A1(n29968), .A2(\xmem_data[98][0] ), .B1(n29967), .B2(
        \xmem_data[99][0] ), .ZN(n29974) );
  AOI22_X1 U32664 ( .A1(n29969), .A2(\xmem_data[100][0] ), .B1(n29896), .B2(
        \xmem_data[101][0] ), .ZN(n29973) );
  AOI22_X1 U32665 ( .A1(n29971), .A2(\xmem_data[102][0] ), .B1(n29970), .B2(
        \xmem_data[103][0] ), .ZN(n29972) );
  NAND4_X1 U32666 ( .A1(n29975), .A2(n29974), .A3(n29973), .A4(n29972), .ZN(
        n30006) );
  AOI22_X1 U32667 ( .A1(n29977), .A2(\xmem_data[104][0] ), .B1(n29976), .B2(
        \xmem_data[105][0] ), .ZN(n29986) );
  AOI22_X1 U32668 ( .A1(n29978), .A2(\xmem_data[106][0] ), .B1(n3194), .B2(
        \xmem_data[107][0] ), .ZN(n29985) );
  AOI22_X1 U32669 ( .A1(n29980), .A2(\xmem_data[108][0] ), .B1(n29979), .B2(
        \xmem_data[109][0] ), .ZN(n29984) );
  AOI22_X1 U32670 ( .A1(n29982), .A2(\xmem_data[110][0] ), .B1(n29981), .B2(
        \xmem_data[111][0] ), .ZN(n29983) );
  NAND4_X1 U32671 ( .A1(n29986), .A2(n29985), .A3(n29984), .A4(n29983), .ZN(
        n30005) );
  AOI22_X1 U32672 ( .A1(n29988), .A2(\xmem_data[112][0] ), .B1(n29987), .B2(
        \xmem_data[113][0] ), .ZN(n29998) );
  AOI22_X1 U32673 ( .A1(n29990), .A2(\xmem_data[114][0] ), .B1(n29989), .B2(
        \xmem_data[115][0] ), .ZN(n29997) );
  AOI22_X1 U32674 ( .A1(n29992), .A2(\xmem_data[116][0] ), .B1(n29991), .B2(
        \xmem_data[117][0] ), .ZN(n29996) );
  AOI22_X1 U32675 ( .A1(n29994), .A2(\xmem_data[118][0] ), .B1(n29993), .B2(
        \xmem_data[119][0] ), .ZN(n29995) );
  NAND4_X1 U32676 ( .A1(n29998), .A2(n29997), .A3(n29996), .A4(n29995), .ZN(
        n30004) );
  AOI22_X1 U32677 ( .A1(n3243), .A2(\xmem_data[120][0] ), .B1(n3242), .B2(
        \xmem_data[121][0] ), .ZN(n30002) );
  AOI22_X1 U32678 ( .A1(n3235), .A2(\xmem_data[122][0] ), .B1(n3238), .B2(
        \xmem_data[123][0] ), .ZN(n30001) );
  AOI22_X1 U32679 ( .A1(n3236), .A2(\xmem_data[124][0] ), .B1(n3225), .B2(
        \xmem_data[125][0] ), .ZN(n30000) );
  AOI22_X1 U32680 ( .A1(n3237), .A2(\xmem_data[126][0] ), .B1(n3234), .B2(
        \xmem_data[127][0] ), .ZN(n29999) );
  NAND4_X1 U32681 ( .A1(n30002), .A2(n30001), .A3(n30000), .A4(n29999), .ZN(
        n30003) );
  INV_X1 U32682 ( .A(n35701), .ZN(n30013) );
  AOI22_X1 U32683 ( .A1(n29481), .A2(\xmem_data[40][0] ), .B1(n29646), .B2(
        \xmem_data[41][0] ), .ZN(n30017) );
  AOI22_X1 U32684 ( .A1(n30171), .A2(\xmem_data[42][0] ), .B1(n29403), .B2(
        \xmem_data[43][0] ), .ZN(n30016) );
  AOI22_X1 U32685 ( .A1(n28751), .A2(\xmem_data[44][0] ), .B1(n30249), .B2(
        \xmem_data[45][0] ), .ZN(n30015) );
  AOI22_X1 U32686 ( .A1(n30304), .A2(\xmem_data[46][0] ), .B1(n27517), .B2(
        \xmem_data[47][0] ), .ZN(n30014) );
  NAND4_X1 U32687 ( .A1(n30017), .A2(n30016), .A3(n30015), .A4(n30014), .ZN(
        n30018) );
  AOI22_X1 U32688 ( .A1(n29481), .A2(\xmem_data[8][0] ), .B1(n29482), .B2(
        \xmem_data[9][0] ), .ZN(n30022) );
  AOI22_X1 U32689 ( .A1(n30171), .A2(\xmem_data[10][0] ), .B1(n28089), .B2(
        \xmem_data[11][0] ), .ZN(n30021) );
  AOI22_X1 U32690 ( .A1(n30665), .A2(\xmem_data[12][0] ), .B1(n27753), .B2(
        \xmem_data[13][0] ), .ZN(n30020) );
  AOI22_X1 U32691 ( .A1(n30304), .A2(\xmem_data[14][0] ), .B1(n16988), .B2(
        \xmem_data[15][0] ), .ZN(n30019) );
  NAND4_X1 U32692 ( .A1(n30022), .A2(n30021), .A3(n30020), .A4(n30019), .ZN(
        n30042) );
  AOI22_X1 U32693 ( .A1(n3210), .A2(\xmem_data[24][0] ), .B1(n30256), .B2(
        \xmem_data[25][0] ), .ZN(n30026) );
  AOI22_X1 U32694 ( .A1(n30048), .A2(\xmem_data[26][0] ), .B1(n20770), .B2(
        \xmem_data[27][0] ), .ZN(n30025) );
  AOI22_X1 U32695 ( .A1(n30199), .A2(\xmem_data[28][0] ), .B1(n3421), .B2(
        \xmem_data[29][0] ), .ZN(n30024) );
  AOI22_X1 U32696 ( .A1(n30200), .A2(\xmem_data[30][0] ), .B1(n3142), .B2(
        \xmem_data[31][0] ), .ZN(n30023) );
  NAND4_X1 U32697 ( .A1(n30026), .A2(n30025), .A3(n30024), .A4(n30023), .ZN(
        n30027) );
  NAND2_X1 U32698 ( .A1(n30027), .A2(n30228), .ZN(n30040) );
  AOI22_X1 U32699 ( .A1(n3211), .A2(\xmem_data[120][0] ), .B1(n30256), .B2(
        \xmem_data[121][0] ), .ZN(n30031) );
  AOI22_X1 U32700 ( .A1(n30258), .A2(\xmem_data[122][0] ), .B1(n30257), .B2(
        \xmem_data[123][0] ), .ZN(n30030) );
  AOI22_X1 U32701 ( .A1(n30260), .A2(\xmem_data[124][0] ), .B1(n3420), .B2(
        \xmem_data[125][0] ), .ZN(n30029) );
  AOI22_X1 U32702 ( .A1(n30200), .A2(\xmem_data[126][0] ), .B1(n3348), .B2(
        \xmem_data[127][0] ), .ZN(n30028) );
  NAND4_X1 U32703 ( .A1(n30031), .A2(n30030), .A3(n30029), .A4(n30028), .ZN(
        n30032) );
  NAND2_X1 U32704 ( .A1(n30032), .A2(n30287), .ZN(n30039) );
  AOI22_X1 U32705 ( .A1(n3210), .A2(\xmem_data[88][0] ), .B1(n30256), .B2(
        \xmem_data[89][0] ), .ZN(n30036) );
  AOI22_X1 U32706 ( .A1(n30258), .A2(\xmem_data[90][0] ), .B1(n30257), .B2(
        \xmem_data[91][0] ), .ZN(n30035) );
  AOI22_X1 U32707 ( .A1(n30260), .A2(\xmem_data[92][0] ), .B1(n3421), .B2(
        \xmem_data[93][0] ), .ZN(n30034) );
  AOI22_X1 U32708 ( .A1(n30320), .A2(\xmem_data[94][0] ), .B1(n3352), .B2(
        \xmem_data[95][0] ), .ZN(n30033) );
  NAND4_X1 U32709 ( .A1(n30036), .A2(n30035), .A3(n30034), .A4(n30033), .ZN(
        n30037) );
  NAND2_X1 U32710 ( .A1(n30037), .A2(n30188), .ZN(n30038) );
  NAND3_X1 U32711 ( .A1(n30040), .A2(n30039), .A3(n30038), .ZN(n30041) );
  AOI22_X1 U32712 ( .A1(n27710), .A2(\xmem_data[0][0] ), .B1(n30182), .B2(
        \xmem_data[1][0] ), .ZN(n30046) );
  AOI22_X1 U32713 ( .A1(n28207), .A2(\xmem_data[2][0] ), .B1(n30278), .B2(
        \xmem_data[3][0] ), .ZN(n30045) );
  AOI22_X1 U32714 ( .A1(n29630), .A2(\xmem_data[4][0] ), .B1(n27833), .B2(
        \xmem_data[5][0] ), .ZN(n30044) );
  AOI22_X1 U32715 ( .A1(n30219), .A2(\xmem_data[6][0] ), .B1(n3131), .B2(
        \xmem_data[7][0] ), .ZN(n30043) );
  NAND4_X1 U32716 ( .A1(n30046), .A2(n30045), .A3(n30044), .A4(n30043), .ZN(
        n30047) );
  AOI22_X1 U32717 ( .A1(n3210), .A2(\xmem_data[56][0] ), .B1(n3193), .B2(
        \xmem_data[57][0] ), .ZN(n30052) );
  AOI22_X1 U32718 ( .A1(n30048), .A2(\xmem_data[58][0] ), .B1(n27717), .B2(
        \xmem_data[59][0] ), .ZN(n30051) );
  AOI22_X1 U32719 ( .A1(n30318), .A2(\xmem_data[60][0] ), .B1(n30317), .B2(
        \xmem_data[61][0] ), .ZN(n30050) );
  AOI22_X1 U32720 ( .A1(n30200), .A2(\xmem_data[62][0] ), .B1(n3153), .B2(
        \xmem_data[63][0] ), .ZN(n30049) );
  NAND4_X1 U32721 ( .A1(n30052), .A2(n30051), .A3(n30050), .A4(n30049), .ZN(
        n30053) );
  NAND4_X1 U32722 ( .A1(n30057), .A2(n30056), .A3(n30055), .A4(n30054), .ZN(
        n30122) );
  AOI22_X1 U32723 ( .A1(n3160), .A2(\xmem_data[112][0] ), .B1(n3185), .B2(
        \xmem_data[113][0] ), .ZN(n30061) );
  AOI22_X1 U32724 ( .A1(n30715), .A2(\xmem_data[114][0] ), .B1(n28754), .B2(
        \xmem_data[115][0] ), .ZN(n30060) );
  AOI22_X1 U32725 ( .A1(n29815), .A2(\xmem_data[116][0] ), .B1(n30170), .B2(
        \xmem_data[117][0] ), .ZN(n30059) );
  AOI22_X1 U32726 ( .A1(n30270), .A2(\xmem_data[118][0] ), .B1(n30269), .B2(
        \xmem_data[119][0] ), .ZN(n30058) );
  NAND4_X1 U32727 ( .A1(n30061), .A2(n30060), .A3(n30059), .A4(n30058), .ZN(
        n30069) );
  AOI22_X1 U32728 ( .A1(n3167), .A2(\xmem_data[48][0] ), .B1(n3190), .B2(
        \xmem_data[49][0] ), .ZN(n30067) );
  AOI22_X1 U32729 ( .A1(n30062), .A2(\xmem_data[50][0] ), .B1(n30309), .B2(
        \xmem_data[51][0] ), .ZN(n30066) );
  AOI22_X1 U32730 ( .A1(n30076), .A2(\xmem_data[52][0] ), .B1(n30716), .B2(
        \xmem_data[53][0] ), .ZN(n30065) );
  AOI22_X1 U32731 ( .A1(n30205), .A2(\xmem_data[54][0] ), .B1(n30311), .B2(
        \xmem_data[55][0] ), .ZN(n30064) );
  NAND4_X1 U32732 ( .A1(n30067), .A2(n30066), .A3(n30065), .A4(n30064), .ZN(
        n30068) );
  AOI22_X1 U32733 ( .A1(n3165), .A2(\xmem_data[16][0] ), .B1(n3191), .B2(
        \xmem_data[17][0] ), .ZN(n30074) );
  AOI22_X1 U32734 ( .A1(n30070), .A2(\xmem_data[18][0] ), .B1(n28147), .B2(
        \xmem_data[19][0] ), .ZN(n30073) );
  AOI22_X1 U32735 ( .A1(n29363), .A2(\xmem_data[20][0] ), .B1(n29640), .B2(
        \xmem_data[21][0] ), .ZN(n30072) );
  AOI22_X1 U32736 ( .A1(n30205), .A2(\xmem_data[22][0] ), .B1(n29379), .B2(
        \xmem_data[23][0] ), .ZN(n30071) );
  NAND4_X1 U32737 ( .A1(n30074), .A2(n30073), .A3(n30072), .A4(n30071), .ZN(
        n30082) );
  AOI22_X1 U32738 ( .A1(n30075), .A2(\xmem_data[82][0] ), .B1(n29439), .B2(
        \xmem_data[83][0] ), .ZN(n30080) );
  AOI22_X1 U32739 ( .A1(n3162), .A2(\xmem_data[80][0] ), .B1(n3190), .B2(
        \xmem_data[81][0] ), .ZN(n30079) );
  AOI22_X1 U32740 ( .A1(n30063), .A2(\xmem_data[84][0] ), .B1(n29487), .B2(
        \xmem_data[85][0] ), .ZN(n30078) );
  AOI22_X1 U32741 ( .A1(n30270), .A2(\xmem_data[86][0] ), .B1(n30269), .B2(
        \xmem_data[87][0] ), .ZN(n30077) );
  NAND4_X1 U32742 ( .A1(n30080), .A2(n30079), .A3(n30078), .A4(n30077), .ZN(
        n30081) );
  AOI22_X1 U32743 ( .A1(n30082), .A2(n30228), .B1(n30081), .B2(n30188), .ZN(
        n30098) );
  AOI22_X1 U32744 ( .A1(n30191), .A2(\xmem_data[72][0] ), .B1(n29646), .B2(
        \xmem_data[73][0] ), .ZN(n30088) );
  AOI22_X1 U32745 ( .A1(n30192), .A2(\xmem_data[74][0] ), .B1(n30083), .B2(
        \xmem_data[75][0] ), .ZN(n30087) );
  AOI22_X1 U32746 ( .A1(n27811), .A2(\xmem_data[76][0] ), .B1(n30090), .B2(
        \xmem_data[77][0] ), .ZN(n30086) );
  AOI22_X1 U32747 ( .A1(n30251), .A2(\xmem_data[78][0] ), .B1(n27455), .B2(
        \xmem_data[79][0] ), .ZN(n30085) );
  NAND4_X1 U32748 ( .A1(n30088), .A2(n30087), .A3(n30086), .A4(n30085), .ZN(
        n30089) );
  NAND2_X1 U32749 ( .A1(n30089), .A2(n30188), .ZN(n30097) );
  AOI22_X1 U32750 ( .A1(n28180), .A2(\xmem_data[104][0] ), .B1(n29704), .B2(
        \xmem_data[105][0] ), .ZN(n30094) );
  AOI22_X1 U32751 ( .A1(n30300), .A2(\xmem_data[106][0] ), .B1(n23792), .B2(
        \xmem_data[107][0] ), .ZN(n30093) );
  AOI22_X1 U32752 ( .A1(n28779), .A2(\xmem_data[108][0] ), .B1(n28684), .B2(
        \xmem_data[109][0] ), .ZN(n30092) );
  AOI22_X1 U32753 ( .A1(n30251), .A2(\xmem_data[110][0] ), .B1(n30303), .B2(
        \xmem_data[111][0] ), .ZN(n30091) );
  NAND4_X1 U32754 ( .A1(n30094), .A2(n30093), .A3(n30092), .A4(n30091), .ZN(
        n30095) );
  NAND2_X1 U32755 ( .A1(n30095), .A2(n30287), .ZN(n30096) );
  NAND4_X1 U32756 ( .A1(n30099), .A2(n30098), .A3(n30097), .A4(n30096), .ZN(
        n30121) );
  AOI22_X1 U32757 ( .A1(n3392), .A2(\xmem_data[34][0] ), .B1(n30278), .B2(
        \xmem_data[35][0] ), .ZN(n30104) );
  AOI22_X1 U32758 ( .A1(n27710), .A2(\xmem_data[32][0] ), .B1(n29432), .B2(
        \xmem_data[33][0] ), .ZN(n30103) );
  AOI22_X1 U32759 ( .A1(n30294), .A2(\xmem_data[36][0] ), .B1(n29495), .B2(
        \xmem_data[37][0] ), .ZN(n30102) );
  AOI22_X1 U32760 ( .A1(n30219), .A2(\xmem_data[38][0] ), .B1(n30295), .B2(
        \xmem_data[39][0] ), .ZN(n30101) );
  NAND4_X1 U32761 ( .A1(n30104), .A2(n30103), .A3(n30102), .A4(n30101), .ZN(
        n30105) );
  AOI22_X1 U32762 ( .A1(n27741), .A2(\xmem_data[96][0] ), .B1(n29672), .B2(
        \xmem_data[97][0] ), .ZN(n30110) );
  AOI22_X1 U32763 ( .A1(n27740), .A2(\xmem_data[98][0] ), .B1(n30292), .B2(
        \xmem_data[99][0] ), .ZN(n30109) );
  AOI22_X1 U32764 ( .A1(n30280), .A2(\xmem_data[100][0] ), .B1(n29495), .B2(
        \xmem_data[101][0] ), .ZN(n30108) );
  AOI22_X1 U32765 ( .A1(n30282), .A2(\xmem_data[102][0] ), .B1(n3137), .B2(
        \xmem_data[103][0] ), .ZN(n30107) );
  NAND4_X1 U32766 ( .A1(n30110), .A2(n30109), .A3(n30108), .A4(n30107), .ZN(
        n30111) );
  AOI22_X1 U32767 ( .A1(n29626), .A2(\xmem_data[64][0] ), .B1(n30222), .B2(
        \xmem_data[65][0] ), .ZN(n30115) );
  AOI22_X1 U32768 ( .A1(n29628), .A2(\xmem_data[66][0] ), .B1(n29627), .B2(
        \xmem_data[67][0] ), .ZN(n30114) );
  AOI22_X1 U32769 ( .A1(n30280), .A2(\xmem_data[68][0] ), .B1(n30217), .B2(
        \xmem_data[69][0] ), .ZN(n30113) );
  AOI22_X1 U32770 ( .A1(n30282), .A2(\xmem_data[70][0] ), .B1(n3138), .B2(
        \xmem_data[71][0] ), .ZN(n30112) );
  NAND4_X1 U32771 ( .A1(n30115), .A2(n30114), .A3(n30113), .A4(n30112), .ZN(
        n30116) );
  NAND3_X1 U32772 ( .A1(n30119), .A2(n30118), .A3(n30117), .ZN(n30120) );
  INV_X1 U32773 ( .A(n35697), .ZN(n30123) );
  OAI21_X1 U32774 ( .B1(n31392), .B2(n31390), .A(n31391), .ZN(n30125) );
  NAND2_X1 U32775 ( .A1(n31392), .A2(n31390), .ZN(n30124) );
  NAND2_X1 U32776 ( .A1(n30125), .A2(n30124), .ZN(n31146) );
  NAND2_X1 U32777 ( .A1(n30126), .A2(n31146), .ZN(n30128) );
  NAND2_X1 U32778 ( .A1(n31143), .A2(n31144), .ZN(n30127) );
  NAND2_X1 U32779 ( .A1(n30128), .A2(n30127), .ZN(n31205) );
  FA_X1 U32780 ( .A(n30131), .B(n30130), .CI(n30129), .CO(n31239), .S(n31624)
         );
  OAI21_X1 U32781 ( .B1(n31414), .B2(n31413), .A(n31412), .ZN(n30132) );
  NAND2_X1 U32782 ( .A1(n30133), .A2(n30132), .ZN(n31767) );
  XNOR2_X1 U32783 ( .A(n30135), .B(n30134), .ZN(n30137) );
  XNOR2_X1 U32784 ( .A(n30137), .B(n30136), .ZN(n31202) );
  NAND2_X1 U32785 ( .A1(n30145), .A2(n30144), .ZN(n30375) );
  FA_X1 U32786 ( .A(n30148), .B(n30147), .CI(n30146), .CO(n30374), .S(n30150)
         );
  NAND2_X1 U32787 ( .A1(n31202), .A2(n31203), .ZN(n30153) );
  FA_X1 U32788 ( .A(n30151), .B(n30149), .CI(n30150), .CO(n31201), .S(n34287)
         );
  OAI21_X1 U32789 ( .B1(n31202), .B2(n31203), .A(n31201), .ZN(n30152) );
  NAND2_X1 U32790 ( .A1(n30152), .A2(n30153), .ZN(n31768) );
  XNOR2_X1 U32791 ( .A(n31767), .B(n31768), .ZN(n30378) );
  FA_X1 U32792 ( .A(n30155), .B(n4012), .CI(n30154), .CO(n31787), .S(n31757)
         );
  XNOR2_X1 U32793 ( .A(n31642), .B(\fmem_data[20][3] ), .ZN(n32518) );
  OAI21_X1 U32794 ( .B1(n32518), .B2(n34495), .A(n30160), .ZN(n30479) );
  XNOR2_X1 U32795 ( .A(n35072), .B(\fmem_data[22][1] ), .ZN(n33948) );
  INV_X1 U32796 ( .A(n34777), .ZN(n30161) );
  NOR2_X1 U32797 ( .A1(n30161), .A2(\fmem_data[22][0] ), .ZN(n30162) );
  OR2_X1 U32798 ( .A1(n33948), .A2(n30162), .ZN(n30478) );
  XNOR2_X1 U32799 ( .A(n35074), .B(\fmem_data[17][1] ), .ZN(n33950) );
  INV_X1 U32800 ( .A(n30163), .ZN(n30480) );
  INV_X1 U32801 ( .A(n30479), .ZN(n30165) );
  INV_X1 U32802 ( .A(n30478), .ZN(n30164) );
  NAND2_X1 U32803 ( .A1(n30165), .A2(n30164), .ZN(n30166) );
  NAND2_X1 U32804 ( .A1(n30480), .A2(n30166), .ZN(n30167) );
  XNOR2_X1 U32805 ( .A(n32442), .B(\fmem_data[1][5] ), .ZN(n32724) );
  OAI22_X1 U32806 ( .A1(n30169), .A2(n34942), .B1(n32724), .B2(n34941), .ZN(
        n30839) );
  AOI22_X1 U32807 ( .A1(n29488), .A2(\xmem_data[84][1] ), .B1(n30266), .B2(
        \xmem_data[85][1] ), .ZN(n30180) );
  AOI22_X1 U32808 ( .A1(n3162), .A2(\xmem_data[80][1] ), .B1(n3187), .B2(
        \xmem_data[81][1] ), .ZN(n30179) );
  AOI22_X1 U32809 ( .A1(n30251), .A2(\xmem_data[78][1] ), .B1(n25607), .B2(
        \xmem_data[79][1] ), .ZN(n30173) );
  AOI22_X1 U32810 ( .A1(n30171), .A2(\xmem_data[74][1] ), .B1(n28233), .B2(
        \xmem_data[75][1] ), .ZN(n30172) );
  NAND2_X1 U32811 ( .A1(n30173), .A2(n30172), .ZN(n30177) );
  AOI22_X1 U32812 ( .A1(n30282), .A2(\xmem_data[70][1] ), .B1(n3138), .B2(
        \xmem_data[71][1] ), .ZN(n30175) );
  AOI22_X1 U32813 ( .A1(n30270), .A2(\xmem_data[86][1] ), .B1(n30269), .B2(
        \xmem_data[87][1] ), .ZN(n30174) );
  NAND2_X1 U32814 ( .A1(n30175), .A2(n30174), .ZN(n30176) );
  NOR2_X1 U32815 ( .A1(n30177), .A2(n30176), .ZN(n30178) );
  NAND3_X1 U32816 ( .A1(n30180), .A2(n30179), .A3(n30178), .ZN(n30187) );
  AOI22_X1 U32817 ( .A1(n28138), .A2(\xmem_data[66][1] ), .B1(n30278), .B2(
        \xmem_data[67][1] ), .ZN(n30181) );
  INV_X1 U32818 ( .A(n30181), .ZN(n30186) );
  AOI22_X1 U32819 ( .A1(n27710), .A2(\xmem_data[64][1] ), .B1(n30106), .B2(
        \xmem_data[65][1] ), .ZN(n30184) );
  AOI22_X1 U32820 ( .A1(n30280), .A2(\xmem_data[68][1] ), .B1(n30696), .B2(
        \xmem_data[69][1] ), .ZN(n30183) );
  NAND2_X1 U32821 ( .A1(n30184), .A2(n30183), .ZN(n30185) );
  NOR3_X1 U32822 ( .A1(n30187), .A2(n30186), .A3(n30185), .ZN(n30189) );
  INV_X1 U32823 ( .A(n30188), .ZN(n30243) );
  NOR2_X1 U32824 ( .A1(n30189), .A2(n30243), .ZN(n30247) );
  AOI22_X1 U32825 ( .A1(n30743), .A2(\xmem_data[8][1] ), .B1(n30730), .B2(
        \xmem_data[9][1] ), .ZN(n30197) );
  AOI22_X1 U32826 ( .A1(n30192), .A2(\xmem_data[10][1] ), .B1(n30943), .B2(
        \xmem_data[11][1] ), .ZN(n30196) );
  AOI22_X1 U32827 ( .A1(n3174), .A2(\xmem_data[12][1] ), .B1(n27753), .B2(
        \xmem_data[13][1] ), .ZN(n30195) );
  AOI22_X1 U32828 ( .A1(n30304), .A2(\xmem_data[14][1] ), .B1(n30892), .B2(
        \xmem_data[15][1] ), .ZN(n30194) );
  NAND4_X1 U32829 ( .A1(n30197), .A2(n30196), .A3(n30195), .A4(n30194), .ZN(
        n30214) );
  AOI22_X1 U32830 ( .A1(n30063), .A2(\xmem_data[20][1] ), .B1(n30685), .B2(
        \xmem_data[21][1] ), .ZN(n30212) );
  AOI22_X1 U32831 ( .A1(n30715), .A2(\xmem_data[18][1] ), .B1(n28147), .B2(
        \xmem_data[19][1] ), .ZN(n30211) );
  AOI22_X1 U32832 ( .A1(n3210), .A2(\xmem_data[24][1] ), .B1(n6247), .B2(
        \xmem_data[25][1] ), .ZN(n30204) );
  AOI22_X1 U32833 ( .A1(n6309), .A2(\xmem_data[26][1] ), .B1(n20567), .B2(
        \xmem_data[27][1] ), .ZN(n30203) );
  AOI22_X1 U32834 ( .A1(n30199), .A2(\xmem_data[28][1] ), .B1(n30259), .B2(
        \xmem_data[29][1] ), .ZN(n30202) );
  AOI22_X1 U32835 ( .A1(n30261), .A2(\xmem_data[30][1] ), .B1(n30864), .B2(
        \xmem_data[31][1] ), .ZN(n30201) );
  NAND4_X1 U32836 ( .A1(n30204), .A2(n30203), .A3(n30202), .A4(n30201), .ZN(
        n30208) );
  AOI22_X1 U32837 ( .A1(n30205), .A2(\xmem_data[22][1] ), .B1(n28202), .B2(
        \xmem_data[23][1] ), .ZN(n30206) );
  INV_X1 U32838 ( .A(n30206), .ZN(n30207) );
  NOR2_X1 U32839 ( .A1(n30208), .A2(n30207), .ZN(n30210) );
  AOI22_X1 U32840 ( .A1(n3163), .A2(\xmem_data[16][1] ), .B1(n3183), .B2(
        \xmem_data[17][1] ), .ZN(n30209) );
  NAND4_X1 U32841 ( .A1(n30212), .A2(n30211), .A3(n30210), .A4(n30209), .ZN(
        n30213) );
  NOR2_X1 U32842 ( .A1(n30213), .A2(n30214), .ZN(n30231) );
  AOI22_X1 U32843 ( .A1(n28700), .A2(\xmem_data[2][1] ), .B1(n30292), .B2(
        \xmem_data[3][1] ), .ZN(n30216) );
  INV_X1 U32844 ( .A(n30216), .ZN(n30227) );
  AOI22_X1 U32845 ( .A1(n30777), .A2(\xmem_data[4][1] ), .B1(n30293), .B2(
        \xmem_data[5][1] ), .ZN(n30221) );
  AOI22_X1 U32846 ( .A1(n30219), .A2(\xmem_data[6][1] ), .B1(n3132), .B2(
        \xmem_data[7][1] ), .ZN(n30220) );
  NAND2_X1 U32847 ( .A1(n30221), .A2(n30220), .ZN(n30226) );
  AOI22_X1 U32848 ( .A1(n29788), .A2(\xmem_data[0][1] ), .B1(n28206), .B2(
        \xmem_data[1][1] ), .ZN(n30224) );
  INV_X1 U32849 ( .A(n30224), .ZN(n30225) );
  NOR3_X1 U32850 ( .A1(n30227), .A2(n30226), .A3(n30225), .ZN(n30230) );
  INV_X1 U32851 ( .A(n30228), .ZN(n30229) );
  AOI21_X1 U32852 ( .B1(n30231), .B2(n30230), .A(n30229), .ZN(n30246) );
  AOI22_X1 U32853 ( .A1(n28146), .A2(\xmem_data[72][1] ), .B1(n27761), .B2(
        \xmem_data[73][1] ), .ZN(n30232) );
  INV_X1 U32854 ( .A(n30232), .ZN(n30242) );
  AOI22_X1 U32855 ( .A1(n3211), .A2(\xmem_data[88][1] ), .B1(n30256), .B2(
        \xmem_data[89][1] ), .ZN(n30236) );
  AOI22_X1 U32856 ( .A1(n30258), .A2(\xmem_data[90][1] ), .B1(n30257), .B2(
        \xmem_data[91][1] ), .ZN(n30235) );
  AOI22_X1 U32857 ( .A1(n30260), .A2(\xmem_data[92][1] ), .B1(n3421), .B2(
        \xmem_data[93][1] ), .ZN(n30234) );
  AOI22_X1 U32858 ( .A1(n30320), .A2(\xmem_data[94][1] ), .B1(n3424), .B2(
        \xmem_data[95][1] ), .ZN(n30233) );
  NAND4_X1 U32859 ( .A1(n30236), .A2(n30235), .A3(n30234), .A4(n30233), .ZN(
        n30241) );
  AOI22_X1 U32860 ( .A1(n30302), .A2(\xmem_data[76][1] ), .B1(n30301), .B2(
        \xmem_data[77][1] ), .ZN(n30239) );
  AOI22_X1 U32861 ( .A1(n30684), .A2(\xmem_data[82][1] ), .B1(n25400), .B2(
        \xmem_data[83][1] ), .ZN(n30238) );
  NAND2_X1 U32862 ( .A1(n30239), .A2(n30238), .ZN(n30240) );
  NOR3_X1 U32863 ( .A1(n30242), .A2(n30241), .A3(n30240), .ZN(n30244) );
  NOR2_X1 U32864 ( .A1(n30244), .A2(n30243), .ZN(n30245) );
  NOR3_X1 U32865 ( .A1(n30247), .A2(n30246), .A3(n30245), .ZN(n30333) );
  AOI22_X1 U32866 ( .A1(n29647), .A2(\xmem_data[104][1] ), .B1(n3369), .B2(
        \xmem_data[105][1] ), .ZN(n30255) );
  AOI22_X1 U32867 ( .A1(n3214), .A2(\xmem_data[106][1] ), .B1(n28152), .B2(
        \xmem_data[107][1] ), .ZN(n30254) );
  AOI22_X1 U32868 ( .A1(n29604), .A2(\xmem_data[108][1] ), .B1(n30193), .B2(
        \xmem_data[109][1] ), .ZN(n30253) );
  AOI22_X1 U32869 ( .A1(n30251), .A2(\xmem_data[110][1] ), .B1(n31354), .B2(
        \xmem_data[111][1] ), .ZN(n30252) );
  AOI22_X1 U32870 ( .A1(n3210), .A2(\xmem_data[120][1] ), .B1(n30256), .B2(
        \xmem_data[121][1] ), .ZN(n30265) );
  AOI22_X1 U32871 ( .A1(n30258), .A2(\xmem_data[122][1] ), .B1(n30257), .B2(
        \xmem_data[123][1] ), .ZN(n30264) );
  AOI22_X1 U32872 ( .A1(n30260), .A2(\xmem_data[124][1] ), .B1(n3421), .B2(
        \xmem_data[125][1] ), .ZN(n30263) );
  AOI22_X1 U32873 ( .A1(n30320), .A2(\xmem_data[126][1] ), .B1(n3433), .B2(
        \xmem_data[127][1] ), .ZN(n30262) );
  NAND4_X1 U32874 ( .A1(n30265), .A2(n30264), .A3(n30263), .A4(n30262), .ZN(
        n30275) );
  AOI22_X1 U32875 ( .A1(n29815), .A2(\xmem_data[116][1] ), .B1(n30170), .B2(
        \xmem_data[117][1] ), .ZN(n30268) );
  AOI22_X1 U32876 ( .A1(n30062), .A2(\xmem_data[114][1] ), .B1(n27855), .B2(
        \xmem_data[115][1] ), .ZN(n30267) );
  NAND2_X1 U32877 ( .A1(n30268), .A2(n30267), .ZN(n30274) );
  AOI22_X1 U32878 ( .A1(n3166), .A2(\xmem_data[112][1] ), .B1(n3186), .B2(
        \xmem_data[113][1] ), .ZN(n30272) );
  AOI22_X1 U32879 ( .A1(n30270), .A2(\xmem_data[118][1] ), .B1(n30269), .B2(
        \xmem_data[119][1] ), .ZN(n30271) );
  NAND2_X1 U32880 ( .A1(n30272), .A2(n30271), .ZN(n30273) );
  NOR3_X1 U32881 ( .A1(n30275), .A2(n30274), .A3(n30273), .ZN(n30276) );
  NAND2_X1 U32882 ( .A1(n30277), .A2(n30276), .ZN(n30289) );
  AOI22_X1 U32883 ( .A1(n27710), .A2(\xmem_data[96][1] ), .B1(n29672), .B2(
        \xmem_data[97][1] ), .ZN(n30286) );
  AOI22_X1 U32884 ( .A1(n28700), .A2(\xmem_data[98][1] ), .B1(n30278), .B2(
        \xmem_data[99][1] ), .ZN(n30285) );
  AOI22_X1 U32885 ( .A1(n30280), .A2(\xmem_data[100][1] ), .B1(n29556), .B2(
        \xmem_data[101][1] ), .ZN(n30284) );
  AOI22_X1 U32886 ( .A1(n30282), .A2(\xmem_data[102][1] ), .B1(n3138), .B2(
        \xmem_data[103][1] ), .ZN(n30283) );
  NAND4_X1 U32887 ( .A1(n30286), .A2(n30285), .A3(n30284), .A4(n30283), .ZN(
        n30288) );
  OAI21_X1 U32888 ( .B1(n30289), .B2(n30288), .A(n30287), .ZN(n30332) );
  AOI22_X1 U32889 ( .A1(n29433), .A2(\xmem_data[32][1] ), .B1(n30290), .B2(
        \xmem_data[33][1] ), .ZN(n30299) );
  AOI22_X1 U32890 ( .A1(n29628), .A2(\xmem_data[34][1] ), .B1(n30292), .B2(
        \xmem_data[35][1] ), .ZN(n30298) );
  AOI22_X1 U32891 ( .A1(n30294), .A2(\xmem_data[36][1] ), .B1(n30776), .B2(
        \xmem_data[37][1] ), .ZN(n30297) );
  AOI22_X1 U32892 ( .A1(n30219), .A2(\xmem_data[38][1] ), .B1(n30295), .B2(
        \xmem_data[39][1] ), .ZN(n30296) );
  NAND4_X1 U32893 ( .A1(n30299), .A2(n30298), .A3(n30297), .A4(n30296), .ZN(
        n30328) );
  AOI22_X1 U32894 ( .A1(n27703), .A2(\xmem_data[40][1] ), .B1(n28665), .B2(
        \xmem_data[41][1] ), .ZN(n30308) );
  AOI22_X1 U32895 ( .A1(n3214), .A2(\xmem_data[42][1] ), .B1(n28051), .B2(
        \xmem_data[43][1] ), .ZN(n30307) );
  AOI22_X1 U32896 ( .A1(n29769), .A2(\xmem_data[44][1] ), .B1(n28110), .B2(
        \xmem_data[45][1] ), .ZN(n30306) );
  AOI22_X1 U32897 ( .A1(n30304), .A2(\xmem_data[46][1] ), .B1(n28053), .B2(
        \xmem_data[47][1] ), .ZN(n30305) );
  NAND4_X1 U32898 ( .A1(n30308), .A2(n30307), .A3(n30306), .A4(n30305), .ZN(
        n30327) );
  AOI22_X1 U32899 ( .A1(n3167), .A2(\xmem_data[48][1] ), .B1(n3186), .B2(
        \xmem_data[49][1] ), .ZN(n30315) );
  AOI22_X1 U32900 ( .A1(n30310), .A2(\xmem_data[50][1] ), .B1(n30309), .B2(
        \xmem_data[51][1] ), .ZN(n30314) );
  AOI22_X1 U32901 ( .A1(n29722), .A2(\xmem_data[52][1] ), .B1(n29640), .B2(
        \xmem_data[53][1] ), .ZN(n30313) );
  AOI22_X1 U32902 ( .A1(n30270), .A2(\xmem_data[54][1] ), .B1(n30311), .B2(
        \xmem_data[55][1] ), .ZN(n30312) );
  NAND4_X1 U32903 ( .A1(n30315), .A2(n30314), .A3(n30313), .A4(n30312), .ZN(
        n30326) );
  AOI22_X1 U32904 ( .A1(n3211), .A2(\xmem_data[56][1] ), .B1(n3193), .B2(
        \xmem_data[57][1] ), .ZN(n30324) );
  AOI22_X1 U32905 ( .A1(n30258), .A2(\xmem_data[58][1] ), .B1(n30674), .B2(
        \xmem_data[59][1] ), .ZN(n30323) );
  AOI22_X1 U32906 ( .A1(n30318), .A2(\xmem_data[60][1] ), .B1(n30317), .B2(
        \xmem_data[61][1] ), .ZN(n30322) );
  AOI22_X1 U32907 ( .A1(n30320), .A2(\xmem_data[62][1] ), .B1(n3153), .B2(
        \xmem_data[63][1] ), .ZN(n30321) );
  NAND4_X1 U32908 ( .A1(n30324), .A2(n30323), .A3(n30322), .A4(n30321), .ZN(
        n30325) );
  NAND2_X1 U32909 ( .A1(n30330), .A2(n30329), .ZN(n30331) );
  XNOR2_X1 U32910 ( .A(n33479), .B(\fmem_data[15][7] ), .ZN(n32108) );
  OAI22_X1 U32911 ( .A1(n32108), .A2(n35696), .B1(n30334), .B2(n35697), .ZN(
        n30838) );
  XNOR2_X1 U32912 ( .A(n32597), .B(\fmem_data[15][5] ), .ZN(n30382) );
  XNOR2_X1 U32913 ( .A(n31513), .B(\fmem_data[15][5] ), .ZN(n34056) );
  OAI22_X1 U32914 ( .A1(n30382), .A2(n34990), .B1(n34989), .B2(n34056), .ZN(
        n30837) );
  OAI21_X1 U32915 ( .B1(n30834), .B2(n30833), .A(n30835), .ZN(n30336) );
  NAND2_X1 U32916 ( .A1(n30834), .A2(n30833), .ZN(n30335) );
  NAND2_X1 U32917 ( .A1(n30336), .A2(n30335), .ZN(n31756) );
  OAI21_X1 U32918 ( .B1(n30339), .B2(n30338), .A(n30337), .ZN(n30341) );
  OAI21_X1 U32919 ( .B1(n31757), .B2(n31756), .A(n31758), .ZN(n30343) );
  NAND2_X1 U32920 ( .A1(n30343), .A2(n30342), .ZN(n31715) );
  FA_X1 U32921 ( .A(n30346), .B(n30345), .CI(n30344), .CO(n31694), .S(n30834)
         );
  INV_X1 U32922 ( .A(n30347), .ZN(n30349) );
  NAND2_X1 U32923 ( .A1(n34503), .A2(n34505), .ZN(n30348) );
  NAND2_X1 U32924 ( .A1(n30349), .A2(n30348), .ZN(n31696) );
  XNOR2_X1 U32925 ( .A(n31694), .B(n31696), .ZN(n30352) );
  XNOR2_X1 U32926 ( .A(n30352), .B(n31695), .ZN(n31929) );
  OR2_X1 U32927 ( .A1(n30354), .A2(n35761), .ZN(n30356) );
  XNOR2_X1 U32928 ( .A(n33573), .B(\fmem_data[28][7] ), .ZN(n31950) );
  OR2_X1 U32929 ( .A1(n31950), .A2(n35760), .ZN(n30355) );
  NAND2_X1 U32930 ( .A1(n30356), .A2(n30355), .ZN(n30405) );
  OAI22_X1 U32931 ( .A1(n30358), .A2(n35497), .B1(n30357), .B2(n35498), .ZN(
        n30404) );
  AOI21_X1 U32932 ( .B1(n30405), .B2(n30404), .A(n30403), .ZN(n30362) );
  NOR2_X1 U32933 ( .A1(n30405), .A2(n30404), .ZN(n30361) );
  NOR2_X1 U32934 ( .A1(n30362), .A2(n30361), .ZN(n31685) );
  AND2_X1 U32935 ( .A1(n34468), .A2(n34470), .ZN(n30363) );
  FA_X1 U32936 ( .A(n30367), .B(n30366), .CI(n30365), .CO(n31868), .S(n31405)
         );
  INV_X1 U32937 ( .A(n31868), .ZN(n30373) );
  XNOR2_X1 U32938 ( .A(n32940), .B(\fmem_data[18][7] ), .ZN(n32008) );
  OAI22_X1 U32939 ( .A1(n32008), .A2(n35704), .B1(n33037), .B2(n35705), .ZN(
        n30989) );
  XNOR2_X1 U32940 ( .A(n32937), .B(\fmem_data[19][7] ), .ZN(n32137) );
  OAI22_X1 U32941 ( .A1(n35656), .A2(n30369), .B1(n32137), .B2(n35655), .ZN(
        n30988) );
  XNOR2_X1 U32942 ( .A(n31664), .B(\fmem_data[22][3] ), .ZN(n32004) );
  OAI22_X1 U32943 ( .A1(n32004), .A2(n34416), .B1(n30370), .B2(n34414), .ZN(
        n30842) );
  XNOR2_X1 U32944 ( .A(n31511), .B(\fmem_data[16][5] ), .ZN(n32006) );
  OAI21_X1 U32945 ( .B1(n30373), .B2(n30372), .A(n30371), .ZN(n31927) );
  XNOR2_X1 U32946 ( .A(n31715), .B(n31716), .ZN(n30377) );
  FA_X1 U32947 ( .A(n30376), .B(n30375), .CI(n30374), .CO(n31714), .S(n31203)
         );
  XNOR2_X1 U32948 ( .A(n30377), .B(n31714), .ZN(n31769) );
  XNOR2_X1 U32949 ( .A(n30378), .B(n31769), .ZN(n31635) );
  XNOR2_X1 U32950 ( .A(n34980), .B(\fmem_data[16][3] ), .ZN(n34037) );
  OAI22_X1 U32951 ( .A1(n30380), .A2(n34501), .B1(n34499), .B2(n34037), .ZN(
        n30453) );
  OR2_X1 U32952 ( .A1(n30382), .A2(n34989), .ZN(n30383) );
  OAI21_X1 U32953 ( .B1(n30384), .B2(n34990), .A(n30383), .ZN(n30808) );
  XNOR2_X1 U32954 ( .A(n33733), .B(\fmem_data[11][7] ), .ZN(n32309) );
  OAI22_X1 U32955 ( .A1(n32309), .A2(n35633), .B1(n30385), .B2(n35634), .ZN(
        n30487) );
  XNOR2_X1 U32956 ( .A(n32554), .B(\fmem_data[26][5] ), .ZN(n32254) );
  OAI22_X1 U32957 ( .A1(n30387), .A2(n35034), .B1(n32254), .B2(n35033), .ZN(
        n30992) );
  OAI21_X1 U32958 ( .B1(n30487), .B2(n30486), .A(n30488), .ZN(n30390) );
  NAND2_X1 U32959 ( .A1(n30487), .A2(n30486), .ZN(n30389) );
  OAI21_X1 U32960 ( .B1(n30809), .B2(n30808), .A(n30811), .ZN(n30391) );
  NAND2_X1 U32961 ( .A1(n30392), .A2(n30391), .ZN(n31752) );
  XNOR2_X1 U32962 ( .A(n32929), .B(\fmem_data[23][7] ), .ZN(n34239) );
  OAI22_X1 U32963 ( .A1(n32141), .A2(n35651), .B1(n34239), .B2(n35652), .ZN(
        n31004) );
  XNOR2_X1 U32964 ( .A(n31672), .B(\fmem_data[18][3] ), .ZN(n33035) );
  OAI22_X1 U32965 ( .A1(n30393), .A2(n33679), .B1(n33681), .B2(n33035), .ZN(
        n30457) );
  OAI22_X1 U32966 ( .A1(n30395), .A2(n35744), .B1(n30394), .B2(n35745), .ZN(
        n30456) );
  INV_X1 U32967 ( .A(n30456), .ZN(n30396) );
  XNOR2_X1 U32968 ( .A(n30457), .B(n30396), .ZN(n31002) );
  INV_X1 U32969 ( .A(n35512), .ZN(n30399) );
  INV_X1 U32970 ( .A(n35508), .ZN(n30400) );
  OAI21_X1 U32971 ( .B1(n31004), .B2(n31002), .A(n31003), .ZN(n30402) );
  NAND2_X1 U32972 ( .A1(n31004), .A2(n31002), .ZN(n30401) );
  XNOR2_X1 U32973 ( .A(n34783), .B(\fmem_data[3][7] ), .ZN(n32652) );
  OAI22_X1 U32974 ( .A1(n30407), .A2(n35638), .B1(n32652), .B2(n35637), .ZN(
        n31009) );
  XNOR2_X1 U32975 ( .A(n33246), .B(\fmem_data[25][5] ), .ZN(n33041) );
  OAI21_X1 U32976 ( .B1(n31009), .B2(n31007), .A(n31006), .ZN(n30410) );
  NAND2_X1 U32977 ( .A1(n31009), .A2(n31007), .ZN(n30409) );
  NAND2_X1 U32978 ( .A1(n30410), .A2(n30409), .ZN(n32350) );
  OAI21_X1 U32979 ( .B1(n32348), .B2(n32347), .A(n32350), .ZN(n30412) );
  NAND2_X1 U32980 ( .A1(n30412), .A2(n30411), .ZN(n31751) );
  XNOR2_X1 U32981 ( .A(n31660), .B(\fmem_data[21][3] ), .ZN(n33158) );
  XNOR2_X1 U32982 ( .A(n33039), .B(\fmem_data[0][3] ), .ZN(n30423) );
  OAI22_X1 U32983 ( .A1(n30416), .A2(n33100), .B1(n30415), .B2(n33098), .ZN(
        n30465) );
  XNOR2_X1 U32984 ( .A(n31452), .B(\fmem_data[10][7] ), .ZN(n33267) );
  OAI22_X1 U32985 ( .A1(n30417), .A2(n35611), .B1(n33267), .B2(n35610), .ZN(
        n31651) );
  XNOR2_X1 U32986 ( .A(n32584), .B(\fmem_data[4][5] ), .ZN(n32318) );
  OAI22_X1 U32987 ( .A1(n30418), .A2(n35011), .B1(n32318), .B2(n35010), .ZN(
        n31650) );
  OAI22_X1 U32988 ( .A1(n30420), .A2(n33105), .B1(n30419), .B2(n33103), .ZN(
        n31649) );
  XNOR2_X1 U32989 ( .A(n31640), .B(n3667), .ZN(n32712) );
  NAND2_X1 U32990 ( .A1(n32712), .A2(n30421), .ZN(n30422) );
  INV_X1 U32991 ( .A(n30824), .ZN(n30427) );
  INV_X1 U32992 ( .A(n30426), .ZN(n30823) );
  NAND2_X1 U32993 ( .A1(n30427), .A2(n30426), .ZN(n30431) );
  NAND2_X1 U32994 ( .A1(n30431), .A2(n30826), .ZN(n30433) );
  NAND2_X1 U32995 ( .A1(n30433), .A2(n30432), .ZN(n30812) );
  INV_X1 U32996 ( .A(n30438), .ZN(n30440) );
  NAND2_X1 U32997 ( .A1(n34462), .A2(n34463), .ZN(n30439) );
  NAND2_X1 U32998 ( .A1(n30440), .A2(n30439), .ZN(n31690) );
  XNOR2_X1 U32999 ( .A(n31691), .B(n31690), .ZN(n30444) );
  NOR2_X1 U33000 ( .A1(n30442), .A2(n30441), .ZN(n30443) );
  XNOR2_X1 U33001 ( .A(n30444), .B(n31689), .ZN(n31726) );
  XNOR2_X1 U33002 ( .A(n31680), .B(n31681), .ZN(n30455) );
  FA_X1 U33003 ( .A(n30454), .B(n30453), .CI(n30452), .CO(n31682), .S(n30809)
         );
  XNOR2_X1 U33004 ( .A(n30455), .B(n31682), .ZN(n31725) );
  OAI22_X1 U33005 ( .A1(n30459), .A2(n35739), .B1(n30458), .B2(n35740), .ZN(
        n30475) );
  OAI21_X1 U33006 ( .B1(n30476), .B2(n30475), .A(n30474), .ZN(n30462) );
  NAND2_X1 U33007 ( .A1(n30462), .A2(n30461), .ZN(n31688) );
  FA_X1 U33008 ( .A(n30467), .B(n30466), .CI(n30465), .CO(n31686), .S(n30814)
         );
  XNOR2_X1 U33009 ( .A(n32039), .B(n32038), .ZN(n30807) );
  XNOR2_X1 U33010 ( .A(n33683), .B(\fmem_data[24][7] ), .ZN(n32666) );
  OAI22_X1 U33011 ( .A1(n32666), .A2(n35489), .B1(n31953), .B2(n35490), .ZN(
        n30484) );
  OAI22_X1 U33012 ( .A1(n32668), .A2(n35708), .B1(n31984), .B2(n35709), .ZN(
        n30482) );
  INV_X1 U33013 ( .A(n30468), .ZN(n30483) );
  OAI21_X1 U33014 ( .B1(n30484), .B2(n30482), .A(n30483), .ZN(n30470) );
  XNOR2_X1 U33015 ( .A(n32586), .B(\fmem_data[12][5] ), .ZN(n32026) );
  OAI22_X1 U33016 ( .A1(n30472), .A2(n33975), .B1(n32026), .B2(n33973), .ZN(
        n31653) );
  XNOR2_X1 U33017 ( .A(n30475), .B(n30474), .ZN(n30477) );
  XNOR2_X1 U33018 ( .A(n30477), .B(n30476), .ZN(n31730) );
  XNOR2_X1 U33019 ( .A(n30479), .B(n30478), .ZN(n30481) );
  XNOR2_X1 U33020 ( .A(n30481), .B(n30480), .ZN(n31875) );
  XNOR2_X1 U33021 ( .A(n30483), .B(n30482), .ZN(n30485) );
  XNOR2_X1 U33022 ( .A(n30485), .B(n30484), .ZN(n31874) );
  XNOR2_X1 U33023 ( .A(n30487), .B(n30486), .ZN(n30489) );
  XNOR2_X1 U33024 ( .A(n30489), .B(n30488), .ZN(n31873) );
  NOR2_X1 U33025 ( .A1(n31860), .A2(n31859), .ZN(n30806) );
  FA_X1 U33026 ( .A(n30492), .B(n30491), .CI(n30490), .CO(n29690), .S(n31160)
         );
  OR2_X1 U33027 ( .A1(n34626), .A2(n3638), .ZN(n30494) );
  OAI22_X1 U33028 ( .A1(n30494), .A2(n35730), .B1(n35729), .B2(n3638), .ZN(
        n30986) );
  AOI22_X1 U33029 ( .A1(n17002), .A2(\xmem_data[32][1] ), .B1(n30495), .B2(
        \xmem_data[33][1] ), .ZN(n30502) );
  AOI22_X1 U33030 ( .A1(n3330), .A2(\xmem_data[34][1] ), .B1(n20781), .B2(
        \xmem_data[35][1] ), .ZN(n30501) );
  AOI22_X1 U33031 ( .A1(n30497), .A2(\xmem_data[36][1] ), .B1(n30496), .B2(
        \xmem_data[37][1] ), .ZN(n30500) );
  AOI22_X1 U33032 ( .A1(n30257), .A2(\xmem_data[38][1] ), .B1(n30498), .B2(
        \xmem_data[39][1] ), .ZN(n30499) );
  NAND4_X1 U33033 ( .A1(n30502), .A2(n30501), .A3(n30500), .A4(n30499), .ZN(
        n30523) );
  AOI22_X1 U33034 ( .A1(n24607), .A2(\xmem_data[40][1] ), .B1(n31346), .B2(
        \xmem_data[41][1] ), .ZN(n30507) );
  AOI22_X1 U33035 ( .A1(n25443), .A2(\xmem_data[42][1] ), .B1(n29286), .B2(
        \xmem_data[43][1] ), .ZN(n30506) );
  AOI22_X1 U33036 ( .A1(n30503), .A2(\xmem_data[44][1] ), .B1(n3218), .B2(
        \xmem_data[45][1] ), .ZN(n30505) );
  AOI22_X1 U33037 ( .A1(n23740), .A2(\xmem_data[46][1] ), .B1(n23739), .B2(
        \xmem_data[47][1] ), .ZN(n30504) );
  NAND4_X1 U33038 ( .A1(n30507), .A2(n30506), .A3(n30505), .A4(n30504), .ZN(
        n30522) );
  AOI22_X1 U33039 ( .A1(n21069), .A2(\xmem_data[48][1] ), .B1(n3256), .B2(
        \xmem_data[49][1] ), .ZN(n30512) );
  AOI22_X1 U33040 ( .A1(n30710), .A2(\xmem_data[50][1] ), .B1(n23771), .B2(
        \xmem_data[51][1] ), .ZN(n30511) );
  AOI22_X1 U33041 ( .A1(n27508), .A2(\xmem_data[52][1] ), .B1(n24158), .B2(
        \xmem_data[53][1] ), .ZN(n30510) );
  AOI22_X1 U33042 ( .A1(n30508), .A2(\xmem_data[54][1] ), .B1(n28515), .B2(
        \xmem_data[55][1] ), .ZN(n30509) );
  NAND4_X1 U33043 ( .A1(n30512), .A2(n30511), .A3(n30510), .A4(n30509), .ZN(
        n30521) );
  AOI22_X1 U33044 ( .A1(n30514), .A2(\xmem_data[56][1] ), .B1(n30513), .B2(
        \xmem_data[57][1] ), .ZN(n30519) );
  AOI22_X1 U33045 ( .A1(n30746), .A2(\xmem_data[58][1] ), .B1(n3208), .B2(
        \xmem_data[59][1] ), .ZN(n30518) );
  AOI22_X1 U33046 ( .A1(n23764), .A2(\xmem_data[60][1] ), .B1(n28492), .B2(
        \xmem_data[61][1] ), .ZN(n30517) );
  AOI22_X1 U33047 ( .A1(n28687), .A2(\xmem_data[62][1] ), .B1(n30515), .B2(
        \xmem_data[63][1] ), .ZN(n30516) );
  NAND4_X1 U33048 ( .A1(n30519), .A2(n30518), .A3(n30517), .A4(n30516), .ZN(
        n30520) );
  OR4_X1 U33049 ( .A1(n30523), .A2(n30522), .A3(n30521), .A4(n30520), .ZN(
        n30566) );
  AOI22_X1 U33050 ( .A1(n31345), .A2(\xmem_data[6][1] ), .B1(n30524), .B2(
        \xmem_data[7][1] ), .ZN(n30532) );
  AOI22_X1 U33051 ( .A1(n3172), .A2(\xmem_data[4][1] ), .B1(n23725), .B2(
        \xmem_data[5][1] ), .ZN(n30526) );
  INV_X1 U33052 ( .A(n30526), .ZN(n30530) );
  AOI22_X1 U33053 ( .A1(n29297), .A2(\xmem_data[2][1] ), .B1(n20781), .B2(
        \xmem_data[3][1] ), .ZN(n30528) );
  NAND2_X1 U33054 ( .A1(n28060), .A2(\xmem_data[1][1] ), .ZN(n30527) );
  NAND2_X1 U33055 ( .A1(n30528), .A2(n30527), .ZN(n30529) );
  NOR2_X1 U33056 ( .A1(n30530), .A2(n30529), .ZN(n30531) );
  NAND2_X1 U33057 ( .A1(n30532), .A2(n30531), .ZN(n30540) );
  AND2_X1 U33058 ( .A1(n3220), .A2(\xmem_data[13][1] ), .ZN(n30533) );
  AOI21_X1 U33059 ( .B1(n28503), .B2(\xmem_data[12][1] ), .A(n30533), .ZN(
        n30538) );
  AOI22_X1 U33060 ( .A1(n3433), .A2(\xmem_data[10][1] ), .B1(n25687), .B2(
        \xmem_data[11][1] ), .ZN(n30537) );
  AOI22_X1 U33061 ( .A1(n28354), .A2(\xmem_data[8][1] ), .B1(n27958), .B2(
        \xmem_data[9][1] ), .ZN(n30536) );
  AOI22_X1 U33062 ( .A1(n20724), .A2(\xmem_data[14][1] ), .B1(n30534), .B2(
        \xmem_data[15][1] ), .ZN(n30535) );
  NAND4_X1 U33063 ( .A1(n30538), .A2(n30537), .A3(n30536), .A4(n30535), .ZN(
        n30539) );
  OR2_X1 U33064 ( .A1(n30540), .A2(n30539), .ZN(n30562) );
  AOI22_X1 U33065 ( .A1(n20541), .A2(\xmem_data[24][1] ), .B1(n30541), .B2(
        \xmem_data[25][1] ), .ZN(n30549) );
  AOI22_X1 U33066 ( .A1(n30948), .A2(\xmem_data[26][1] ), .B1(n30542), .B2(
        \xmem_data[27][1] ), .ZN(n30548) );
  AOI22_X1 U33067 ( .A1(n17020), .A2(\xmem_data[28][1] ), .B1(n30544), .B2(
        \xmem_data[29][1] ), .ZN(n30547) );
  AOI22_X1 U33068 ( .A1(n30950), .A2(\xmem_data[30][1] ), .B1(n30545), .B2(
        \xmem_data[31][1] ), .ZN(n30546) );
  NAND4_X1 U33069 ( .A1(n30549), .A2(n30548), .A3(n30547), .A4(n30546), .ZN(
        n30560) );
  AOI22_X1 U33070 ( .A1(n28475), .A2(\xmem_data[16][1] ), .B1(n30550), .B2(
        \xmem_data[17][1] ), .ZN(n30556) );
  AOI22_X1 U33071 ( .A1(n3280), .A2(\xmem_data[18][1] ), .B1(n29103), .B2(
        \xmem_data[19][1] ), .ZN(n30555) );
  AOI22_X1 U33072 ( .A1(n30551), .A2(\xmem_data[20][1] ), .B1(n30854), .B2(
        \xmem_data[21][1] ), .ZN(n30554) );
  AOI22_X1 U33073 ( .A1(n25708), .A2(\xmem_data[22][1] ), .B1(n30552), .B2(
        \xmem_data[23][1] ), .ZN(n30553) );
  NAND4_X1 U33074 ( .A1(n30556), .A2(n30555), .A3(n30554), .A4(n30553), .ZN(
        n30559) );
  AND2_X1 U33075 ( .A1(n30557), .A2(\xmem_data[0][1] ), .ZN(n30558) );
  OR3_X1 U33076 ( .A1(n30560), .A2(n30559), .A3(n30558), .ZN(n30561) );
  OR2_X1 U33077 ( .A1(n30562), .A2(n30561), .ZN(n30564) );
  AOI22_X1 U33078 ( .A1(n30566), .A2(n30565), .B1(n30564), .B2(n30563), .ZN(
        n30631) );
  AOI22_X1 U33079 ( .A1(n20593), .A2(\xmem_data[64][1] ), .B1(n21051), .B2(
        \xmem_data[65][1] ), .ZN(n30570) );
  AOI22_X1 U33080 ( .A1(n30600), .A2(\xmem_data[66][1] ), .B1(n30599), .B2(
        \xmem_data[67][1] ), .ZN(n30569) );
  AOI22_X1 U33081 ( .A1(n3171), .A2(\xmem_data[68][1] ), .B1(n27526), .B2(
        \xmem_data[69][1] ), .ZN(n30568) );
  AOI22_X1 U33082 ( .A1(n30257), .A2(\xmem_data[70][1] ), .B1(n30601), .B2(
        \xmem_data[71][1] ), .ZN(n30567) );
  NAND4_X1 U33083 ( .A1(n30570), .A2(n30569), .A3(n30568), .A4(n30567), .ZN(
        n30587) );
  AOI22_X1 U33084 ( .A1(n30592), .A2(\xmem_data[76][1] ), .B1(n3217), .B2(
        \xmem_data[77][1] ), .ZN(n30575) );
  AOI22_X1 U33085 ( .A1(n3348), .A2(\xmem_data[74][1] ), .B1(n30589), .B2(
        \xmem_data[75][1] ), .ZN(n30574) );
  AOI22_X1 U33086 ( .A1(n30588), .A2(\xmem_data[72][1] ), .B1(n30571), .B2(
        \xmem_data[73][1] ), .ZN(n30573) );
  AOI22_X1 U33087 ( .A1(n30593), .A2(\xmem_data[78][1] ), .B1(n24207), .B2(
        \xmem_data[79][1] ), .ZN(n30572) );
  NAND4_X1 U33088 ( .A1(n30575), .A2(n30574), .A3(n30573), .A4(n30572), .ZN(
        n30586) );
  AOI22_X1 U33089 ( .A1(n30606), .A2(\xmem_data[80][1] ), .B1(n20806), .B2(
        \xmem_data[81][1] ), .ZN(n30579) );
  AOI22_X1 U33090 ( .A1(n3140), .A2(\xmem_data[82][1] ), .B1(n28045), .B2(
        \xmem_data[83][1] ), .ZN(n30578) );
  AOI22_X1 U33091 ( .A1(n30607), .A2(\xmem_data[84][1] ), .B1(n3358), .B2(
        \xmem_data[85][1] ), .ZN(n30577) );
  AOI22_X1 U33092 ( .A1(n30608), .A2(\xmem_data[86][1] ), .B1(n22702), .B2(
        \xmem_data[87][1] ), .ZN(n30576) );
  NAND4_X1 U33093 ( .A1(n30579), .A2(n30578), .A3(n30577), .A4(n30576), .ZN(
        n30585) );
  AOI22_X1 U33094 ( .A1(n30614), .A2(\xmem_data[88][1] ), .B1(n30613), .B2(
        \xmem_data[89][1] ), .ZN(n30583) );
  AOI22_X1 U33095 ( .A1(n29396), .A2(\xmem_data[90][1] ), .B1(n30615), .B2(
        \xmem_data[91][1] ), .ZN(n30582) );
  AOI22_X1 U33096 ( .A1(n24214), .A2(\xmem_data[92][1] ), .B1(n28058), .B2(
        \xmem_data[93][1] ), .ZN(n30581) );
  AOI22_X1 U33097 ( .A1(n30617), .A2(\xmem_data[94][1] ), .B1(n30616), .B2(
        \xmem_data[95][1] ), .ZN(n30580) );
  NAND4_X1 U33098 ( .A1(n30583), .A2(n30582), .A3(n30581), .A4(n30580), .ZN(
        n30584) );
  OR4_X1 U33099 ( .A1(n30587), .A2(n30586), .A3(n30585), .A4(n30584), .ZN(
        n30629) );
  AOI22_X1 U33100 ( .A1(n30588), .A2(\xmem_data[104][1] ), .B1(n3203), .B2(
        \xmem_data[105][1] ), .ZN(n30597) );
  AOI22_X1 U33101 ( .A1(n3348), .A2(\xmem_data[106][1] ), .B1(n30589), .B2(
        \xmem_data[107][1] ), .ZN(n30596) );
  AND2_X1 U33102 ( .A1(n3222), .A2(\xmem_data[109][1] ), .ZN(n30591) );
  AOI21_X1 U33103 ( .B1(n30592), .B2(\xmem_data[108][1] ), .A(n30591), .ZN(
        n30595) );
  AOI22_X1 U33104 ( .A1(n30593), .A2(\xmem_data[110][1] ), .B1(n30963), .B2(
        \xmem_data[111][1] ), .ZN(n30594) );
  NAND4_X1 U33105 ( .A1(n30597), .A2(n30596), .A3(n30595), .A4(n30594), .ZN(
        n30625) );
  AOI22_X1 U33106 ( .A1(n3177), .A2(\xmem_data[96][1] ), .B1(n25716), .B2(
        \xmem_data[97][1] ), .ZN(n30605) );
  AOI22_X1 U33107 ( .A1(n30600), .A2(\xmem_data[98][1] ), .B1(n30599), .B2(
        \xmem_data[99][1] ), .ZN(n30604) );
  AOI22_X1 U33108 ( .A1(n3171), .A2(\xmem_data[100][1] ), .B1(n27981), .B2(
        \xmem_data[101][1] ), .ZN(n30603) );
  AOI22_X1 U33109 ( .A1(n30674), .A2(\xmem_data[102][1] ), .B1(n30601), .B2(
        \xmem_data[103][1] ), .ZN(n30602) );
  NAND4_X1 U33110 ( .A1(n30605), .A2(n30604), .A3(n30603), .A4(n30602), .ZN(
        n30624) );
  AOI22_X1 U33111 ( .A1(n30606), .A2(\xmem_data[112][1] ), .B1(n27550), .B2(
        \xmem_data[113][1] ), .ZN(n30612) );
  AOI22_X1 U33112 ( .A1(n27905), .A2(\xmem_data[114][1] ), .B1(n25514), .B2(
        \xmem_data[115][1] ), .ZN(n30611) );
  AOI22_X1 U33113 ( .A1(n30607), .A2(\xmem_data[116][1] ), .B1(n20546), .B2(
        \xmem_data[117][1] ), .ZN(n30610) );
  AOI22_X1 U33114 ( .A1(n30608), .A2(\xmem_data[118][1] ), .B1(n22740), .B2(
        \xmem_data[119][1] ), .ZN(n30609) );
  NAND4_X1 U33115 ( .A1(n30612), .A2(n30611), .A3(n30610), .A4(n30609), .ZN(
        n30623) );
  AOI22_X1 U33116 ( .A1(n30614), .A2(\xmem_data[120][1] ), .B1(n30613), .B2(
        \xmem_data[121][1] ), .ZN(n30621) );
  AOI22_X1 U33117 ( .A1(n25461), .A2(\xmem_data[122][1] ), .B1(n30615), .B2(
        \xmem_data[123][1] ), .ZN(n30620) );
  AOI22_X1 U33118 ( .A1(n24214), .A2(\xmem_data[124][1] ), .B1(n31329), .B2(
        \xmem_data[125][1] ), .ZN(n30619) );
  AOI22_X1 U33119 ( .A1(n30617), .A2(\xmem_data[126][1] ), .B1(n30616), .B2(
        \xmem_data[127][1] ), .ZN(n30618) );
  NAND4_X1 U33120 ( .A1(n30621), .A2(n30620), .A3(n30619), .A4(n30618), .ZN(
        n30622) );
  OR4_X1 U33121 ( .A1(n30625), .A2(n30624), .A3(n30623), .A4(n30622), .ZN(
        n30627) );
  AOI22_X1 U33122 ( .A1(n30629), .A2(n30628), .B1(n30627), .B2(n30626), .ZN(
        n30630) );
  XNOR2_X1 U33123 ( .A(n32953), .B(\fmem_data[26][7] ), .ZN(n34034) );
  XNOR2_X1 U33124 ( .A(n36111), .B(\fmem_data[26][7] ), .ZN(n30632) );
  OAI22_X1 U33125 ( .A1(n34034), .A2(n35712), .B1(n30632), .B2(n35711), .ZN(
        n30985) );
  AOI22_X1 U33126 ( .A1(n29590), .A2(\xmem_data[112][0] ), .B1(n29646), .B2(
        \xmem_data[113][0] ), .ZN(n30639) );
  AOI22_X1 U33127 ( .A1(n30664), .A2(\xmem_data[114][0] ), .B1(n30663), .B2(
        \xmem_data[115][0] ), .ZN(n30638) );
  AOI22_X1 U33128 ( .A1(n3174), .A2(\xmem_data[116][0] ), .B1(n30249), .B2(
        \xmem_data[117][0] ), .ZN(n30637) );
  AOI22_X1 U33129 ( .A1(n30667), .A2(\xmem_data[118][0] ), .B1(n28091), .B2(
        \xmem_data[119][0] ), .ZN(n30636) );
  NAND4_X1 U33130 ( .A1(n30639), .A2(n30638), .A3(n30637), .A4(n30636), .ZN(
        n30653) );
  AOI22_X1 U33131 ( .A1(n30673), .A2(\xmem_data[96][0] ), .B1(n30672), .B2(
        \xmem_data[97][0] ), .ZN(n30643) );
  AOI22_X1 U33132 ( .A1(n30675), .A2(\xmem_data[98][0] ), .B1(n30674), .B2(
        \xmem_data[99][0] ), .ZN(n30642) );
  AOI22_X1 U33133 ( .A1(n30677), .A2(\xmem_data[100][0] ), .B1(n30676), .B2(
        \xmem_data[101][0] ), .ZN(n30641) );
  AOI22_X1 U33134 ( .A1(n30678), .A2(\xmem_data[102][0] ), .B1(n3434), .B2(
        \xmem_data[103][0] ), .ZN(n30640) );
  NAND4_X1 U33135 ( .A1(n30643), .A2(n30642), .A3(n30641), .A4(n30640), .ZN(
        n30652) );
  AOI22_X1 U33136 ( .A1(n30764), .A2(\xmem_data[122][0] ), .B1(n28687), .B2(
        \xmem_data[123][0] ), .ZN(n30650) );
  AOI22_X1 U33137 ( .A1(n3166), .A2(\xmem_data[120][0] ), .B1(n3187), .B2(
        \xmem_data[121][0] ), .ZN(n30649) );
  AOI22_X1 U33138 ( .A1(n28173), .A2(\xmem_data[124][0] ), .B1(n29487), .B2(
        \xmem_data[125][0] ), .ZN(n30648) );
  AOI22_X1 U33139 ( .A1(n30646), .A2(\xmem_data[126][0] ), .B1(n30645), .B2(
        \xmem_data[127][0] ), .ZN(n30647) );
  NAND4_X1 U33140 ( .A1(n30650), .A2(n30649), .A3(n30648), .A4(n30647), .ZN(
        n30651) );
  OR3_X1 U33141 ( .A1(n30653), .A2(n30652), .A3(n30651), .ZN(n30661) );
  AOI22_X1 U33142 ( .A1(n29433), .A2(\xmem_data[104][0] ), .B1(n30654), .B2(
        \xmem_data[105][0] ), .ZN(n30658) );
  AOI22_X1 U33143 ( .A1(n30279), .A2(\xmem_data[106][0] ), .B1(n23770), .B2(
        \xmem_data[107][0] ), .ZN(n30657) );
  AOI22_X1 U33144 ( .A1(n30697), .A2(\xmem_data[108][0] ), .B1(n3170), .B2(
        \xmem_data[109][0] ), .ZN(n30656) );
  AOI22_X1 U33145 ( .A1(n30699), .A2(\xmem_data[110][0] ), .B1(n30698), .B2(
        \xmem_data[111][0] ), .ZN(n30655) );
  NAND4_X1 U33146 ( .A1(n30658), .A2(n30657), .A3(n30656), .A4(n30655), .ZN(
        n30660) );
  OAI21_X1 U33147 ( .B1(n30661), .B2(n30660), .A(n30659), .ZN(n30788) );
  AOI22_X1 U33148 ( .A1(n27703), .A2(\xmem_data[80][0] ), .B1(n29347), .B2(
        \xmem_data[81][0] ), .ZN(n30671) );
  AOI22_X1 U33149 ( .A1(n30664), .A2(\xmem_data[82][0] ), .B1(n30663), .B2(
        \xmem_data[83][0] ), .ZN(n30670) );
  AOI22_X1 U33150 ( .A1(n3173), .A2(\xmem_data[84][0] ), .B1(n30193), .B2(
        \xmem_data[85][0] ), .ZN(n30669) );
  AOI22_X1 U33151 ( .A1(n30667), .A2(\xmem_data[86][0] ), .B1(n3465), .B2(
        \xmem_data[87][0] ), .ZN(n30668) );
  NAND4_X1 U33152 ( .A1(n30671), .A2(n30670), .A3(n30669), .A4(n30668), .ZN(
        n30694) );
  AOI22_X1 U33153 ( .A1(n30673), .A2(\xmem_data[64][0] ), .B1(n30672), .B2(
        \xmem_data[65][0] ), .ZN(n30682) );
  AOI22_X1 U33154 ( .A1(n30675), .A2(\xmem_data[66][0] ), .B1(n30674), .B2(
        \xmem_data[67][0] ), .ZN(n30681) );
  AOI22_X1 U33155 ( .A1(n30677), .A2(\xmem_data[68][0] ), .B1(n30676), .B2(
        \xmem_data[69][0] ), .ZN(n30680) );
  AOI22_X1 U33156 ( .A1(n30678), .A2(\xmem_data[70][0] ), .B1(n3153), .B2(
        \xmem_data[71][0] ), .ZN(n30679) );
  NAND4_X1 U33157 ( .A1(n30682), .A2(n30681), .A3(n30680), .A4(n30679), .ZN(
        n30693) );
  AND2_X1 U33158 ( .A1(n25400), .A2(\xmem_data[91][0] ), .ZN(n30683) );
  AOI21_X1 U33159 ( .B1(n30684), .B2(\xmem_data[90][0] ), .A(n30683), .ZN(
        n30691) );
  AOI22_X1 U33160 ( .A1(n3163), .A2(\xmem_data[88][0] ), .B1(n3189), .B2(
        \xmem_data[89][0] ), .ZN(n30690) );
  AOI22_X1 U33161 ( .A1(n28173), .A2(\xmem_data[92][0] ), .B1(n30716), .B2(
        \xmem_data[93][0] ), .ZN(n30689) );
  AOI22_X1 U33162 ( .A1(n30687), .A2(\xmem_data[94][0] ), .B1(n30686), .B2(
        \xmem_data[95][0] ), .ZN(n30688) );
  NAND4_X1 U33163 ( .A1(n30691), .A2(n30690), .A3(n30689), .A4(n30688), .ZN(
        n30692) );
  OR3_X1 U33164 ( .A1(n30694), .A2(n30693), .A3(n30692), .ZN(n30706) );
  AOI22_X1 U33165 ( .A1(n29433), .A2(\xmem_data[72][0] ), .B1(n30106), .B2(
        \xmem_data[73][0] ), .ZN(n30703) );
  AOI22_X1 U33166 ( .A1(n29699), .A2(\xmem_data[74][0] ), .B1(n30593), .B2(
        \xmem_data[75][0] ), .ZN(n30702) );
  AOI22_X1 U33167 ( .A1(n30697), .A2(\xmem_data[76][0] ), .B1(n29798), .B2(
        \xmem_data[77][0] ), .ZN(n30701) );
  AOI22_X1 U33168 ( .A1(n30699), .A2(\xmem_data[78][0] ), .B1(n30698), .B2(
        \xmem_data[79][0] ), .ZN(n30700) );
  NAND4_X1 U33169 ( .A1(n30703), .A2(n30702), .A3(n30701), .A4(n30700), .ZN(
        n30705) );
  OAI21_X1 U33170 ( .B1(n30706), .B2(n30705), .A(n30704), .ZN(n30787) );
  AOI22_X1 U33171 ( .A1(n29433), .A2(\xmem_data[8][0] ), .B1(n30707), .B2(
        \xmem_data[9][0] ), .ZN(n30714) );
  AOI22_X1 U33172 ( .A1(n28138), .A2(\xmem_data[10][0] ), .B1(n30292), .B2(
        \xmem_data[11][0] ), .ZN(n30713) );
  AOI22_X1 U33173 ( .A1(n28219), .A2(\xmem_data[12][0] ), .B1(n29556), .B2(
        \xmem_data[13][0] ), .ZN(n30712) );
  AOI22_X1 U33174 ( .A1(n3224), .A2(\xmem_data[14][0] ), .B1(n30710), .B2(
        \xmem_data[15][0] ), .ZN(n30711) );
  NAND4_X1 U33175 ( .A1(n30714), .A2(n30713), .A3(n30712), .A4(n30711), .ZN(
        n30740) );
  AOI22_X1 U33176 ( .A1(n3168), .A2(\xmem_data[24][0] ), .B1(n3189), .B2(
        \xmem_data[25][0] ), .ZN(n30721) );
  AOI22_X1 U33177 ( .A1(n30715), .A2(\xmem_data[26][0] ), .B1(n29639), .B2(
        \xmem_data[27][0] ), .ZN(n30720) );
  AOI22_X1 U33178 ( .A1(n29488), .A2(\xmem_data[28][0] ), .B1(n29721), .B2(
        \xmem_data[29][0] ), .ZN(n30719) );
  AOI22_X1 U33179 ( .A1(n30767), .A2(\xmem_data[30][0] ), .B1(n29816), .B2(
        \xmem_data[31][0] ), .ZN(n30718) );
  NAND4_X1 U33180 ( .A1(n30721), .A2(n30720), .A3(n30719), .A4(n30718), .ZN(
        n30739) );
  AOI22_X1 U33181 ( .A1(n7041), .A2(\xmem_data[0][0] ), .B1(n7042), .B2(
        \xmem_data[1][0] ), .ZN(n30729) );
  AOI22_X1 U33182 ( .A1(n30722), .A2(\xmem_data[2][0] ), .B1(n28036), .B2(
        \xmem_data[3][0] ), .ZN(n30728) );
  AOI22_X1 U33183 ( .A1(n30724), .A2(\xmem_data[4][0] ), .B1(n30723), .B2(
        \xmem_data[5][0] ), .ZN(n30727) );
  AOI22_X1 U33184 ( .A1(n30725), .A2(\xmem_data[6][0] ), .B1(n3414), .B2(
        \xmem_data[7][0] ), .ZN(n30726) );
  NAND4_X1 U33185 ( .A1(n30729), .A2(n30728), .A3(n30727), .A4(n30726), .ZN(
        n30738) );
  AOI22_X1 U33186 ( .A1(n29481), .A2(\xmem_data[16][0] ), .B1(n29389), .B2(
        \xmem_data[17][0] ), .ZN(n30736) );
  AOI22_X1 U33187 ( .A1(n30731), .A2(\xmem_data[18][0] ), .B1(n20716), .B2(
        \xmem_data[19][0] ), .ZN(n30735) );
  AOI22_X1 U33188 ( .A1(n30665), .A2(\xmem_data[20][0] ), .B1(n30634), .B2(
        \xmem_data[21][0] ), .ZN(n30734) );
  AOI22_X1 U33189 ( .A1(n30732), .A2(\xmem_data[22][0] ), .B1(n21048), .B2(
        \xmem_data[23][0] ), .ZN(n30733) );
  NAND4_X1 U33190 ( .A1(n30736), .A2(n30735), .A3(n30734), .A4(n30733), .ZN(
        n30737) );
  OR4_X1 U33191 ( .A1(n30740), .A2(n30739), .A3(n30738), .A4(n30737), .ZN(
        n30742) );
  NAND2_X1 U33192 ( .A1(n30742), .A2(n30741), .ZN(n30786) );
  AOI22_X1 U33193 ( .A1(n29446), .A2(\xmem_data[48][0] ), .B1(n28238), .B2(
        \xmem_data[49][0] ), .ZN(n30751) );
  AOI22_X1 U33194 ( .A1(n26543), .A2(\xmem_data[50][0] ), .B1(n30744), .B2(
        \xmem_data[51][0] ), .ZN(n30750) );
  AOI22_X1 U33195 ( .A1(n29769), .A2(\xmem_data[52][0] ), .B1(n30084), .B2(
        \xmem_data[53][0] ), .ZN(n30749) );
  AOI22_X1 U33196 ( .A1(n30747), .A2(\xmem_data[54][0] ), .B1(n28053), .B2(
        \xmem_data[55][0] ), .ZN(n30748) );
  NAND4_X1 U33197 ( .A1(n30751), .A2(n30750), .A3(n30749), .A4(n30748), .ZN(
        n30774) );
  AOI22_X1 U33198 ( .A1(n30753), .A2(\xmem_data[32][0] ), .B1(n30752), .B2(
        \xmem_data[33][0] ), .ZN(n30763) );
  AOI22_X1 U33199 ( .A1(n30755), .A2(\xmem_data[34][0] ), .B1(n30754), .B2(
        \xmem_data[35][0] ), .ZN(n30762) );
  AOI22_X1 U33200 ( .A1(n30757), .A2(\xmem_data[36][0] ), .B1(n30756), .B2(
        \xmem_data[37][0] ), .ZN(n30761) );
  AOI22_X1 U33201 ( .A1(n30759), .A2(\xmem_data[38][0] ), .B1(n3144), .B2(
        \xmem_data[39][0] ), .ZN(n30760) );
  NAND4_X1 U33202 ( .A1(n30763), .A2(n30762), .A3(n30761), .A4(n30760), .ZN(
        n30773) );
  AOI22_X1 U33203 ( .A1(n3163), .A2(\xmem_data[56][0] ), .B1(n3187), .B2(
        \xmem_data[57][0] ), .ZN(n30771) );
  AOI22_X1 U33204 ( .A1(n30764), .A2(\xmem_data[58][0] ), .B1(n24115), .B2(
        \xmem_data[59][0] ), .ZN(n30770) );
  AOI22_X1 U33205 ( .A1(n29363), .A2(\xmem_data[60][0] ), .B1(n29640), .B2(
        \xmem_data[61][0] ), .ZN(n30769) );
  AOI22_X1 U33206 ( .A1(n30767), .A2(\xmem_data[62][0] ), .B1(n29573), .B2(
        \xmem_data[63][0] ), .ZN(n30768) );
  NAND4_X1 U33207 ( .A1(n30771), .A2(n30770), .A3(n30769), .A4(n30768), .ZN(
        n30772) );
  OR3_X1 U33208 ( .A1(n30774), .A2(n30773), .A3(n30772), .ZN(n30784) );
  AOI22_X1 U33209 ( .A1(n28136), .A2(\xmem_data[40][0] ), .B1(n30707), .B2(
        \xmem_data[41][0] ), .ZN(n30781) );
  AOI22_X1 U33210 ( .A1(n29423), .A2(\xmem_data[42][0] ), .B1(n30964), .B2(
        \xmem_data[43][0] ), .ZN(n30780) );
  AOI22_X1 U33211 ( .A1(n30777), .A2(\xmem_data[44][0] ), .B1(n29708), .B2(
        \xmem_data[45][0] ), .ZN(n30779) );
  AOI22_X1 U33212 ( .A1(n3224), .A2(\xmem_data[46][0] ), .B1(n27905), .B2(
        \xmem_data[47][0] ), .ZN(n30778) );
  NAND4_X1 U33213 ( .A1(n30781), .A2(n30780), .A3(n30779), .A4(n30778), .ZN(
        n30783) );
  OAI21_X1 U33214 ( .B1(n30784), .B2(n30783), .A(n30782), .ZN(n30785) );
  INV_X1 U33215 ( .A(n35652), .ZN(n30789) );
  AND2_X1 U33216 ( .A1(n3116), .A2(n30789), .ZN(n31191) );
  XNOR2_X1 U33217 ( .A(n31800), .B(\fmem_data[29][1] ), .ZN(n32731) );
  OR2_X1 U33218 ( .A1(n32731), .A2(n3575), .ZN(n30790) );
  OAI21_X1 U33219 ( .B1(n32243), .B2(n36120), .A(n30790), .ZN(n31190) );
  NAND2_X1 U33220 ( .A1(n31191), .A2(n31190), .ZN(n30793) );
  XNOR2_X1 U33221 ( .A(n32321), .B(\fmem_data[17][3] ), .ZN(n32134) );
  OAI21_X1 U33222 ( .B1(n31190), .B2(n31191), .A(n31192), .ZN(n30792) );
  NAND2_X1 U33223 ( .A1(n30793), .A2(n30792), .ZN(n31158) );
  FA_X1 U33224 ( .A(n30798), .B(n30797), .CI(n30796), .CO(n30802), .S(n31890)
         );
  INV_X1 U33225 ( .A(n35634), .ZN(n30799) );
  AND2_X1 U33226 ( .A1(n36313), .A2(n30799), .ZN(n31909) );
  XNOR2_X1 U33227 ( .A(n31512), .B(\fmem_data[17][5] ), .ZN(n34044) );
  OAI22_X1 U33228 ( .A1(n32531), .A2(n34043), .B1(n34044), .B2(n34045), .ZN(
        n31908) );
  FA_X1 U33229 ( .A(n30803), .B(n30802), .CI(n30801), .CO(n30148), .S(n31181)
         );
  INV_X1 U33230 ( .A(n31861), .ZN(n30805) );
  NAND2_X1 U33231 ( .A1(n31860), .A2(n31859), .ZN(n30804) );
  OAI21_X1 U33232 ( .B1(n30806), .B2(n30805), .A(n30804), .ZN(n32037) );
  XNOR2_X1 U33233 ( .A(n30807), .B(n32037), .ZN(n32461) );
  XNOR2_X1 U33234 ( .A(n30811), .B(n30810), .ZN(n31762) );
  FA_X1 U33235 ( .A(n30814), .B(n30813), .CI(n30812), .CO(n31750), .S(n31761)
         );
  OAI22_X1 U33236 ( .A1(n32539), .A2(n35181), .B1(n30815), .B2(n35182), .ZN(
        n31118) );
  XNOR2_X1 U33237 ( .A(n31662), .B(\fmem_data[12][1] ), .ZN(n32587) );
  INV_X1 U33238 ( .A(n31878), .ZN(n30822) );
  XNOR2_X1 U33239 ( .A(n35316), .B(\fmem_data[15][1] ), .ZN(n33929) );
  XNOR2_X1 U33240 ( .A(n35030), .B(\fmem_data[15][1] ), .ZN(n32212) );
  NOR2_X1 U33241 ( .A1(n31877), .A2(n31876), .ZN(n30821) );
  NAND2_X1 U33242 ( .A1(n31876), .A2(n31877), .ZN(n30820) );
  OAI21_X1 U33243 ( .B1(n30822), .B2(n30821), .A(n30820), .ZN(n31001) );
  XNOR2_X1 U33244 ( .A(n30824), .B(n30823), .ZN(n30825) );
  INV_X1 U33245 ( .A(n30827), .ZN(n31738) );
  INV_X1 U33246 ( .A(n30828), .ZN(n30830) );
  NAND2_X1 U33247 ( .A1(n34734), .A2(n3572), .ZN(n30829) );
  NAND2_X1 U33248 ( .A1(n30830), .A2(n30829), .ZN(n31737) );
  XNOR2_X1 U33249 ( .A(n34334), .B(\fmem_data[27][7] ), .ZN(n32289) );
  OAI22_X1 U33250 ( .A1(n32289), .A2(n35641), .B1(n30831), .B2(n35642), .ZN(
        n31736) );
  XNOR2_X1 U33251 ( .A(n30834), .B(n30833), .ZN(n30836) );
  FA_X1 U33252 ( .A(n30839), .B(n30838), .CI(n30837), .CO(n30835), .S(n31180)
         );
  FA_X1 U33253 ( .A(n30842), .B(n30841), .CI(n30840), .CO(n31866), .S(n31179)
         );
  FA_X1 U33254 ( .A(n30845), .B(n30843), .CI(n30844), .CO(n30366), .S(n31149)
         );
  XNOR2_X1 U33255 ( .A(n30846), .B(\fmem_data[13][3] ), .ZN(n32542) );
  OAI22_X1 U33256 ( .A1(n32542), .A2(n33570), .B1(n30847), .B2(n33568), .ZN(
        n31139) );
  AOI22_X1 U33257 ( .A1(n31327), .A2(\xmem_data[6][0] ), .B1(n25423), .B2(
        \xmem_data[7][0] ), .ZN(n30848) );
  AOI22_X1 U33258 ( .A1(n30849), .A2(\xmem_data[16][0] ), .B1(n30598), .B2(
        \xmem_data[17][0] ), .ZN(n30853) );
  AOI22_X1 U33259 ( .A1(n20950), .A2(\xmem_data[18][0] ), .B1(n14975), .B2(
        \xmem_data[19][0] ), .ZN(n30852) );
  AOI22_X1 U33260 ( .A1(n24166), .A2(\xmem_data[20][0] ), .B1(n29017), .B2(
        \xmem_data[21][0] ), .ZN(n30851) );
  AOI22_X1 U33261 ( .A1(n29298), .A2(\xmem_data[22][0] ), .B1(n28035), .B2(
        \xmem_data[23][0] ), .ZN(n30850) );
  NAND4_X1 U33262 ( .A1(n30853), .A2(n30852), .A3(n30851), .A4(n30850), .ZN(
        n30859) );
  AOI22_X1 U33263 ( .A1(n24438), .A2(\xmem_data[0][0] ), .B1(n27903), .B2(
        \xmem_data[1][0] ), .ZN(n30857) );
  AOI22_X1 U33264 ( .A1(n23813), .A2(\xmem_data[4][0] ), .B1(n30854), .B2(
        \xmem_data[5][0] ), .ZN(n30856) );
  NAND2_X1 U33265 ( .A1(n20808), .A2(\xmem_data[2][0] ), .ZN(n30855) );
  NAND3_X1 U33266 ( .A1(n30857), .A2(n30856), .A3(n30855), .ZN(n30858) );
  OR3_X1 U33267 ( .A1(n30860), .A2(n30859), .A3(n30858), .ZN(n30870) );
  AOI22_X1 U33268 ( .A1(n30862), .A2(\xmem_data[24][0] ), .B1(n30861), .B2(
        \xmem_data[25][0] ), .ZN(n30868) );
  AOI22_X1 U33269 ( .A1(n30864), .A2(\xmem_data[26][0] ), .B1(n30863), .B2(
        \xmem_data[27][0] ), .ZN(n30867) );
  AOI22_X1 U33270 ( .A1(n21066), .A2(\xmem_data[28][0] ), .B1(n3218), .B2(
        \xmem_data[29][0] ), .ZN(n30866) );
  AOI22_X1 U33271 ( .A1(n25612), .A2(\xmem_data[30][0] ), .B1(n28319), .B2(
        \xmem_data[31][0] ), .ZN(n30865) );
  NAND4_X1 U33272 ( .A1(n30868), .A2(n30867), .A3(n30866), .A4(n30865), .ZN(
        n30869) );
  NOR2_X1 U33273 ( .A1(n30870), .A2(n30869), .ZN(n30881) );
  AOI22_X1 U33274 ( .A1(n30514), .A2(\xmem_data[8][0] ), .B1(n20544), .B2(
        \xmem_data[9][0] ), .ZN(n30876) );
  AOI22_X1 U33275 ( .A1(n30666), .A2(\xmem_data[10][0] ), .B1(n27516), .B2(
        \xmem_data[11][0] ), .ZN(n30875) );
  AOI22_X1 U33276 ( .A1(n24593), .A2(\xmem_data[12][0] ), .B1(n14970), .B2(
        \xmem_data[13][0] ), .ZN(n30874) );
  AOI22_X1 U33277 ( .A1(n30872), .A2(\xmem_data[14][0] ), .B1(n30871), .B2(
        \xmem_data[15][0] ), .ZN(n30873) );
  NAND4_X1 U33278 ( .A1(n30876), .A2(n30875), .A3(n30874), .A4(n30873), .ZN(
        n30878) );
  NOR2_X1 U33279 ( .A1(n30878), .A2(n3736), .ZN(n30880) );
  AOI21_X1 U33280 ( .B1(n30881), .B2(n30880), .A(n30879), .ZN(n30921) );
  AOI22_X1 U33281 ( .A1(n30883), .A2(\xmem_data[32][0] ), .B1(n30882), .B2(
        \xmem_data[33][0] ), .ZN(n30890) );
  AOI22_X1 U33282 ( .A1(n3281), .A2(\xmem_data[34][0] ), .B1(n28007), .B2(
        \xmem_data[35][0] ), .ZN(n30889) );
  AOI22_X1 U33283 ( .A1(n30885), .A2(\xmem_data[36][0] ), .B1(n30884), .B2(
        \xmem_data[37][0] ), .ZN(n30888) );
  AOI22_X1 U33284 ( .A1(n30886), .A2(\xmem_data[38][0] ), .B1(n20958), .B2(
        \xmem_data[39][0] ), .ZN(n30887) );
  NAND4_X1 U33285 ( .A1(n30890), .A2(n30889), .A3(n30888), .A4(n30887), .ZN(
        n30917) );
  AOI22_X1 U33286 ( .A1(n25710), .A2(\xmem_data[40][0] ), .B1(n20584), .B2(
        \xmem_data[41][0] ), .ZN(n30897) );
  AOI22_X1 U33287 ( .A1(n27755), .A2(\xmem_data[42][0] ), .B1(n24457), .B2(
        \xmem_data[43][0] ), .ZN(n30896) );
  AOI22_X1 U33288 ( .A1(n25635), .A2(\xmem_data[44][0] ), .B1(n31270), .B2(
        \xmem_data[45][0] ), .ZN(n30895) );
  AOI22_X1 U33289 ( .A1(n30893), .A2(\xmem_data[46][0] ), .B1(n27523), .B2(
        \xmem_data[47][0] ), .ZN(n30894) );
  NAND4_X1 U33290 ( .A1(n30897), .A2(n30896), .A3(n30895), .A4(n30894), .ZN(
        n30916) );
  AOI22_X1 U33291 ( .A1(n3325), .A2(\xmem_data[48][0] ), .B1(n30898), .B2(
        \xmem_data[49][0] ), .ZN(n30905) );
  AOI22_X1 U33292 ( .A1(n3301), .A2(\xmem_data[50][0] ), .B1(n28495), .B2(
        \xmem_data[51][0] ), .ZN(n30904) );
  AOI22_X1 U33293 ( .A1(n25582), .A2(\xmem_data[52][0] ), .B1(n28500), .B2(
        \xmem_data[53][0] ), .ZN(n30903) );
  AOI22_X1 U33294 ( .A1(n30901), .A2(\xmem_data[54][0] ), .B1(n30900), .B2(
        \xmem_data[55][0] ), .ZN(n30902) );
  NAND4_X1 U33295 ( .A1(n30905), .A2(n30904), .A3(n30903), .A4(n30902), .ZN(
        n30915) );
  AOI22_X1 U33296 ( .A1(n30906), .A2(\xmem_data[60][0] ), .B1(n3221), .B2(
        \xmem_data[61][0] ), .ZN(n30913) );
  AOI22_X1 U33297 ( .A1(n3352), .A2(\xmem_data[58][0] ), .B1(n25485), .B2(
        \xmem_data[59][0] ), .ZN(n30912) );
  AOI22_X1 U33298 ( .A1(n30909), .A2(\xmem_data[56][0] ), .B1(n30908), .B2(
        \xmem_data[57][0] ), .ZN(n30911) );
  AOI22_X1 U33299 ( .A1(n28367), .A2(\xmem_data[62][0] ), .B1(n29255), .B2(
        \xmem_data[63][0] ), .ZN(n30910) );
  NAND4_X1 U33300 ( .A1(n30913), .A2(n30912), .A3(n30911), .A4(n30910), .ZN(
        n30914) );
  OR4_X1 U33301 ( .A1(n30917), .A2(n30916), .A3(n30915), .A4(n30914), .ZN(
        n30919) );
  AND2_X1 U33302 ( .A1(n30919), .A2(n30918), .ZN(n30920) );
  NOR2_X1 U33303 ( .A1(n30921), .A2(n30920), .ZN(n30978) );
  AOI22_X1 U33304 ( .A1(n24438), .A2(\xmem_data[96][0] ), .B1(n22711), .B2(
        \xmem_data[97][0] ), .ZN(n30925) );
  AOI22_X1 U33305 ( .A1(n3128), .A2(\xmem_data[98][0] ), .B1(n28045), .B2(
        \xmem_data[99][0] ), .ZN(n30924) );
  AOI22_X1 U33306 ( .A1(n27551), .A2(\xmem_data[100][0] ), .B1(n27988), .B2(
        \xmem_data[101][0] ), .ZN(n30923) );
  AOI22_X1 U33307 ( .A1(n30943), .A2(\xmem_data[102][0] ), .B1(n13168), .B2(
        \xmem_data[103][0] ), .ZN(n30922) );
  NAND4_X1 U33308 ( .A1(n30925), .A2(n30924), .A3(n30923), .A4(n30922), .ZN(
        n30941) );
  AOI22_X1 U33309 ( .A1(n3176), .A2(\xmem_data[104][0] ), .B1(n28517), .B2(
        \xmem_data[105][0] ), .ZN(n30929) );
  AOI22_X1 U33310 ( .A1(n3465), .A2(\xmem_data[106][0] ), .B1(n27989), .B2(
        \xmem_data[107][0] ), .ZN(n30928) );
  AOI22_X1 U33311 ( .A1(n30949), .A2(\xmem_data[108][0] ), .B1(n31355), .B2(
        \xmem_data[109][0] ), .ZN(n30927) );
  AOI22_X1 U33312 ( .A1(n30950), .A2(\xmem_data[110][0] ), .B1(n24709), .B2(
        \xmem_data[111][0] ), .ZN(n30926) );
  NAND4_X1 U33313 ( .A1(n30929), .A2(n30928), .A3(n30927), .A4(n30926), .ZN(
        n30940) );
  AOI22_X1 U33314 ( .A1(n30956), .A2(\xmem_data[112][0] ), .B1(n30955), .B2(
        \xmem_data[113][0] ), .ZN(n30933) );
  AOI22_X1 U33315 ( .A1(n3308), .A2(\xmem_data[114][0] ), .B1(n20507), .B2(
        \xmem_data[115][0] ), .ZN(n30932) );
  AOI22_X1 U33316 ( .A1(n3179), .A2(\xmem_data[116][0] ), .B1(n28500), .B2(
        \xmem_data[117][0] ), .ZN(n30931) );
  AOI22_X1 U33317 ( .A1(n27498), .A2(\xmem_data[118][0] ), .B1(n24524), .B2(
        \xmem_data[119][0] ), .ZN(n30930) );
  NAND4_X1 U33318 ( .A1(n30933), .A2(n30932), .A3(n30931), .A4(n30930), .ZN(
        n30939) );
  AOI22_X1 U33319 ( .A1(n20953), .A2(\xmem_data[120][0] ), .B1(n28317), .B2(
        \xmem_data[121][0] ), .ZN(n30937) );
  AOI22_X1 U33320 ( .A1(n3333), .A2(\xmem_data[122][0] ), .B1(n24172), .B2(
        \xmem_data[123][0] ), .ZN(n30936) );
  AOI22_X1 U33321 ( .A1(n30962), .A2(\xmem_data[124][0] ), .B1(n3220), .B2(
        \xmem_data[125][0] ), .ZN(n30935) );
  AOI22_X1 U33322 ( .A1(n30964), .A2(\xmem_data[126][0] ), .B1(n30963), .B2(
        \xmem_data[127][0] ), .ZN(n30934) );
  NAND4_X1 U33323 ( .A1(n30937), .A2(n30936), .A3(n30935), .A4(n30934), .ZN(
        n30938) );
  OR4_X1 U33324 ( .A1(n30941), .A2(n30940), .A3(n30939), .A4(n30938), .ZN(
        n30975) );
  AOI22_X1 U33325 ( .A1(n25416), .A2(\xmem_data[64][0] ), .B1(n13444), .B2(
        \xmem_data[65][0] ), .ZN(n30947) );
  AOI22_X1 U33326 ( .A1(n3129), .A2(\xmem_data[66][0] ), .B1(n29103), .B2(
        \xmem_data[67][0] ), .ZN(n30946) );
  AOI22_X1 U33327 ( .A1(n27551), .A2(\xmem_data[68][0] ), .B1(n27943), .B2(
        \xmem_data[69][0] ), .ZN(n30945) );
  AOI22_X1 U33328 ( .A1(n30943), .A2(\xmem_data[70][0] ), .B1(n13168), .B2(
        \xmem_data[71][0] ), .ZN(n30944) );
  NAND4_X1 U33329 ( .A1(n30947), .A2(n30946), .A3(n30945), .A4(n30944), .ZN(
        n30972) );
  AOI22_X1 U33330 ( .A1(n23763), .A2(\xmem_data[72][0] ), .B1(n20798), .B2(
        \xmem_data[73][0] ), .ZN(n30954) );
  AOI22_X1 U33331 ( .A1(n29807), .A2(\xmem_data[74][0] ), .B1(n13188), .B2(
        \xmem_data[75][0] ), .ZN(n30953) );
  AOI22_X1 U33332 ( .A1(n30949), .A2(\xmem_data[76][0] ), .B1(n17043), .B2(
        \xmem_data[77][0] ), .ZN(n30952) );
  AOI22_X1 U33333 ( .A1(n30950), .A2(\xmem_data[78][0] ), .B1(n24592), .B2(
        \xmem_data[79][0] ), .ZN(n30951) );
  NAND4_X1 U33334 ( .A1(n30954), .A2(n30953), .A3(n30952), .A4(n30951), .ZN(
        n30971) );
  AOI22_X1 U33335 ( .A1(n30956), .A2(\xmem_data[80][0] ), .B1(n30955), .B2(
        \xmem_data[81][0] ), .ZN(n30960) );
  AOI22_X1 U33336 ( .A1(n29379), .A2(\xmem_data[82][0] ), .B1(n27975), .B2(
        \xmem_data[83][0] ), .ZN(n30959) );
  AOI22_X1 U33337 ( .A1(n22684), .A2(\xmem_data[84][0] ), .B1(n27526), .B2(
        \xmem_data[85][0] ), .ZN(n30958) );
  AOI22_X1 U33338 ( .A1(n14982), .A2(\xmem_data[86][0] ), .B1(n20769), .B2(
        \xmem_data[87][0] ), .ZN(n30957) );
  NAND4_X1 U33339 ( .A1(n30960), .A2(n30959), .A3(n30958), .A4(n30957), .ZN(
        n30970) );
  AOI22_X1 U33340 ( .A1(n3380), .A2(\xmem_data[88][0] ), .B1(n25357), .B2(
        \xmem_data[89][0] ), .ZN(n30968) );
  AOI22_X1 U33341 ( .A1(n3333), .A2(\xmem_data[90][0] ), .B1(n3247), .B2(
        \xmem_data[91][0] ), .ZN(n30967) );
  AOI22_X1 U33342 ( .A1(n30962), .A2(\xmem_data[92][0] ), .B1(n3219), .B2(
        \xmem_data[93][0] ), .ZN(n30966) );
  AOI22_X1 U33343 ( .A1(n30964), .A2(\xmem_data[94][0] ), .B1(n30963), .B2(
        \xmem_data[95][0] ), .ZN(n30965) );
  NAND4_X1 U33344 ( .A1(n30968), .A2(n30967), .A3(n30966), .A4(n30965), .ZN(
        n30969) );
  OR4_X1 U33345 ( .A1(n30972), .A2(n30971), .A3(n30970), .A4(n30969), .ZN(
        n30973) );
  AOI22_X1 U33346 ( .A1(n30976), .A2(n30975), .B1(n30974), .B2(n30973), .ZN(
        n30977) );
  INV_X1 U33347 ( .A(n35611), .ZN(n30979) );
  XNOR2_X1 U33348 ( .A(n3359), .B(\fmem_data[2][1] ), .ZN(n32527) );
  XNOR2_X1 U33349 ( .A(n31705), .B(\fmem_data[17][1] ), .ZN(n33949) );
  OAI22_X1 U33350 ( .A1(n32544), .A2(n34529), .B1(n33949), .B2(n3566), .ZN(
        n31119) );
  XNOR2_X1 U33351 ( .A(n31638), .B(\fmem_data[24][3] ), .ZN(n32717) );
  XNOR2_X1 U33352 ( .A(n3454), .B(\fmem_data[19][3] ), .ZN(n32728) );
  OAI22_X1 U33353 ( .A1(n30984), .A2(n34472), .B1(n32728), .B2(n34474), .ZN(
        n31742) );
  FA_X1 U33354 ( .A(n30987), .B(n30986), .CI(n30985), .CO(n31741), .S(n31159)
         );
  FA_X1 U33355 ( .A(n30990), .B(n30989), .CI(n30988), .CO(n31867), .S(n31153)
         );
  FA_X1 U33356 ( .A(n30993), .B(n30992), .CI(n30991), .CO(n30488), .S(n31157)
         );
  FA_X1 U33357 ( .A(n30996), .B(n30995), .CI(n30994), .CO(n31003), .S(n31156)
         );
  FA_X1 U33358 ( .A(n31001), .B(n31000), .CI(n30999), .CO(n31760), .S(n32100)
         );
  XNOR2_X1 U33359 ( .A(n31003), .B(n31002), .ZN(n31005) );
  XNOR2_X1 U33360 ( .A(n31005), .B(n31004), .ZN(n31872) );
  FA_X1 U33361 ( .A(n31012), .B(n31011), .CI(n31010), .CO(n29525), .S(n31115)
         );
  XNOR2_X1 U33362 ( .A(n32064), .B(\fmem_data[0][3] ), .ZN(n32536) );
  XNOR2_X1 U33363 ( .A(n31125), .B(\fmem_data[0][3] ), .ZN(n32714) );
  AOI22_X1 U33364 ( .A1(n31255), .A2(\xmem_data[16][1] ), .B1(n31254), .B2(
        \xmem_data[17][1] ), .ZN(n31018) );
  AOI22_X1 U33365 ( .A1(n3206), .A2(\xmem_data[18][1] ), .B1(n25581), .B2(
        \xmem_data[19][1] ), .ZN(n31017) );
  AOI22_X1 U33366 ( .A1(n3338), .A2(\xmem_data[20][1] ), .B1(n24167), .B2(
        \xmem_data[21][1] ), .ZN(n31016) );
  AOI22_X1 U33367 ( .A1(n29151), .A2(\xmem_data[22][1] ), .B1(n31256), .B2(
        \xmem_data[23][1] ), .ZN(n31015) );
  NAND4_X1 U33368 ( .A1(n31018), .A2(n31017), .A3(n31016), .A4(n31015), .ZN(
        n31021) );
  AOI22_X1 U33369 ( .A1(n21308), .A2(\xmem_data[28][1] ), .B1(n27437), .B2(
        \xmem_data[29][1] ), .ZN(n31019) );
  AOI22_X1 U33370 ( .A1(n31348), .A2(\xmem_data[30][1] ), .B1(n3220), .B2(
        \xmem_data[31][1] ), .ZN(n31024) );
  AOI22_X1 U33371 ( .A1(n3380), .A2(\xmem_data[26][1] ), .B1(n31262), .B2(
        \xmem_data[27][1] ), .ZN(n31023) );
  AOI22_X1 U33372 ( .A1(n30257), .A2(\xmem_data[24][1] ), .B1(n31261), .B2(
        \xmem_data[25][1] ), .ZN(n31022) );
  AOI22_X1 U33373 ( .A1(n28367), .A2(\xmem_data[0][1] ), .B1(n20500), .B2(
        \xmem_data[1][1] ), .ZN(n31026) );
  AOI22_X1 U33374 ( .A1(n31276), .A2(\xmem_data[6][1] ), .B1(n28415), .B2(
        \xmem_data[7][1] ), .ZN(n31028) );
  NAND2_X1 U33375 ( .A1(n29762), .A2(\xmem_data[4][1] ), .ZN(n31027) );
  NAND2_X1 U33376 ( .A1(n31028), .A2(n31027), .ZN(n31031) );
  AOI22_X1 U33377 ( .A1(n20994), .A2(\xmem_data[2][1] ), .B1(n31275), .B2(
        \xmem_data[3][1] ), .ZN(n31029) );
  INV_X1 U33378 ( .A(n31029), .ZN(n31030) );
  OR3_X1 U33379 ( .A1(n31032), .A2(n31031), .A3(n31030), .ZN(n31038) );
  AOI22_X1 U33380 ( .A1(n27453), .A2(\xmem_data[8][1] ), .B1(n24448), .B2(
        \xmem_data[9][1] ), .ZN(n31036) );
  AOI22_X1 U33381 ( .A1(n31268), .A2(\xmem_data[10][1] ), .B1(n25709), .B2(
        \xmem_data[11][1] ), .ZN(n31035) );
  AOI22_X1 U33382 ( .A1(n30543), .A2(\xmem_data[12][1] ), .B1(n31269), .B2(
        \xmem_data[13][1] ), .ZN(n31034) );
  AOI22_X1 U33383 ( .A1(n22676), .A2(\xmem_data[14][1] ), .B1(n31270), .B2(
        \xmem_data[15][1] ), .ZN(n31033) );
  NAND4_X1 U33384 ( .A1(n31036), .A2(n31035), .A3(n31034), .A4(n31033), .ZN(
        n31037) );
  OR2_X1 U33385 ( .A1(n31038), .A2(n31037), .ZN(n31039) );
  NOR2_X1 U33386 ( .A1(n31040), .A2(n31039), .ZN(n31043) );
  NAND2_X1 U33387 ( .A1(n28343), .A2(\xmem_data[5][1] ), .ZN(n31042) );
  AOI21_X1 U33388 ( .B1(n31043), .B2(n31042), .A(n31041), .ZN(n31044) );
  INV_X1 U33389 ( .A(n31044), .ZN(n31110) );
  AOI22_X1 U33390 ( .A1(n31368), .A2(\xmem_data[96][1] ), .B1(n31367), .B2(
        \xmem_data[97][1] ), .ZN(n31048) );
  AOI22_X1 U33391 ( .A1(n20725), .A2(\xmem_data[98][1] ), .B1(n24564), .B2(
        \xmem_data[99][1] ), .ZN(n31047) );
  AOI22_X1 U33392 ( .A1(n30698), .A2(\xmem_data[100][1] ), .B1(n29306), .B2(
        \xmem_data[101][1] ), .ZN(n31046) );
  AOI22_X1 U33393 ( .A1(n30607), .A2(\xmem_data[102][1] ), .B1(n28415), .B2(
        \xmem_data[103][1] ), .ZN(n31045) );
  NAND4_X1 U33394 ( .A1(n31048), .A2(n31047), .A3(n31046), .A4(n31045), .ZN(
        n31064) );
  AOI22_X1 U33395 ( .A1(n31353), .A2(\xmem_data[104][1] ), .B1(n25423), .B2(
        \xmem_data[105][1] ), .ZN(n31052) );
  AOI22_X1 U33396 ( .A1(n28298), .A2(\xmem_data[106][1] ), .B1(n28052), .B2(
        \xmem_data[107][1] ), .ZN(n31051) );
  AOI22_X1 U33397 ( .A1(n31354), .A2(\xmem_data[108][1] ), .B1(n27864), .B2(
        \xmem_data[109][1] ), .ZN(n31050) );
  AOI22_X1 U33398 ( .A1(n21007), .A2(\xmem_data[110][1] ), .B1(n31355), .B2(
        \xmem_data[111][1] ), .ZN(n31049) );
  NAND4_X1 U33399 ( .A1(n31052), .A2(n31051), .A3(n31050), .A4(n31049), .ZN(
        n31063) );
  AOI22_X1 U33400 ( .A1(n17044), .A2(\xmem_data[112][1] ), .B1(n31360), .B2(
        \xmem_data[113][1] ), .ZN(n31056) );
  AOI22_X1 U33401 ( .A1(n29240), .A2(\xmem_data[114][1] ), .B1(n31361), .B2(
        \xmem_data[115][1] ), .ZN(n31055) );
  AOI22_X1 U33402 ( .A1(n29573), .A2(\xmem_data[116][1] ), .B1(n31362), .B2(
        \xmem_data[117][1] ), .ZN(n31054) );
  AOI22_X1 U33403 ( .A1(n27542), .A2(\xmem_data[118][1] ), .B1(n17049), .B2(
        \xmem_data[119][1] ), .ZN(n31053) );
  NAND4_X1 U33404 ( .A1(n31056), .A2(n31055), .A3(n31054), .A4(n31053), .ZN(
        n31062) );
  AOI22_X1 U33405 ( .A1(n31345), .A2(\xmem_data[120][1] ), .B1(n31344), .B2(
        \xmem_data[121][1] ), .ZN(n31060) );
  AOI22_X1 U33406 ( .A1(n25408), .A2(\xmem_data[122][1] ), .B1(n31346), .B2(
        \xmem_data[123][1] ), .ZN(n31059) );
  AOI22_X1 U33407 ( .A1(n3332), .A2(\xmem_data[124][1] ), .B1(n31347), .B2(
        \xmem_data[125][1] ), .ZN(n31058) );
  AOI22_X1 U33408 ( .A1(n31348), .A2(\xmem_data[126][1] ), .B1(n3217), .B2(
        \xmem_data[127][1] ), .ZN(n31057) );
  NAND4_X1 U33409 ( .A1(n31060), .A2(n31059), .A3(n31058), .A4(n31057), .ZN(
        n31061) );
  OR4_X1 U33410 ( .A1(n31064), .A2(n31063), .A3(n31062), .A4(n31061), .ZN(
        n31086) );
  AOI22_X1 U33411 ( .A1(n31368), .A2(\xmem_data[64][1] ), .B1(n31367), .B2(
        \xmem_data[65][1] ), .ZN(n31068) );
  AOI22_X1 U33412 ( .A1(n3342), .A2(\xmem_data[66][1] ), .B1(n28342), .B2(
        \xmem_data[67][1] ), .ZN(n31067) );
  AOI22_X1 U33413 ( .A1(n23742), .A2(\xmem_data[68][1] ), .B1(n25514), .B2(
        \xmem_data[69][1] ), .ZN(n31066) );
  AOI22_X1 U33414 ( .A1(n24638), .A2(\xmem_data[70][1] ), .B1(n3358), .B2(
        \xmem_data[71][1] ), .ZN(n31065) );
  NAND4_X1 U33415 ( .A1(n31068), .A2(n31067), .A3(n31066), .A4(n31065), .ZN(
        n31084) );
  AOI22_X1 U33416 ( .A1(n31353), .A2(\xmem_data[72][1] ), .B1(n22675), .B2(
        \xmem_data[73][1] ), .ZN(n31072) );
  AOI22_X1 U33417 ( .A1(n3175), .A2(\xmem_data[74][1] ), .B1(n25572), .B2(
        \xmem_data[75][1] ), .ZN(n31071) );
  AOI22_X1 U33418 ( .A1(n25607), .A2(\xmem_data[76][1] ), .B1(n20543), .B2(
        \xmem_data[77][1] ), .ZN(n31070) );
  AOI22_X1 U33419 ( .A1(n20542), .A2(\xmem_data[78][1] ), .B1(n31355), .B2(
        \xmem_data[79][1] ), .ZN(n31069) );
  NAND4_X1 U33420 ( .A1(n31072), .A2(n31071), .A3(n31070), .A4(n31069), .ZN(
        n31083) );
  AOI22_X1 U33421 ( .A1(n28302), .A2(\xmem_data[80][1] ), .B1(n31360), .B2(
        \xmem_data[81][1] ), .ZN(n31076) );
  AOI22_X1 U33422 ( .A1(n24647), .A2(\xmem_data[82][1] ), .B1(n31361), .B2(
        \xmem_data[83][1] ), .ZN(n31075) );
  AOI22_X1 U33423 ( .A1(n20817), .A2(\xmem_data[84][1] ), .B1(n31362), .B2(
        \xmem_data[85][1] ), .ZN(n31074) );
  AOI22_X1 U33424 ( .A1(n25582), .A2(\xmem_data[86][1] ), .B1(n28292), .B2(
        \xmem_data[87][1] ), .ZN(n31073) );
  NAND4_X1 U33425 ( .A1(n31076), .A2(n31075), .A3(n31074), .A4(n31073), .ZN(
        n31082) );
  AOI22_X1 U33426 ( .A1(n31345), .A2(\xmem_data[88][1] ), .B1(n31344), .B2(
        \xmem_data[89][1] ), .ZN(n31080) );
  AOI22_X1 U33427 ( .A1(n24526), .A2(\xmem_data[90][1] ), .B1(n31346), .B2(
        \xmem_data[91][1] ), .ZN(n31079) );
  AOI22_X1 U33428 ( .A1(n3433), .A2(\xmem_data[92][1] ), .B1(n31347), .B2(
        \xmem_data[93][1] ), .ZN(n31078) );
  AOI22_X1 U33429 ( .A1(n31348), .A2(\xmem_data[94][1] ), .B1(n3222), .B2(
        \xmem_data[95][1] ), .ZN(n31077) );
  NAND4_X1 U33430 ( .A1(n31080), .A2(n31079), .A3(n31078), .A4(n31077), .ZN(
        n31081) );
  OR4_X1 U33431 ( .A1(n31084), .A2(n31083), .A3(n31082), .A4(n31081), .ZN(
        n31085) );
  AOI22_X1 U33432 ( .A1(n31376), .A2(n31086), .B1(n31342), .B2(n31085), .ZN(
        n31109) );
  AOI22_X1 U33433 ( .A1(n24632), .A2(\xmem_data[32][1] ), .B1(n22667), .B2(
        \xmem_data[33][1] ), .ZN(n31090) );
  AOI22_X1 U33434 ( .A1(n17010), .A2(\xmem_data[34][1] ), .B1(n28342), .B2(
        \xmem_data[35][1] ), .ZN(n31089) );
  AOI22_X1 U33435 ( .A1(n20808), .A2(\xmem_data[36][1] ), .B1(n27547), .B2(
        \xmem_data[37][1] ), .ZN(n31088) );
  AOI22_X1 U33436 ( .A1(n31321), .A2(\xmem_data[38][1] ), .B1(n13475), .B2(
        \xmem_data[39][1] ), .ZN(n31087) );
  NAND4_X1 U33437 ( .A1(n31090), .A2(n31089), .A3(n31088), .A4(n31087), .ZN(
        n31106) );
  AOI22_X1 U33438 ( .A1(n31327), .A2(\xmem_data[40][1] ), .B1(n31326), .B2(
        \xmem_data[41][1] ), .ZN(n31094) );
  AOI22_X1 U33439 ( .A1(n28980), .A2(\xmem_data[42][1] ), .B1(n23715), .B2(
        \xmem_data[43][1] ), .ZN(n31093) );
  AOI22_X1 U33440 ( .A1(n31328), .A2(\xmem_data[44][1] ), .B1(n24457), .B2(
        \xmem_data[45][1] ), .ZN(n31092) );
  AOI22_X1 U33441 ( .A1(n31330), .A2(\xmem_data[46][1] ), .B1(n31329), .B2(
        \xmem_data[47][1] ), .ZN(n31091) );
  NAND4_X1 U33442 ( .A1(n31094), .A2(n31093), .A3(n31092), .A4(n31091), .ZN(
        n31105) );
  AOI22_X1 U33443 ( .A1(n21008), .A2(\xmem_data[48][1] ), .B1(n25399), .B2(
        \xmem_data[49][1] ), .ZN(n31098) );
  AOI22_X1 U33444 ( .A1(n28493), .A2(\xmem_data[50][1] ), .B1(n24117), .B2(
        \xmem_data[51][1] ), .ZN(n31097) );
  AOI22_X1 U33445 ( .A1(n31315), .A2(\xmem_data[52][1] ), .B1(n31314), .B2(
        \xmem_data[53][1] ), .ZN(n31096) );
  AOI22_X1 U33446 ( .A1(n31316), .A2(\xmem_data[54][1] ), .B1(n27463), .B2(
        \xmem_data[55][1] ), .ZN(n31095) );
  NAND4_X1 U33447 ( .A1(n31098), .A2(n31097), .A3(n31096), .A4(n31095), .ZN(
        n31104) );
  AOI22_X1 U33448 ( .A1(n31308), .A2(\xmem_data[56][1] ), .B1(n20769), .B2(
        \xmem_data[57][1] ), .ZN(n31102) );
  AOI22_X1 U33449 ( .A1(n3380), .A2(\xmem_data[58][1] ), .B1(n31309), .B2(
        \xmem_data[59][1] ), .ZN(n31101) );
  AOI22_X1 U33450 ( .A1(n23754), .A2(\xmem_data[60][1] ), .B1(n28501), .B2(
        \xmem_data[61][1] ), .ZN(n31100) );
  AOI22_X1 U33451 ( .A1(n24631), .A2(\xmem_data[62][1] ), .B1(n3217), .B2(
        \xmem_data[63][1] ), .ZN(n31099) );
  NAND4_X1 U33452 ( .A1(n31102), .A2(n31101), .A3(n31100), .A4(n31099), .ZN(
        n31103) );
  OR4_X1 U33453 ( .A1(n31106), .A2(n31105), .A3(n31104), .A4(n31103), .ZN(
        n31107) );
  NAND2_X1 U33454 ( .A1(n31107), .A2(n31340), .ZN(n31108) );
  XNOR2_X1 U33455 ( .A(n34610), .B(\fmem_data[12][5] ), .ZN(n32135) );
  OAI22_X1 U33456 ( .A1(n32135), .A2(n33973), .B1(n33974), .B2(n33975), .ZN(
        n31914) );
  XNOR2_X1 U33457 ( .A(n31592), .B(\fmem_data[29][3] ), .ZN(n32529) );
  XNOR2_X1 U33458 ( .A(n32242), .B(\fmem_data[29][3] ), .ZN(n33965) );
  OAI21_X1 U33459 ( .B1(n31913), .B2(n31914), .A(n31915), .ZN(n31112) );
  NAND2_X1 U33460 ( .A1(n31112), .A2(n31111), .ZN(n31113) );
  FA_X1 U33461 ( .A(n31115), .B(n31114), .CI(n31113), .CO(n31870), .S(n32475)
         );
  FA_X1 U33462 ( .A(n31118), .B(n31117), .CI(n31116), .CO(n31878), .S(n32055)
         );
  FA_X1 U33463 ( .A(n31121), .B(n31120), .CI(n31119), .CO(n31147), .S(n32054)
         );
  XNOR2_X1 U33464 ( .A(n36312), .B(\fmem_data[10][5] ), .ZN(n31124) );
  XNOR2_X1 U33465 ( .A(n31128), .B(n31127), .ZN(n31130) );
  XNOR2_X1 U33466 ( .A(n31130), .B(n31129), .ZN(n32473) );
  FA_X1 U33467 ( .A(n31133), .B(n31132), .CI(n31131), .CO(n31413), .S(n32468)
         );
  FA_X1 U33468 ( .A(n31136), .B(n31135), .CI(n31134), .CO(n31143), .S(n32087)
         );
  FA_X1 U33469 ( .A(n31139), .B(n31138), .CI(n31137), .CO(n31148), .S(n32086)
         );
  FA_X1 U33470 ( .A(n31142), .B(n31141), .CI(n31140), .CO(n31189), .S(n32085)
         );
  XNOR2_X1 U33471 ( .A(n31144), .B(n31143), .ZN(n31145) );
  XNOR2_X1 U33472 ( .A(n31146), .B(n31145), .ZN(n32478) );
  FA_X1 U33473 ( .A(n31149), .B(n31148), .CI(n31147), .CO(n31178), .S(n32476)
         );
  OAI21_X1 U33474 ( .B1(n32477), .B2(n32478), .A(n32476), .ZN(n31151) );
  NAND2_X1 U33475 ( .A1(n32477), .A2(n3393), .ZN(n31150) );
  NAND2_X1 U33476 ( .A1(n31151), .A2(n31150), .ZN(n32103) );
  FA_X1 U33477 ( .A(n31154), .B(n31153), .CI(n31152), .CO(n31930), .S(n32102)
         );
  FA_X1 U33478 ( .A(n31157), .B(n31156), .CI(n31155), .CO(n31152), .S(n31438)
         );
  FA_X1 U33479 ( .A(n31160), .B(n31159), .CI(n31158), .CO(n31183), .S(n31437)
         );
  XNOR2_X1 U33480 ( .A(n31161), .B(\fmem_data[22][1] ), .ZN(n33809) );
  XNOR2_X1 U33481 ( .A(n32005), .B(\fmem_data[16][3] ), .ZN(n31453) );
  OAI22_X1 U33482 ( .A1(n31165), .A2(n35006), .B1(n31164), .B2(n35007), .ZN(
        n32082) );
  XNOR2_X1 U33483 ( .A(n36101), .B(\fmem_data[24][5] ), .ZN(n31166) );
  OAI22_X1 U33484 ( .A1(n31167), .A2(n34039), .B1(n31166), .B2(n34041), .ZN(
        n32491) );
  OR2_X1 U33485 ( .A1(n36313), .A2(n3697), .ZN(n31170) );
  XNOR2_X1 U33486 ( .A(n32727), .B(\fmem_data[19][1] ), .ZN(n32426) );
  OAI22_X1 U33487 ( .A1(n32426), .A2(n36226), .B1(n31171), .B2(n3633), .ZN(
        n32495) );
  XNOR2_X1 U33488 ( .A(n36315), .B(\fmem_data[3][5] ), .ZN(n31175) );
  OAI22_X1 U33489 ( .A1(n31175), .A2(n34918), .B1(n31174), .B2(n34919), .ZN(
        n32493) );
  OAI21_X1 U33490 ( .B1(n32495), .B2(n32492), .A(n32493), .ZN(n31177) );
  NAND2_X1 U33491 ( .A1(n31177), .A2(n31176), .ZN(n32483) );
  FA_X1 U33492 ( .A(n31180), .B(n31179), .CI(n31178), .CO(n31931), .S(n32499)
         );
  FA_X1 U33493 ( .A(n31183), .B(n31182), .CI(n31181), .CO(n31861), .S(n32500)
         );
  FA_X1 U33494 ( .A(n31186), .B(n31185), .CI(n31184), .CO(n31404), .S(n31435)
         );
  FA_X1 U33495 ( .A(n31189), .B(n31187), .CI(n31188), .CO(n31210), .S(n31434)
         );
  XNOR2_X1 U33496 ( .A(n31191), .B(n31190), .ZN(n31193) );
  XNOR2_X1 U33497 ( .A(n32427), .B(\fmem_data[8][3] ), .ZN(n34209) );
  XNOR2_X1 U33498 ( .A(n36314), .B(n3488), .ZN(n31194) );
  OAI22_X1 U33499 ( .A1(n33880), .A2(n34944), .B1(n31194), .B2(n34945), .ZN(
        n31496) );
  XNOR2_X1 U33500 ( .A(n36228), .B(\fmem_data[20][5] ), .ZN(n31195) );
  XNOR2_X1 U33501 ( .A(n3116), .B(\fmem_data[23][5] ), .ZN(n31197) );
  XNOR2_X1 U33502 ( .A(n3451), .B(\fmem_data[3][3] ), .ZN(n33895) );
  XNOR2_X1 U33503 ( .A(n33720), .B(\fmem_data[3][3] ), .ZN(n34421) );
  OR2_X1 U33504 ( .A1(n3116), .A2(n3687), .ZN(n31198) );
  OAI21_X1 U33505 ( .B1(n32499), .B2(n32500), .A(n32501), .ZN(n31200) );
  NAND2_X1 U33506 ( .A1(n31200), .A2(n31199), .ZN(n32466) );
  XNOR2_X1 U33507 ( .A(n31635), .B(n31634), .ZN(n31418) );
  XNOR2_X1 U33508 ( .A(n31201), .B(n31202), .ZN(n31204) );
  XNOR2_X1 U33509 ( .A(n31204), .B(n31203), .ZN(n31421) );
  FA_X1 U33510 ( .A(n31207), .B(n31206), .CI(n31205), .CO(n31240), .S(n31432)
         );
  XNOR2_X1 U33511 ( .A(n31209), .B(n31208), .ZN(n31211) );
  XNOR2_X1 U33512 ( .A(n31211), .B(n31210), .ZN(n31431) );
  FA_X1 U33513 ( .A(n31214), .B(n31213), .CI(n31212), .CO(n31187), .S(n31440)
         );
  FA_X1 U33514 ( .A(n31217), .B(n31216), .CI(n31215), .CO(n31128), .S(n31439)
         );
  OR2_X1 U33515 ( .A1(n31440), .A2(n31439), .ZN(n31222) );
  XNOR2_X1 U33516 ( .A(n31219), .B(\fmem_data[26][1] ), .ZN(n32555) );
  XNOR2_X1 U33517 ( .A(n31220), .B(\fmem_data[26][1] ), .ZN(n33640) );
  OAI22_X1 U33518 ( .A1(n32555), .A2(n33725), .B1(n33640), .B2(n3678), .ZN(
        n31558) );
  XNOR2_X1 U33519 ( .A(n32165), .B(\fmem_data[2][1] ), .ZN(n32788) );
  XNOR2_X1 U33520 ( .A(n31221), .B(\fmem_data[2][1] ), .ZN(n32526) );
  OAI22_X1 U33521 ( .A1(n32788), .A2(n34343), .B1(n3578), .B2(n32526), .ZN(
        n31557) );
  XNOR2_X1 U33522 ( .A(n33553), .B(\fmem_data[5][3] ), .ZN(n32424) );
  XNOR2_X1 U33523 ( .A(n32419), .B(\fmem_data[5][3] ), .ZN(n33852) );
  OAI22_X1 U33524 ( .A1(n32424), .A2(n33851), .B1(n33852), .B2(n33850), .ZN(
        n31556) );
  XNOR2_X1 U33525 ( .A(n33019), .B(\fmem_data[23][3] ), .ZN(n34020) );
  XNOR2_X1 U33526 ( .A(n32929), .B(\fmem_data[23][3] ), .ZN(n34413) );
  NAND2_X1 U33527 ( .A1(n31222), .A2(n31441), .ZN(n31224) );
  NAND2_X1 U33528 ( .A1(n31224), .A2(n31223), .ZN(n31601) );
  XNOR2_X1 U33529 ( .A(n36339), .B(\fmem_data[15][5] ), .ZN(n31226) );
  XNOR2_X1 U33530 ( .A(n33479), .B(\fmem_data[15][5] ), .ZN(n33940) );
  OAI22_X1 U33531 ( .A1(n31226), .A2(n34989), .B1(n33940), .B2(n34990), .ZN(
        n31608) );
  XNOR2_X1 U33532 ( .A(n32440), .B(\fmem_data[7][3] ), .ZN(n33992) );
  XNOR2_X1 U33533 ( .A(n3313), .B(\fmem_data[7][3] ), .ZN(n32604) );
  FA_X1 U33534 ( .A(n31229), .B(n31228), .CI(n31227), .CO(n31184), .S(n31548)
         );
  XNOR2_X1 U33535 ( .A(n32444), .B(\fmem_data[27][3] ), .ZN(n33996) );
  XNOR2_X1 U33536 ( .A(n32978), .B(\fmem_data[27][3] ), .ZN(n34426) );
  OAI22_X1 U33537 ( .A1(n34463), .A2(n33996), .B1(n34462), .B2(n34426), .ZN(
        n31615) );
  XNOR2_X1 U33538 ( .A(n36313), .B(\fmem_data[11][5] ), .ZN(n31230) );
  OAI22_X1 U33539 ( .A1(n31231), .A2(n34932), .B1(n31230), .B2(n34933), .ZN(
        n31614) );
  INV_X1 U33540 ( .A(n33963), .ZN(n31232) );
  XNOR2_X1 U33541 ( .A(n31233), .B(\fmem_data[5][1] ), .ZN(n34022) );
  OAI22_X1 U33542 ( .A1(n32420), .A2(n34483), .B1(n34022), .B2(n3576), .ZN(
        n31530) );
  FA_X1 U33543 ( .A(n31236), .B(n31235), .CI(n31234), .CO(n31407), .S(n31600)
         );
  OAI21_X1 U33544 ( .B1(n31601), .B2(n31602), .A(n31600), .ZN(n31238) );
  NAND2_X1 U33545 ( .A1(n31238), .A2(n31237), .ZN(n31430) );
  FA_X1 U33546 ( .A(n31241), .B(n31240), .CI(n31239), .CO(n31412), .S(n31426)
         );
  XNOR2_X1 U33547 ( .A(n31980), .B(\fmem_data[27][1] ), .ZN(n34190) );
  XNOR2_X1 U33548 ( .A(n3278), .B(\fmem_data[27][1] ), .ZN(n32445) );
  OAI22_X1 U33549 ( .A1(n34190), .A2(n3482), .B1(n32445), .B2(n36240), .ZN(
        n31564) );
  XNOR2_X1 U33550 ( .A(n32256), .B(\fmem_data[23][1] ), .ZN(n32417) );
  OAI22_X1 U33551 ( .A1(n33905), .A2(n3662), .B1(n32417), .B2(n36241), .ZN(
        n31611) );
  XNOR2_X1 U33552 ( .A(n31246), .B(\fmem_data[11][1] ), .ZN(n33946) );
  XNOR2_X1 U33553 ( .A(n3316), .B(\fmem_data[11][1] ), .ZN(n33778) );
  XNOR2_X1 U33554 ( .A(n36316), .B(\fmem_data[27][5] ), .ZN(n31249) );
  XNOR2_X1 U33555 ( .A(n32438), .B(\fmem_data[31][3] ), .ZN(n33907) );
  AOI22_X1 U33556 ( .A1(n27396), .A2(\xmem_data[4][0] ), .B1(n28343), .B2(
        \xmem_data[5][0] ), .ZN(n31253) );
  INV_X1 U33557 ( .A(n31253), .ZN(n31286) );
  AOI22_X1 U33558 ( .A1(n31255), .A2(\xmem_data[16][0] ), .B1(n31254), .B2(
        \xmem_data[17][0] ), .ZN(n31260) );
  AOI22_X1 U33559 ( .A1(n30956), .A2(\xmem_data[18][0] ), .B1(n28494), .B2(
        \xmem_data[19][0] ), .ZN(n31259) );
  AOI22_X1 U33560 ( .A1(n3269), .A2(\xmem_data[20][0] ), .B1(n29245), .B2(
        \xmem_data[21][0] ), .ZN(n31258) );
  AOI22_X1 U33561 ( .A1(n24467), .A2(\xmem_data[22][0] ), .B1(n31256), .B2(
        \xmem_data[23][0] ), .ZN(n31257) );
  NAND4_X1 U33562 ( .A1(n31260), .A2(n31259), .A3(n31258), .A4(n31257), .ZN(
        n31283) );
  AOI22_X1 U33563 ( .A1(n30901), .A2(\xmem_data[24][0] ), .B1(n31261), .B2(
        \xmem_data[25][0] ), .ZN(n31267) );
  AOI22_X1 U33564 ( .A1(n3380), .A2(\xmem_data[26][0] ), .B1(n31262), .B2(
        \xmem_data[27][0] ), .ZN(n31266) );
  AOI22_X1 U33565 ( .A1(n3142), .A2(\xmem_data[28][0] ), .B1(n27501), .B2(
        \xmem_data[29][0] ), .ZN(n31265) );
  AOI22_X1 U33566 ( .A1(n25508), .A2(\xmem_data[30][0] ), .B1(n3220), .B2(
        \xmem_data[31][0] ), .ZN(n31264) );
  NAND4_X1 U33567 ( .A1(n31267), .A2(n31266), .A3(n31265), .A4(n31264), .ZN(
        n31282) );
  AOI22_X1 U33568 ( .A1(n28152), .A2(\xmem_data[8][0] ), .B1(n24212), .B2(
        \xmem_data[9][0] ), .ZN(n31274) );
  AOI22_X1 U33569 ( .A1(n31268), .A2(\xmem_data[10][0] ), .B1(n28052), .B2(
        \xmem_data[11][0] ), .ZN(n31273) );
  AOI22_X1 U33570 ( .A1(n16988), .A2(\xmem_data[12][0] ), .B1(n31269), .B2(
        \xmem_data[13][0] ), .ZN(n31272) );
  AOI22_X1 U33571 ( .A1(n29010), .A2(\xmem_data[14][0] ), .B1(n31270), .B2(
        \xmem_data[15][0] ), .ZN(n31271) );
  NAND4_X1 U33572 ( .A1(n31274), .A2(n31273), .A3(n31272), .A4(n31271), .ZN(
        n31281) );
  AOI22_X1 U33573 ( .A1(n23741), .A2(\xmem_data[2][0] ), .B1(n31275), .B2(
        \xmem_data[3][0] ), .ZN(n31279) );
  AOI22_X1 U33574 ( .A1(n31276), .A2(\xmem_data[6][0] ), .B1(n14933), .B2(
        \xmem_data[7][0] ), .ZN(n31278) );
  AOI22_X1 U33575 ( .A1(n29789), .A2(\xmem_data[0][0] ), .B1(n20500), .B2(
        \xmem_data[1][0] ), .ZN(n31277) );
  NAND3_X1 U33576 ( .A1(n31279), .A2(n31278), .A3(n31277), .ZN(n31280) );
  OR4_X1 U33577 ( .A1(n31283), .A2(n31282), .A3(n31281), .A4(n31280), .ZN(
        n31285) );
  OAI21_X1 U33578 ( .B1(n31286), .B2(n31285), .A(n31284), .ZN(n31381) );
  AOI22_X1 U33579 ( .A1(n31345), .A2(\xmem_data[88][0] ), .B1(n31344), .B2(
        \xmem_data[89][0] ), .ZN(n31291) );
  AOI22_X1 U33580 ( .A1(n20710), .A2(\xmem_data[90][0] ), .B1(n31346), .B2(
        \xmem_data[91][0] ), .ZN(n31290) );
  AOI22_X1 U33581 ( .A1(n3142), .A2(\xmem_data[92][0] ), .B1(n31347), .B2(
        \xmem_data[93][0] ), .ZN(n31289) );
  AND2_X1 U33582 ( .A1(n3221), .A2(\xmem_data[95][0] ), .ZN(n31287) );
  AOI21_X1 U33583 ( .B1(n31348), .B2(\xmem_data[94][0] ), .A(n31287), .ZN(
        n31288) );
  NAND4_X1 U33584 ( .A1(n31291), .A2(n31290), .A3(n31289), .A4(n31288), .ZN(
        n31307) );
  AOI22_X1 U33585 ( .A1(n31353), .A2(\xmem_data[72][0] ), .B1(n28515), .B2(
        \xmem_data[73][0] ), .ZN(n31295) );
  AOI22_X1 U33586 ( .A1(n3176), .A2(\xmem_data[74][0] ), .B1(n29046), .B2(
        \xmem_data[75][0] ), .ZN(n31294) );
  AOI22_X1 U33587 ( .A1(n25461), .A2(\xmem_data[76][0] ), .B1(n13188), .B2(
        \xmem_data[77][0] ), .ZN(n31293) );
  AOI22_X1 U33588 ( .A1(n25434), .A2(\xmem_data[78][0] ), .B1(n31355), .B2(
        \xmem_data[79][0] ), .ZN(n31292) );
  NAND4_X1 U33589 ( .A1(n31295), .A2(n31294), .A3(n31293), .A4(n31292), .ZN(
        n31306) );
  AOI22_X1 U33590 ( .A1(n17044), .A2(\xmem_data[80][0] ), .B1(n31360), .B2(
        \xmem_data[81][0] ), .ZN(n31299) );
  AOI22_X1 U33591 ( .A1(n27524), .A2(\xmem_data[82][0] ), .B1(n31361), .B2(
        \xmem_data[83][0] ), .ZN(n31298) );
  AOI22_X1 U33592 ( .A1(n28701), .A2(\xmem_data[84][0] ), .B1(n31362), .B2(
        \xmem_data[85][0] ), .ZN(n31297) );
  AOI22_X1 U33593 ( .A1(n20782), .A2(\xmem_data[86][0] ), .B1(n28500), .B2(
        \xmem_data[87][0] ), .ZN(n31296) );
  NAND4_X1 U33594 ( .A1(n31299), .A2(n31298), .A3(n31297), .A4(n31296), .ZN(
        n31305) );
  AOI22_X1 U33595 ( .A1(n31368), .A2(\xmem_data[64][0] ), .B1(n31367), .B2(
        \xmem_data[65][0] ), .ZN(n31303) );
  AOI22_X1 U33596 ( .A1(n24565), .A2(\xmem_data[66][0] ), .B1(n22711), .B2(
        \xmem_data[67][0] ), .ZN(n31302) );
  AOI22_X1 U33597 ( .A1(n3128), .A2(\xmem_data[68][0] ), .B1(n28007), .B2(
        \xmem_data[69][0] ), .ZN(n31301) );
  AOI22_X1 U33598 ( .A1(n27447), .A2(\xmem_data[70][0] ), .B1(n20546), .B2(
        \xmem_data[71][0] ), .ZN(n31300) );
  NAND4_X1 U33599 ( .A1(n31303), .A2(n31302), .A3(n31301), .A4(n31300), .ZN(
        n31304) );
  OR4_X1 U33600 ( .A1(n31307), .A2(n31306), .A3(n31305), .A4(n31304), .ZN(
        n31343) );
  AOI22_X1 U33601 ( .A1(n31308), .A2(\xmem_data[56][0] ), .B1(n24686), .B2(
        \xmem_data[57][0] ), .ZN(n31313) );
  AOI22_X1 U33602 ( .A1(n24688), .A2(\xmem_data[58][0] ), .B1(n31309), .B2(
        \xmem_data[59][0] ), .ZN(n31312) );
  AOI22_X1 U33603 ( .A1(n3387), .A2(\xmem_data[60][0] ), .B1(n13468), .B2(
        \xmem_data[61][0] ), .ZN(n31311) );
  AOI22_X1 U33604 ( .A1(n25508), .A2(\xmem_data[62][0] ), .B1(n3217), .B2(
        \xmem_data[63][0] ), .ZN(n31310) );
  NAND4_X1 U33605 ( .A1(n31313), .A2(n31312), .A3(n31311), .A4(n31310), .ZN(
        n31339) );
  AOI22_X1 U33606 ( .A1(n23722), .A2(\xmem_data[48][0] ), .B1(n30515), .B2(
        \xmem_data[49][0] ), .ZN(n31320) );
  AOI22_X1 U33607 ( .A1(n21010), .A2(\xmem_data[50][0] ), .B1(n28429), .B2(
        \xmem_data[51][0] ), .ZN(n31319) );
  AOI22_X1 U33608 ( .A1(n31315), .A2(\xmem_data[52][0] ), .B1(n31314), .B2(
        \xmem_data[53][0] ), .ZN(n31318) );
  AOI22_X1 U33609 ( .A1(n31316), .A2(\xmem_data[54][0] ), .B1(n25723), .B2(
        \xmem_data[55][0] ), .ZN(n31317) );
  NAND4_X1 U33610 ( .A1(n31320), .A2(n31319), .A3(n31318), .A4(n31317), .ZN(
        n31337) );
  AOI22_X1 U33611 ( .A1(n25414), .A2(\xmem_data[32][0] ), .B1(n22710), .B2(
        \xmem_data[33][0] ), .ZN(n31325) );
  AOI22_X1 U33612 ( .A1(n28475), .A2(\xmem_data[34][0] ), .B1(n30882), .B2(
        \xmem_data[35][0] ), .ZN(n31324) );
  AOI22_X1 U33613 ( .A1(n27396), .A2(\xmem_data[36][0] ), .B1(n24657), .B2(
        \xmem_data[37][0] ), .ZN(n31323) );
  AOI22_X1 U33614 ( .A1(n31321), .A2(\xmem_data[38][0] ), .B1(n13475), .B2(
        \xmem_data[39][0] ), .ZN(n31322) );
  NAND4_X1 U33615 ( .A1(n31325), .A2(n31324), .A3(n31323), .A4(n31322), .ZN(
        n31336) );
  AOI22_X1 U33616 ( .A1(n31327), .A2(\xmem_data[40][0] ), .B1(n31326), .B2(
        \xmem_data[41][0] ), .ZN(n31334) );
  AOI22_X1 U33617 ( .A1(n24131), .A2(\xmem_data[42][0] ), .B1(n25382), .B2(
        \xmem_data[43][0] ), .ZN(n31333) );
  AOI22_X1 U33618 ( .A1(n31328), .A2(\xmem_data[44][0] ), .B1(n23716), .B2(
        \xmem_data[45][0] ), .ZN(n31332) );
  AOI22_X1 U33619 ( .A1(n31330), .A2(\xmem_data[46][0] ), .B1(n31329), .B2(
        \xmem_data[47][0] ), .ZN(n31331) );
  NAND4_X1 U33620 ( .A1(n31334), .A2(n31333), .A3(n31332), .A4(n31331), .ZN(
        n31335) );
  OR3_X1 U33621 ( .A1(n31337), .A2(n31336), .A3(n31335), .ZN(n31338) );
  OR2_X1 U33622 ( .A1(n31339), .A2(n31338), .ZN(n31341) );
  AOI22_X1 U33623 ( .A1(n31343), .A2(n31342), .B1(n31341), .B2(n31340), .ZN(
        n31380) );
  AOI22_X1 U33624 ( .A1(n31345), .A2(\xmem_data[120][0] ), .B1(n31344), .B2(
        \xmem_data[121][0] ), .ZN(n31352) );
  AOI22_X1 U33625 ( .A1(n29124), .A2(\xmem_data[122][0] ), .B1(n31346), .B2(
        \xmem_data[123][0] ), .ZN(n31351) );
  AOI22_X1 U33626 ( .A1(n25725), .A2(\xmem_data[124][0] ), .B1(n31347), .B2(
        \xmem_data[125][0] ), .ZN(n31350) );
  AOI22_X1 U33627 ( .A1(n31348), .A2(\xmem_data[126][0] ), .B1(n3222), .B2(
        \xmem_data[127][0] ), .ZN(n31349) );
  NAND4_X1 U33628 ( .A1(n31352), .A2(n31351), .A3(n31350), .A4(n31349), .ZN(
        n31378) );
  AOI22_X1 U33629 ( .A1(n31353), .A2(\xmem_data[104][0] ), .B1(n27452), .B2(
        \xmem_data[105][0] ), .ZN(n31359) );
  AOI22_X1 U33630 ( .A1(n28298), .A2(\xmem_data[106][0] ), .B1(n30613), .B2(
        \xmem_data[107][0] ), .ZN(n31358) );
  AOI22_X1 U33631 ( .A1(n30948), .A2(\xmem_data[108][0] ), .B1(n27989), .B2(
        \xmem_data[109][0] ), .ZN(n31357) );
  AOI22_X1 U33632 ( .A1(n29317), .A2(\xmem_data[110][0] ), .B1(n31355), .B2(
        \xmem_data[111][0] ), .ZN(n31356) );
  NAND4_X1 U33633 ( .A1(n31359), .A2(n31358), .A3(n31357), .A4(n31356), .ZN(
        n31375) );
  AOI22_X1 U33634 ( .A1(n20815), .A2(\xmem_data[112][0] ), .B1(n31360), .B2(
        \xmem_data[113][0] ), .ZN(n31366) );
  AOI22_X1 U33635 ( .A1(n3205), .A2(\xmem_data[114][0] ), .B1(n31361), .B2(
        \xmem_data[115][0] ), .ZN(n31365) );
  AOI22_X1 U33636 ( .A1(n30311), .A2(\xmem_data[116][0] ), .B1(n31362), .B2(
        \xmem_data[117][0] ), .ZN(n31364) );
  AOI22_X1 U33637 ( .A1(n25582), .A2(\xmem_data[118][0] ), .B1(n25406), .B2(
        \xmem_data[119][0] ), .ZN(n31363) );
  NAND4_X1 U33638 ( .A1(n31366), .A2(n31365), .A3(n31364), .A4(n31363), .ZN(
        n31374) );
  AOI22_X1 U33639 ( .A1(n31368), .A2(\xmem_data[96][0] ), .B1(n31367), .B2(
        \xmem_data[97][0] ), .ZN(n31372) );
  AOI22_X1 U33640 ( .A1(n24141), .A2(\xmem_data[98][0] ), .B1(n22711), .B2(
        \xmem_data[99][0] ), .ZN(n31371) );
  AOI22_X1 U33641 ( .A1(n30295), .A2(\xmem_data[100][0] ), .B1(n28510), .B2(
        \xmem_data[101][0] ), .ZN(n31370) );
  AOI22_X1 U33642 ( .A1(n20961), .A2(\xmem_data[102][0] ), .B1(n3357), .B2(
        \xmem_data[103][0] ), .ZN(n31369) );
  NAND4_X1 U33643 ( .A1(n31372), .A2(n31371), .A3(n31370), .A4(n31369), .ZN(
        n31373) );
  OR3_X1 U33644 ( .A1(n31375), .A2(n31374), .A3(n31373), .ZN(n31377) );
  OAI21_X1 U33645 ( .B1(n31378), .B2(n31377), .A(n31376), .ZN(n31379) );
  INV_X1 U33646 ( .A(n33975), .ZN(n31382) );
  XNOR2_X1 U33647 ( .A(n32283), .B(\fmem_data[18][1] ), .ZN(n32437) );
  XNOR2_X1 U33648 ( .A(n3442), .B(\fmem_data[18][1] ), .ZN(n33792) );
  OAI22_X1 U33649 ( .A1(n32437), .A2(n36104), .B1(n33792), .B2(n3580), .ZN(
        n31523) );
  OAI22_X1 U33650 ( .A1(n32422), .A2(n33796), .B1(n3456), .B2(n33797), .ZN(
        n31524) );
  OAI21_X1 U33651 ( .B1(n31522), .B2(n31523), .A(n31524), .ZN(n31385) );
  NAND2_X1 U33652 ( .A1(n31385), .A2(n31384), .ZN(n31554) );
  XNOR2_X1 U33653 ( .A(n3272), .B(\fmem_data[31][1] ), .ZN(n34112) );
  XNOR2_X1 U33654 ( .A(n3320), .B(\fmem_data[31][1] ), .ZN(n32439) );
  FA_X1 U33655 ( .A(n31389), .B(n31388), .CI(n31387), .CO(n31186), .S(n31463)
         );
  XNOR2_X1 U33656 ( .A(n32936), .B(\fmem_data[19][3] ), .ZN(n32595) );
  OAI22_X1 U33657 ( .A1(n34192), .A2(n34472), .B1(n32595), .B2(n34474), .ZN(
        n31578) );
  XNOR2_X1 U33658 ( .A(n32616), .B(\fmem_data[9][3] ), .ZN(n33876) );
  OR2_X1 U33659 ( .A1(n36316), .A2(n3636), .ZN(n31397) );
  OAI22_X1 U33660 ( .A1(n31398), .A2(n34835), .B1(n34836), .B2(n3648), .ZN(
        n31571) );
  XNOR2_X1 U33661 ( .A(n32953), .B(\fmem_data[26][3] ), .ZN(n32434) );
  OAI22_X1 U33662 ( .A1(n32434), .A2(n32779), .B1(n32780), .B2(n31399), .ZN(
        n31521) );
  INV_X1 U33663 ( .A(n33328), .ZN(n31400) );
  INV_X1 U33664 ( .A(n33105), .ZN(n31401) );
  XNOR2_X1 U33665 ( .A(n33027), .B(\fmem_data[7][1] ), .ZN(n33989) );
  XNOR2_X1 U33666 ( .A(n32174), .B(\fmem_data[7][1] ), .ZN(n32441) );
  OAI22_X1 U33667 ( .A1(n33989), .A2(n3581), .B1(n32441), .B2(n36218), .ZN(
        n31569) );
  XNOR2_X1 U33668 ( .A(n3366), .B(\fmem_data[3][1] ), .ZN(n33872) );
  XNOR2_X1 U33669 ( .A(n3262), .B(\fmem_data[3][1] ), .ZN(n32561) );
  OAI22_X1 U33670 ( .A1(n33872), .A2(n3582), .B1(n32561), .B2(n36199), .ZN(
        n31568) );
  XNOR2_X1 U33671 ( .A(n32603), .B(\fmem_data[7][5] ), .ZN(n34072) );
  XNOR2_X1 U33672 ( .A(n36311), .B(\fmem_data[7][5] ), .ZN(n31403) );
  OAI22_X1 U33673 ( .A1(n34072), .A2(n34835), .B1(n31403), .B2(n34836), .ZN(
        n31567) );
  FA_X1 U33674 ( .A(n31406), .B(n31405), .CI(n31404), .CO(n31132), .S(n31629)
         );
  FA_X1 U33675 ( .A(n31409), .B(n31408), .CI(n31407), .CO(n31131), .S(n31628)
         );
  OAI21_X1 U33676 ( .B1(n31427), .B2(n31426), .A(n31428), .ZN(n31411) );
  NAND2_X1 U33677 ( .A1(n31411), .A2(n31410), .ZN(n31420) );
  XNOR2_X1 U33678 ( .A(n31415), .B(n31414), .ZN(n31419) );
  OAI21_X1 U33679 ( .B1(n31421), .B2(n31420), .A(n31419), .ZN(n31417) );
  NAND2_X1 U33680 ( .A1(n31421), .A2(n31420), .ZN(n31416) );
  NAND2_X1 U33681 ( .A1(n31417), .A2(n31416), .ZN(n31633) );
  XNOR2_X1 U33682 ( .A(n31418), .B(n31633), .ZN(n33405) );
  XNOR2_X1 U33683 ( .A(n31420), .B(n31419), .ZN(n31422) );
  XNOR2_X1 U33684 ( .A(n31422), .B(n31421), .ZN(n33411) );
  FA_X1 U33685 ( .A(n31424), .B(n31425), .CI(n31423), .CO(n35438), .S(n33410)
         );
  XNOR2_X1 U33686 ( .A(n31427), .B(n31426), .ZN(n31429) );
  XNOR2_X1 U33687 ( .A(n31429), .B(n31428), .ZN(n33418) );
  FA_X1 U33688 ( .A(n31432), .B(n31431), .CI(n31430), .CO(n31427), .S(n33525)
         );
  FA_X1 U33689 ( .A(n31434), .B(n31435), .CI(n31433), .CO(n32501), .S(n33424)
         );
  FA_X1 U33690 ( .A(n31438), .B(n31437), .CI(n31436), .CO(n32101), .S(n33423)
         );
  XNOR2_X1 U33691 ( .A(n31440), .B(n31439), .ZN(n31442) );
  XNOR2_X1 U33692 ( .A(n31442), .B(n31441), .ZN(n33427) );
  XNOR2_X1 U33693 ( .A(n32513), .B(\fmem_data[25][3] ), .ZN(n32079) );
  OAI22_X1 U33694 ( .A1(n31445), .A2(n35011), .B1(n31444), .B2(n35010), .ZN(
        n31918) );
  INV_X1 U33695 ( .A(n33250), .ZN(n31447) );
  INV_X1 U33696 ( .A(n34206), .ZN(n31448) );
  INV_X1 U33697 ( .A(n33174), .ZN(n31449) );
  XNOR2_X1 U33698 ( .A(n31452), .B(\fmem_data[10][1] ), .ZN(n34532) );
  XNOR2_X1 U33699 ( .A(n33754), .B(\fmem_data[0][3] ), .ZN(n34538) );
  INV_X1 U33700 ( .A(n32975), .ZN(n31455) );
  INV_X1 U33701 ( .A(n32974), .ZN(n31454) );
  NAND2_X1 U33702 ( .A1(n31455), .A2(n31454), .ZN(n31456) );
  NAND2_X1 U33703 ( .A1(n32977), .A2(n31456), .ZN(n31458) );
  NAND2_X1 U33704 ( .A1(n31458), .A2(n31457), .ZN(n33432) );
  FA_X1 U33705 ( .A(n31461), .B(n31460), .CI(n31459), .CO(n32053), .S(n33431)
         );
  FA_X1 U33706 ( .A(n31464), .B(n31463), .CI(n31462), .CO(n31622), .S(n33425)
         );
  XNOR2_X1 U33707 ( .A(n31466), .B(n31465), .ZN(n31468) );
  XNOR2_X1 U33708 ( .A(n31468), .B(n31467), .ZN(n33669) );
  XNOR2_X1 U33709 ( .A(n33754), .B(\fmem_data[0][5] ), .ZN(n32563) );
  XNOR2_X1 U33710 ( .A(n36296), .B(\fmem_data[0][5] ), .ZN(n31469) );
  FA_X1 U33711 ( .A(n31472), .B(n31471), .CI(n31470), .CO(n31480), .S(n33674)
         );
  XNOR2_X1 U33712 ( .A(n34859), .B(\fmem_data[25][1] ), .ZN(n32148) );
  OAI22_X1 U33713 ( .A1(n31473), .A2(n34045), .B1(n34043), .B2(n3626), .ZN(
        n33890) );
  XNOR2_X1 U33714 ( .A(n33889), .B(n33890), .ZN(n31475) );
  XNOR2_X1 U33715 ( .A(n36110), .B(\fmem_data[25][5] ), .ZN(n31474) );
  XNOR2_X1 U33716 ( .A(n32078), .B(\fmem_data[25][5] ), .ZN(n34048) );
  OAI22_X1 U33717 ( .A1(n31474), .A2(n34985), .B1(n34048), .B2(n34986), .ZN(
        n33891) );
  XNOR2_X1 U33718 ( .A(n31475), .B(n33891), .ZN(n33675) );
  OAI21_X1 U33719 ( .B1(n33673), .B2(n33674), .A(n33675), .ZN(n31477) );
  NAND2_X1 U33720 ( .A1(n33674), .A2(n33673), .ZN(n31476) );
  NAND2_X1 U33721 ( .A1(n31477), .A2(n31476), .ZN(n33631) );
  FA_X1 U33722 ( .A(n31480), .B(n31479), .CI(n31478), .CO(n28406), .S(n33632)
         );
  XNOR2_X1 U33723 ( .A(n33631), .B(n33632), .ZN(n31485) );
  XNOR2_X1 U33724 ( .A(n31485), .B(n33630), .ZN(n33668) );
  FA_X1 U33725 ( .A(n31488), .B(n31487), .CI(n31486), .CO(n33672), .S(n33567)
         );
  XNOR2_X1 U33726 ( .A(n31489), .B(\fmem_data[21][1] ), .ZN(n34024) );
  INV_X1 U33727 ( .A(n33100), .ZN(n31490) );
  XNOR2_X1 U33728 ( .A(n32513), .B(\fmem_data[25][1] ), .ZN(n31500) );
  OR2_X1 U33729 ( .A1(n36313), .A2(n3657), .ZN(n31493) );
  OAI22_X1 U33730 ( .A1(n31493), .A2(n34533), .B1(n34429), .B2(n3657), .ZN(
        n33718) );
  FA_X1 U33731 ( .A(n31497), .B(n31496), .CI(n31495), .CO(n31605), .S(n33540)
         );
  INV_X1 U33732 ( .A(n32780), .ZN(n31498) );
  INV_X1 U33733 ( .A(n33059), .ZN(n31499) );
  OR2_X1 U33734 ( .A1(n33471), .A2(n33470), .ZN(n31501) );
  XNOR2_X1 U33735 ( .A(n32078), .B(\fmem_data[25][1] ), .ZN(n33449) );
  OAI22_X1 U33736 ( .A1(n33449), .A2(n34440), .B1(n31500), .B2(n3483), .ZN(
        n33473) );
  NAND2_X1 U33737 ( .A1(n31501), .A2(n33473), .ZN(n31503) );
  NAND2_X1 U33738 ( .A1(n33471), .A2(n33470), .ZN(n31502) );
  NAND2_X1 U33739 ( .A1(n31503), .A2(n31502), .ZN(n33490) );
  XNOR2_X1 U33740 ( .A(n31946), .B(\fmem_data[22][3] ), .ZN(n34417) );
  OAI22_X1 U33741 ( .A1(n31504), .A2(n34416), .B1(n34417), .B2(n34414), .ZN(
        n33491) );
  FA_X1 U33742 ( .A(n31510), .B(n31509), .CI(n31508), .CO(n33584), .S(n33563)
         );
  XNOR2_X1 U33743 ( .A(n32005), .B(\fmem_data[16][1] ), .ZN(n33557) );
  XNOR2_X1 U33744 ( .A(n32321), .B(\fmem_data[17][1] ), .ZN(n33834) );
  XNOR2_X1 U33745 ( .A(n33939), .B(\fmem_data[15][1] ), .ZN(n33480) );
  XNOR2_X1 U33746 ( .A(n3425), .B(\fmem_data[15][1] ), .ZN(n32598) );
  OAI21_X1 U33747 ( .B1(n33542), .B2(n33540), .A(n33541), .ZN(n31515) );
  NAND2_X1 U33748 ( .A1(n33542), .A2(n33540), .ZN(n31514) );
  NAND2_X1 U33749 ( .A1(n31515), .A2(n31514), .ZN(n33667) );
  INV_X1 U33750 ( .A(n33614), .ZN(n31599) );
  FA_X1 U33751 ( .A(n31518), .B(n31517), .CI(n31516), .CO(n31604), .S(n33536)
         );
  XNOR2_X1 U33752 ( .A(n31523), .B(n31522), .ZN(n31525) );
  XNOR2_X1 U33753 ( .A(n31525), .B(n31524), .ZN(n33438) );
  INV_X1 U33754 ( .A(n33873), .ZN(n31527) );
  INV_X1 U33755 ( .A(n33568), .ZN(n31528) );
  INV_X1 U33756 ( .A(n34431), .ZN(n31529) );
  XNOR2_X1 U33757 ( .A(n32235), .B(\fmem_data[12][1] ), .ZN(n34733) );
  FA_X1 U33758 ( .A(n31532), .B(n31531), .CI(n31530), .CO(n31613), .S(n33506)
         );
  XNOR2_X1 U33759 ( .A(n36112), .B(\fmem_data[12][3] ), .ZN(n31533) );
  INV_X1 U33760 ( .A(n33797), .ZN(n31534) );
  INV_X1 U33761 ( .A(n34537), .ZN(n31535) );
  INV_X1 U33762 ( .A(n34497), .ZN(n31536) );
  INV_X1 U33763 ( .A(n33596), .ZN(n31537) );
  INV_X1 U33764 ( .A(n34201), .ZN(n31538) );
  AND2_X1 U33765 ( .A1(n34615), .A2(n31538), .ZN(n34479) );
  XNOR2_X1 U33766 ( .A(n36244), .B(\fmem_data[14][3] ), .ZN(n31543) );
  XNOR2_X1 U33767 ( .A(n3376), .B(\fmem_data[11][1] ), .ZN(n32930) );
  XNOR2_X1 U33768 ( .A(n32023), .B(\fmem_data[11][1] ), .ZN(n33777) );
  OAI22_X1 U33769 ( .A1(n36196), .A2(n32930), .B1(n33777), .B2(n3577), .ZN(
        n33550) );
  OAI21_X1 U33770 ( .B1(n33548), .B2(n33547), .A(n33550), .ZN(n31546) );
  NAND2_X1 U33771 ( .A1(n33548), .A2(n33547), .ZN(n31545) );
  NAND2_X1 U33772 ( .A1(n31546), .A2(n31545), .ZN(n33504) );
  FA_X1 U33773 ( .A(n31549), .B(n31548), .CI(n31547), .CO(n31602), .S(n33477)
         );
  FA_X1 U33774 ( .A(n31552), .B(n31551), .CI(n31550), .CO(n31623), .S(n33476)
         );
  FA_X1 U33775 ( .A(n31555), .B(n31554), .CI(n31553), .CO(n31464), .S(n33533)
         );
  FA_X1 U33776 ( .A(n31558), .B(n31556), .CI(n31557), .CO(n31574), .S(n32995)
         );
  XNOR2_X1 U33777 ( .A(n31655), .B(\fmem_data[30][1] ), .ZN(n32573) );
  XNOR2_X1 U33778 ( .A(n32615), .B(\fmem_data[24][1] ), .ZN(n31910) );
  OAI21_X1 U33779 ( .B1(n32995), .B2(n32992), .A(n32993), .ZN(n31559) );
  NAND2_X1 U33780 ( .A1(n31560), .A2(n31559), .ZN(n33532) );
  FA_X1 U33781 ( .A(n31563), .B(n31562), .CI(n31561), .CO(n31550), .S(n33531)
         );
  FA_X1 U33782 ( .A(n31566), .B(n31565), .CI(n31564), .CO(n31552), .S(n33530)
         );
  FA_X1 U33783 ( .A(n31569), .B(n31567), .CI(n31568), .CO(n31618), .S(n33529)
         );
  FA_X1 U33784 ( .A(n31572), .B(n31571), .CI(n31570), .CO(n31619), .S(n33528)
         );
  FA_X1 U33785 ( .A(n31575), .B(n31574), .CI(n31573), .CO(n31441), .S(n33515)
         );
  FA_X1 U33786 ( .A(n31578), .B(n31577), .CI(n31576), .CO(n31620), .S(n33514)
         );
  XNOR2_X1 U33787 ( .A(n32898), .B(\fmem_data[8][3] ), .ZN(n33832) );
  XNOR2_X1 U33788 ( .A(n34626), .B(\fmem_data[8][3] ), .ZN(n31579) );
  OAI22_X1 U33789 ( .A1(n33832), .A2(n34206), .B1(n31579), .B2(n34208), .ZN(
        n33501) );
  INV_X1 U33790 ( .A(n33855), .ZN(n31580) );
  INV_X1 U33791 ( .A(n33681), .ZN(n31581) );
  INV_X1 U33792 ( .A(n33850), .ZN(n31582) );
  XNOR2_X1 U33793 ( .A(n31992), .B(\fmem_data[22][1] ), .ZN(n33810) );
  NOR2_X1 U33794 ( .A1(n31588), .A2(n3693), .ZN(n31584) );
  NOR2_X1 U33795 ( .A1(n31585), .A2(n3693), .ZN(n31583) );
  NOR2_X1 U33796 ( .A1(n31584), .A2(n31583), .ZN(n31590) );
  INV_X1 U33797 ( .A(n31585), .ZN(n31586) );
  NOR2_X1 U33798 ( .A1(n31586), .A2(\fmem_data[22][1] ), .ZN(n31587) );
  NAND2_X1 U33799 ( .A1(n31588), .A2(n31587), .ZN(n31589) );
  NAND2_X1 U33800 ( .A1(n31590), .A2(n31589), .ZN(n34776) );
  OR2_X1 U33801 ( .A1(n36299), .A2(n3627), .ZN(n31591) );
  OAI22_X1 U33802 ( .A1(n31591), .A2(n34501), .B1(n34499), .B2(n3627), .ZN(
        n33486) );
  OAI22_X1 U33803 ( .A1(n33580), .A2(n3575), .B1(n32928), .B2(n36120), .ZN(
        n33487) );
  XNOR2_X1 U33804 ( .A(n32131), .B(\fmem_data[4][1] ), .ZN(n32980) );
  OAI21_X1 U33805 ( .B1(n33486), .B2(n33487), .A(n33485), .ZN(n31594) );
  NAND2_X1 U33806 ( .A1(n31594), .A2(n31593), .ZN(n33441) );
  XNOR2_X1 U33807 ( .A(n31957), .B(\fmem_data[6][1] ), .ZN(n33812) );
  XNOR2_X1 U33808 ( .A(n32117), .B(\fmem_data[6][1] ), .ZN(n32883) );
  NOR2_X1 U33809 ( .A1(n33613), .A2(n33612), .ZN(n31598) );
  NAND2_X1 U33810 ( .A1(n33613), .A2(n33612), .ZN(n31597) );
  OAI21_X1 U33811 ( .B1(n31598), .B2(n31599), .A(n31597), .ZN(n33523) );
  XNOR2_X1 U33812 ( .A(n31601), .B(n31600), .ZN(n31603) );
  XNOR2_X1 U33813 ( .A(n31603), .B(n31602), .ZN(n33611) );
  FA_X1 U33814 ( .A(n31606), .B(n31605), .CI(n31604), .CO(n31433), .S(n33539)
         );
  FA_X1 U33815 ( .A(n31609), .B(n31608), .CI(n31607), .CO(n31549), .S(n33510)
         );
  FA_X1 U33816 ( .A(n31612), .B(n31611), .CI(n31610), .CO(n31551), .S(n33509)
         );
  FA_X1 U33817 ( .A(n31615), .B(n31614), .CI(n31613), .CO(n31547), .S(n33511)
         );
  OAI21_X1 U33818 ( .B1(n33509), .B2(n33510), .A(n33511), .ZN(n31617) );
  NAND2_X1 U33819 ( .A1(n33510), .A2(n33509), .ZN(n31616) );
  NAND2_X1 U33820 ( .A1(n31617), .A2(n31616), .ZN(n33538) );
  FA_X1 U33821 ( .A(n31620), .B(n31619), .CI(n31618), .CO(n31621), .S(n33537)
         );
  FA_X1 U33822 ( .A(n31623), .B(n31622), .CI(n31621), .CO(n31630), .S(n33609)
         );
  XNOR2_X1 U33823 ( .A(n31625), .B(n31624), .ZN(n31627) );
  XNOR2_X1 U33824 ( .A(n31627), .B(n31626), .ZN(n33619) );
  FA_X1 U33825 ( .A(n31630), .B(n31629), .CI(n31628), .CO(n31428), .S(n33618)
         );
  OAI21_X1 U33826 ( .B1(n33406), .B2(n33405), .A(n33407), .ZN(n31632) );
  NAND2_X1 U33827 ( .A1(n33406), .A2(n33405), .ZN(n31631) );
  NAND2_X1 U33828 ( .A1(n31632), .A2(n31631), .ZN(n35454) );
  OAI21_X1 U33829 ( .B1(n31635), .B2(n31634), .A(n31633), .ZN(n31637) );
  NAND2_X1 U33830 ( .A1(n31635), .A2(n31634), .ZN(n31636) );
  NAND2_X1 U33831 ( .A1(n31637), .A2(n31636), .ZN(n35434) );
  XNOR2_X1 U33832 ( .A(n35240), .B(\fmem_data[3][5] ), .ZN(n34917) );
  XNOR2_X1 U33833 ( .A(n32188), .B(\fmem_data[3][5] ), .ZN(n33029) );
  OAI22_X1 U33834 ( .A1(n34917), .A2(n34919), .B1(n33029), .B2(n34918), .ZN(
        n31707) );
  XNOR2_X1 U33835 ( .A(n35238), .B(\fmem_data[11][5] ), .ZN(n34931) );
  XNOR2_X1 U33836 ( .A(n35112), .B(\fmem_data[11][5] ), .ZN(n31978) );
  OAI22_X1 U33837 ( .A1(n34931), .A2(n34932), .B1(n31978), .B2(n34933), .ZN(
        n31711) );
  AOI21_X1 U33838 ( .B1(n31645), .B2(n31646), .A(n31644), .ZN(n31648) );
  NOR2_X1 U33839 ( .A1(n31646), .A2(n31645), .ZN(n31647) );
  NOR2_X1 U33840 ( .A1(n31648), .A2(n31647), .ZN(n31710) );
  FA_X1 U33841 ( .A(n31651), .B(n31650), .CI(n31649), .CO(n31729), .S(n30813)
         );
  FA_X1 U33842 ( .A(n31654), .B(n31653), .CI(n31652), .CO(n31728), .S(n31731)
         );
  XNOR2_X1 U33843 ( .A(n31657), .B(\fmem_data[28][7] ), .ZN(n35400) );
  XNOR2_X1 U33844 ( .A(n31895), .B(\fmem_data[4][7] ), .ZN(n33306) );
  XNOR2_X1 U33845 ( .A(n31663), .B(\fmem_data[12][7] ), .ZN(n35123) );
  XNOR2_X1 U33846 ( .A(n35355), .B(\fmem_data[10][5] ), .ZN(n35087) );
  XNOR2_X1 U33847 ( .A(n35140), .B(\fmem_data[7][5] ), .ZN(n33028) );
  XNOR2_X1 U33848 ( .A(n35359), .B(\fmem_data[7][5] ), .ZN(n34837) );
  OAI22_X1 U33849 ( .A1(n33028), .A2(n34836), .B1(n34835), .B2(n34837), .ZN(
        n31699) );
  XNOR2_X1 U33850 ( .A(n35405), .B(\fmem_data[5][5] ), .ZN(n33310) );
  AOI21_X1 U33851 ( .B1(n33859), .B2(n33857), .A(n33310), .ZN(n31667) );
  XNOR2_X1 U33852 ( .A(n31669), .B(\fmem_data[13][7] ), .ZN(n35105) );
  XNOR2_X1 U33853 ( .A(n31670), .B(\fmem_data[26][7] ), .ZN(n35107) );
  OAI22_X1 U33854 ( .A1(n31671), .A2(n35711), .B1(n35107), .B2(n35712), .ZN(
        n35119) );
  XNOR2_X1 U33855 ( .A(n3371), .B(\fmem_data[18][7] ), .ZN(n31819) );
  XNOR2_X1 U33856 ( .A(n3356), .B(\fmem_data[18][7] ), .ZN(n35109) );
  XNOR2_X1 U33857 ( .A(n35397), .B(\fmem_data[16][5] ), .ZN(n33329) );
  XNOR2_X1 U33858 ( .A(n35399), .B(\fmem_data[28][5] ), .ZN(n33323) );
  FA_X1 U33859 ( .A(n31677), .B(n31678), .CI(n31679), .CO(n35407), .S(n31790)
         );
  OAI21_X1 U33860 ( .B1(n31682), .B2(n31681), .A(n31680), .ZN(n31684) );
  NAND2_X1 U33861 ( .A1(n31682), .A2(n31681), .ZN(n31683) );
  NAND2_X1 U33862 ( .A1(n31684), .A2(n31683), .ZN(n31749) );
  FA_X1 U33863 ( .A(n3492), .B(n31685), .CI(n3728), .CO(n31748), .S(n31928) );
  FA_X1 U33864 ( .A(n31688), .B(n31687), .CI(n31686), .CO(n31747), .S(n31724)
         );
  OAI21_X1 U33865 ( .B1(n31695), .B2(n31696), .A(n31694), .ZN(n31698) );
  NAND2_X1 U33866 ( .A1(n31698), .A2(n31697), .ZN(n31720) );
  FA_X1 U33867 ( .A(n31701), .B(n31700), .CI(n31699), .CO(n35253), .S(n31721)
         );
  OAI21_X1 U33868 ( .B1(n31722), .B2(n31720), .A(n31721), .ZN(n31703) );
  NAND2_X1 U33869 ( .A1(n31722), .A2(n31720), .ZN(n31702) );
  NAND2_X1 U33870 ( .A1(n31703), .A2(n31702), .ZN(n35292) );
  XNOR2_X1 U33871 ( .A(n35293), .B(n35292), .ZN(n31713) );
  AOI21_X1 U33872 ( .B1(n33643), .B2(n33642), .A(n33385), .ZN(n31706) );
  FA_X1 U33873 ( .A(n31709), .B(n31708), .CI(n31707), .CO(n35311), .S(n31746)
         );
  FA_X1 U33874 ( .A(n31712), .B(n31710), .CI(n31711), .CO(n35310), .S(n31745)
         );
  XNOR2_X1 U33875 ( .A(n31713), .B(n35291), .ZN(n35300) );
  OAI21_X1 U33876 ( .B1(n31719), .B2(n31718), .A(n31717), .ZN(n35299) );
  XNOR2_X1 U33877 ( .A(n31721), .B(n31720), .ZN(n31723) );
  XNOR2_X1 U33878 ( .A(n31723), .B(n31722), .ZN(n35055) );
  FA_X1 U33879 ( .A(n31726), .B(n31725), .CI(n31724), .CO(n35054), .S(n32038)
         );
  FA_X1 U33880 ( .A(n31729), .B(n31728), .CI(n31727), .CO(n31744), .S(n31755)
         );
  FA_X1 U33881 ( .A(n31732), .B(n31731), .CI(n31730), .CO(n31754), .S(n31860)
         );
  FA_X1 U33882 ( .A(n31735), .B(n31734), .CI(n31733), .CO(n31680), .S(n31865)
         );
  OAI21_X1 U33883 ( .B1(n31738), .B2(n31737), .A(n31736), .ZN(n31740) );
  NAND2_X1 U33884 ( .A1(n31738), .A2(n31737), .ZN(n31739) );
  NAND2_X1 U33885 ( .A1(n31740), .A2(n31739), .ZN(n31864) );
  FA_X1 U33886 ( .A(n31743), .B(n31742), .CI(n31741), .CO(n31863), .S(n31154)
         );
  FA_X1 U33887 ( .A(n31746), .B(n31745), .CI(n31744), .CO(n35309), .S(n35049)
         );
  FA_X1 U33888 ( .A(n31749), .B(n31748), .CI(n31747), .CO(n35293), .S(n35048)
         );
  FA_X1 U33889 ( .A(n31752), .B(n31751), .CI(n31750), .CO(n35047), .S(n32039)
         );
  FA_X1 U33890 ( .A(n31755), .B(n31754), .CI(n31753), .CO(n35053), .S(n31857)
         );
  XNOR2_X1 U33891 ( .A(n31757), .B(n31756), .ZN(n31759) );
  XNOR2_X1 U33892 ( .A(n31759), .B(n31758), .ZN(n31856) );
  FA_X1 U33893 ( .A(n31761), .B(n31762), .CI(n31760), .CO(n31855), .S(n32277)
         );
  OAI21_X1 U33894 ( .B1(n31857), .B2(n31856), .A(n31855), .ZN(n31764) );
  NAND2_X1 U33895 ( .A1(n31764), .A2(n31763), .ZN(n32048) );
  OAI21_X1 U33896 ( .B1(n32050), .B2(n32049), .A(n32048), .ZN(n31766) );
  NAND2_X1 U33897 ( .A1(n32050), .A2(n32049), .ZN(n31765) );
  NAND2_X1 U33898 ( .A1(n31766), .A2(n31765), .ZN(n35428) );
  OAI21_X1 U33899 ( .B1(n31768), .B2(n31769), .A(n31767), .ZN(n31771) );
  NAND2_X1 U33900 ( .A1(n31771), .A2(n31770), .ZN(n35427) );
  XNOR2_X1 U33901 ( .A(n35434), .B(n35435), .ZN(n31854) );
  NAND2_X1 U33902 ( .A1(n31774), .A2(n31773), .ZN(n31776) );
  OAI21_X1 U33903 ( .B1(n31774), .B2(n31773), .A(n31772), .ZN(n31775) );
  NAND2_X1 U33904 ( .A1(n31776), .A2(n31775), .ZN(n35432) );
  FA_X1 U33905 ( .A(n31778), .B(n31779), .CI(n31777), .CO(n35350), .S(n31786)
         );
  FA_X1 U33906 ( .A(n31782), .B(n31780), .CI(n31781), .CO(n35349), .S(n31794)
         );
  FA_X1 U33907 ( .A(n31785), .B(n31784), .CI(n31783), .CO(n35348), .S(n31805)
         );
  FA_X1 U33908 ( .A(n31788), .B(n31787), .CI(n31786), .CO(n35416), .S(n31812)
         );
  FA_X1 U33909 ( .A(n31789), .B(n31791), .CI(n31790), .CO(n35415), .S(n31811)
         );
  FA_X1 U33910 ( .A(n31794), .B(n31793), .CI(n31792), .CO(n35420), .S(n31847)
         );
  FA_X1 U33911 ( .A(n31797), .B(n31796), .CI(n31795), .CO(n35347), .S(n31788)
         );
  XNOR2_X1 U33912 ( .A(n31800), .B(\fmem_data[29][7] ), .ZN(n35358) );
  XNOR2_X1 U33913 ( .A(n35120), .B(\fmem_data[6][5] ), .ZN(n33368) );
  XNOR2_X1 U33914 ( .A(n35403), .B(\fmem_data[21][5] ), .ZN(n33304) );
  AOI21_X1 U33915 ( .B1(n34195), .B2(n34194), .A(n33304), .ZN(n31802) );
  INV_X1 U33916 ( .A(n31802), .ZN(n35344) );
  XNOR2_X1 U33917 ( .A(n35395), .B(\fmem_data[24][5] ), .ZN(n33371) );
  OAI21_X1 U33918 ( .B1(n31807), .B2(n31806), .A(n31805), .ZN(n31809) );
  NAND2_X1 U33919 ( .A1(n31809), .A2(n31808), .ZN(n35418) );
  FA_X1 U33920 ( .A(n31812), .B(n31811), .CI(n31810), .CO(n35421), .S(n31773)
         );
  XNOR2_X1 U33921 ( .A(n35102), .B(\fmem_data[14][5] ), .ZN(n33101) );
  AOI21_X1 U33922 ( .B1(n33100), .B2(n33098), .A(n33101), .ZN(n31814) );
  XNOR2_X1 U33923 ( .A(n32188), .B(\fmem_data[3][7] ), .ZN(n35241) );
  OAI22_X1 U33924 ( .A1(n31815), .A2(n35637), .B1(n35241), .B2(n35638), .ZN(
        n35161) );
  XNOR2_X1 U33925 ( .A(n33214), .B(\fmem_data[24][7] ), .ZN(n35396) );
  XNOR2_X1 U33926 ( .A(n31818), .B(\fmem_data[19][7] ), .ZN(n33134) );
  OAI22_X1 U33927 ( .A1(n35271), .A2(n35656), .B1(n33134), .B2(n35655), .ZN(
        n35165) );
  OAI22_X1 U33928 ( .A1(n31820), .A2(n35704), .B1(n35705), .B2(n31819), .ZN(
        n34866) );
  XNOR2_X1 U33929 ( .A(n35108), .B(\fmem_data[18][5] ), .ZN(n35008) );
  OAI22_X1 U33930 ( .A1(n35008), .A2(n35006), .B1(n31821), .B2(n35007), .ZN(
        n34865) );
  XNOR2_X1 U33931 ( .A(n35324), .B(\fmem_data[4][5] ), .ZN(n35009) );
  OAI22_X1 U33932 ( .A1(n35009), .A2(n35011), .B1(n31822), .B2(n35010), .ZN(
        n34864) );
  XNOR2_X1 U33933 ( .A(n33039), .B(\fmem_data[0][7] ), .ZN(n35402) );
  XNOR2_X1 U33934 ( .A(n35340), .B(\fmem_data[20][5] ), .ZN(n35038) );
  XNOR2_X1 U33935 ( .A(n35178), .B(\fmem_data[20][5] ), .ZN(n33252) );
  OAI22_X1 U33936 ( .A1(n35036), .A2(n35038), .B1(n33252), .B2(n35037), .ZN(
        n34883) );
  XNOR2_X1 U33937 ( .A(n35326), .B(\fmem_data[25][5] ), .ZN(n34984) );
  FA_X1 U33938 ( .A(n31829), .B(n31830), .CI(n31828), .CO(n35124), .S(n35175)
         );
  AOI21_X1 U33939 ( .B1(n33963), .B2(n33961), .A(n33130), .ZN(n31831) );
  INV_X1 U33940 ( .A(n31831), .ZN(n35126) );
  FA_X1 U33941 ( .A(n31835), .B(n31834), .CI(n31833), .CO(n35411), .S(n31844)
         );
  XNOR2_X1 U33942 ( .A(n35410), .B(n35411), .ZN(n31842) );
  NOR2_X1 U33943 ( .A1(n31838), .A2(n31837), .ZN(n31841) );
  OAI21_X1 U33944 ( .B1(n31841), .B2(n31840), .A(n31839), .ZN(n35412) );
  XNOR2_X1 U33945 ( .A(n31842), .B(n35412), .ZN(n35190) );
  FA_X1 U33946 ( .A(n31845), .B(n31844), .CI(n31843), .CO(n35189), .S(n31853)
         );
  OAI21_X1 U33947 ( .B1(n31848), .B2(n31847), .A(n31846), .ZN(n31850) );
  NAND2_X1 U33948 ( .A1(n31848), .A2(n31847), .ZN(n31849) );
  NAND2_X1 U33949 ( .A1(n31850), .A2(n31849), .ZN(n35425) );
  FA_X1 U33950 ( .A(n31853), .B(n31852), .CI(n31851), .CO(n35424), .S(n35216)
         );
  XNOR2_X1 U33951 ( .A(n31854), .B(n35433), .ZN(n35455) );
  XNOR2_X1 U33952 ( .A(n31856), .B(n31855), .ZN(n31858) );
  XNOR2_X1 U33953 ( .A(n31858), .B(n31857), .ZN(n32462) );
  XNOR2_X1 U33954 ( .A(n31860), .B(n31859), .ZN(n31862) );
  XNOR2_X1 U33955 ( .A(n31862), .B(n31861), .ZN(n32471) );
  FA_X1 U33956 ( .A(n31865), .B(n31864), .CI(n31863), .CO(n31753), .S(n31926)
         );
  XNOR2_X1 U33957 ( .A(n31867), .B(n31866), .ZN(n31869) );
  XNOR2_X1 U33958 ( .A(n31869), .B(n31868), .ZN(n31925) );
  FA_X1 U33959 ( .A(n31872), .B(n31871), .CI(n31870), .CO(n31924), .S(n32099)
         );
  FA_X1 U33960 ( .A(n31875), .B(n31874), .CI(n31873), .CO(n31859), .S(n32498)
         );
  XNOR2_X1 U33961 ( .A(n31877), .B(n31876), .ZN(n31879) );
  XNOR2_X1 U33962 ( .A(n31879), .B(n31878), .ZN(n32094) );
  XNOR2_X1 U33963 ( .A(n31882), .B(\fmem_data[21][1] ), .ZN(n34023) );
  OAI22_X1 U33964 ( .A1(n34023), .A2(n34613), .B1(n31883), .B2(n3570), .ZN(
        n31906) );
  OAI22_X1 U33965 ( .A1(n33860), .A2(n33857), .B1(n31884), .B2(n33859), .ZN(
        n31905) );
  XNOR2_X1 U33966 ( .A(n31885), .B(\fmem_data[5][1] ), .ZN(n34021) );
  OAI22_X1 U33967 ( .A1(n34021), .A2(n34483), .B1(n31886), .B2(n3576), .ZN(
        n31904) );
  FA_X1 U33968 ( .A(n31891), .B(n31890), .CI(n31889), .CO(n31182), .S(n32092)
         );
  XNOR2_X1 U33969 ( .A(n35280), .B(\fmem_data[1][1] ), .ZN(n34078) );
  XNOR2_X1 U33970 ( .A(n31893), .B(\fmem_data[27][3] ), .ZN(n33995) );
  OAI22_X1 U33971 ( .A1(n31894), .A2(n34463), .B1(n34462), .B2(n33995), .ZN(
        n32157) );
  XNOR2_X1 U33972 ( .A(n31895), .B(\fmem_data[4][1] ), .ZN(n32585) );
  OAI22_X1 U33973 ( .A1(n31896), .A2(n3569), .B1(n32585), .B2(n34598), .ZN(
        n31903) );
  XNOR2_X1 U33974 ( .A(n31897), .B(\fmem_data[28][3] ), .ZN(n33856) );
  OAI22_X1 U33975 ( .A1(n33856), .A2(n33853), .B1(n31898), .B2(n33855), .ZN(
        n31902) );
  XNOR2_X1 U33976 ( .A(n31900), .B(\fmem_data[20][3] ), .ZN(n32517) );
  OAI22_X1 U33977 ( .A1(n32128), .A2(n34495), .B1(n32517), .B2(n34497), .ZN(
        n31901) );
  FA_X1 U33978 ( .A(n31903), .B(n31902), .CI(n31901), .CO(n32156), .S(n32267)
         );
  FA_X1 U33979 ( .A(n31906), .B(n31905), .CI(n31904), .CO(n32160), .S(n32266)
         );
  FA_X1 U33980 ( .A(n31909), .B(n31908), .CI(n31907), .CO(n31889), .S(n32265)
         );
  XNOR2_X1 U33981 ( .A(n32442), .B(\fmem_data[1][3] ), .ZN(n33993) );
  OAI22_X1 U33982 ( .A1(n32594), .A2(n34466), .B1(n33993), .B2(n34779), .ZN(
        n32486) );
  XNOR2_X1 U33983 ( .A(n31914), .B(n31913), .ZN(n31916) );
  XNOR2_X1 U33984 ( .A(n31916), .B(n31915), .ZN(n32481) );
  FA_X1 U33985 ( .A(n31919), .B(n31918), .CI(n31917), .CO(n32480), .S(n33433)
         );
  OAI21_X1 U33986 ( .B1(n32089), .B2(n32088), .A(n32090), .ZN(n31921) );
  NAND2_X1 U33987 ( .A1(n31921), .A2(n31920), .ZN(n32496) );
  OAI21_X1 U33988 ( .B1(n32469), .B2(n32471), .A(n32470), .ZN(n31922) );
  NAND2_X1 U33989 ( .A1(n31923), .A2(n31922), .ZN(n32463) );
  FA_X1 U33990 ( .A(n31926), .B(n31925), .CI(n31924), .CO(n32044), .S(n32469)
         );
  FA_X1 U33991 ( .A(n31929), .B(n31928), .CI(n31927), .CO(n31716), .S(n32043)
         );
  XNOR2_X1 U33992 ( .A(n32044), .B(n32043), .ZN(n31933) );
  FA_X1 U33993 ( .A(n31932), .B(n31931), .CI(n31930), .CO(n32042), .S(n32276)
         );
  XNOR2_X1 U33994 ( .A(n31933), .B(n32042), .ZN(n32465) );
  OAI21_X1 U33995 ( .B1(n32462), .B2(n32463), .A(n32465), .ZN(n31935) );
  NAND2_X1 U33996 ( .A1(n32462), .A2(n32463), .ZN(n31934) );
  NAND2_X1 U33997 ( .A1(n31935), .A2(n31934), .ZN(n35063) );
  OAI22_X1 U33998 ( .A1(n31937), .A2(n35641), .B1(n31936), .B2(n35642), .ZN(
        n33112) );
  OAI22_X1 U33999 ( .A1(n31939), .A2(n35618), .B1(n31938), .B2(n35619), .ZN(
        n33111) );
  OAI22_X1 U34000 ( .A1(n34235), .A2(n34908), .B1(n31941), .B2(n34909), .ZN(
        n33110) );
  OAI22_X1 U34001 ( .A1(n31945), .A2(n33603), .B1(n31944), .B2(n33741), .ZN(
        n32300) );
  XNOR2_X1 U34002 ( .A(n31946), .B(\fmem_data[22][7] ), .ZN(n34102) );
  OAI22_X1 U34003 ( .A1(n34102), .A2(n35584), .B1(n31947), .B2(n35585), .ZN(
        n32299) );
  OAI22_X1 U34004 ( .A1(n31949), .A2(n33690), .B1(n31948), .B2(n34736), .ZN(
        n32711) );
  XNOR2_X1 U34005 ( .A(n34630), .B(\fmem_data[14][7] ), .ZN(n34097) );
  OAI22_X1 U34006 ( .A1(n34097), .A2(n35576), .B1(n31952), .B2(n35577), .ZN(
        n32709) );
  INV_X1 U34007 ( .A(n31956), .ZN(n32186) );
  INV_X1 U34008 ( .A(n31960), .ZN(n32184) );
  FA_X1 U34009 ( .A(n31963), .B(n31962), .CI(n31961), .CO(n31691), .S(n32352)
         );
  INV_X1 U34010 ( .A(n31967), .ZN(n32172) );
  AOI21_X1 U34011 ( .B1(n34483), .B2(n3576), .A(n31968), .ZN(n31969) );
  XNOR2_X1 U34012 ( .A(n32727), .B(\fmem_data[19][7] ), .ZN(n33135) );
  OAI22_X1 U34013 ( .A1(n31979), .A2(n34933), .B1(n34932), .B2(n31978), .ZN(
        n33107) );
  OAI22_X1 U34014 ( .A1(n33168), .A2(n34904), .B1(n31981), .B2(n34903), .ZN(
        n33125) );
  OAI22_X1 U34015 ( .A1(n31983), .A2(n35637), .B1(n31982), .B2(n35638), .ZN(
        n33124) );
  OAI22_X1 U34016 ( .A1(n31987), .A2(n35037), .B1(n31986), .B2(n35036), .ZN(
        n32649) );
  OAI22_X1 U34017 ( .A1(n31989), .A2(n35581), .B1(n35580), .B2(n31988), .ZN(
        n32648) );
  AOI21_X1 U34018 ( .B1(n3573), .B2(n36298), .A(n31990), .ZN(n31991) );
  INV_X1 U34019 ( .A(n31991), .ZN(n32647) );
  XNOR2_X1 U34020 ( .A(n31996), .B(\fmem_data[8][3] ), .ZN(n33061) );
  OAI22_X1 U34021 ( .A1(n31998), .A2(n34437), .B1(n31997), .B2(n34435), .ZN(
        n33074) );
  OAI22_X1 U34022 ( .A1(n35088), .A2(n32000), .B1(n31999), .B2(n35089), .ZN(
        n33073) );
  OAI22_X1 U34023 ( .A1(n32004), .A2(n34414), .B1(n32003), .B2(n34416), .ZN(
        n32521) );
  FA_X1 U34024 ( .A(n32011), .B(n32010), .CI(n32009), .CO(n33024), .S(n32721)
         );
  OAI22_X1 U34025 ( .A1(n32013), .A2(n34497), .B1(n32012), .B2(n34495), .ZN(
        n33023) );
  XNOR2_X1 U34026 ( .A(n32014), .B(\fmem_data[2][3] ), .ZN(n32642) );
  OAI22_X1 U34027 ( .A1(n33796), .A2(n32642), .B1(n32015), .B2(n33797), .ZN(
        n33022) );
  OAI22_X1 U34028 ( .A1(n32019), .A2(n35722), .B1(n35721), .B2(n32018), .ZN(
        n33049) );
  XNOR2_X1 U34029 ( .A(n32554), .B(\fmem_data[26][7] ), .ZN(n34033) );
  XNOR2_X1 U34030 ( .A(n32023), .B(\fmem_data[11][5] ), .ZN(n33971) );
  OAI22_X1 U34031 ( .A1(n32024), .A2(n34932), .B1(n33971), .B2(n34933), .ZN(
        n32360) );
  OAI22_X1 U34032 ( .A1(n33976), .A2(n33973), .B1(n32026), .B2(n33975), .ZN(
        n32358) );
  INV_X1 U34033 ( .A(n32358), .ZN(n32031) );
  INV_X1 U34034 ( .A(n36100), .ZN(n32027) );
  NOR2_X1 U34035 ( .A1(n32027), .A2(\fmem_data[24][0] ), .ZN(n32028) );
  OR2_X1 U34036 ( .A1(n32029), .A2(n32028), .ZN(n32357) );
  INV_X1 U34037 ( .A(n32357), .ZN(n32030) );
  NAND2_X1 U34038 ( .A1(n32031), .A2(n32030), .ZN(n32032) );
  NAND2_X1 U34039 ( .A1(n32360), .A2(n32032), .ZN(n32034) );
  NAND2_X1 U34040 ( .A1(n32034), .A2(n32033), .ZN(n33220) );
  OAI21_X1 U34041 ( .B1(n32039), .B2(n32038), .A(n32037), .ZN(n32041) );
  NAND2_X1 U34042 ( .A1(n32039), .A2(n32038), .ZN(n32040) );
  NAND2_X1 U34043 ( .A1(n32041), .A2(n32040), .ZN(n34971) );
  XNOR2_X1 U34044 ( .A(n34970), .B(n34971), .ZN(n32047) );
  NAND2_X1 U34045 ( .A1(n32046), .A2(n32045), .ZN(n34969) );
  XNOR2_X1 U34046 ( .A(n32047), .B(n34969), .ZN(n35062) );
  XNOR2_X1 U34047 ( .A(n35063), .B(n35062), .ZN(n32052) );
  XNOR2_X1 U34048 ( .A(n32049), .B(n32048), .ZN(n32051) );
  XNOR2_X1 U34049 ( .A(n32051), .B(n32050), .ZN(n35064) );
  XNOR2_X1 U34050 ( .A(n32052), .B(n35064), .ZN(n33404) );
  FA_X1 U34051 ( .A(n32055), .B(n32054), .CI(n32053), .CO(n32474), .S(n33003)
         );
  XNOR2_X1 U34052 ( .A(n3295), .B(\fmem_data[13][1] ), .ZN(n34741) );
  OAI22_X1 U34053 ( .A1(n32056), .A2(n3571), .B1(n34741), .B2(n34742), .ZN(
        n32967) );
  OR2_X1 U34054 ( .A1(n32059), .A2(n3647), .ZN(n32061) );
  XNOR2_X1 U34055 ( .A(n32127), .B(\fmem_data[20][1] ), .ZN(n33552) );
  OR2_X1 U34056 ( .A1(n33552), .A2(n36227), .ZN(n32060) );
  NAND2_X1 U34057 ( .A1(n32061), .A2(n32060), .ZN(n32965) );
  OAI21_X1 U34058 ( .B1(n32967), .B2(n32966), .A(n32965), .ZN(n32063) );
  NAND2_X1 U34059 ( .A1(n32063), .A2(n32062), .ZN(n32945) );
  XNOR2_X1 U34060 ( .A(n32064), .B(\fmem_data[0][1] ), .ZN(n33578) );
  OAI22_X1 U34061 ( .A1(n33578), .A2(n3564), .B1(n33755), .B2(n36295), .ZN(
        n32935) );
  OAI22_X1 U34062 ( .A1(n32067), .A2(n34201), .B1(n32066), .B2(n34199), .ZN(
        n32934) );
  XNOR2_X1 U34063 ( .A(n33749), .B(\fmem_data[13][3] ), .ZN(n33571) );
  OAI21_X1 U34064 ( .B1(n32945), .B2(n32944), .A(n32946), .ZN(n32074) );
  NAND2_X1 U34065 ( .A1(n32074), .A2(n32073), .ZN(n32927) );
  INV_X1 U34066 ( .A(n34986), .ZN(n32076) );
  INV_X1 U34067 ( .A(n35034), .ZN(n32077) );
  XNOR2_X1 U34068 ( .A(n32078), .B(\fmem_data[25][3] ), .ZN(n32606) );
  OAI22_X1 U34069 ( .A1(n32606), .A2(n33057), .B1(n32079), .B2(n33059), .ZN(
        n32414) );
  FA_X1 U34070 ( .A(n32084), .B(n32083), .CI(n32082), .CO(n32485), .S(n32925)
         );
  FA_X1 U34071 ( .A(n32087), .B(n32086), .CI(n32085), .CO(n32477), .S(n33001)
         );
  INV_X1 U34072 ( .A(n32920), .ZN(n32097) );
  XNOR2_X1 U34073 ( .A(n32089), .B(n32088), .ZN(n32091) );
  XNOR2_X1 U34074 ( .A(n32091), .B(n32090), .ZN(n32919) );
  FA_X1 U34075 ( .A(n32094), .B(n32093), .CI(n32092), .CO(n32497), .S(n32918)
         );
  NOR2_X1 U34076 ( .A1(n32919), .A2(n32918), .ZN(n32096) );
  OAI21_X1 U34077 ( .B1(n32097), .B2(n32096), .A(n32095), .ZN(n32913) );
  FA_X1 U34078 ( .A(n32100), .B(n32099), .CI(n32098), .CO(n32275), .S(n32912)
         );
  FA_X1 U34079 ( .A(n32103), .B(n32102), .CI(n32101), .CO(n32467), .S(n32911)
         );
  OAI21_X1 U34080 ( .B1(n32913), .B2(n32912), .A(n32911), .ZN(n32105) );
  NAND2_X1 U34081 ( .A1(n32913), .A2(n32912), .ZN(n32104) );
  NAND2_X1 U34082 ( .A1(n32105), .A2(n32104), .ZN(n33006) );
  XNOR2_X1 U34083 ( .A(n3313), .B(\fmem_data[7][5] ), .ZN(n34071) );
  OAI22_X1 U34084 ( .A1(n32107), .A2(n34835), .B1(n34071), .B2(n34836), .ZN(
        n32315) );
  XNOR2_X1 U34085 ( .A(n36339), .B(\fmem_data[15][7] ), .ZN(n32109) );
  OAI22_X1 U34086 ( .A1(n32109), .A2(n35696), .B1(n32108), .B2(n35697), .ZN(
        n32314) );
  XNOR2_X1 U34087 ( .A(n3320), .B(\fmem_data[31][3] ), .ZN(n33906) );
  OAI22_X1 U34088 ( .A1(n32111), .A2(n34470), .B1(n33906), .B2(n34468), .ZN(
        n32303) );
  XNOR2_X1 U34089 ( .A(n35112), .B(\fmem_data[11][1] ), .ZN(n33945) );
  OAI22_X1 U34090 ( .A1(n32112), .A2(n3577), .B1(n33945), .B2(n36196), .ZN(
        n32302) );
  INV_X1 U34091 ( .A(n35585), .ZN(n32113) );
  INV_X1 U34092 ( .A(n35577), .ZN(n32114) );
  XNOR2_X1 U34093 ( .A(n32117), .B(\fmem_data[6][3] ), .ZN(n33597) );
  OAI22_X1 U34094 ( .A1(n32118), .A2(n33596), .B1(n33597), .B2(n33598), .ZN(
        n32684) );
  INV_X1 U34095 ( .A(n33828), .ZN(n32119) );
  INV_X1 U34096 ( .A(n33859), .ZN(n32121) );
  XNOR2_X1 U34097 ( .A(n32124), .B(\fmem_data[22][3] ), .ZN(n34415) );
  OAI22_X1 U34098 ( .A1(n32126), .A2(n3574), .B1(n32428), .B2(n34625), .ZN(
        n32797) );
  XNOR2_X1 U34099 ( .A(n32131), .B(\fmem_data[4][3] ), .ZN(n32689) );
  XNOR2_X1 U34100 ( .A(n36337), .B(\fmem_data[19][7] ), .ZN(n32138) );
  OAI22_X1 U34101 ( .A1(n32138), .A2(n35655), .B1(n32137), .B2(n35656), .ZN(
        n32632) );
  XNOR2_X1 U34102 ( .A(n33743), .B(\fmem_data[9][5] ), .ZN(n32227) );
  OR2_X1 U34103 ( .A1(n36316), .A2(n3698), .ZN(n32140) );
  XNOR2_X1 U34104 ( .A(n3116), .B(\fmem_data[23][7] ), .ZN(n32142) );
  OAI22_X1 U34105 ( .A1(n32142), .A2(n35651), .B1(n32141), .B2(n35652), .ZN(
        n32201) );
  OAI22_X1 U34106 ( .A1(n32144), .A2(n32779), .B1(n32143), .B2(n32780), .ZN(
        n32661) );
  XNOR2_X1 U34107 ( .A(n32145), .B(\fmem_data[18][1] ), .ZN(n33793) );
  OAI22_X1 U34108 ( .A1(n33793), .A2(n36104), .B1(n32146), .B2(n3580), .ZN(
        n32660) );
  OAI22_X1 U34109 ( .A1(n32148), .A2(n34440), .B1(n3483), .B2(n32147), .ZN(
        n32659) );
  OAI22_X1 U34110 ( .A1(n32150), .A2(n34909), .B1(n32149), .B2(n34908), .ZN(
        n32199) );
  OR2_X1 U34111 ( .A1(n3116), .A2(n3668), .ZN(n32155) );
  XNOR2_X1 U34112 ( .A(n32808), .B(n32807), .ZN(n32170) );
  FA_X1 U34113 ( .A(n32158), .B(n32157), .CI(n32156), .CO(n32339), .S(n32089)
         );
  FA_X1 U34114 ( .A(n32161), .B(n32160), .CI(n32159), .CO(n32337), .S(n32093)
         );
  XNOR2_X1 U34115 ( .A(n32163), .B(\fmem_data[26][1] ), .ZN(n33641) );
  OAI22_X1 U34116 ( .A1(n33641), .A2(n33725), .B1(n3678), .B2(n32164), .ZN(
        n32611) );
  XNOR2_X1 U34117 ( .A(n32165), .B(\fmem_data[2][3] ), .ZN(n33798) );
  OAI22_X1 U34118 ( .A1(n33798), .A2(n33796), .B1(n32166), .B2(n33797), .ZN(
        n32610) );
  XNOR2_X1 U34119 ( .A(n34862), .B(\fmem_data[16][1] ), .ZN(n34026) );
  OAI22_X1 U34120 ( .A1(n34026), .A2(n36298), .B1(n32167), .B2(n3573), .ZN(
        n32609) );
  XNOR2_X1 U34121 ( .A(n35145), .B(\fmem_data[27][1] ), .ZN(n34189) );
  XNOR2_X1 U34122 ( .A(n32337), .B(n32338), .ZN(n32169) );
  XNOR2_X1 U34123 ( .A(n32339), .B(n32169), .ZN(n32806) );
  XNOR2_X1 U34124 ( .A(n32170), .B(n32806), .ZN(n32917) );
  FA_X1 U34125 ( .A(n32173), .B(n32172), .CI(n32171), .CO(n32351), .S(n32356)
         );
  XNOR2_X1 U34126 ( .A(n32174), .B(\fmem_data[7][3] ), .ZN(n33991) );
  OAI22_X1 U34127 ( .A1(n32175), .A2(n34505), .B1(n33991), .B2(n34503), .ZN(
        n32333) );
  XNOR2_X1 U34128 ( .A(n35110), .B(\fmem_data[31][1] ), .ZN(n34111) );
  OAI22_X1 U34129 ( .A1(n32178), .A2(n3931), .B1(n34111), .B2(n36216), .ZN(
        n32331) );
  XNOR2_X1 U34130 ( .A(n35140), .B(\fmem_data[7][1] ), .ZN(n33990) );
  OAI22_X1 U34131 ( .A1(n33990), .A2(n36218), .B1(n32181), .B2(n3581), .ZN(
        n32335) );
  OAI22_X1 U34132 ( .A1(n32183), .A2(n34923), .B1(n32182), .B2(n34922), .ZN(
        n32334) );
  FA_X1 U34133 ( .A(n32186), .B(n32185), .CI(n32184), .CO(n32353), .S(n32282)
         );
  XNOR2_X1 U34134 ( .A(n32188), .B(\fmem_data[3][1] ), .ZN(n33871) );
  OAI22_X1 U34135 ( .A1(n32189), .A2(n3582), .B1(n33871), .B2(n36199), .ZN(
        n32634) );
  XNOR2_X1 U34136 ( .A(n33484), .B(\fmem_data[31][5] ), .ZN(n33879) );
  OAI22_X1 U34137 ( .A1(n34944), .A2(n32190), .B1(n33879), .B2(n34945), .ZN(
        n32633) );
  XNOR2_X1 U34138 ( .A(n35114), .B(\fmem_data[23][1] ), .ZN(n33904) );
  OAI22_X1 U34139 ( .A1(n32191), .A2(n3662), .B1(n33904), .B2(n36241), .ZN(
        n32219) );
  XNOR2_X1 U34140 ( .A(n36311), .B(\fmem_data[7][7] ), .ZN(n32192) );
  OAI22_X1 U34141 ( .A1(n32193), .A2(n35619), .B1(n32192), .B2(n35618), .ZN(
        n32218) );
  XNOR2_X1 U34142 ( .A(n32194), .B(\fmem_data[3][3] ), .ZN(n33894) );
  OAI22_X1 U34143 ( .A1(n32195), .A2(n34420), .B1(n33894), .B2(n34418), .ZN(
        n32217) );
  FA_X1 U34144 ( .A(n32198), .B(n32197), .CI(n32196), .CO(n32338), .S(n32705)
         );
  FA_X1 U34145 ( .A(n32201), .B(n32200), .CI(n32199), .CO(n32305), .S(n32703)
         );
  XNOR2_X1 U34146 ( .A(n33939), .B(\fmem_data[15][3] ), .ZN(n32602) );
  OAI22_X1 U34147 ( .A1(n32205), .A2(n34364), .B1(n34363), .B2(n32602), .ZN(
        n32413) );
  OAI21_X1 U34148 ( .B1(n32411), .B2(n32410), .A(n32413), .ZN(n32207) );
  NAND2_X1 U34149 ( .A1(n32207), .A2(n32206), .ZN(n32272) );
  FA_X1 U34150 ( .A(n32210), .B(n32209), .CI(n32208), .CO(n32274), .S(n32926)
         );
  XNOR2_X1 U34151 ( .A(n32211), .B(\fmem_data[15][1] ), .ZN(n34403) );
  OAI21_X1 U34152 ( .B1(n32272), .B2(n32274), .A(n32271), .ZN(n32214) );
  NAND2_X1 U34153 ( .A1(n32214), .A2(n32213), .ZN(n32704) );
  OAI21_X1 U34154 ( .B1(n32705), .B2(n32703), .A(n32704), .ZN(n32216) );
  NAND2_X1 U34155 ( .A1(n32216), .A2(n32215), .ZN(n32367) );
  FA_X1 U34156 ( .A(n32219), .B(n32218), .CI(n32217), .CO(n32280), .S(n32372)
         );
  INV_X1 U34157 ( .A(n35615), .ZN(n32220) );
  OAI22_X1 U34158 ( .A1(n34196), .A2(n34194), .B1(n32221), .B2(n34195), .ZN(
        n32263) );
  INV_X1 U34159 ( .A(n32222), .ZN(n32224) );
  XNOR2_X1 U34160 ( .A(n32224), .B(n32223), .ZN(n32262) );
  XNOR2_X1 U34161 ( .A(n32228), .B(\fmem_data[5][3] ), .ZN(n33849) );
  FA_X1 U34162 ( .A(n32232), .B(n32231), .CI(n32230), .CO(n32301), .S(n32268)
         );
  XNOR2_X1 U34163 ( .A(n3376), .B(\fmem_data[11][3] ), .ZN(n34428) );
  OAI22_X1 U34164 ( .A1(n34533), .A2(n32234), .B1(n34428), .B2(n34429), .ZN(
        n32448) );
  INV_X1 U34165 ( .A(n32702), .ZN(n32248) );
  XNOR2_X1 U34166 ( .A(n33227), .B(\fmem_data[14][1] ), .ZN(n32601) );
  XNOR2_X1 U34167 ( .A(n32242), .B(\fmem_data[29][1] ), .ZN(n33579) );
  OAI22_X1 U34168 ( .A1(n32243), .A2(n3575), .B1(n33579), .B2(n36120), .ZN(
        n32627) );
  NOR2_X1 U34169 ( .A1(n32700), .A2(n32699), .ZN(n32247) );
  NAND2_X1 U34170 ( .A1(n32700), .A2(n32699), .ZN(n32246) );
  OAI21_X1 U34171 ( .B1(n32248), .B2(n32247), .A(n32246), .ZN(n32370) );
  FA_X1 U34172 ( .A(n32251), .B(n32250), .CI(n32249), .CO(n32304), .S(n32375)
         );
  INV_X1 U34173 ( .A(n35709), .ZN(n32252) );
  INV_X1 U34174 ( .A(n35753), .ZN(n32253) );
  XNOR2_X1 U34175 ( .A(n32953), .B(\fmem_data[26][5] ), .ZN(n33786) );
  OAI22_X1 U34176 ( .A1(n33786), .A2(n35033), .B1(n32254), .B2(n35034), .ZN(
        n32656) );
  XNOR2_X1 U34177 ( .A(n32256), .B(\fmem_data[23][3] ), .ZN(n34019) );
  OAI22_X1 U34178 ( .A1(n32257), .A2(n34412), .B1(n34019), .B2(n34410), .ZN(
        n32361) );
  FA_X1 U34179 ( .A(n32264), .B(n32263), .CI(n32262), .CO(n32364), .S(n32270)
         );
  FA_X1 U34180 ( .A(n32267), .B(n32266), .CI(n32265), .CO(n32088), .S(n33000)
         );
  FA_X1 U34181 ( .A(n32270), .B(n32269), .CI(n32268), .CO(n32371), .S(n32999)
         );
  XNOR2_X1 U34182 ( .A(n32272), .B(n32271), .ZN(n32273) );
  XNOR2_X1 U34183 ( .A(n32274), .B(n32273), .ZN(n32998) );
  FA_X1 U34184 ( .A(n32276), .B(n32277), .CI(n32275), .CO(n32460), .S(n33008)
         );
  OAI21_X1 U34185 ( .B1(n33006), .B2(n33007), .A(n33008), .ZN(n32279) );
  NAND2_X1 U34186 ( .A1(n33006), .A2(n33007), .ZN(n32278) );
  NAND2_X1 U34187 ( .A1(n32279), .A2(n32278), .ZN(n32507) );
  FA_X1 U34188 ( .A(n32282), .B(n32281), .CI(n32280), .CO(n32383), .S(n32368)
         );
  XNOR2_X1 U34189 ( .A(n32283), .B(\fmem_data[18][3] ), .ZN(n33646) );
  OAI22_X1 U34190 ( .A1(n33646), .A2(n33679), .B1(n32284), .B2(n33681), .ZN(
        n32664) );
  INV_X1 U34191 ( .A(n35516), .ZN(n32285) );
  XNOR2_X1 U34192 ( .A(n33554), .B(\fmem_data[2][5] ), .ZN(n33848) );
  OAI22_X1 U34193 ( .A1(n33848), .A2(n35018), .B1(n32286), .B2(n35019), .ZN(
        n32662) );
  XNOR2_X1 U34194 ( .A(n36316), .B(n3698), .ZN(n32288) );
  NAND2_X1 U34195 ( .A1(n32288), .A2(n32287), .ZN(n32296) );
  OR2_X1 U34196 ( .A1(n32289), .A2(n35642), .ZN(n32295) );
  NAND3_X1 U34197 ( .A1(n32296), .A2(n32295), .A3(n32293), .ZN(n32294) );
  NAND2_X1 U34198 ( .A1(n32328), .A2(n32294), .ZN(n32298) );
  NAND2_X1 U34199 ( .A1(n32296), .A2(n32295), .ZN(n32329) );
  NAND2_X1 U34200 ( .A1(n32329), .A2(n32327), .ZN(n32297) );
  NAND2_X1 U34201 ( .A1(n32298), .A2(n32297), .ZN(n32326) );
  FA_X1 U34202 ( .A(n3707), .B(n32300), .CI(n32299), .CO(n33083), .S(n32325)
         );
  FA_X1 U34203 ( .A(n32303), .B(n32302), .CI(n32301), .CO(n32324), .S(n32408)
         );
  FA_X1 U34204 ( .A(n32306), .B(n32305), .CI(n32304), .CO(n32381), .S(n32807)
         );
  OAI22_X1 U34205 ( .A1(n32308), .A2(n34903), .B1(n32307), .B2(n34904), .ZN(
        n32638) );
  XNOR2_X1 U34206 ( .A(n36313), .B(\fmem_data[11][7] ), .ZN(n32310) );
  OAI22_X1 U34207 ( .A1(n32310), .A2(n35633), .B1(n32309), .B2(n35634), .ZN(
        n32637) );
  FA_X1 U34208 ( .A(n32313), .B(n32312), .CI(n32311), .CO(n32636), .S(n32269)
         );
  FA_X1 U34209 ( .A(n32316), .B(n32315), .CI(n32314), .CO(n32342), .S(n32409)
         );
  XNOR2_X1 U34210 ( .A(n32319), .B(\fmem_data[29][3] ), .ZN(n33966) );
  OAI22_X1 U34211 ( .A1(n33966), .A2(n34424), .B1(n32320), .B2(n34422), .ZN(
        n33067) );
  XNOR2_X1 U34212 ( .A(n32342), .B(n32343), .ZN(n32323) );
  XNOR2_X1 U34213 ( .A(n32344), .B(n32323), .ZN(n32399) );
  FA_X1 U34214 ( .A(n32326), .B(n32325), .CI(n32324), .CO(n32382), .S(n32398)
         );
  FA_X1 U34215 ( .A(n32333), .B(n32332), .CI(n32331), .CO(n32355), .S(n32405)
         );
  FA_X1 U34216 ( .A(n32336), .B(n32335), .CI(n32334), .CO(n32354), .S(n32404)
         );
  OAI21_X1 U34217 ( .B1(n32338), .B2(n32339), .A(n32337), .ZN(n32341) );
  NAND2_X1 U34218 ( .A1(n32339), .A2(n32338), .ZN(n32340) );
  NAND2_X1 U34219 ( .A1(n32341), .A2(n32340), .ZN(n32389) );
  OAI21_X1 U34220 ( .B1(n32344), .B2(n32343), .A(n32342), .ZN(n32346) );
  NAND2_X1 U34221 ( .A1(n32344), .A2(n32343), .ZN(n32345) );
  NAND2_X1 U34222 ( .A1(n32346), .A2(n32345), .ZN(n32388) );
  XNOR2_X1 U34223 ( .A(n32348), .B(n32347), .ZN(n32349) );
  XNOR2_X1 U34224 ( .A(n32350), .B(n32349), .ZN(n32387) );
  FA_X1 U34225 ( .A(n32353), .B(n32352), .CI(n32351), .CO(n33117), .S(n32386)
         );
  FA_X1 U34226 ( .A(n32356), .B(n32355), .CI(n32354), .CO(n32385), .S(n32369)
         );
  FA_X1 U34227 ( .A(n32363), .B(n32362), .CI(n32361), .CO(n32377), .S(n32374)
         );
  FA_X1 U34228 ( .A(n32366), .B(n32365), .CI(n32364), .CO(n32376), .S(n32373)
         );
  FA_X1 U34229 ( .A(n32369), .B(n32368), .CI(n32367), .CO(n32392), .S(n32916)
         );
  FA_X1 U34230 ( .A(n32372), .B(n32371), .CI(n32370), .CO(n32402), .S(n32858)
         );
  FA_X1 U34231 ( .A(n32375), .B(n32374), .CI(n32373), .CO(n32400), .S(n32857)
         );
  FA_X1 U34232 ( .A(n32378), .B(n32377), .CI(n32376), .CO(n32384), .S(n32401)
         );
  OAI21_X1 U34233 ( .B1(n32402), .B2(n32400), .A(n32401), .ZN(n32380) );
  NAND2_X1 U34234 ( .A1(n32402), .A2(n32400), .ZN(n32379) );
  NAND2_X1 U34235 ( .A1(n32380), .A2(n32379), .ZN(n32391) );
  XNOR2_X1 U34236 ( .A(n33094), .B(n33095), .ZN(n32390) );
  FA_X1 U34237 ( .A(n32383), .B(n32382), .CI(n32381), .CO(n33149), .S(n32396)
         );
  FA_X1 U34238 ( .A(n32386), .B(n32385), .CI(n32384), .CO(n33148), .S(n32393)
         );
  FA_X1 U34239 ( .A(n32389), .B(n32388), .CI(n32387), .CO(n33147), .S(n32394)
         );
  XNOR2_X1 U34240 ( .A(n32390), .B(n33093), .ZN(n32508) );
  FA_X1 U34241 ( .A(n32393), .B(n32392), .CI(n32391), .CO(n33094), .S(n32512)
         );
  FA_X1 U34242 ( .A(n32396), .B(n32395), .CI(n32394), .CO(n33095), .S(n32511)
         );
  FA_X1 U34243 ( .A(n32399), .B(n32398), .CI(n32397), .CO(n32395), .S(n32852)
         );
  XNOR2_X1 U34244 ( .A(n32401), .B(n32400), .ZN(n32403) );
  XNOR2_X1 U34245 ( .A(n32403), .B(n32402), .ZN(n32851) );
  FA_X1 U34246 ( .A(n32406), .B(n32405), .CI(n32404), .CO(n32397), .S(n32855)
         );
  FA_X1 U34247 ( .A(n32409), .B(n32408), .CI(n32407), .CO(n32808), .S(n32854)
         );
  XNOR2_X1 U34248 ( .A(n32413), .B(n32412), .ZN(n32906) );
  FA_X1 U34249 ( .A(n32416), .B(n32415), .CI(n32414), .CO(n32209), .S(n32875)
         );
  XNOR2_X1 U34250 ( .A(n33019), .B(\fmem_data[23][1] ), .ZN(n34360) );
  XNOR2_X1 U34251 ( .A(n33551), .B(\fmem_data[20][3] ), .ZN(n34498) );
  OAI22_X1 U34252 ( .A1(n34498), .A2(n34495), .B1(n32418), .B2(n34497), .ZN(
        n32873) );
  XNOR2_X1 U34253 ( .A(n32419), .B(\fmem_data[5][1] ), .ZN(n34482) );
  XNOR2_X1 U34254 ( .A(n3353), .B(\fmem_data[2][3] ), .ZN(n32421) );
  OAI22_X1 U34255 ( .A1(n32422), .A2(n33797), .B1(n33796), .B2(n32421), .ZN(
        n34792) );
  OAI22_X1 U34256 ( .A1(n33748), .A2(n34625), .B1(n32428), .B2(n3574), .ZN(
        n32866) );
  OAI21_X1 U34257 ( .B1(n32869), .B2(n32867), .A(n32866), .ZN(n32430) );
  NAND2_X1 U34258 ( .A1(n32869), .A2(n32867), .ZN(n32429) );
  NAND2_X1 U34259 ( .A1(n32430), .A2(n32429), .ZN(n32904) );
  INV_X1 U34260 ( .A(n32861), .ZN(n32456) );
  OR2_X1 U34261 ( .A1(n34626), .A2(n3700), .ZN(n32432) );
  OAI22_X1 U34262 ( .A1(n32432), .A2(n34206), .B1(n34208), .B2(n3700), .ZN(
        n32896) );
  XNOR2_X1 U34263 ( .A(n36111), .B(\fmem_data[26][3] ), .ZN(n32433) );
  OAI22_X1 U34264 ( .A1(n32434), .A2(n32780), .B1(n32433), .B2(n32779), .ZN(
        n32895) );
  OR2_X1 U34265 ( .A1(n36296), .A2(n3667), .ZN(n32436) );
  OAI22_X1 U34266 ( .A1(n32436), .A2(n34537), .B1(n34535), .B2(n3667), .ZN(
        n32893) );
  XNOR2_X1 U34267 ( .A(n32596), .B(\fmem_data[18][1] ), .ZN(n32941) );
  OAI22_X1 U34268 ( .A1(n32437), .A2(n3580), .B1(n32941), .B2(n36104), .ZN(
        n32892) );
  XNOR2_X1 U34269 ( .A(n32440), .B(\fmem_data[7][1] ), .ZN(n33700) );
  OAI22_X1 U34270 ( .A1(n33700), .A2(n36218), .B1(n32441), .B2(n3581), .ZN(
        n32844) );
  XNOR2_X1 U34271 ( .A(n32444), .B(\fmem_data[27][1] ), .ZN(n33736) );
  OAI22_X1 U34272 ( .A1(n33736), .A2(n36240), .B1(n32445), .B2(n3482), .ZN(
        n32842) );
  FA_X1 U34273 ( .A(n32448), .B(n32447), .CI(n32446), .CO(n32702), .S(n34763)
         );
  OAI21_X1 U34274 ( .B1(n34762), .B2(n34761), .A(n34763), .ZN(n32450) );
  NAND2_X1 U34275 ( .A1(n32450), .A2(n32449), .ZN(n32860) );
  FA_X1 U34276 ( .A(n32453), .B(n32452), .CI(n32451), .CO(n32407), .S(n32859)
         );
  NOR2_X1 U34277 ( .A1(n32860), .A2(n32859), .ZN(n32455) );
  NAND2_X1 U34278 ( .A1(n32860), .A2(n32859), .ZN(n32454) );
  OAI21_X1 U34279 ( .B1(n32456), .B2(n32455), .A(n32454), .ZN(n32853) );
  OAI21_X1 U34280 ( .B1(n32507), .B2(n32508), .A(n32506), .ZN(n32458) );
  NAND2_X1 U34281 ( .A1(n32507), .A2(n32508), .ZN(n32457) );
  NAND2_X1 U34282 ( .A1(n32458), .A2(n32457), .ZN(n33403) );
  FA_X1 U34283 ( .A(n32461), .B(n32460), .CI(n32459), .CO(n31634), .S(n33413)
         );
  XNOR2_X1 U34284 ( .A(n32463), .B(n32462), .ZN(n32464) );
  XNOR2_X1 U34285 ( .A(n32465), .B(n32464), .ZN(n33412) );
  FA_X1 U34286 ( .A(n32468), .B(n32467), .CI(n32466), .CO(n32459), .S(n33012)
         );
  XNOR2_X1 U34287 ( .A(n32470), .B(n32469), .ZN(n32472) );
  XNOR2_X1 U34288 ( .A(n32472), .B(n32471), .ZN(n33011) );
  FA_X1 U34289 ( .A(n32475), .B(n32474), .CI(n32473), .CO(n32098), .S(n32924)
         );
  XNOR2_X1 U34290 ( .A(n32477), .B(n32476), .ZN(n32479) );
  XNOR2_X1 U34291 ( .A(n32479), .B(n3393), .ZN(n32923) );
  FA_X1 U34292 ( .A(n32482), .B(n32481), .CI(n32480), .CO(n32090), .S(n33430)
         );
  FA_X1 U34293 ( .A(n32485), .B(n32484), .CI(n32483), .CO(n31436), .S(n33429)
         );
  FA_X1 U34294 ( .A(n32488), .B(n32487), .CI(n32486), .CO(n32482), .S(n33436)
         );
  FA_X1 U34295 ( .A(n32491), .B(n32490), .CI(n32489), .CO(n32484), .S(n33435)
         );
  XNOR2_X1 U34296 ( .A(n32493), .B(n32492), .ZN(n32494) );
  XNOR2_X1 U34297 ( .A(n32495), .B(n32494), .ZN(n33434) );
  FA_X1 U34298 ( .A(n32498), .B(n32497), .CI(n32496), .CO(n32470), .S(n33420)
         );
  OAI21_X1 U34299 ( .B1(n33413), .B2(n33412), .A(n33414), .ZN(n32504) );
  NAND2_X1 U34300 ( .A1(n33413), .A2(n33412), .ZN(n32503) );
  NAND2_X1 U34301 ( .A1(n32504), .A2(n32503), .ZN(n33402) );
  XNOR2_X1 U34302 ( .A(n35455), .B(n35456), .ZN(n32505) );
  XNOR2_X1 U34303 ( .A(n35454), .B(n32505), .ZN(n36440) );
  XNOR2_X1 U34304 ( .A(n32507), .B(n32506), .ZN(n32509) );
  XNOR2_X1 U34305 ( .A(n32509), .B(n32508), .ZN(n36033) );
  FA_X1 U34306 ( .A(n32512), .B(n32511), .CI(n32510), .CO(n32506), .S(n36037)
         );
  FA_X1 U34307 ( .A(n32521), .B(n32520), .CI(n32519), .CO(n32722), .S(n32762)
         );
  OAI22_X1 U34308 ( .A1(n32529), .A2(n34422), .B1(n34423), .B2(n34424), .ZN(
        n32775) );
  XNOR2_X1 U34309 ( .A(n33751), .B(\fmem_data[17][5] ), .ZN(n32530) );
  OAI22_X1 U34310 ( .A1(n32531), .A2(n34045), .B1(n32530), .B2(n34043), .ZN(
        n32548) );
  INV_X1 U34311 ( .A(n34045), .ZN(n32532) );
  INV_X1 U34312 ( .A(n35003), .ZN(n32533) );
  INV_X1 U34313 ( .A(n35011), .ZN(n32534) );
  AND2_X1 U34314 ( .A1(n34599), .A2(n32534), .ZN(n32618) );
  OAI21_X1 U34315 ( .B1(n32791), .B2(n32792), .A(n32793), .ZN(n32538) );
  NAND2_X1 U34316 ( .A1(n32538), .A2(n32537), .ZN(n32761) );
  XNOR2_X1 U34317 ( .A(n33800), .B(\fmem_data[13][5] ), .ZN(n32540) );
  OAI22_X1 U34318 ( .A1(n32540), .A2(n35181), .B1(n32539), .B2(n35182), .ZN(
        n32568) );
  XNOR2_X1 U34319 ( .A(n32541), .B(\fmem_data[13][3] ), .ZN(n33569) );
  OAI22_X1 U34320 ( .A1(n32542), .A2(n33568), .B1(n33569), .B2(n33570), .ZN(
        n32567) );
  XNOR2_X1 U34321 ( .A(n32568), .B(n32567), .ZN(n32545) );
  OAI22_X1 U34322 ( .A1(n33833), .A2(n34529), .B1(n32544), .B2(n3566), .ZN(
        n32566) );
  FA_X1 U34323 ( .A(n32548), .B(n32547), .CI(n32546), .CO(n32793), .S(n34725)
         );
  OR2_X1 U34324 ( .A1(n34623), .A2(n3701), .ZN(n32549) );
  OAI22_X1 U34325 ( .A1(n32549), .A2(n33850), .B1(n33851), .B2(n3701), .ZN(
        n32889) );
  OAI22_X1 U34326 ( .A1(n32550), .A2(n33681), .B1(n33679), .B2(n3664), .ZN(
        n32888) );
  OR2_X1 U34327 ( .A1(n34612), .A2(n3646), .ZN(n32553) );
  OAI22_X1 U34328 ( .A1(n32553), .A2(n33596), .B1(n33598), .B2(n3646), .ZN(
        n34748) );
  XNOR2_X1 U34329 ( .A(n32554), .B(\fmem_data[26][1] ), .ZN(n33724) );
  OAI22_X1 U34330 ( .A1(n32555), .A2(n3678), .B1(n33724), .B2(n33725), .ZN(
        n34747) );
  INV_X1 U34331 ( .A(n32557), .ZN(n32556) );
  NAND2_X1 U34332 ( .A1(n32556), .A2(\fmem_data[3][1] ), .ZN(n32559) );
  NAND3_X1 U34333 ( .A1(n3275), .A2(n32557), .A3(n3695), .ZN(n32558) );
  OAI211_X1 U34334 ( .C1(n3274), .C2(n3695), .A(n32559), .B(n32558), .ZN(
        n33721) );
  OAI22_X1 U34335 ( .A1(n33721), .A2(n36199), .B1(n32561), .B2(n3582), .ZN(
        n32839) );
  OAI21_X1 U34336 ( .B1(n32568), .B2(n32567), .A(n32566), .ZN(n32570) );
  NAND2_X1 U34337 ( .A1(n32570), .A2(n32569), .ZN(n32745) );
  OAI22_X1 U34338 ( .A1(n32574), .A2(n3560), .B1(n32573), .B2(n34788), .ZN(
        n32799) );
  INV_X1 U34339 ( .A(n35041), .ZN(n32577) );
  INV_X1 U34340 ( .A(n34039), .ZN(n32578) );
  INV_X1 U34341 ( .A(n35182), .ZN(n32579) );
  XNOR2_X1 U34342 ( .A(n34624), .B(\fmem_data[28][5] ), .ZN(n32580) );
  OAI22_X1 U34343 ( .A1(n32581), .A2(n33828), .B1(n32580), .B2(n33827), .ZN(
        n32623) );
  XNOR2_X1 U34344 ( .A(n32736), .B(n32735), .ZN(n32591) );
  XNOR2_X1 U34345 ( .A(n32586), .B(\fmem_data[12][1] ), .ZN(n33780) );
  OAI22_X1 U34346 ( .A1(n32587), .A2(n3572), .B1(n33780), .B2(n34734), .ZN(
        n32773) );
  INV_X1 U34347 ( .A(n35019), .ZN(n32588) );
  INV_X1 U34348 ( .A(n33643), .ZN(n32589) );
  INV_X1 U34349 ( .A(n35036), .ZN(n32590) );
  XNOR2_X1 U34350 ( .A(n32591), .B(n32737), .ZN(n32826) );
  NAND2_X1 U34351 ( .A1(n32593), .A2(n32592), .ZN(n34802) );
  XNOR2_X1 U34352 ( .A(n32937), .B(\fmem_data[19][3] ), .ZN(n34473) );
  OAI22_X1 U34353 ( .A1(n32595), .A2(n34472), .B1(n34473), .B2(n34474), .ZN(
        n34731) );
  XNOR2_X1 U34354 ( .A(n32940), .B(\fmem_data[18][3] ), .ZN(n33682) );
  XNOR2_X1 U34355 ( .A(n32596), .B(\fmem_data[18][3] ), .ZN(n33645) );
  OAI22_X1 U34356 ( .A1(n34402), .A2(n3568), .B1(n32598), .B2(n36223), .ZN(
        n34527) );
  XNOR2_X1 U34357 ( .A(n33225), .B(\fmem_data[16][1] ), .ZN(n34025) );
  XNOR2_X1 U34358 ( .A(n32600), .B(\fmem_data[14][1] ), .ZN(n33593) );
  XNOR2_X1 U34359 ( .A(n32603), .B(\fmem_data[7][3] ), .ZN(n34506) );
  OAI22_X1 U34360 ( .A1(n34506), .A2(n34503), .B1(n32604), .B2(n34505), .ZN(
        n32871) );
  XNOR2_X1 U34361 ( .A(n36110), .B(\fmem_data[25][3] ), .ZN(n32607) );
  OAI22_X1 U34362 ( .A1(n32607), .A2(n33057), .B1(n32606), .B2(n33059), .ZN(
        n34540) );
  FA_X1 U34363 ( .A(n32611), .B(n32610), .CI(n32609), .CO(n32197), .S(n32672)
         );
  XNOR2_X1 U34364 ( .A(n32616), .B(\fmem_data[9][1] ), .ZN(n34478) );
  XNOR2_X1 U34365 ( .A(n32617), .B(\fmem_data[9][1] ), .ZN(n34197) );
  OAI22_X1 U34366 ( .A1(n34478), .A2(n34476), .B1(n34197), .B2(n3579), .ZN(
        n34775) );
  FA_X1 U34367 ( .A(n32620), .B(n32619), .CI(n32618), .CO(n32547), .S(n34774)
         );
  FA_X1 U34368 ( .A(n32624), .B(n32623), .CI(n32622), .CO(n32735), .S(n34759)
         );
  FA_X1 U34369 ( .A(n32627), .B(n32626), .CI(n32625), .CO(n32699), .S(n34758)
         );
  NAND2_X1 U34370 ( .A1(n32629), .A2(n32628), .ZN(n34801) );
  FA_X1 U34371 ( .A(n32632), .B(n32631), .CI(n32630), .CO(n32306), .S(n32676)
         );
  FA_X1 U34372 ( .A(n32635), .B(n32634), .CI(n32633), .CO(n32281), .S(n32675)
         );
  FA_X1 U34373 ( .A(n32638), .B(n32637), .CI(n32636), .CO(n32344), .S(n32677)
         );
  OAI21_X1 U34374 ( .B1(n32676), .B2(n32675), .A(n32677), .ZN(n32640) );
  NAND2_X1 U34375 ( .A1(n32676), .A2(n32675), .ZN(n32639) );
  NAND2_X1 U34376 ( .A1(n32640), .A2(n32639), .ZN(n32816) );
  OAI22_X1 U34377 ( .A1(n32642), .A2(n33797), .B1(n33796), .B2(n32641), .ZN(
        n33077) );
  OAI22_X1 U34378 ( .A1(n32644), .A2(n33853), .B1(n32643), .B2(n33855), .ZN(
        n33076) );
  OAI22_X1 U34379 ( .A1(n32646), .A2(n33249), .B1(n32645), .B2(n33250), .ZN(
        n33075) );
  FA_X1 U34380 ( .A(n32649), .B(n32647), .CI(n32648), .CO(n33025), .S(n33277)
         );
  XNOR2_X1 U34381 ( .A(n36315), .B(\fmem_data[3][7] ), .ZN(n32653) );
  OAI22_X1 U34382 ( .A1(n32653), .A2(n35637), .B1(n32652), .B2(n35638), .ZN(
        n32749) );
  INV_X1 U34383 ( .A(n36311), .ZN(n36122) );
  NAND2_X1 U34384 ( .A1(n36122), .A2(\fmem_data[7][7] ), .ZN(n32654) );
  OAI22_X1 U34385 ( .A1(n32654), .A2(n35619), .B1(n35618), .B2(n3490), .ZN(
        n32748) );
  XNOR2_X1 U34386 ( .A(n32655), .B(n33275), .ZN(n32815) );
  FA_X1 U34387 ( .A(n32658), .B(n32657), .CI(n32656), .CO(n32363), .S(n32681)
         );
  FA_X1 U34388 ( .A(n32661), .B(n32660), .CI(n32659), .CO(n32200), .S(n32680)
         );
  FA_X1 U34389 ( .A(n32664), .B(n32663), .CI(n32662), .CO(n32328), .S(n32679)
         );
  OR2_X1 U34390 ( .A1(n36313), .A2(n3663), .ZN(n32669) );
  FA_X1 U34391 ( .A(n32672), .B(n32671), .CI(n32670), .CO(n32770), .S(n32829)
         );
  XNOR2_X1 U34392 ( .A(n32676), .B(n32675), .ZN(n32678) );
  XNOR2_X1 U34393 ( .A(n32678), .B(n32677), .ZN(n32821) );
  FA_X1 U34394 ( .A(n32681), .B(n32680), .CI(n32679), .CO(n32769), .S(n32865)
         );
  FA_X1 U34395 ( .A(n32684), .B(n32683), .CI(n32682), .CO(n32453), .S(n34753)
         );
  XNOR2_X1 U34396 ( .A(n32686), .B(n32685), .ZN(n32688) );
  XNOR2_X1 U34397 ( .A(n32688), .B(n32687), .ZN(n34729) );
  FA_X1 U34398 ( .A(n32693), .B(n32692), .CI(n32691), .CO(n32624), .S(n34727)
         );
  FA_X1 U34399 ( .A(n32696), .B(n32695), .CI(n32694), .CO(n32700), .S(n34754)
         );
  OAI21_X1 U34400 ( .B1(n34753), .B2(n34752), .A(n34754), .ZN(n32698) );
  NAND2_X1 U34401 ( .A1(n32698), .A2(n32697), .ZN(n32864) );
  XNOR2_X1 U34402 ( .A(n32700), .B(n32699), .ZN(n32701) );
  XNOR2_X1 U34403 ( .A(n32702), .B(n32701), .ZN(n32863) );
  XNOR2_X1 U34404 ( .A(n32704), .B(n32703), .ZN(n32706) );
  XNOR2_X1 U34405 ( .A(n32706), .B(n32705), .ZN(n32819) );
  OAI21_X1 U34406 ( .B1(n34808), .B2(n34806), .A(n34807), .ZN(n32707) );
  NAND2_X1 U34407 ( .A1(n32708), .A2(n32707), .ZN(n33294) );
  FA_X1 U34408 ( .A(n32710), .B(n32711), .CI(n32709), .CO(n33082), .S(n33210)
         );
  NAND2_X1 U34409 ( .A1(n32712), .A2(n31535), .ZN(n32713) );
  OAI21_X1 U34410 ( .B1(n34535), .B2(n32714), .A(n32713), .ZN(n32744) );
  XNOR2_X1 U34411 ( .A(n36312), .B(\fmem_data[10][7] ), .ZN(n32715) );
  XNOR2_X1 U34412 ( .A(n34531), .B(\fmem_data[10][7] ), .ZN(n33268) );
  OAI22_X1 U34413 ( .A1(n32717), .A2(n34431), .B1(n32716), .B2(n34433), .ZN(
        n32742) );
  FA_X1 U34414 ( .A(n32720), .B(n32719), .CI(n32718), .CO(n33208), .S(n32768)
         );
  FA_X1 U34415 ( .A(n32723), .B(n32722), .CI(n32721), .CO(n32812), .S(n34675)
         );
  XNOR2_X1 U34416 ( .A(n32727), .B(\fmem_data[19][3] ), .ZN(n34191) );
  OAI22_X1 U34417 ( .A1(n34191), .A2(n34474), .B1(n32728), .B2(n34472), .ZN(
        n32758) );
  OAI21_X1 U34418 ( .B1(n32737), .B2(n32736), .A(n32735), .ZN(n32739) );
  NAND2_X1 U34419 ( .A1(n32739), .A2(n32738), .ZN(n34397) );
  OAI21_X1 U34420 ( .B1(n34396), .B2(n34395), .A(n34397), .ZN(n32741) );
  NAND2_X1 U34421 ( .A1(n34396), .A2(n34395), .ZN(n32740) );
  NAND2_X1 U34422 ( .A1(n32741), .A2(n32740), .ZN(n34674) );
  FA_X1 U34423 ( .A(n32744), .B(n32743), .CI(n32742), .CO(n33209), .S(n32767)
         );
  FA_X1 U34424 ( .A(n32747), .B(n32746), .CI(n32745), .CO(n32766), .S(n32825)
         );
  FA_X1 U34425 ( .A(n32750), .B(n32748), .CI(n32749), .CO(n33275), .S(n32765)
         );
  FA_X1 U34426 ( .A(n32760), .B(n32759), .CI(n32758), .CO(n33155), .S(n34396)
         );
  XNOR2_X1 U34427 ( .A(n33290), .B(n33289), .ZN(n32764) );
  FA_X1 U34428 ( .A(n32763), .B(n32762), .CI(n32761), .CO(n33288), .S(n34803)
         );
  XNOR2_X1 U34429 ( .A(n32764), .B(n33288), .ZN(n34718) );
  XNOR2_X1 U34430 ( .A(n32769), .B(n32768), .ZN(n32771) );
  XNOR2_X1 U34431 ( .A(n32771), .B(n32770), .ZN(n32823) );
  FA_X1 U34432 ( .A(n32774), .B(n32773), .CI(n32772), .CO(n32737), .S(n34517)
         );
  FA_X1 U34433 ( .A(n32777), .B(n32776), .CI(n32775), .CO(n32792), .S(n34516)
         );
  XNOR2_X1 U34434 ( .A(n3365), .B(\fmem_data[9][3] ), .ZN(n32782) );
  OAI22_X1 U34435 ( .A1(n32783), .A2(n33873), .B1(n32782), .B2(n33875), .ZN(
        n34765) );
  FA_X1 U34436 ( .A(n32786), .B(n32785), .CI(n32784), .CO(n32772), .S(n32846)
         );
  XNOR2_X1 U34437 ( .A(n32787), .B(\fmem_data[2][1] ), .ZN(n34342) );
  OAI22_X1 U34438 ( .A1(n34343), .A2(n34342), .B1(n32788), .B2(n3578), .ZN(
        n34770) );
  OR2_X1 U34439 ( .A1(n36101), .A2(n3605), .ZN(n32789) );
  FA_X1 U34440 ( .A(n32797), .B(n32796), .CI(n32795), .CO(n32452), .S(n32835)
         );
  FA_X1 U34441 ( .A(n32800), .B(n32798), .CI(n32799), .CO(n32736), .S(n32834)
         );
  FA_X1 U34442 ( .A(n32803), .B(n32802), .CI(n32801), .CO(n32451), .S(n32833)
         );
  OAI21_X1 U34443 ( .B1(n34722), .B2(n34720), .A(n34721), .ZN(n32805) );
  NAND2_X1 U34444 ( .A1(n34722), .A2(n34720), .ZN(n32804) );
  NAND2_X1 U34445 ( .A1(n32805), .A2(n32804), .ZN(n32822) );
  OAI21_X1 U34446 ( .B1(n32808), .B2(n32807), .A(n32806), .ZN(n32810) );
  NAND2_X1 U34447 ( .A1(n32808), .A2(n32807), .ZN(n32809) );
  NAND2_X1 U34448 ( .A1(n32810), .A2(n32809), .ZN(n33089) );
  FA_X1 U34449 ( .A(n32813), .B(n32812), .CI(n32811), .CO(n33084), .S(n33090)
         );
  XNOR2_X1 U34450 ( .A(n33089), .B(n33090), .ZN(n32817) );
  FA_X1 U34451 ( .A(n32816), .B(n32815), .CI(n32814), .CO(n33088), .S(n34806)
         );
  XNOR2_X1 U34452 ( .A(n32817), .B(n33088), .ZN(n33293) );
  XNOR2_X1 U34453 ( .A(n33295), .B(n33293), .ZN(n32818) );
  XNOR2_X1 U34454 ( .A(n33294), .B(n32818), .ZN(n36036) );
  FA_X1 U34455 ( .A(n32821), .B(n32820), .CI(n32819), .CO(n34807), .S(n36267)
         );
  FA_X1 U34456 ( .A(n32824), .B(n32823), .CI(n32822), .CO(n34717), .S(n36266)
         );
  XNOR2_X1 U34457 ( .A(n32828), .B(n32827), .ZN(n36078) );
  XNOR2_X1 U34458 ( .A(n32830), .B(n32829), .ZN(n32832) );
  XNOR2_X1 U34459 ( .A(n32832), .B(n32831), .ZN(n36080) );
  FA_X1 U34460 ( .A(n32835), .B(n32834), .CI(n32833), .CO(n34721), .S(n36162)
         );
  FA_X1 U34461 ( .A(n32838), .B(n32837), .CI(n32836), .CO(n32831), .S(n36161)
         );
  FA_X1 U34462 ( .A(n32841), .B(n32840), .CI(n32839), .CO(n34724), .S(n36169)
         );
  FA_X1 U34463 ( .A(n32844), .B(n32843), .CI(n32842), .CO(n34761), .S(n36168)
         );
  FA_X1 U34464 ( .A(n32847), .B(n32846), .CI(n32845), .CO(n34515), .S(n36167)
         );
  OAI21_X1 U34465 ( .B1(n36078), .B2(n36080), .A(n36079), .ZN(n32849) );
  NAND2_X1 U34466 ( .A1(n32849), .A2(n32848), .ZN(n36265) );
  FA_X1 U34467 ( .A(n32852), .B(n32851), .CI(n32850), .CO(n32510), .S(n36153)
         );
  FA_X1 U34468 ( .A(n32855), .B(n32854), .CI(n32853), .CO(n32850), .S(n36270)
         );
  FA_X1 U34469 ( .A(n32858), .B(n32857), .CI(n32856), .CO(n32915), .S(n36269)
         );
  XNOR2_X1 U34470 ( .A(n32860), .B(n32859), .ZN(n32862) );
  XNOR2_X1 U34471 ( .A(n32862), .B(n32861), .ZN(n36182) );
  FA_X1 U34472 ( .A(n32865), .B(n32864), .CI(n32863), .CO(n32820), .S(n36181)
         );
  FA_X1 U34473 ( .A(n32872), .B(n32871), .CI(n32870), .CO(n32836), .S(n36171)
         );
  FA_X1 U34474 ( .A(n32875), .B(n32874), .CI(n32873), .CO(n32905), .S(n36170)
         );
  OAI21_X1 U34475 ( .B1(n36172), .B2(n36171), .A(n36170), .ZN(n32877) );
  NAND2_X1 U34476 ( .A1(n32877), .A2(n32876), .ZN(n36185) );
  FA_X1 U34477 ( .A(n32880), .B(n32879), .CI(n32878), .CO(n34762), .S(n36176)
         );
  INV_X1 U34478 ( .A(n34505), .ZN(n32881) );
  OAI22_X1 U34479 ( .A1(n33757), .A2(n34017), .B1(n32883), .B2(n3559), .ZN(
        n36205) );
  INV_X1 U34480 ( .A(n34463), .ZN(n32884) );
  AND2_X1 U34481 ( .A1(n36316), .A2(n32884), .ZN(n36206) );
  OAI21_X1 U34482 ( .B1(n36204), .B2(n36205), .A(n36206), .ZN(n32886) );
  NAND2_X1 U34483 ( .A1(n32886), .A2(n32885), .ZN(n36135) );
  FA_X1 U34484 ( .A(n32889), .B(n32888), .CI(n32887), .CO(n32841), .S(n36134)
         );
  INV_X1 U34485 ( .A(n34412), .ZN(n32890) );
  AND2_X1 U34486 ( .A1(n3116), .A2(n32890), .ZN(n36258) );
  INV_X1 U34487 ( .A(n34364), .ZN(n32891) );
  FA_X1 U34488 ( .A(n32894), .B(n32893), .CI(n32892), .CO(n32879), .S(n36195)
         );
  FA_X1 U34489 ( .A(n32897), .B(n32896), .CI(n32895), .CO(n32880), .S(n36194)
         );
  XNOR2_X1 U34490 ( .A(n32899), .B(\fmem_data[8][1] ), .ZN(n33747) );
  INV_X1 U34491 ( .A(n34420), .ZN(n32900) );
  INV_X1 U34492 ( .A(n34472), .ZN(n32901) );
  OAI21_X1 U34493 ( .B1(n36176), .B2(n36175), .A(n36174), .ZN(n32903) );
  NAND2_X1 U34494 ( .A1(n32903), .A2(n32902), .ZN(n36184) );
  FA_X1 U34495 ( .A(n32906), .B(n32905), .CI(n32904), .CO(n32861), .S(n36183)
         );
  OAI21_X1 U34496 ( .B1(n36037), .B2(n36036), .A(n36038), .ZN(n32910) );
  NAND2_X1 U34497 ( .A1(n36037), .A2(n36036), .ZN(n32909) );
  NAND2_X1 U34498 ( .A1(n32910), .A2(n32909), .ZN(n36032) );
  XNOR2_X1 U34499 ( .A(n32912), .B(n32911), .ZN(n32914) );
  XNOR2_X1 U34500 ( .A(n32914), .B(n32913), .ZN(n36159) );
  FA_X1 U34501 ( .A(n32917), .B(n32916), .CI(n32915), .CO(n33007), .S(n36158)
         );
  XNOR2_X1 U34502 ( .A(n32919), .B(n32918), .ZN(n32921) );
  XNOR2_X1 U34503 ( .A(n32921), .B(n32920), .ZN(n36374) );
  FA_X1 U34504 ( .A(n32924), .B(n32923), .CI(n32922), .CO(n33421), .S(n36373)
         );
  FA_X1 U34505 ( .A(n32927), .B(n32926), .CI(n32925), .CO(n33002), .S(n36284)
         );
  OAI22_X1 U34506 ( .A1(n36121), .A2(n36120), .B1(n32928), .B2(n3575), .ZN(
        n36259) );
  XNOR2_X1 U34507 ( .A(n32929), .B(\fmem_data[23][1] ), .ZN(n34359) );
  XNOR2_X1 U34508 ( .A(n34361), .B(n3735), .ZN(n36242) );
  XNOR2_X1 U34509 ( .A(n33733), .B(\fmem_data[11][1] ), .ZN(n36197) );
  OAI22_X1 U34510 ( .A1(n3577), .A2(n32930), .B1(n36197), .B2(n36196), .ZN(
        n36261) );
  OAI21_X1 U34511 ( .B1(n36259), .B2(n36260), .A(n36261), .ZN(n32932) );
  NAND2_X1 U34512 ( .A1(n32932), .A2(n32931), .ZN(n36294) );
  FA_X1 U34513 ( .A(n32935), .B(n32934), .CI(n32933), .CO(n32944), .S(n36293)
         );
  XNOR2_X1 U34514 ( .A(n32937), .B(\fmem_data[19][1] ), .ZN(n36225) );
  OAI22_X1 U34515 ( .A1(n34345), .A2(n3633), .B1(n36225), .B2(n36226), .ZN(
        n36306) );
  XNOR2_X1 U34516 ( .A(n32938), .B(\fmem_data[1][1] ), .ZN(n33689) );
  OAI21_X1 U34517 ( .B1(n36306), .B2(n36305), .A(n36304), .ZN(n32943) );
  NAND2_X1 U34518 ( .A1(n32943), .A2(n32942), .ZN(n36292) );
  XNOR2_X1 U34519 ( .A(n32945), .B(n32944), .ZN(n32947) );
  XNOR2_X1 U34520 ( .A(n32947), .B(n32946), .ZN(n36409) );
  NAND2_X1 U34521 ( .A1(n34529), .A2(n32948), .ZN(n36327) );
  NAND2_X1 U34522 ( .A1(n36100), .A2(n32949), .ZN(n36326) );
  NAND2_X1 U34523 ( .A1(n34742), .A2(n32950), .ZN(n36325) );
  OR2_X1 U34524 ( .A1(n36228), .A2(n4018), .ZN(n32951) );
  NAND2_X1 U34525 ( .A1(n36227), .A2(n32951), .ZN(n36324) );
  NAND2_X1 U34526 ( .A1(n34625), .A2(n32952), .ZN(n36323) );
  XNOR2_X1 U34527 ( .A(n32953), .B(\fmem_data[26][1] ), .ZN(n33726) );
  OAI22_X1 U34528 ( .A1(n33726), .A2(n3678), .B1(n36111), .B2(n33725), .ZN(
        n36322) );
  NAND2_X1 U34529 ( .A1(n34476), .A2(n32954), .ZN(n36342) );
  NAND2_X1 U34530 ( .A1(n36104), .A2(n32955), .ZN(n36341) );
  NAND2_X1 U34531 ( .A1(n34483), .A2(n32956), .ZN(n36340) );
  INV_X1 U34532 ( .A(n36290), .ZN(n32971) );
  FA_X1 U34533 ( .A(n32959), .B(n32958), .CI(n32957), .CO(n33500), .S(n36351)
         );
  XNOR2_X1 U34534 ( .A(n33789), .B(\fmem_data[30][1] ), .ZN(n34789) );
  FA_X1 U34535 ( .A(n32962), .B(n32961), .CI(n32960), .CO(n33497), .S(n36352)
         );
  OAI21_X1 U34536 ( .B1(n36351), .B2(n36350), .A(n36352), .ZN(n32963) );
  NAND2_X1 U34537 ( .A1(n32964), .A2(n32963), .ZN(n36288) );
  XNOR2_X1 U34538 ( .A(n32966), .B(n32965), .ZN(n32968) );
  XNOR2_X1 U34539 ( .A(n32968), .B(n32967), .ZN(n36289) );
  NOR2_X1 U34540 ( .A1(n36288), .A2(n36289), .ZN(n32970) );
  OAI21_X1 U34541 ( .B1(n32971), .B2(n32970), .A(n32969), .ZN(n36411) );
  OAI21_X1 U34542 ( .B1(n36410), .B2(n36409), .A(n36411), .ZN(n32973) );
  NAND2_X1 U34543 ( .A1(n36409), .A2(n36410), .ZN(n32972) );
  NAND2_X1 U34544 ( .A1(n32973), .A2(n32972), .ZN(n36286) );
  XNOR2_X1 U34545 ( .A(n3260), .B(\fmem_data[27][1] ), .ZN(n33735) );
  XNOR2_X1 U34546 ( .A(n34334), .B(\fmem_data[27][1] ), .ZN(n36239) );
  OAI22_X1 U34547 ( .A1(n3482), .A2(n33735), .B1(n36239), .B2(n36240), .ZN(
        n36252) );
  XNOR2_X1 U34548 ( .A(n33803), .B(\fmem_data[24][1] ), .ZN(n34771) );
  OAI22_X2 U34549 ( .A1(n36102), .A2(n36100), .B1(n34771), .B2(n3565), .ZN(
        n36254) );
  NAND2_X1 U34550 ( .A1(n36252), .A2(n36254), .ZN(n32983) );
  OAI22_X1 U34551 ( .A1(n34600), .A2(n34598), .B1(n32980), .B2(n3569), .ZN(
        n36253) );
  NAND2_X1 U34552 ( .A1(n36252), .A2(n36253), .ZN(n32982) );
  NAND2_X1 U34553 ( .A1(n36254), .A2(n36253), .ZN(n32981) );
  NAND3_X1 U34554 ( .A1(n32983), .A2(n32982), .A3(n32981), .ZN(n36358) );
  FA_X1 U34555 ( .A(n32986), .B(n32985), .CI(n32984), .CO(n32946), .S(n36357)
         );
  FA_X1 U34556 ( .A(n32989), .B(n32988), .CI(n32987), .CO(n32977), .S(n36359)
         );
  OAI21_X1 U34557 ( .B1(n36358), .B2(n36357), .A(n36359), .ZN(n32991) );
  NAND2_X1 U34558 ( .A1(n36358), .A2(n36357), .ZN(n32990) );
  NAND2_X1 U34559 ( .A1(n32991), .A2(n32990), .ZN(n36320) );
  OAI21_X1 U34560 ( .B1(n36284), .B2(n36286), .A(n36285), .ZN(n32997) );
  NAND2_X1 U34561 ( .A1(n36284), .A2(n36286), .ZN(n32996) );
  NAND2_X1 U34562 ( .A1(n32997), .A2(n32996), .ZN(n36283) );
  FA_X1 U34563 ( .A(n33000), .B(n32999), .CI(n32998), .CO(n32856), .S(n36282)
         );
  FA_X1 U34564 ( .A(n33003), .B(n33002), .CI(n33001), .CO(n32920), .S(n36281)
         );
  OAI21_X1 U34565 ( .B1(n36374), .B2(n36373), .A(n36376), .ZN(n33005) );
  NAND2_X1 U34566 ( .A1(n36374), .A2(n36373), .ZN(n33004) );
  NAND2_X1 U34567 ( .A1(n33005), .A2(n33004), .ZN(n36157) );
  XNOR2_X1 U34568 ( .A(n33007), .B(n33006), .ZN(n33009) );
  FA_X1 U34569 ( .A(n33012), .B(n33011), .CI(n33010), .CO(n33414), .S(n36151)
         );
  OAI21_X1 U34570 ( .B1(n36150), .B2(n36149), .A(n36151), .ZN(n33014) );
  NAND2_X1 U34571 ( .A1(n36150), .A2(n36149), .ZN(n33013) );
  NAND2_X1 U34572 ( .A1(n33014), .A2(n33013), .ZN(n36034) );
  OAI21_X1 U34573 ( .B1(n36032), .B2(n36033), .A(n36034), .ZN(n33015) );
  NAND2_X1 U34574 ( .A1(n33015), .A2(n33016), .ZN(n36027) );
  INV_X1 U34575 ( .A(n33018), .ZN(n33144) );
  FA_X1 U34576 ( .A(n33023), .B(n33022), .CI(n33021), .CO(n33142), .S(n33222)
         );
  FA_X1 U34577 ( .A(n33026), .B(n33025), .CI(n33024), .CO(n33121), .S(n32813)
         );
  OAI22_X1 U34578 ( .A1(n33030), .A2(n34918), .B1(n33029), .B2(n34919), .ZN(
        n33137) );
  OAI22_X1 U34579 ( .A1(n33034), .A2(n35006), .B1(n33033), .B2(n35007), .ZN(
        n33065) );
  OAI22_X1 U34580 ( .A1(n33036), .A2(n33681), .B1(n33035), .B2(n33679), .ZN(
        n33064) );
  OAI22_X1 U34581 ( .A1(n33042), .A2(n34986), .B1(n33041), .B2(n34985), .ZN(
        n33080) );
  OAI22_X1 U34582 ( .A1(n33044), .A2(n33873), .B1(n33043), .B2(n33875), .ZN(
        n33079) );
  OAI22_X1 U34583 ( .A1(n33046), .A2(n35034), .B1(n33045), .B2(n35033), .ZN(
        n33078) );
  FA_X1 U34584 ( .A(n33049), .B(n33048), .CI(n33047), .CO(n33362), .S(n33221)
         );
  XNOR2_X1 U34585 ( .A(n33055), .B(\fmem_data[4][3] ), .ZN(n33175) );
  OAI22_X1 U34586 ( .A1(n33056), .A2(n33174), .B1(n33175), .B2(n33176), .ZN(
        n33238) );
  OAI22_X1 U34587 ( .A1(n33060), .A2(n33059), .B1(n33058), .B2(n33057), .ZN(
        n33237) );
  OAI22_X1 U34588 ( .A1(n33062), .A2(n34206), .B1(n34208), .B2(n33061), .ZN(
        n33236) );
  FA_X1 U34589 ( .A(n33065), .B(n33064), .CI(n33063), .CO(n33376), .S(n33070)
         );
  FA_X1 U34590 ( .A(n33068), .B(n33067), .CI(n33066), .CO(n33069), .S(n32343)
         );
  FA_X1 U34591 ( .A(n33071), .B(n33070), .CI(n33069), .CO(n33389), .S(n33284)
         );
  FA_X1 U34592 ( .A(n33072), .B(n33073), .CI(n33074), .CO(n33213), .S(n32723)
         );
  FA_X1 U34593 ( .A(n33077), .B(n33076), .CI(n33075), .CO(n33212), .S(n33278)
         );
  FA_X1 U34594 ( .A(n33080), .B(n33079), .CI(n33078), .CO(n33374), .S(n33211)
         );
  FA_X1 U34595 ( .A(n33083), .B(n33081), .CI(n33082), .CO(n33118), .S(n33282)
         );
  XNOR2_X1 U34596 ( .A(n33085), .B(n33084), .ZN(n33087) );
  XNOR2_X1 U34597 ( .A(n33087), .B(n33086), .ZN(n33153) );
  NAND2_X1 U34598 ( .A1(n33092), .A2(n33091), .ZN(n33152) );
  OAI21_X1 U34599 ( .B1(n33095), .B2(n33094), .A(n33093), .ZN(n33097) );
  NAND2_X1 U34600 ( .A1(n33095), .A2(n33094), .ZN(n33096) );
  NAND2_X1 U34601 ( .A1(n33097), .A2(n33096), .ZN(n35057) );
  XNOR2_X1 U34602 ( .A(n35058), .B(n35057), .ZN(n33151) );
  FA_X1 U34603 ( .A(n33109), .B(n33108), .CI(n33107), .CO(n34976), .S(n33115)
         );
  XNOR2_X1 U34604 ( .A(n34975), .B(n34976), .ZN(n33113) );
  FA_X1 U34605 ( .A(n33112), .B(n33111), .CI(n33110), .CO(n34977), .S(n33119)
         );
  XNOR2_X1 U34606 ( .A(n33113), .B(n34977), .ZN(n35052) );
  FA_X1 U34607 ( .A(n33116), .B(n33115), .CI(n33114), .CO(n35051), .S(n33085)
         );
  FA_X1 U34608 ( .A(n33119), .B(n33118), .CI(n33117), .CO(n35050), .S(n33086)
         );
  FA_X1 U34609 ( .A(n33122), .B(n33121), .CI(n33120), .CO(n34999), .S(n33399)
         );
  FA_X1 U34610 ( .A(n33125), .B(n33124), .CI(n33123), .CO(n34997), .S(n33114)
         );
  XNOR2_X1 U34611 ( .A(n35073), .B(\fmem_data[22][5] ), .ZN(n33223) );
  XNOR2_X1 U34612 ( .A(n35357), .B(\fmem_data[29][5] ), .ZN(n35086) );
  OAI22_X1 U34613 ( .A1(n33135), .A2(n35655), .B1(n33134), .B2(n35656), .ZN(
        n35044) );
  XNOR2_X1 U34614 ( .A(n34999), .B(n34998), .ZN(n33146) );
  FA_X1 U34615 ( .A(n33138), .B(n33137), .CI(n33136), .CO(n35027), .S(n33120)
         );
  FA_X1 U34616 ( .A(n33141), .B(n33140), .CI(n33139), .CO(n35026), .S(n33116)
         );
  XNOR2_X1 U34617 ( .A(n35027), .B(n35026), .ZN(n33145) );
  FA_X1 U34618 ( .A(n33144), .B(n33143), .CI(n33142), .CO(n35025), .S(n33122)
         );
  XNOR2_X1 U34619 ( .A(n33145), .B(n35025), .ZN(n35000) );
  XNOR2_X1 U34620 ( .A(n33146), .B(n35000), .ZN(n34959) );
  XNOR2_X1 U34621 ( .A(n34960), .B(n34959), .ZN(n33150) );
  FA_X1 U34622 ( .A(n33149), .B(n33148), .CI(n33147), .CO(n34958), .S(n33093)
         );
  XNOR2_X1 U34623 ( .A(n33151), .B(n35059), .ZN(n34964) );
  FA_X1 U34624 ( .A(n33154), .B(n33153), .CI(n33152), .CO(n35058), .S(n34816)
         );
  FA_X1 U34625 ( .A(n33157), .B(n33156), .CI(n33155), .CO(n34679), .S(n33289)
         );
  OAI22_X1 U34626 ( .A1(n33159), .A2(n34199), .B1(n33158), .B2(n34201), .ZN(
        n33202) );
  INV_X1 U34627 ( .A(n34598), .ZN(n33160) );
  NOR2_X1 U34628 ( .A1(n33160), .A2(\fmem_data[4][0] ), .ZN(n33161) );
  OR2_X1 U34629 ( .A1(n33162), .A2(n33161), .ZN(n33201) );
  FA_X1 U34630 ( .A(n33173), .B(n33172), .CI(n33171), .CO(n34221), .S(n32763)
         );
  OAI22_X1 U34631 ( .A1(n33177), .A2(n33176), .B1(n33175), .B2(n33174), .ZN(
        n33262) );
  AOI21_X1 U34632 ( .B1(n34440), .B2(n3483), .A(n33178), .ZN(n33179) );
  INV_X1 U34633 ( .A(n33179), .ZN(n33261) );
  OAI22_X1 U34634 ( .A1(n33924), .A2(n35515), .B1(n33182), .B2(n35516), .ZN(
        n33193) );
  OAI22_X1 U34635 ( .A1(n33190), .A2(n34779), .B1(n33189), .B2(n34466), .ZN(
        n33230) );
  FA_X1 U34636 ( .A(n33193), .B(n33192), .CI(n33191), .CO(n33229), .S(n34219)
         );
  INV_X1 U34637 ( .A(n36227), .ZN(n33194) );
  NOR2_X1 U34638 ( .A1(n33194), .A2(\fmem_data[20][0] ), .ZN(n33195) );
  INV_X1 U34639 ( .A(n33198), .ZN(n33259) );
  XNOR2_X1 U34640 ( .A(n33202), .B(n33201), .ZN(n33204) );
  XNOR2_X1 U34641 ( .A(n33204), .B(n33203), .ZN(n34217) );
  FA_X1 U34642 ( .A(n33207), .B(n33206), .CI(n33205), .CO(n34216), .S(n34395)
         );
  FA_X1 U34643 ( .A(n33210), .B(n33209), .CI(n33208), .CO(n33285), .S(n34676)
         );
  FA_X1 U34644 ( .A(n33213), .B(n33212), .CI(n33211), .CO(n33337), .S(n33283)
         );
  XNOR2_X1 U34645 ( .A(n33214), .B(\fmem_data[24][5] ), .ZN(n33370) );
  OAI22_X1 U34646 ( .A1(n33217), .A2(n35701), .B1(n33216), .B2(n35700), .ZN(
        n33301) );
  OAI22_X1 U34647 ( .A1(n33219), .A2(n34923), .B1(n33218), .B2(n34922), .ZN(
        n33300) );
  FA_X1 U34648 ( .A(n33222), .B(n33221), .CI(n33220), .CO(n33335), .S(n32811)
         );
  XNOR2_X1 U34649 ( .A(n33225), .B(\fmem_data[16][7] ), .ZN(n34863) );
  FA_X1 U34650 ( .A(n33231), .B(n33230), .CI(n33229), .CO(n33350), .S(n33287)
         );
  FA_X1 U34651 ( .A(n33237), .B(n33238), .CI(n33236), .CO(n33331), .S(n33071)
         );
  FA_X1 U34652 ( .A(n33245), .B(n33244), .CI(n33243), .CO(n33353), .S(n34678)
         );
  XNOR2_X1 U34653 ( .A(n33246), .B(\fmem_data[25][7] ), .ZN(n34860) );
  INV_X1 U34654 ( .A(n33251), .ZN(n33378) );
  XNOR2_X1 U34655 ( .A(n33394), .B(n33393), .ZN(n33281) );
  FA_X1 U34656 ( .A(n32753), .B(n33255), .CI(n33254), .CO(n33340), .S(n33156)
         );
  FA_X1 U34657 ( .A(n3705), .B(n33259), .CI(n33258), .CO(n33338), .S(n34218)
         );
  FA_X1 U34658 ( .A(n33262), .B(n33261), .CI(n33260), .CO(n33346), .S(n34220)
         );
  AOI21_X1 U34659 ( .B1(n34625), .B2(n3574), .A(n33263), .ZN(n33264) );
  INV_X1 U34660 ( .A(n33264), .ZN(n34096) );
  AOI21_X1 U34661 ( .B1(n36104), .B2(n3580), .A(n33265), .ZN(n33266) );
  INV_X1 U34662 ( .A(n33266), .ZN(n34095) );
  OAI22_X1 U34663 ( .A1(n33268), .A2(n35610), .B1(n33267), .B2(n35611), .ZN(
        n34094) );
  OR2_X1 U34664 ( .A1(n33277), .A2(n33278), .ZN(n33276) );
  NAND2_X1 U34665 ( .A1(n33276), .A2(n33275), .ZN(n33280) );
  NAND2_X1 U34666 ( .A1(n33280), .A2(n33279), .ZN(n34671) );
  XNOR2_X1 U34667 ( .A(n33281), .B(n33392), .ZN(n33360) );
  FA_X1 U34668 ( .A(n33283), .B(n33284), .CI(n33282), .CO(n33397), .S(n34703)
         );
  FA_X1 U34669 ( .A(n33287), .B(n33286), .CI(n33285), .CO(n33357), .S(n34702)
         );
  OAI21_X1 U34670 ( .B1(n33290), .B2(n33289), .A(n33288), .ZN(n33292) );
  NAND2_X1 U34671 ( .A1(n33292), .A2(n33291), .ZN(n34701) );
  OAI21_X1 U34672 ( .B1(n33294), .B2(n33295), .A(n33293), .ZN(n33297) );
  NAND2_X1 U34673 ( .A1(n33295), .A2(n33294), .ZN(n33296) );
  NAND2_X1 U34674 ( .A1(n33297), .A2(n33296), .ZN(n34815) );
  OAI21_X1 U34675 ( .B1(n34816), .B2(n34814), .A(n34815), .ZN(n33299) );
  NAND2_X1 U34676 ( .A1(n34816), .A2(n34814), .ZN(n33298) );
  NAND2_X1 U34677 ( .A1(n33299), .A2(n33298), .ZN(n34965) );
  FA_X1 U34678 ( .A(n33302), .B(n33301), .CI(n33300), .CO(n34916), .S(n33336)
         );
  OAI22_X1 U34679 ( .A1(n33323), .A2(n33828), .B1(n33322), .B2(n33827), .ZN(
        n34831) );
  OAI22_X1 U34680 ( .A1(n33329), .A2(n33328), .B1(n33327), .B2(n33326), .ZN(
        n34832) );
  XNOR2_X1 U34681 ( .A(n34826), .B(n34825), .ZN(n33334) );
  FA_X1 U34682 ( .A(n33333), .B(n33332), .CI(n33331), .CO(n34824), .S(n33349)
         );
  XNOR2_X1 U34683 ( .A(n33334), .B(n34824), .ZN(n34852) );
  FA_X1 U34684 ( .A(n33337), .B(n33336), .CI(n33335), .CO(n34851), .S(n33356)
         );
  FA_X1 U34685 ( .A(n33340), .B(n33339), .CI(n33338), .CO(n34693), .S(n34673)
         );
  FA_X1 U34686 ( .A(n33343), .B(n33342), .CI(n33341), .CO(n35081), .S(n34691)
         );
  FA_X1 U34687 ( .A(n33346), .B(n33345), .CI(n33344), .CO(n34692), .S(n34672)
         );
  FA_X1 U34688 ( .A(n33351), .B(n33350), .CI(n33349), .CO(n34847), .S(n33394)
         );
  XNOR2_X1 U34689 ( .A(n34848), .B(n34847), .ZN(n33355) );
  FA_X1 U34690 ( .A(n33354), .B(n33353), .CI(n33352), .CO(n34846), .S(n33393)
         );
  XNOR2_X1 U34691 ( .A(n33355), .B(n34846), .ZN(n34892) );
  FA_X1 U34692 ( .A(n33358), .B(n33357), .CI(n33356), .CO(n34891), .S(n33361)
         );
  FA_X1 U34693 ( .A(n33361), .B(n33360), .CI(n33359), .CO(n34894), .S(n34814)
         );
  XNOR2_X1 U34694 ( .A(n34896), .B(n34894), .ZN(n33400) );
  INV_X1 U34695 ( .A(n33362), .ZN(n33367) );
  NOR2_X1 U34696 ( .A1(n33364), .A2(n33363), .ZN(n33366) );
  NAND2_X1 U34697 ( .A1(n33364), .A2(n33363), .ZN(n33365) );
  OAI21_X1 U34698 ( .B1(n33367), .B2(n33366), .A(n33365), .ZN(n34845) );
  OAI22_X1 U34699 ( .A1(n33369), .A2(n33954), .B1(n33956), .B2(n33368), .ZN(
        n34938) );
  FA_X1 U34700 ( .A(n33376), .B(n33375), .CI(n33374), .CO(n34843), .S(n33391)
         );
  FA_X1 U34701 ( .A(n33379), .B(n33378), .CI(n33377), .CO(n34901), .S(n33352)
         );
  FA_X1 U34702 ( .A(n33382), .B(n33381), .CI(n33380), .CO(n34900), .S(n33351)
         );
  FA_X1 U34703 ( .A(n33391), .B(n33390), .CI(n33389), .CO(n34951), .S(n33398)
         );
  FA_X1 U34704 ( .A(n33397), .B(n33398), .CI(n33399), .CO(n34955), .S(n33154)
         );
  XNOR2_X1 U34705 ( .A(n33400), .B(n34895), .ZN(n34966) );
  XNOR2_X1 U34706 ( .A(n34965), .B(n34966), .ZN(n33401) );
  XNOR2_X1 U34707 ( .A(n34964), .B(n33401), .ZN(n36026) );
  FA_X1 U34708 ( .A(n33404), .B(n33403), .CI(n33402), .CO(n35456), .S(n36025)
         );
  NOR2_X1 U34709 ( .A1(n36440), .A2(n36439), .ZN(n34823) );
  XNOR2_X1 U34710 ( .A(n33406), .B(n33405), .ZN(n33408) );
  XNOR2_X1 U34711 ( .A(n33408), .B(n33407), .ZN(n36649) );
  FA_X1 U34712 ( .A(n33411), .B(n33410), .CI(n33409), .CO(n33407), .S(n36639)
         );
  XNOR2_X1 U34713 ( .A(n33413), .B(n33412), .ZN(n33415) );
  XNOR2_X1 U34714 ( .A(n33415), .B(n33414), .ZN(n36637) );
  FA_X1 U34715 ( .A(n33417), .B(n33418), .CI(n33416), .CO(n33409), .S(n36628)
         );
  FA_X1 U34716 ( .A(n33421), .B(n33420), .CI(n33419), .CO(n33010), .S(n36379)
         );
  FA_X1 U34717 ( .A(n33424), .B(n33423), .CI(n33422), .CO(n33524), .S(n36277)
         );
  FA_X1 U34718 ( .A(n33427), .B(n33426), .CI(n33425), .CO(n33422), .S(n36280)
         );
  FA_X1 U34719 ( .A(n33430), .B(n33429), .CI(n33428), .CO(n32922), .S(n36279)
         );
  FA_X1 U34720 ( .A(n33433), .B(n33432), .CI(n33431), .CO(n33426), .S(n36368)
         );
  FA_X1 U34721 ( .A(n33436), .B(n33435), .CI(n33434), .CO(n33428), .S(n36367)
         );
  FA_X1 U34722 ( .A(n33439), .B(n33438), .CI(n33437), .CO(n33535), .S(n36470)
         );
  FA_X1 U34723 ( .A(n33442), .B(n33441), .CI(n33440), .CO(n33513), .S(n36469)
         );
  FA_X1 U34724 ( .A(n33445), .B(n33444), .CI(n33443), .CO(n33440), .S(n36402)
         );
  FA_X1 U34725 ( .A(n33448), .B(n33447), .CI(n33446), .CO(n32989), .S(n36334)
         );
  OAI22_X1 U34726 ( .A1(n33449), .A2(n3483), .B1(n36110), .B2(n34440), .ZN(
        n36345) );
  NAND2_X1 U34727 ( .A1(n33725), .A2(n33450), .ZN(n36344) );
  XNOR2_X1 U34728 ( .A(n33451), .B(\fmem_data[9][1] ), .ZN(n33744) );
  OAI22_X1 U34729 ( .A1(n33744), .A2(n3579), .B1(n34476), .B2(n3365), .ZN(
        n36343) );
  OAI21_X1 U34730 ( .B1(n36345), .B2(n36344), .A(n36343), .ZN(n33453) );
  NAND2_X1 U34731 ( .A1(n36345), .A2(n36344), .ZN(n33452) );
  NAND2_X1 U34732 ( .A1(n33453), .A2(n33452), .ZN(n36335) );
  NAND3_X1 U34733 ( .A1(n3389), .A2(n33454), .A3(n3945), .ZN(n33457) );
  OR2_X1 U34734 ( .A1(n3389), .A2(n3945), .ZN(n33456) );
  NAND3_X1 U34735 ( .A1(n33458), .A2(n33457), .A3(n33456), .ZN(n36219) );
  XNOR2_X1 U34736 ( .A(n3313), .B(\fmem_data[7][1] ), .ZN(n33699) );
  OAI22_X1 U34737 ( .A1(n36219), .A2(n36218), .B1(n3581), .B2(n33699), .ZN(
        n36333) );
  OAI21_X1 U34738 ( .B1(n36334), .B2(n36335), .A(n36333), .ZN(n33461) );
  NAND2_X1 U34739 ( .A1(n36334), .A2(n36335), .ZN(n33460) );
  NAND2_X1 U34740 ( .A1(n33461), .A2(n33460), .ZN(n36403) );
  FA_X1 U34741 ( .A(n33464), .B(n33463), .CI(n33462), .CO(n33494), .S(n36356)
         );
  NAND3_X1 U34742 ( .A1(n33466), .A2(n33465), .A3(\fmem_data[4][1] ), .ZN(
        n33467) );
  NAND2_X1 U34743 ( .A1(n34598), .A2(n33467), .ZN(n36303) );
  OR2_X1 U34744 ( .A1(n34612), .A2(n3682), .ZN(n33468) );
  NAND2_X1 U34745 ( .A1(n34017), .A2(n33468), .ZN(n36302) );
  NAND2_X1 U34746 ( .A1(n34745), .A2(n33469), .ZN(n36301) );
  NOR2_X1 U34747 ( .A1(n33475), .A2(n33474), .ZN(n36468) );
  FA_X1 U34748 ( .A(n33478), .B(n33477), .CI(n33476), .CO(n33613), .S(n36389)
         );
  XNOR2_X1 U34749 ( .A(n33479), .B(\fmem_data[15][1] ), .ZN(n36222) );
  OAI22_X1 U34750 ( .A1(n36222), .A2(n36223), .B1(n3568), .B2(n33480), .ZN(
        n36349) );
  NAND2_X1 U34751 ( .A1(n34440), .A2(n33481), .ZN(n36310) );
  OAI21_X1 U34752 ( .B1(n36296), .B2(n4020), .A(n36295), .ZN(n36309) );
  NAND2_X1 U34753 ( .A1(n34343), .A2(n33482), .ZN(n36308) );
  XNOR2_X1 U34754 ( .A(n33483), .B(\fmem_data[31][1] ), .ZN(n36211) );
  XNOR2_X1 U34755 ( .A(n33484), .B(\fmem_data[31][1] ), .ZN(n33701) );
  OAI22_X1 U34756 ( .A1(n36211), .A2(n36216), .B1(n33701), .B2(n3931), .ZN(
        n36347) );
  XNOR2_X1 U34757 ( .A(n33486), .B(n33485), .ZN(n33488) );
  XNOR2_X1 U34758 ( .A(n33488), .B(n33487), .ZN(n36407) );
  XNOR2_X1 U34759 ( .A(n33490), .B(n33489), .ZN(n33492) );
  XNOR2_X1 U34760 ( .A(n33492), .B(n33491), .ZN(n36406) );
  FA_X1 U34761 ( .A(n33495), .B(n33494), .CI(n33493), .CO(n33505), .S(n36400)
         );
  FA_X1 U34762 ( .A(n33498), .B(n33497), .CI(n33496), .CO(n33437), .S(n36398)
         );
  FA_X1 U34763 ( .A(n33501), .B(n33500), .CI(n33499), .CO(n33442), .S(n36399)
         );
  OAI21_X1 U34764 ( .B1(n36400), .B2(n36398), .A(n36399), .ZN(n33503) );
  NAND2_X1 U34765 ( .A1(n36400), .A2(n36398), .ZN(n33502) );
  NAND2_X1 U34766 ( .A1(n33503), .A2(n33502), .ZN(n36413) );
  FA_X1 U34767 ( .A(n33506), .B(n33505), .CI(n33504), .CO(n33534), .S(n36415)
         );
  OAI21_X1 U34768 ( .B1(n36414), .B2(n36413), .A(n36415), .ZN(n33508) );
  NAND2_X1 U34769 ( .A1(n36414), .A2(n36413), .ZN(n33507) );
  NAND2_X1 U34770 ( .A1(n33508), .A2(n33507), .ZN(n36393) );
  XNOR2_X1 U34771 ( .A(n33510), .B(n33509), .ZN(n33512) );
  XNOR2_X1 U34772 ( .A(n33512), .B(n33511), .ZN(n36392) );
  FA_X1 U34773 ( .A(n33515), .B(n33514), .CI(n33513), .CO(n33518), .S(n36391)
         );
  OAI21_X1 U34774 ( .B1(n36393), .B2(n36392), .A(n36391), .ZN(n33517) );
  NAND2_X1 U34775 ( .A1(n33517), .A2(n33516), .ZN(n36388) );
  FA_X1 U34776 ( .A(n33520), .B(n33519), .CI(n33518), .CO(n33612), .S(n36387)
         );
  OAI21_X1 U34777 ( .B1(n36389), .B2(n36388), .A(n36387), .ZN(n33522) );
  NAND2_X1 U34778 ( .A1(n33522), .A2(n33521), .ZN(n36275) );
  FA_X1 U34779 ( .A(n33525), .B(n33524), .CI(n33523), .CO(n33417), .S(n36380)
         );
  OAI21_X1 U34780 ( .B1(n36379), .B2(n36381), .A(n36380), .ZN(n33527) );
  NAND2_X1 U34781 ( .A1(n36381), .A2(n36379), .ZN(n33526) );
  NAND2_X1 U34782 ( .A1(n33527), .A2(n33526), .ZN(n36627) );
  FA_X1 U34783 ( .A(n33530), .B(n33529), .CI(n33528), .CO(n33519), .S(n36397)
         );
  FA_X1 U34784 ( .A(n33533), .B(n33532), .CI(n33531), .CO(n33520), .S(n36396)
         );
  FA_X1 U34785 ( .A(n33539), .B(n33538), .CI(n33537), .CO(n33610), .S(n36419)
         );
  FA_X1 U34786 ( .A(n33546), .B(n33545), .CI(n33544), .CO(n33562), .S(n36484)
         );
  XNOR2_X1 U34787 ( .A(n33548), .B(n33547), .ZN(n33549) );
  XNOR2_X1 U34788 ( .A(n33550), .B(n33549), .ZN(n36482) );
  XNOR2_X1 U34789 ( .A(n33551), .B(\fmem_data[20][1] ), .ZN(n36229) );
  XNOR2_X1 U34790 ( .A(n33553), .B(\fmem_data[5][1] ), .ZN(n34484) );
  XNOR2_X1 U34791 ( .A(n33554), .B(\fmem_data[2][1] ), .ZN(n34344) );
  OAI22_X1 U34792 ( .A1(n34344), .A2(n3578), .B1(n3353), .B2(n34343), .ZN(
        n36329) );
  OAI22_X1 U34793 ( .A1(n36300), .A2(n36298), .B1(n33557), .B2(n3573), .ZN(
        n36471) );
  OAI21_X1 U34794 ( .B1(n36472), .B2(n36473), .A(n36471), .ZN(n33559) );
  NAND2_X1 U34795 ( .A1(n33559), .A2(n33558), .ZN(n36483) );
  FA_X1 U34796 ( .A(n33564), .B(n33563), .CI(n33562), .CO(n33541), .S(n36466)
         );
  FA_X1 U34797 ( .A(n33567), .B(n33566), .CI(n33565), .CO(n33542), .S(n36465)
         );
  OAI22_X1 U34798 ( .A1(n33571), .A2(n33570), .B1(n33569), .B2(n33568), .ZN(
        n33589) );
  INV_X1 U34799 ( .A(n35089), .ZN(n33572) );
  OAI22_X1 U34800 ( .A1(n33580), .A2(n36120), .B1(n33579), .B2(n3575), .ZN(
        n33696) );
  FA_X1 U34801 ( .A(n33586), .B(n33585), .CI(n33584), .CO(n31466), .S(n33661)
         );
  FA_X1 U34802 ( .A(n33589), .B(n33588), .CI(n33587), .CO(n33639), .S(n33769)
         );
  XNOR2_X1 U34803 ( .A(n36312), .B(\fmem_data[10][3] ), .ZN(n33591) );
  XNOR2_X1 U34804 ( .A(n33592), .B(\fmem_data[14][1] ), .ZN(n34738) );
  OAI22_X1 U34805 ( .A1(n33593), .A2(n3563), .B1(n34738), .B2(n34739), .ZN(
        n33715) );
  OAI21_X1 U34806 ( .B1(n36490), .B2(n36492), .A(n36489), .ZN(n33606) );
  NAND2_X1 U34807 ( .A1(n33606), .A2(n33605), .ZN(n36421) );
  OAI21_X1 U34808 ( .B1(n36420), .B2(n36419), .A(n36421), .ZN(n33608) );
  NAND2_X1 U34809 ( .A1(n33608), .A2(n33607), .ZN(n36385) );
  FA_X1 U34810 ( .A(n33611), .B(n33610), .CI(n33609), .CO(n33620), .S(n36383)
         );
  XNOR2_X1 U34811 ( .A(n33612), .B(n33613), .ZN(n33615) );
  XNOR2_X1 U34812 ( .A(n33615), .B(n33614), .ZN(n36384) );
  OAI21_X1 U34813 ( .B1(n36385), .B2(n36383), .A(n36384), .ZN(n33617) );
  NAND2_X1 U34814 ( .A1(n36385), .A2(n36383), .ZN(n33616) );
  NAND2_X1 U34815 ( .A1(n33617), .A2(n33616), .ZN(n36616) );
  FA_X1 U34816 ( .A(n33618), .B(n33619), .CI(n33620), .CO(n33416), .S(n36617)
         );
  FA_X1 U34817 ( .A(n33623), .B(n33622), .CI(n33621), .CO(n31625), .S(n34292)
         );
  FA_X1 U34818 ( .A(n33626), .B(n33625), .CI(n33624), .CO(n31626), .S(n34294)
         );
  XNOR2_X1 U34819 ( .A(n34292), .B(n34294), .ZN(n33656) );
  FA_X1 U34820 ( .A(n33629), .B(n33628), .CI(n33627), .CO(n34151), .S(n34174)
         );
  OAI21_X1 U34821 ( .B1(n33632), .B2(n33631), .A(n33630), .ZN(n33634) );
  NAND2_X1 U34822 ( .A1(n33634), .A2(n33633), .ZN(n34173) );
  XNOR2_X1 U34823 ( .A(n34174), .B(n34173), .ZN(n33655) );
  FA_X1 U34824 ( .A(n33637), .B(n33635), .CI(n33636), .CO(n33627), .S(n33665)
         );
  FA_X1 U34825 ( .A(n33639), .B(n3494), .CI(n33638), .CO(n33663), .S(n33662)
         );
  OAI22_X1 U34826 ( .A1(n33641), .A2(n3678), .B1(n33640), .B2(n33725), .ZN(
        n34067) );
  OR2_X1 U34827 ( .A1(n36296), .A2(n3629), .ZN(n33644) );
  OAI22_X1 U34828 ( .A1(n33644), .A2(n33643), .B1(n33642), .B2(n3629), .ZN(
        n34066) );
  INV_X1 U34829 ( .A(n34942), .ZN(n33647) );
  FA_X1 U34830 ( .A(n33652), .B(n33651), .CI(n33650), .CO(n34366), .S(n33767)
         );
  NAND2_X1 U34831 ( .A1(n33654), .A2(n33653), .ZN(n34172) );
  XNOR2_X1 U34832 ( .A(n33655), .B(n34172), .ZN(n34293) );
  XNOR2_X1 U34833 ( .A(n33656), .B(n34293), .ZN(n36425) );
  FA_X1 U34834 ( .A(n33659), .B(n33658), .CI(n33657), .CO(n33624), .S(n33917)
         );
  FA_X1 U34835 ( .A(n33662), .B(n33661), .CI(n33660), .CO(n33916), .S(n36489)
         );
  XNOR2_X1 U34836 ( .A(n33664), .B(n33663), .ZN(n33666) );
  XNOR2_X1 U34837 ( .A(n33666), .B(n33665), .ZN(n33915) );
  FA_X1 U34838 ( .A(n33669), .B(n33668), .CI(n33667), .CO(n33614), .S(n36455)
         );
  FA_X1 U34839 ( .A(n33672), .B(n33671), .CI(n33670), .CO(n31467), .S(n33819)
         );
  XNOR2_X1 U34840 ( .A(n33674), .B(n33673), .ZN(n33676) );
  OAI22_X1 U34841 ( .A1(n33682), .A2(n33681), .B1(n33680), .B2(n33679), .ZN(
        n33762) );
  XNOR2_X1 U34842 ( .A(n33683), .B(\fmem_data[24][3] ), .ZN(n34434) );
  FA_X1 U34843 ( .A(n33687), .B(n33686), .CI(n33685), .CO(n33670), .S(n33710)
         );
  XNOR2_X1 U34844 ( .A(n36315), .B(\fmem_data[3][3] ), .ZN(n33692) );
  XNOR2_X1 U34845 ( .A(n34783), .B(\fmem_data[3][3] ), .ZN(n34419) );
  OAI22_X1 U34846 ( .A1(n33692), .A2(n34418), .B1(n34419), .B2(n34420), .ZN(
        n33764) );
  OAI21_X1 U34847 ( .B1(n33711), .B2(n33710), .A(n33712), .ZN(n33694) );
  NAND2_X1 U34848 ( .A1(n33711), .A2(n33710), .ZN(n33693) );
  NAND2_X1 U34849 ( .A1(n33694), .A2(n33693), .ZN(n33817) );
  FA_X1 U34850 ( .A(n33697), .B(n33696), .CI(n33695), .CO(n33638), .S(n33836)
         );
  OR2_X1 U34851 ( .A1(n36315), .A2(n3642), .ZN(n33698) );
  OAI22_X1 U34852 ( .A1(n33698), .A2(n34420), .B1(n34418), .B2(n3642), .ZN(
        n33737) );
  OAI21_X1 U34853 ( .B1(n33737), .B2(n33738), .A(n33739), .ZN(n33704) );
  NAND2_X1 U34854 ( .A1(n33704), .A2(n33703), .ZN(n33835) );
  XNOR2_X1 U34855 ( .A(n33836), .B(n33835), .ZN(n33709) );
  INV_X1 U34856 ( .A(n34919), .ZN(n33705) );
  INV_X1 U34857 ( .A(n34835), .ZN(n33706) );
  AND2_X1 U34858 ( .A1(n36311), .A2(n33706), .ZN(n33821) );
  XNOR2_X1 U34859 ( .A(n33822), .B(n33821), .ZN(n33708) );
  INV_X1 U34860 ( .A(n34903), .ZN(n33707) );
  AND2_X1 U34861 ( .A1(n36316), .A2(n33707), .ZN(n33820) );
  XNOR2_X1 U34862 ( .A(n33708), .B(n33820), .ZN(n33837) );
  XNOR2_X1 U34863 ( .A(n33709), .B(n33837), .ZN(n36507) );
  XNOR2_X1 U34864 ( .A(n33711), .B(n33710), .ZN(n33713) );
  XNOR2_X1 U34865 ( .A(n33713), .B(n33712), .ZN(n36509) );
  FA_X1 U34866 ( .A(n33716), .B(n33715), .CI(n33714), .CO(n33768), .S(n36516)
         );
  FA_X1 U34867 ( .A(n33719), .B(n33718), .CI(n33717), .CO(n33565), .S(n36515)
         );
  XNOR2_X1 U34868 ( .A(n33720), .B(\fmem_data[3][1] ), .ZN(n34784) );
  OAI22_X1 U34869 ( .A1(n33721), .A2(n3582), .B1(n34784), .B2(n36199), .ZN(
        n34354) );
  OAI22_X1 U34870 ( .A1(n33722), .A2(n34505), .B1(n34503), .B2(n3685), .ZN(
        n34355) );
  XNOR2_X1 U34871 ( .A(n34354), .B(n34355), .ZN(n33728) );
  INV_X1 U34872 ( .A(n34435), .ZN(n33723) );
  OAI22_X1 U34873 ( .A1(n33726), .A2(n33725), .B1(n33724), .B2(n3678), .ZN(
        n34605) );
  INV_X1 U34874 ( .A(n34422), .ZN(n33727) );
  XNOR2_X1 U34875 ( .A(n33728), .B(n34353), .ZN(n36514) );
  OAI21_X1 U34876 ( .B1(n36507), .B2(n36509), .A(n36508), .ZN(n33730) );
  NAND2_X1 U34877 ( .A1(n33730), .A2(n33729), .ZN(n36462) );
  XNOR2_X1 U34878 ( .A(n36339), .B(\fmem_data[15][3] ), .ZN(n33732) );
  OAI22_X1 U34879 ( .A1(n33732), .A2(n34363), .B1(n33731), .B2(n34364), .ZN(
        n33816) );
  XNOR2_X1 U34880 ( .A(n36313), .B(\fmem_data[11][3] ), .ZN(n33734) );
  OAI22_X1 U34881 ( .A1(n33734), .A2(n34429), .B1(n34430), .B2(n34533), .ZN(
        n33815) );
  XNOR2_X1 U34882 ( .A(n33738), .B(n33737), .ZN(n33740) );
  XNOR2_X1 U34883 ( .A(n33740), .B(n33739), .ZN(n36601) );
  INV_X1 U34884 ( .A(n33741), .ZN(n33742) );
  XNOR2_X1 U34885 ( .A(n33743), .B(\fmem_data[9][1] ), .ZN(n34477) );
  OAI22_X1 U34886 ( .A1(n34477), .A2(n3579), .B1(n34476), .B2(n33744), .ZN(
        n34608) );
  INV_X1 U34887 ( .A(n34414), .ZN(n33745) );
  INV_X1 U34888 ( .A(n36505), .ZN(n33772) );
  XNOR2_X1 U34889 ( .A(n33749), .B(\fmem_data[13][1] ), .ZN(n34743) );
  OAI22_X1 U34890 ( .A1(n34743), .A2(n3571), .B1(n34742), .B2(n33800), .ZN(
        n36534) );
  OAI21_X1 U34891 ( .B1(n36534), .B2(n36533), .A(n36535), .ZN(n33753) );
  NAND2_X1 U34892 ( .A1(n33753), .A2(n33752), .ZN(n36479) );
  XNOR2_X1 U34893 ( .A(n33756), .B(\fmem_data[28][1] ), .ZN(n34746) );
  FA_X1 U34894 ( .A(n33763), .B(n33762), .CI(n33761), .CO(n33711), .S(n36487)
         );
  FA_X1 U34895 ( .A(n33766), .B(n33765), .CI(n33764), .CO(n33712), .S(n36486)
         );
  FA_X1 U34896 ( .A(n33769), .B(n33768), .CI(n33767), .CO(n33660), .S(n36503)
         );
  NOR2_X1 U34897 ( .A1(n36504), .A2(n36503), .ZN(n33771) );
  OAI21_X1 U34898 ( .B1(n33772), .B2(n33771), .A(n33770), .ZN(n36464) );
  OAI21_X1 U34899 ( .B1(n36461), .B2(n36462), .A(n36464), .ZN(n33774) );
  NAND2_X1 U34900 ( .A1(n36462), .A2(n36461), .ZN(n33773) );
  NAND2_X1 U34901 ( .A1(n33774), .A2(n33773), .ZN(n36454) );
  OAI21_X1 U34902 ( .B1(n36456), .B2(n36455), .A(n36454), .ZN(n33776) );
  NAND2_X1 U34903 ( .A1(n33776), .A2(n33775), .ZN(n36424) );
  INV_X1 U34904 ( .A(n34909), .ZN(n33779) );
  AND2_X1 U34905 ( .A1(n3116), .A2(n33779), .ZN(n33805) );
  OAI21_X1 U34906 ( .B1(n33807), .B2(n33805), .A(n33806), .ZN(n33783) );
  NAND2_X1 U34907 ( .A1(n33807), .A2(n33805), .ZN(n33782) );
  NAND2_X1 U34908 ( .A1(n33783), .A2(n33782), .ZN(n33908) );
  OAI22_X1 U34909 ( .A1(n33784), .A2(n35041), .B1(n35040), .B2(n3608), .ZN(
        n33901) );
  OAI22_X1 U34910 ( .A1(n34626), .A2(n33785), .B1(n35004), .B2(n3594), .ZN(
        n33900) );
  XNOR2_X1 U34911 ( .A(n33901), .B(n33900), .ZN(n33788) );
  XNOR2_X1 U34912 ( .A(n36111), .B(\fmem_data[26][5] ), .ZN(n33787) );
  XNOR2_X1 U34913 ( .A(n33788), .B(n33899), .ZN(n33911) );
  XNOR2_X1 U34914 ( .A(n33911), .B(n33910), .ZN(n33791) );
  XNOR2_X1 U34915 ( .A(n33908), .B(n33791), .ZN(n36062) );
  OAI22_X1 U34916 ( .A1(n33793), .A2(n3580), .B1(n33792), .B2(n36104), .ZN(
        n33870) );
  OAI22_X1 U34917 ( .A1(n33798), .A2(n33797), .B1(n3456), .B2(n33796), .ZN(
        n33983) );
  OR2_X1 U34918 ( .A1(n36101), .A2(n3651), .ZN(n33799) );
  OAI22_X1 U34919 ( .A1(n33801), .A2(n35182), .B1(n35181), .B2(n3612), .ZN(
        n33981) );
  XNOR2_X1 U34920 ( .A(n33982), .B(n33981), .ZN(n33802) );
  XNOR2_X1 U34921 ( .A(n3319), .B(n33802), .ZN(n33998) );
  OAI22_X1 U34922 ( .A1(n33804), .A2(n34431), .B1(n34432), .B2(n34433), .ZN(
        n33997) );
  XNOR2_X1 U34923 ( .A(n33808), .B(n33807), .ZN(n34574) );
  OAI22_X1 U34924 ( .A1(n33810), .A2(n34777), .B1(n33809), .B2(n3567), .ZN(
        n33842) );
  OAI22_X1 U34925 ( .A1(n33812), .A2(n34017), .B1(n33811), .B2(n3559), .ZN(
        n33841) );
  INV_X1 U34926 ( .A(n34990), .ZN(n33813) );
  FA_X1 U34927 ( .A(n33816), .B(n33815), .CI(n33814), .CO(n34572), .S(n36602)
         );
  INV_X1 U34928 ( .A(n34570), .ZN(n33865) );
  FA_X1 U34929 ( .A(n33819), .B(n33818), .CI(n33817), .CO(n34568), .S(n36461)
         );
  OAI21_X1 U34930 ( .B1(n33822), .B2(n33821), .A(n33820), .ZN(n33824) );
  OR2_X1 U34931 ( .A1(n34623), .A2(n3635), .ZN(n33825) );
  OAI22_X1 U34932 ( .A1(n33825), .A2(n33859), .B1(n33857), .B2(n3635), .ZN(
        n34107) );
  OAI22_X1 U34933 ( .A1(n36105), .A2(n33826), .B1(n35007), .B2(n3649), .ZN(
        n34106) );
  OR2_X1 U34934 ( .A1(n34624), .A2(n3650), .ZN(n33829) );
  OAI22_X1 U34935 ( .A1(n33829), .A2(n33828), .B1(n33827), .B2(n3650), .ZN(
        n34105) );
  INV_X1 U34936 ( .A(n34923), .ZN(n33830) );
  OAI22_X1 U34937 ( .A1(n33834), .A2(n34529), .B1(n33833), .B2(n3566), .ZN(
        n34507) );
  OAI21_X1 U34938 ( .B1(n33837), .B2(n33836), .A(n33835), .ZN(n33839) );
  NAND2_X1 U34939 ( .A1(n34639), .A2(n34640), .ZN(n33862) );
  FA_X1 U34940 ( .A(n33842), .B(n33841), .CI(n33840), .CO(n33883), .S(n34573)
         );
  XNOR2_X1 U34941 ( .A(n33844), .B(\fmem_data[9][5] ), .ZN(n33845) );
  OAI22_X1 U34942 ( .A1(n33846), .A2(n35041), .B1(n33845), .B2(n35040), .ZN(
        n33897) );
  XNOR2_X1 U34943 ( .A(n3354), .B(\fmem_data[2][5] ), .ZN(n33847) );
  OAI22_X1 U34944 ( .A1(n33848), .A2(n35019), .B1(n33847), .B2(n35018), .ZN(
        n33896) );
  OAI22_X1 U34945 ( .A1(n33852), .A2(n33851), .B1(n33850), .B2(n33849), .ZN(
        n34215) );
  OAI21_X1 U34946 ( .B1(n34639), .B2(n34640), .A(n34641), .ZN(n33861) );
  NAND2_X1 U34947 ( .A1(n33862), .A2(n33861), .ZN(n34569) );
  NOR2_X1 U34948 ( .A1(n34568), .A2(n34569), .ZN(n33864) );
  OAI21_X1 U34949 ( .B1(n33865), .B2(n33864), .A(n33863), .ZN(n34299) );
  OAI22_X1 U34950 ( .A1(n33867), .A2(n36221), .B1(n33866), .B2(n3558), .ZN(
        n34141) );
  FA_X1 U34951 ( .A(n33870), .B(n33869), .CI(n33868), .CO(n34140), .S(n33999)
         );
  OAI22_X1 U34952 ( .A1(n36199), .A2(n33872), .B1(n3582), .B2(n33871), .ZN(
        n34139) );
  OAI22_X1 U34953 ( .A1(n33876), .A2(n33875), .B1(n33874), .B2(n33873), .ZN(
        n34015) );
  OAI22_X1 U34954 ( .A1(n33880), .A2(n34945), .B1(n33879), .B2(n34944), .ZN(
        n34013) );
  FA_X1 U34955 ( .A(n33883), .B(n33882), .CI(n33881), .CO(n34331), .S(n34641)
         );
  FA_X1 U34956 ( .A(n33888), .B(n33887), .CI(n33886), .CO(n34149), .S(n34155)
         );
  XNOR2_X1 U34957 ( .A(n34156), .B(n34155), .ZN(n33914) );
  NAND2_X1 U34958 ( .A1(n33891), .A2(n33890), .ZN(n33892) );
  OAI22_X1 U34959 ( .A1(n33895), .A2(n34418), .B1(n33894), .B2(n34420), .ZN(
        n34090) );
  FA_X1 U34960 ( .A(n33898), .B(n33897), .CI(n33896), .CO(n34089), .S(n33882)
         );
  OAI21_X1 U34961 ( .B1(n33901), .B2(n33900), .A(n33899), .ZN(n33903) );
  NAND2_X1 U34962 ( .A1(n33903), .A2(n33902), .ZN(n34085) );
  OAI22_X1 U34963 ( .A1(n33905), .A2(n36241), .B1(n3662), .B2(n33904), .ZN(
        n34084) );
  OAI22_X1 U34964 ( .A1(n33907), .A2(n34468), .B1(n33906), .B2(n34470), .ZN(
        n34083) );
  OR2_X1 U34965 ( .A1(n33910), .A2(n33911), .ZN(n33909) );
  NAND2_X1 U34966 ( .A1(n33909), .A2(n33908), .ZN(n33913) );
  NAND2_X1 U34967 ( .A1(n33913), .A2(n33912), .ZN(n34324) );
  XNOR2_X1 U34968 ( .A(n33914), .B(n34154), .ZN(n34298) );
  FA_X1 U34969 ( .A(n33917), .B(n33916), .CI(n33915), .CO(n34297), .S(n36456)
         );
  OAI21_X1 U34970 ( .B1(n36616), .B2(n36617), .A(n36618), .ZN(n33919) );
  NAND2_X1 U34971 ( .A1(n36617), .A2(n36616), .ZN(n33918) );
  NAND2_X1 U34972 ( .A1(n33919), .A2(n33918), .ZN(n36629) );
  OAI21_X1 U34973 ( .B1(n36628), .B2(n36627), .A(n36629), .ZN(n33921) );
  NAND2_X1 U34974 ( .A1(n36628), .A2(n36627), .ZN(n33920) );
  NAND2_X1 U34975 ( .A1(n33921), .A2(n33920), .ZN(n36638) );
  OAI21_X1 U34976 ( .B1(n36639), .B2(n36637), .A(n36638), .ZN(n33923) );
  NAND2_X1 U34977 ( .A1(n33923), .A2(n33922), .ZN(n36648) );
  XNOR2_X1 U34978 ( .A(n36112), .B(\fmem_data[12][7] ), .ZN(n33925) );
  XNOR2_X1 U34979 ( .A(n34227), .B(n34228), .ZN(n33935) );
  FA_X1 U34980 ( .A(n33934), .B(n33933), .CI(n33932), .CO(n34224), .S(n34229)
         );
  XNOR2_X1 U34981 ( .A(n33935), .B(n34229), .ZN(n34254) );
  FA_X1 U34982 ( .A(n33938), .B(n33937), .CI(n33936), .CO(n34227), .S(n34123)
         );
  XNOR2_X1 U34983 ( .A(n33939), .B(\fmem_data[15][5] ), .ZN(n34057) );
  OAI22_X1 U34984 ( .A1(n33940), .A2(n34989), .B1(n34057), .B2(n34990), .ZN(
        n34118) );
  XNOR2_X1 U34985 ( .A(n33942), .B(n33941), .ZN(n33944) );
  XNOR2_X1 U34986 ( .A(n33944), .B(n33943), .ZN(n34117) );
  OAI22_X1 U34987 ( .A1(n33946), .A2(n36196), .B1(n33945), .B2(n3577), .ZN(
        n34116) );
  OAI21_X1 U34988 ( .B1(n34123), .B2(n34122), .A(n34121), .ZN(n33953) );
  NAND2_X1 U34989 ( .A1(n33953), .A2(n33952), .ZN(n34253) );
  OAI22_X1 U34990 ( .A1(n33957), .A2(n33956), .B1(n33955), .B2(n33954), .ZN(
        n34002) );
  INV_X1 U34991 ( .A(n35761), .ZN(n33958) );
  INV_X1 U34992 ( .A(n35705), .ZN(n33959) );
  INV_X1 U34993 ( .A(n35498), .ZN(n33960) );
  OAI22_X1 U34994 ( .A1(n33972), .A2(n34933), .B1(n33971), .B2(n34932), .ZN(
        n34008) );
  OAI21_X1 U34995 ( .B1(n34008), .B2(n34006), .A(n34007), .ZN(n33980) );
  NAND2_X1 U34996 ( .A1(n34008), .A2(n34006), .ZN(n33979) );
  NAND2_X1 U34997 ( .A1(n33980), .A2(n33979), .ZN(n34274) );
  OAI21_X1 U34998 ( .B1(n33983), .B2(n33982), .A(n33981), .ZN(n33985) );
  NAND2_X1 U34999 ( .A1(n3319), .A2(n33982), .ZN(n33984) );
  NAND2_X1 U35000 ( .A1(n33985), .A2(n33984), .ZN(n34088) );
  FA_X1 U35001 ( .A(n33988), .B(n33987), .CI(n33986), .CO(n34087), .S(n33671)
         );
  OAI22_X1 U35002 ( .A1(n33990), .A2(n3581), .B1(n33989), .B2(n36218), .ZN(
        n34086) );
  OAI22_X1 U35003 ( .A1(n33992), .A2(n34503), .B1(n33991), .B2(n34505), .ZN(
        n34064) );
  OAI22_X1 U35004 ( .A1(n33996), .A2(n34462), .B1(n33995), .B2(n34463), .ZN(
        n34062) );
  FA_X1 U35005 ( .A(n33999), .B(n33998), .CI(n33997), .CO(n34317), .S(n36061)
         );
  FA_X1 U35006 ( .A(n34002), .B(n34001), .CI(n34000), .CO(n34276), .S(n34132)
         );
  FA_X1 U35007 ( .A(n34005), .B(n34004), .CI(n34003), .CO(n34030), .S(n34131)
         );
  XNOR2_X1 U35008 ( .A(n34007), .B(n34006), .ZN(n34009) );
  XNOR2_X1 U35009 ( .A(n34009), .B(n34008), .ZN(n34130) );
  FA_X1 U35010 ( .A(n34012), .B(n34011), .CI(n34010), .CO(n34029), .S(n34146)
         );
  FA_X1 U35011 ( .A(n34015), .B(n34014), .CI(n34013), .CO(n34145), .S(n34330)
         );
  OAI22_X1 U35012 ( .A1(n34020), .A2(n34410), .B1(n34019), .B2(n34412), .ZN(
        n34315) );
  OAI22_X1 U35013 ( .A1(n34022), .A2(n34483), .B1(n3576), .B2(n34021), .ZN(
        n34406) );
  OAI22_X1 U35014 ( .A1(n34024), .A2(n34613), .B1(n3570), .B2(n34023), .ZN(
        n34405) );
  OAI22_X1 U35015 ( .A1(n34026), .A2(n3573), .B1(n34025), .B2(n36298), .ZN(
        n34404) );
  OAI21_X1 U35016 ( .B1(n34451), .B2(n34450), .A(n34452), .ZN(n34028) );
  NAND2_X1 U35017 ( .A1(n34451), .A2(n34450), .ZN(n34027) );
  NAND2_X1 U35018 ( .A1(n34028), .A2(n34027), .ZN(n34446) );
  OAI22_X1 U35019 ( .A1(n34038), .A2(n34499), .B1(n34501), .B2(n34037), .ZN(
        n34243) );
  XNOR2_X1 U35020 ( .A(n34264), .B(n34263), .ZN(n34058) );
  OR2_X1 U35021 ( .A1(n34047), .A2(n34986), .ZN(n34050) );
  OR2_X1 U35022 ( .A1(n34048), .A2(n34985), .ZN(n34049) );
  INV_X1 U35023 ( .A(n35745), .ZN(n34051) );
  INV_X1 U35024 ( .A(n35712), .ZN(n34052) );
  OR2_X1 U35025 ( .A1(n34210), .A2(n34211), .ZN(n34053) );
  NAND2_X1 U35026 ( .A1(n3323), .A2(n34053), .ZN(n34055) );
  NAND2_X1 U35027 ( .A1(n34211), .A2(n34210), .ZN(n34054) );
  NAND2_X1 U35028 ( .A1(n34055), .A2(n34054), .ZN(n34204) );
  OAI22_X1 U35029 ( .A1(n34057), .A2(n34989), .B1(n34990), .B2(n34056), .ZN(
        n34203) );
  XNOR2_X1 U35030 ( .A(n34058), .B(n34261), .ZN(n34187) );
  FA_X1 U35031 ( .A(n34061), .B(n34060), .CI(n34059), .CO(n34275), .S(n34127)
         );
  FA_X1 U35032 ( .A(n34064), .B(n34063), .CI(n34062), .CO(n34126), .S(n34318)
         );
  FA_X1 U35033 ( .A(n34067), .B(n34066), .CI(n34065), .CO(n34313), .S(n34368)
         );
  FA_X1 U35034 ( .A(n34070), .B(n34069), .CI(n34068), .CO(n34001), .S(n34312)
         );
  OAI22_X1 U35035 ( .A1(n34072), .A2(n34836), .B1(n34071), .B2(n34835), .ZN(
        n34311) );
  OAI21_X1 U35036 ( .B1(n34447), .B2(n34446), .A(n34448), .ZN(n34074) );
  NAND2_X1 U35037 ( .A1(n34447), .A2(n34446), .ZN(n34073) );
  NAND2_X1 U35038 ( .A1(n34074), .A2(n34073), .ZN(n34381) );
  INV_X1 U35039 ( .A(n34381), .ZN(n34162) );
  FA_X1 U35040 ( .A(n34077), .B(n34076), .CI(n34075), .CO(n34255), .S(n34248)
         );
  FA_X1 U35041 ( .A(n34082), .B(n34081), .CI(n34080), .CO(n34246), .S(n34121)
         );
  FA_X1 U35042 ( .A(n34085), .B(n34084), .CI(n34083), .CO(n34305), .S(n34325)
         );
  FA_X1 U35043 ( .A(n34088), .B(n34087), .CI(n34086), .CO(n34304), .S(n34319)
         );
  FA_X1 U35044 ( .A(n34091), .B(n34090), .CI(n34089), .CO(n34306), .S(n34326)
         );
  OAI21_X1 U35045 ( .B1(n34305), .B2(n34304), .A(n34306), .ZN(n34093) );
  NAND2_X1 U35046 ( .A1(n34305), .A2(n34304), .ZN(n34092) );
  NAND2_X1 U35047 ( .A1(n34093), .A2(n34092), .ZN(n34184) );
  FA_X1 U35048 ( .A(n34096), .B(n34095), .CI(n34094), .CO(n33345), .S(n34251)
         );
  XNOR2_X1 U35049 ( .A(n36244), .B(\fmem_data[14][7] ), .ZN(n34098) );
  OAI22_X1 U35050 ( .A1(n34098), .A2(n35576), .B1(n34097), .B2(n35577), .ZN(
        n34135) );
  XNOR2_X1 U35051 ( .A(n36243), .B(\fmem_data[22][7] ), .ZN(n34101) );
  OAI22_X1 U35052 ( .A1(n34102), .A2(n35585), .B1(n35584), .B2(n34101), .ZN(
        n34133) );
  FA_X1 U35053 ( .A(n34104), .B(n33272), .CI(n34103), .CO(n33344), .S(n34249)
         );
  FA_X1 U35054 ( .A(n34107), .B(n34106), .CI(n34105), .CO(n34138), .S(n34114)
         );
  FA_X1 U35055 ( .A(n34110), .B(n34109), .CI(n34108), .CO(n26379), .S(n34137)
         );
  OAI22_X1 U35056 ( .A1(n34112), .A2(n36216), .B1(n34111), .B2(n3931), .ZN(
        n34136) );
  FA_X1 U35057 ( .A(n34115), .B(n34114), .CI(n34113), .CO(n34322), .S(n34639)
         );
  FA_X1 U35058 ( .A(n34118), .B(n34117), .CI(n34116), .CO(n34122), .S(n34320)
         );
  OAI21_X1 U35059 ( .B1(n34321), .B2(n34322), .A(n34320), .ZN(n34120) );
  NAND2_X1 U35060 ( .A1(n34321), .A2(n34322), .ZN(n34119) );
  NAND2_X1 U35061 ( .A1(n34120), .A2(n34119), .ZN(n34455) );
  XNOR2_X1 U35062 ( .A(n34122), .B(n34121), .ZN(n34124) );
  XNOR2_X1 U35063 ( .A(n34124), .B(n34123), .ZN(n34454) );
  FA_X1 U35064 ( .A(n34127), .B(n34126), .CI(n34125), .CO(n34186), .S(n34456)
         );
  OAI21_X1 U35065 ( .B1(n34455), .B2(n34454), .A(n34456), .ZN(n34129) );
  NAND2_X1 U35066 ( .A1(n34455), .A2(n34454), .ZN(n34128) );
  NAND2_X1 U35067 ( .A1(n34129), .A2(n34128), .ZN(n34377) );
  FA_X1 U35068 ( .A(n34132), .B(n34131), .CI(n34130), .CO(n34280), .S(n34450)
         );
  FA_X1 U35069 ( .A(n34134), .B(n34135), .CI(n34133), .CO(n34250), .S(n34300)
         );
  FA_X1 U35070 ( .A(n34138), .B(n34137), .CI(n34136), .CO(n34301), .S(n34321)
         );
  FA_X1 U35071 ( .A(n34141), .B(n34140), .CI(n34139), .CO(n34302), .S(n34332)
         );
  OAI21_X1 U35072 ( .B1(n34300), .B2(n34301), .A(n34302), .ZN(n34143) );
  NAND2_X1 U35073 ( .A1(n34143), .A2(n34142), .ZN(n34279) );
  FA_X1 U35074 ( .A(n34146), .B(n34145), .CI(n34144), .CO(n34278), .S(n34452)
         );
  INV_X1 U35075 ( .A(n34382), .ZN(n34161) );
  NOR2_X1 U35076 ( .A1(n34382), .A2(n34381), .ZN(n34160) );
  XNOR2_X1 U35077 ( .A(n34148), .B(n34147), .ZN(n34150) );
  XNOR2_X1 U35078 ( .A(n34150), .B(n34149), .ZN(n34291) );
  FA_X1 U35079 ( .A(n34153), .B(n34152), .CI(n34151), .CO(n34181), .S(n34290)
         );
  OAI21_X1 U35080 ( .B1(n34155), .B2(n34156), .A(n34154), .ZN(n34158) );
  NAND2_X1 U35081 ( .A1(n34156), .A2(n34155), .ZN(n34157) );
  NAND2_X1 U35082 ( .A1(n34158), .A2(n34157), .ZN(n34289) );
  INV_X1 U35083 ( .A(n34383), .ZN(n34159) );
  OAI22_X1 U35084 ( .A1(n34162), .A2(n34161), .B1(n34160), .B2(n34159), .ZN(
        n35449) );
  FA_X1 U35085 ( .A(n34165), .B(n34164), .CI(n34163), .CO(n27314), .S(n34285)
         );
  FA_X1 U35086 ( .A(n34168), .B(n34167), .CI(n34166), .CO(n34180), .S(n34374)
         );
  FA_X1 U35087 ( .A(n34171), .B(n34170), .CI(n34169), .CO(n34163), .S(n34373)
         );
  OAI21_X1 U35088 ( .B1(n34174), .B2(n34173), .A(n34172), .ZN(n34175) );
  NAND2_X1 U35089 ( .A1(n34176), .A2(n34175), .ZN(n34372) );
  OAI21_X1 U35090 ( .B1(n34374), .B2(n34373), .A(n34372), .ZN(n34178) );
  NAND2_X1 U35091 ( .A1(n34178), .A2(n34177), .ZN(n34284) );
  XNOR2_X1 U35092 ( .A(n34180), .B(n34179), .ZN(n34182) );
  XNOR2_X1 U35093 ( .A(n34182), .B(n34181), .ZN(n34283) );
  FA_X1 U35094 ( .A(n34185), .B(n34183), .CI(n34184), .CO(n34700), .S(n34378)
         );
  FA_X1 U35095 ( .A(n34188), .B(n34187), .CI(n34186), .CO(n34699), .S(n34448)
         );
  OAI22_X1 U35096 ( .A1(n34192), .A2(n34474), .B1(n34191), .B2(n34472), .ZN(
        n34309) );
  XNOR2_X1 U35097 ( .A(n34615), .B(\fmem_data[21][5] ), .ZN(n34193) );
  OAI22_X1 U35098 ( .A1(n34196), .A2(n34195), .B1(n34194), .B2(n34193), .ZN(
        n34409) );
  OAI22_X1 U35099 ( .A1(n34198), .A2(n3579), .B1(n34197), .B2(n34476), .ZN(
        n34408) );
  OAI22_X1 U35100 ( .A1(n34202), .A2(n34201), .B1(n34200), .B2(n34199), .ZN(
        n34407) );
  FA_X1 U35101 ( .A(n34205), .B(n34204), .CI(n34203), .CO(n34261), .S(n34393)
         );
  FA_X1 U35102 ( .A(n34215), .B(n34214), .CI(n34213), .CO(n34399), .S(n33881)
         );
  FA_X1 U35103 ( .A(n34218), .B(n34217), .CI(n34216), .CO(n33286), .S(n34386)
         );
  FA_X1 U35104 ( .A(n34221), .B(n34220), .CI(n34219), .CO(n34677), .S(n34385)
         );
  OAI21_X1 U35105 ( .B1(n34387), .B2(n34386), .A(n34385), .ZN(n34223) );
  NAND2_X1 U35106 ( .A1(n34387), .A2(n34386), .ZN(n34222) );
  NAND2_X1 U35107 ( .A1(n34223), .A2(n34222), .ZN(n34698) );
  FA_X1 U35108 ( .A(n34226), .B(n34225), .CI(n34224), .CO(n12717), .S(n34658)
         );
  OAI21_X1 U35109 ( .B1(n34229), .B2(n34228), .A(n34227), .ZN(n34231) );
  NAND2_X1 U35110 ( .A1(n34229), .A2(n34228), .ZN(n34230) );
  NAND2_X1 U35111 ( .A1(n34231), .A2(n34230), .ZN(n34657) );
  FA_X1 U35112 ( .A(n34238), .B(n34237), .CI(n34236), .CO(n34662), .S(n34031)
         );
  FA_X1 U35113 ( .A(n34245), .B(n34244), .CI(n34243), .CO(n34665), .S(n34264)
         );
  FA_X1 U35114 ( .A(n34246), .B(n34247), .CI(n34248), .CO(n34660), .S(n34185)
         );
  FA_X1 U35115 ( .A(n34251), .B(n34250), .CI(n34249), .CO(n34659), .S(n34183)
         );
  FA_X1 U35116 ( .A(n34254), .B(n34253), .CI(n34252), .CO(n34653), .S(n34447)
         );
  FA_X1 U35117 ( .A(n34257), .B(n34256), .CI(n34255), .CO(n18727), .S(n34683)
         );
  FA_X1 U35118 ( .A(n34260), .B(n34259), .CI(n34258), .CO(n12727), .S(n34682)
         );
  XNOR2_X1 U35119 ( .A(n34683), .B(n34682), .ZN(n34267) );
  OR2_X1 U35120 ( .A1(n34264), .A2(n34263), .ZN(n34262) );
  NAND2_X1 U35121 ( .A1(n34262), .A2(n34261), .ZN(n34266) );
  NAND2_X1 U35122 ( .A1(n34266), .A2(n34265), .ZN(n34681) );
  XNOR2_X1 U35123 ( .A(n34267), .B(n34681), .ZN(n34697) );
  FA_X1 U35124 ( .A(n34270), .B(n34269), .CI(n34268), .CO(n12725), .S(n34688)
         );
  FA_X1 U35125 ( .A(n34273), .B(n34272), .CI(n34271), .CO(n12724), .S(n34687)
         );
  XNOR2_X1 U35126 ( .A(n34688), .B(n34687), .ZN(n34277) );
  FA_X1 U35127 ( .A(n34276), .B(n34275), .CI(n34274), .CO(n34686), .S(n34252)
         );
  XNOR2_X1 U35128 ( .A(n34277), .B(n34686), .ZN(n34696) );
  FA_X1 U35129 ( .A(n34280), .B(n34279), .CI(n34278), .CO(n34695), .S(n34376)
         );
  OAI21_X1 U35130 ( .B1(n34715), .B2(n34714), .A(n34713), .ZN(n34282) );
  NAND2_X1 U35131 ( .A1(n34282), .A2(n34281), .ZN(n35447) );
  FA_X1 U35132 ( .A(n34285), .B(n34284), .CI(n34283), .CO(n35448), .S(n34550)
         );
  FA_X1 U35133 ( .A(n34288), .B(n34287), .CI(n34286), .CO(n31423), .S(n34549)
         );
  FA_X1 U35134 ( .A(n34290), .B(n34291), .CI(n34289), .CO(n34383), .S(n34553)
         );
  OAI21_X1 U35135 ( .B1(n34294), .B2(n34293), .A(n34292), .ZN(n34296) );
  NAND2_X1 U35136 ( .A1(n34294), .A2(n34293), .ZN(n34295) );
  NAND2_X1 U35137 ( .A1(n34296), .A2(n34295), .ZN(n34552) );
  FA_X1 U35138 ( .A(n34298), .B(n34299), .CI(n34297), .CO(n34551), .S(n36423)
         );
  XNOR2_X1 U35139 ( .A(n34301), .B(n34300), .ZN(n34303) );
  XNOR2_X1 U35140 ( .A(n34303), .B(n34302), .ZN(n34391) );
  XNOR2_X1 U35141 ( .A(n34305), .B(n34304), .ZN(n34307) );
  XNOR2_X1 U35142 ( .A(n34307), .B(n34306), .ZN(n34390) );
  FA_X1 U35143 ( .A(n34309), .B(n34310), .CI(n34308), .CO(n34394), .S(n34329)
         );
  FA_X1 U35144 ( .A(n34313), .B(n34312), .CI(n34311), .CO(n34125), .S(n34328)
         );
  FA_X1 U35145 ( .A(n34316), .B(n34315), .CI(n34314), .CO(n34144), .S(n34327)
         );
  FA_X1 U35146 ( .A(n34319), .B(n34318), .CI(n34317), .CO(n34451), .S(n36069)
         );
  XNOR2_X1 U35147 ( .A(n34321), .B(n34320), .ZN(n34323) );
  XNOR2_X1 U35148 ( .A(n34323), .B(n34322), .ZN(n36068) );
  FA_X1 U35149 ( .A(n34326), .B(n34325), .CI(n34324), .CO(n34154), .S(n36067)
         );
  FA_X1 U35150 ( .A(n34329), .B(n34328), .CI(n34327), .CO(n34389), .S(n34567)
         );
  XNOR2_X1 U35151 ( .A(n34331), .B(n34330), .ZN(n34333) );
  XNOR2_X1 U35152 ( .A(n34333), .B(n34332), .ZN(n34566) );
  XNOR2_X1 U35153 ( .A(n36316), .B(\fmem_data[27][3] ), .ZN(n34335) );
  XNOR2_X1 U35154 ( .A(n34334), .B(\fmem_data[27][3] ), .ZN(n34427) );
  OAI22_X1 U35155 ( .A1(n34335), .A2(n34462), .B1(n34427), .B2(n34463), .ZN(
        n34633) );
  OR2_X1 U35156 ( .A1(n3116), .A2(n3674), .ZN(n34336) );
  INV_X1 U35157 ( .A(n34501), .ZN(n34339) );
  INV_X1 U35158 ( .A(n34340), .ZN(n34341) );
  OAI22_X1 U35159 ( .A1(n34344), .A2(n34343), .B1(n34342), .B2(n3578), .ZN(
        n34619) );
  FA_X1 U35160 ( .A(n34349), .B(n34348), .CI(n34347), .CO(n34601), .S(n36600)
         );
  INV_X1 U35161 ( .A(n36058), .ZN(n34371) );
  FA_X1 U35162 ( .A(n34352), .B(n34351), .CI(n34350), .CO(n34367), .S(n34577)
         );
  NOR2_X1 U35163 ( .A1(n34355), .A2(n34354), .ZN(n34358) );
  INV_X1 U35164 ( .A(n34353), .ZN(n34357) );
  OAI21_X1 U35165 ( .B1(n34358), .B2(n34357), .A(n34356), .ZN(n34576) );
  OAI22_X1 U35166 ( .A1(n34360), .A2(n3662), .B1(n34359), .B2(n36241), .ZN(
        n36093) );
  XNOR2_X1 U35167 ( .A(n3116), .B(\fmem_data[23][3] ), .ZN(n34362) );
  OAI22_X1 U35168 ( .A1(n34411), .A2(n34412), .B1(n34410), .B2(n34362), .ZN(
        n36092) );
  FA_X1 U35169 ( .A(n34368), .B(n34367), .CI(n34366), .CO(n33664), .S(n36056)
         );
  NOR2_X1 U35170 ( .A1(n36057), .A2(n36056), .ZN(n34370) );
  OAI21_X1 U35171 ( .B1(n34371), .B2(n34370), .A(n34369), .ZN(n34565) );
  XNOR2_X1 U35172 ( .A(n34373), .B(n34372), .ZN(n34375) );
  FA_X1 U35173 ( .A(n34378), .B(n34377), .CI(n34376), .CO(n34382), .S(n34555)
         );
  OAI21_X1 U35174 ( .B1(n34556), .B2(n34554), .A(n34555), .ZN(n34380) );
  NAND2_X1 U35175 ( .A1(n34556), .A2(n34554), .ZN(n34379) );
  NAND2_X1 U35176 ( .A1(n34380), .A2(n34379), .ZN(n34650) );
  XNOR2_X1 U35177 ( .A(n34382), .B(n34381), .ZN(n34384) );
  XNOR2_X1 U35178 ( .A(n34384), .B(n34383), .ZN(n34649) );
  XNOR2_X1 U35179 ( .A(n34386), .B(n34385), .ZN(n34388) );
  XNOR2_X1 U35180 ( .A(n34388), .B(n34387), .ZN(n34709) );
  FA_X1 U35181 ( .A(n34390), .B(n34391), .CI(n34389), .CO(n34708), .S(n34560)
         );
  FA_X1 U35182 ( .A(n34393), .B(n34394), .CI(n34392), .CO(n34387), .S(n34800)
         );
  XNOR2_X1 U35183 ( .A(n34396), .B(n34395), .ZN(n34398) );
  FA_X1 U35184 ( .A(n34401), .B(n34400), .CI(n34399), .CO(n34392), .S(n34458)
         );
  FA_X1 U35185 ( .A(n34406), .B(n34405), .CI(n34404), .CO(n34314), .S(n34493)
         );
  FA_X1 U35186 ( .A(n34407), .B(n34408), .CI(n34409), .CO(n34308), .S(n34492)
         );
  OAI22_X1 U35187 ( .A1(n34421), .A2(n34420), .B1(n34419), .B2(n34418), .ZN(
        n34489) );
  OAI22_X1 U35188 ( .A1(n34427), .A2(n34462), .B1(n34463), .B2(n34426), .ZN(
        n34511) );
  OAI22_X1 U35189 ( .A1(n34430), .A2(n34429), .B1(n34428), .B2(n34533), .ZN(
        n34510) );
  OAI21_X1 U35190 ( .B1(n34519), .B2(n34520), .A(n34518), .ZN(n34443) );
  NAND2_X1 U35191 ( .A1(n34443), .A2(n34442), .ZN(n34460) );
  OAI21_X1 U35192 ( .B1(n34458), .B2(n34459), .A(n34460), .ZN(n34445) );
  NAND2_X1 U35193 ( .A1(n34445), .A2(n34444), .ZN(n34798) );
  XNOR2_X1 U35194 ( .A(n34446), .B(n34447), .ZN(n34449) );
  XNOR2_X1 U35195 ( .A(n34451), .B(n34450), .ZN(n34453) );
  XNOR2_X1 U35196 ( .A(n34453), .B(n34452), .ZN(n34562) );
  XNOR2_X1 U35197 ( .A(n34454), .B(n34455), .ZN(n34457) );
  XNOR2_X1 U35198 ( .A(n34457), .B(n34456), .ZN(n34561) );
  XNOR2_X1 U35199 ( .A(n34459), .B(n34458), .ZN(n34461) );
  XNOR2_X1 U35200 ( .A(n34461), .B(n34460), .ZN(n36070) );
  OR2_X1 U35201 ( .A1(n36316), .A2(n3643), .ZN(n34464) );
  XNOR2_X1 U35202 ( .A(n36337), .B(\fmem_data[19][3] ), .ZN(n34475) );
  OAI22_X1 U35203 ( .A1(n34475), .A2(n34474), .B1(n34473), .B2(n34472), .ZN(
        n34579) );
  INV_X1 U35204 ( .A(n34479), .ZN(n34481) );
  XNOR2_X1 U35205 ( .A(n34481), .B(n34480), .ZN(n34587) );
  OAI22_X1 U35206 ( .A1(n34484), .A2(n34483), .B1(n34482), .B2(n3576), .ZN(
        n34586) );
  OAI21_X1 U35207 ( .B1(n34579), .B2(n34578), .A(n34580), .ZN(n34488) );
  NAND2_X1 U35208 ( .A1(n34579), .A2(n34578), .ZN(n34487) );
  NAND2_X1 U35209 ( .A1(n34488), .A2(n34487), .ZN(n34635) );
  FA_X1 U35210 ( .A(n34491), .B(n34490), .CI(n34489), .CO(n34519), .S(n34634)
         );
  FA_X1 U35211 ( .A(n34494), .B(n34493), .CI(n34492), .CO(n34459), .S(n36063)
         );
  OAI22_X1 U35212 ( .A1(n34498), .A2(n34497), .B1(n34496), .B2(n34495), .ZN(
        n34584) );
  FA_X1 U35213 ( .A(n34509), .B(n34508), .CI(n34507), .CO(n34113), .S(n36083)
         );
  FA_X1 U35214 ( .A(n34512), .B(n34511), .CI(n34510), .CO(n34520), .S(n36082)
         );
  OAI21_X1 U35215 ( .B1(n36065), .B2(n36063), .A(n36064), .ZN(n34514) );
  NAND2_X1 U35216 ( .A1(n36065), .A2(n36063), .ZN(n34513) );
  NAND2_X1 U35217 ( .A1(n34514), .A2(n34513), .ZN(n36071) );
  FA_X1 U35218 ( .A(n34517), .B(n34516), .CI(n34515), .CO(n34722), .S(n36126)
         );
  XNOR2_X1 U35219 ( .A(n34519), .B(n34518), .ZN(n34521) );
  XNOR2_X1 U35220 ( .A(n34521), .B(n34520), .ZN(n36125) );
  FA_X1 U35221 ( .A(n34524), .B(n34523), .CI(n34522), .CO(n34518), .S(n36129)
         );
  FA_X1 U35222 ( .A(n34527), .B(n34526), .CI(n34525), .CO(n32837), .S(n36128)
         );
  XNOR2_X1 U35223 ( .A(n34531), .B(\fmem_data[10][1] ), .ZN(n36103) );
  OAI22_X1 U35224 ( .A1(n36103), .A2(n36114), .B1(n34532), .B2(n3561), .ZN(
        n36117) );
  INV_X1 U35225 ( .A(n34533), .ZN(n34534) );
  AND2_X1 U35226 ( .A1(n36313), .A2(n34534), .ZN(n36116) );
  XNOR2_X1 U35227 ( .A(n36296), .B(\fmem_data[0][3] ), .ZN(n34536) );
  FA_X1 U35228 ( .A(n34541), .B(n34540), .CI(n34539), .CO(n32870), .S(n36107)
         );
  OAI21_X1 U35229 ( .B1(n36070), .B2(n36071), .A(n36072), .ZN(n34543) );
  NAND2_X1 U35230 ( .A1(n34543), .A2(n34542), .ZN(n34563) );
  OAI21_X1 U35231 ( .B1(n3391), .B2(n34561), .A(n34563), .ZN(n34545) );
  NAND2_X1 U35232 ( .A1(n3391), .A2(n34561), .ZN(n34544) );
  NAND2_X1 U35233 ( .A1(n34545), .A2(n34544), .ZN(n36048) );
  OAI21_X1 U35234 ( .B1(n36050), .B2(n36049), .A(n36048), .ZN(n34547) );
  NAND2_X1 U35235 ( .A1(n34547), .A2(n34546), .ZN(n34648) );
  FA_X1 U35236 ( .A(n34550), .B(n34549), .CI(n34548), .CO(n35467), .S(n36631)
         );
  FA_X1 U35237 ( .A(n34553), .B(n34552), .CI(n34551), .CO(n34548), .S(n36620)
         );
  XNOR2_X1 U35238 ( .A(n34555), .B(n34554), .ZN(n34557) );
  XNOR2_X1 U35239 ( .A(n34557), .B(n3463), .ZN(n36622) );
  FA_X1 U35240 ( .A(n34559), .B(n34560), .CI(n34558), .CO(n34556), .S(n36453)
         );
  XNOR2_X1 U35241 ( .A(n34562), .B(n34561), .ZN(n34564) );
  XNOR2_X1 U35242 ( .A(n34564), .B(n34563), .ZN(n36452) );
  FA_X1 U35243 ( .A(n34567), .B(n34566), .CI(n34565), .CO(n34558), .S(n36460)
         );
  XNOR2_X1 U35244 ( .A(n34569), .B(n34568), .ZN(n34571) );
  XNOR2_X1 U35245 ( .A(n34571), .B(n34570), .ZN(n36459) );
  FA_X1 U35246 ( .A(n34574), .B(n34573), .CI(n34572), .CO(n36060), .S(n36596)
         );
  FA_X1 U35247 ( .A(n34577), .B(n34576), .CI(n34575), .CO(n36057), .S(n36595)
         );
  FA_X1 U35248 ( .A(n34584), .B(n34583), .CI(n34582), .CO(n36084), .S(n36604)
         );
  FA_X1 U35249 ( .A(n34587), .B(n34586), .CI(n34585), .CO(n34580), .S(n36553)
         );
  NOR2_X1 U35250 ( .A1(n34588), .A2(n3693), .ZN(n34591) );
  NOR2_X1 U35251 ( .A1(n34589), .A2(n3693), .ZN(n34590) );
  NOR2_X1 U35252 ( .A1(n34591), .A2(n34590), .ZN(n34592) );
  NAND2_X1 U35253 ( .A1(n34593), .A2(n34592), .ZN(n34778) );
  NAND2_X1 U35254 ( .A1(n34739), .A2(n34594), .ZN(n36567) );
  NAND2_X1 U35255 ( .A1(n36120), .A2(n34595), .ZN(n36566) );
  NAND2_X1 U35256 ( .A1(n34777), .A2(n34597), .ZN(n36570) );
  INV_X1 U35257 ( .A(n36498), .ZN(n34645) );
  FA_X1 U35258 ( .A(n34603), .B(n34602), .CI(n34601), .CO(n36058), .S(n36606)
         );
  FA_X1 U35259 ( .A(n34606), .B(n34605), .CI(n34604), .CO(n34353), .S(n36542)
         );
  FA_X1 U35260 ( .A(n34609), .B(n34608), .CI(n34607), .CO(n34349), .S(n36541)
         );
  OAI22_X1 U35261 ( .A1(n36112), .A2(n34734), .B1(n34735), .B2(n3572), .ZN(
        n36539) );
  AND2_X1 U35262 ( .A1(n3353), .A2(\fmem_data[2][0] ), .ZN(n36559) );
  INV_X1 U35263 ( .A(n34613), .ZN(n34614) );
  XNOR2_X1 U35264 ( .A(n34618), .B(n34617), .ZN(n36537) );
  FA_X1 U35265 ( .A(n34621), .B(n34620), .CI(n34619), .CO(n36089), .S(n36556)
         );
  NAND2_X1 U35266 ( .A1(n36298), .A2(n34622), .ZN(n36519) );
  NAND2_X1 U35267 ( .A1(n34788), .A2(n34628), .ZN(n36529) );
  NAND2_X1 U35268 ( .A1(n34734), .A2(n34629), .ZN(n36528) );
  XNOR2_X1 U35269 ( .A(n34630), .B(\fmem_data[14][1] ), .ZN(n34740) );
  FA_X1 U35270 ( .A(n34633), .B(n34632), .CI(n34631), .CO(n34603), .S(n36511)
         );
  FA_X1 U35271 ( .A(n34636), .B(n34635), .CI(n34634), .CO(n36065), .S(n36608)
         );
  OAI21_X1 U35272 ( .B1(n36606), .B2(n36607), .A(n36608), .ZN(n34638) );
  NAND2_X1 U35273 ( .A1(n36607), .A2(n36606), .ZN(n34637) );
  NAND2_X1 U35274 ( .A1(n34638), .A2(n34637), .ZN(n36497) );
  XNOR2_X1 U35275 ( .A(n34640), .B(n34639), .ZN(n34642) );
  XNOR2_X1 U35276 ( .A(n34642), .B(n34641), .ZN(n36496) );
  NOR2_X1 U35277 ( .A1(n36497), .A2(n36496), .ZN(n34644) );
  NAND2_X1 U35278 ( .A1(n36497), .A2(n36496), .ZN(n34643) );
  OAI21_X1 U35279 ( .B1(n34645), .B2(n34644), .A(n34643), .ZN(n36458) );
  OAI21_X1 U35280 ( .B1(n36620), .B2(n36622), .A(n36621), .ZN(n34647) );
  NAND2_X1 U35281 ( .A1(n36620), .A2(n36622), .ZN(n34646) );
  NAND2_X1 U35282 ( .A1(n34647), .A2(n34646), .ZN(n36632) );
  NAND2_X1 U35283 ( .A1(n36631), .A2(n36632), .ZN(n34652) );
  FA_X1 U35284 ( .A(n34650), .B(n34649), .CI(n34648), .CO(n35466), .S(n36633)
         );
  OAI21_X1 U35285 ( .B1(n36631), .B2(n36632), .A(n36633), .ZN(n34651) );
  NAND2_X1 U35286 ( .A1(n34651), .A2(n34652), .ZN(n36642) );
  FA_X1 U35287 ( .A(n34655), .B(n34654), .CI(n34653), .CO(n35219), .S(n34714)
         );
  FA_X1 U35288 ( .A(n34658), .B(n34657), .CI(n34656), .CO(n34855), .S(n34655)
         );
  FA_X1 U35289 ( .A(n34661), .B(n34660), .CI(n34659), .CO(n34856), .S(n34654)
         );
  XNOR2_X1 U35290 ( .A(n34855), .B(n34856), .ZN(n34670) );
  FA_X1 U35291 ( .A(n34664), .B(n34663), .CI(n34662), .CO(n34886), .S(n34656)
         );
  FA_X1 U35292 ( .A(n34667), .B(n34666), .CI(n34665), .CO(n34885), .S(n34661)
         );
  FA_X1 U35293 ( .A(n3704), .B(n34669), .CI(n34668), .CO(n35082), .S(n34884)
         );
  XNOR2_X1 U35294 ( .A(n34670), .B(n34854), .ZN(n35220) );
  XNOR2_X1 U35295 ( .A(n35219), .B(n35220), .ZN(n34680) );
  FA_X1 U35296 ( .A(n34673), .B(n34672), .CI(n34671), .CO(n33392), .S(n34706)
         );
  FA_X1 U35297 ( .A(n34676), .B(n34675), .CI(n34674), .CO(n34705), .S(n34719)
         );
  FA_X1 U35298 ( .A(n34677), .B(n34678), .CI(n34679), .CO(n33358), .S(n34704)
         );
  XNOR2_X1 U35299 ( .A(n34680), .B(n35218), .ZN(n35452) );
  XNOR2_X1 U35300 ( .A(n34692), .B(n34691), .ZN(n34694) );
  XNOR2_X1 U35301 ( .A(n34694), .B(n34693), .ZN(n34888) );
  FA_X1 U35302 ( .A(n34697), .B(n34696), .CI(n34695), .CO(n35227), .S(n34713)
         );
  FA_X1 U35303 ( .A(n34700), .B(n34699), .CI(n34698), .CO(n35226), .S(n34715)
         );
  FA_X1 U35304 ( .A(n34703), .B(n34702), .CI(n34701), .CO(n33359), .S(n34712)
         );
  FA_X1 U35305 ( .A(n34704), .B(n34705), .CI(n34706), .CO(n35218), .S(n34711)
         );
  FA_X1 U35306 ( .A(n34708), .B(n34709), .CI(n34707), .CO(n34710), .S(n36050)
         );
  FA_X1 U35307 ( .A(n34712), .B(n34711), .CI(n34710), .CO(n35450), .S(n36041)
         );
  XNOR2_X1 U35308 ( .A(n34714), .B(n34713), .ZN(n34716) );
  XNOR2_X1 U35309 ( .A(n34716), .B(n34715), .ZN(n36040) );
  FA_X1 U35310 ( .A(n34719), .B(n34718), .CI(n34717), .CO(n33295), .S(n36044)
         );
  XNOR2_X1 U35311 ( .A(n34721), .B(n34720), .ZN(n34723) );
  XNOR2_X1 U35312 ( .A(n34723), .B(n34722), .ZN(n36075) );
  FA_X1 U35313 ( .A(n34726), .B(n34725), .CI(n34724), .CO(n32827), .S(n36165)
         );
  FA_X1 U35314 ( .A(n34729), .B(n34728), .CI(n34727), .CO(n34752), .S(n36132)
         );
  FA_X1 U35315 ( .A(n34732), .B(n34730), .CI(n34731), .CO(n32838), .S(n36131)
         );
  OAI22_X1 U35316 ( .A1(n34735), .A2(n34734), .B1(n3572), .B2(n34733), .ZN(
        n36096) );
  INV_X1 U35317 ( .A(n34736), .ZN(n34737) );
  OAI22_X1 U35318 ( .A1(n34740), .A2(n34739), .B1(n34738), .B2(n3563), .ZN(
        n36094) );
  OAI22_X1 U35319 ( .A1(n34746), .A2(n34745), .B1(n34744), .B2(n3562), .ZN(
        n36098) );
  FA_X1 U35321 ( .A(n34749), .B(n34748), .CI(n34747), .CO(n32840), .S(n36136)
         );
  OAI21_X1 U35322 ( .B1(n36139), .B2(n36137), .A(n36136), .ZN(n34751) );
  NAND2_X1 U35323 ( .A1(n34751), .A2(n34750), .ZN(n36130) );
  XNOR2_X1 U35324 ( .A(n34753), .B(n34752), .ZN(n34755) );
  XNOR2_X1 U35325 ( .A(n34755), .B(n34754), .ZN(n36163) );
  OAI21_X1 U35326 ( .B1(n36165), .B2(n36164), .A(n36163), .ZN(n34757) );
  NAND2_X1 U35327 ( .A1(n36164), .A2(n36165), .ZN(n34756) );
  NAND2_X1 U35328 ( .A1(n34757), .A2(n34756), .ZN(n36074) );
  FA_X1 U35329 ( .A(n34760), .B(n34759), .CI(n34758), .CO(n32830), .S(n36186)
         );
  XNOR2_X1 U35330 ( .A(n34762), .B(n34761), .ZN(n34764) );
  XNOR2_X1 U35331 ( .A(n34764), .B(n34763), .ZN(n36187) );
  FA_X1 U35332 ( .A(n34767), .B(n34766), .CI(n34765), .CO(n32847), .S(n36142)
         );
  FA_X1 U35333 ( .A(n34770), .B(n34769), .CI(n34768), .CO(n32845), .S(n36141)
         );
  FA_X1 U35334 ( .A(n34775), .B(n34774), .CI(n34773), .CO(n34760), .S(n36191)
         );
  OAI22_X1 U35335 ( .A1(n34778), .A2(n34777), .B1(n34776), .B2(n3567), .ZN(
        n36246) );
  INV_X1 U35336 ( .A(n36246), .ZN(n34782) );
  INV_X1 U35337 ( .A(n34779), .ZN(n34780) );
  INV_X1 U35338 ( .A(n36247), .ZN(n34781) );
  NAND2_X1 U35339 ( .A1(n34782), .A2(n34781), .ZN(n34785) );
  XNOR2_X1 U35340 ( .A(n34783), .B(\fmem_data[3][1] ), .ZN(n36119) );
  OAI22_X1 U35341 ( .A1(n34784), .A2(n3582), .B1(n36119), .B2(n36199), .ZN(
        n36248) );
  NAND2_X1 U35342 ( .A1(n34785), .A2(n36248), .ZN(n34787) );
  NAND2_X1 U35343 ( .A1(n36247), .A2(n36246), .ZN(n34786) );
  NAND2_X1 U35344 ( .A1(n34787), .A2(n34786), .ZN(n36235) );
  FA_X1 U35345 ( .A(n34793), .B(n34792), .CI(n34791), .CO(n32869), .S(n36233)
         );
  OAI21_X1 U35346 ( .B1(n36186), .B2(n36187), .A(n36188), .ZN(n34795) );
  NAND2_X1 U35347 ( .A1(n34795), .A2(n34794), .ZN(n36076) );
  OAI21_X1 U35348 ( .B1(n36074), .B2(n36075), .A(n36076), .ZN(n34797) );
  NAND2_X1 U35349 ( .A1(n36075), .A2(n36074), .ZN(n34796) );
  NAND2_X1 U35350 ( .A1(n34797), .A2(n34796), .ZN(n36055) );
  FA_X1 U35351 ( .A(n34799), .B(n34800), .CI(n34798), .CO(n34707), .S(n36052)
         );
  FA_X1 U35352 ( .A(n34803), .B(n34802), .CI(n34801), .CO(n34808), .S(n36053)
         );
  OAI21_X1 U35353 ( .B1(n36055), .B2(n36052), .A(n36053), .ZN(n34805) );
  NAND2_X1 U35354 ( .A1(n36055), .A2(n36052), .ZN(n34804) );
  NAND2_X1 U35355 ( .A1(n34805), .A2(n34804), .ZN(n36045) );
  XNOR2_X1 U35356 ( .A(n34807), .B(n34806), .ZN(n34809) );
  XNOR2_X1 U35357 ( .A(n34809), .B(n34808), .ZN(n36047) );
  OAI21_X1 U35358 ( .B1(n36044), .B2(n36045), .A(n36047), .ZN(n34811) );
  NAND2_X1 U35359 ( .A1(n36044), .A2(n36045), .ZN(n34810) );
  NAND2_X1 U35360 ( .A1(n34811), .A2(n34810), .ZN(n36042) );
  OAI21_X1 U35361 ( .B1(n36041), .B2(n36040), .A(n36042), .ZN(n34813) );
  NAND2_X1 U35362 ( .A1(n36041), .A2(n36040), .ZN(n34812) );
  NAND2_X1 U35363 ( .A1(n34813), .A2(n34812), .ZN(n35471) );
  XNOR2_X1 U35364 ( .A(n35470), .B(n35471), .ZN(n34818) );
  XNOR2_X1 U35365 ( .A(n34815), .B(n34814), .ZN(n34817) );
  XNOR2_X1 U35366 ( .A(n34818), .B(n35469), .ZN(n36644) );
  OAI21_X1 U35367 ( .B1(n36641), .B2(n36642), .A(n36644), .ZN(n34820) );
  NAND2_X1 U35368 ( .A1(n3284), .A2(n36642), .ZN(n34819) );
  NAND2_X1 U35369 ( .A1(n34820), .A2(n34819), .ZN(n36647) );
  INV_X1 U35370 ( .A(n36442), .ZN(n34822) );
  NAND2_X1 U35371 ( .A1(n36440), .A2(n36439), .ZN(n34821) );
  OAI21_X1 U35372 ( .B1(n34823), .B2(n34822), .A(n34821), .ZN(n36024) );
  OAI21_X1 U35373 ( .B1(n34832), .B2(n34831), .A(n34830), .ZN(n34834) );
  NAND2_X1 U35374 ( .A1(n34834), .A2(n34833), .ZN(n35079) );
  NAND2_X1 U35375 ( .A1(n34842), .A2(n34841), .ZN(n35078) );
  FA_X1 U35376 ( .A(n34845), .B(n34844), .CI(n34843), .CO(n35369), .S(n34953)
         );
  OAI21_X1 U35377 ( .B1(n34848), .B2(n34847), .A(n34846), .ZN(n34850) );
  NAND2_X1 U35378 ( .A1(n34848), .A2(n34847), .ZN(n34849) );
  NAND2_X1 U35379 ( .A1(n34850), .A2(n34849), .ZN(n35379) );
  FA_X1 U35380 ( .A(n34853), .B(n34852), .CI(n34851), .CO(n35378), .S(n34893)
         );
  OAI21_X1 U35381 ( .B1(n34855), .B2(n34856), .A(n34854), .ZN(n34858) );
  NAND2_X1 U35382 ( .A1(n34858), .A2(n34857), .ZN(n35225) );
  OAI22_X1 U35383 ( .A1(n34983), .A2(n35745), .B1(n35744), .B2(n34860), .ZN(
        n35144) );
  XNOR2_X1 U35384 ( .A(n35338), .B(\fmem_data[9][5] ), .ZN(n35039) );
  XNOR2_X1 U35385 ( .A(n34862), .B(\fmem_data[16][7] ), .ZN(n34981) );
  OAI22_X1 U35386 ( .A1(n34863), .A2(n35752), .B1(n34981), .B2(n35753), .ZN(
        n35142) );
  FA_X1 U35387 ( .A(n34866), .B(n34865), .CI(n34864), .CO(n35164), .S(n35185)
         );
  XNOR2_X1 U35388 ( .A(n35184), .B(n35185), .ZN(n34874) );
  INV_X1 U35389 ( .A(n34870), .ZN(n34867) );
  NAND2_X1 U35390 ( .A1(n34867), .A2(n14573), .ZN(n34868) );
  NAND2_X1 U35391 ( .A1(n34869), .A2(n34868), .ZN(n34873) );
  NAND2_X1 U35392 ( .A1(n34871), .A2(n34870), .ZN(n34872) );
  NAND2_X1 U35393 ( .A1(n34873), .A2(n34872), .ZN(n35186) );
  XNOR2_X1 U35394 ( .A(n34874), .B(n35186), .ZN(n35200) );
  FA_X1 U35395 ( .A(n34877), .B(n34876), .CI(n34875), .CO(n35149), .S(n12720)
         );
  FA_X1 U35396 ( .A(n34880), .B(n34879), .CI(n34878), .CO(n35148), .S(n18725)
         );
  FA_X1 U35397 ( .A(n34883), .B(n34882), .CI(n34881), .CO(n35132), .S(n35147)
         );
  XNOR2_X1 U35398 ( .A(n35200), .B(n35199), .ZN(n34887) );
  FA_X1 U35399 ( .A(n34886), .B(n34885), .CI(n34884), .CO(n35198), .S(n34854)
         );
  XNOR2_X1 U35400 ( .A(n34887), .B(n35198), .ZN(n35224) );
  FA_X1 U35401 ( .A(n34890), .B(n34889), .CI(n34888), .CO(n35223), .S(n35228)
         );
  FA_X1 U35402 ( .A(n34893), .B(n34892), .CI(n34891), .CO(n35381), .S(n34896)
         );
  OAI21_X1 U35403 ( .B1(n34895), .B2(n34896), .A(n34894), .ZN(n34898) );
  NAND2_X1 U35404 ( .A1(n34898), .A2(n34897), .ZN(n35230) );
  FA_X1 U35405 ( .A(n34901), .B(n34900), .CI(n34899), .CO(n35354), .S(n34952)
         );
  INV_X1 U35406 ( .A(n34902), .ZN(n34906) );
  INV_X1 U35407 ( .A(n34910), .ZN(n35245) );
  FA_X1 U35408 ( .A(n34913), .B(n34912), .CI(n34911), .CO(n35244), .S(n34899)
         );
  FA_X1 U35409 ( .A(n34916), .B(n34915), .CI(n34914), .CO(n35352), .S(n34853)
         );
  AOI21_X1 U35410 ( .B1(n34919), .B2(n34918), .A(n34917), .ZN(n34920) );
  INV_X1 U35411 ( .A(n34920), .ZN(n35363) );
  AOI21_X1 U35412 ( .B1(n34923), .B2(n34922), .A(n34921), .ZN(n34924) );
  INV_X1 U35413 ( .A(n34924), .ZN(n35362) );
  XNOR2_X1 U35414 ( .A(n35363), .B(n35362), .ZN(n34928) );
  FA_X1 U35415 ( .A(n34927), .B(n34926), .CI(n34925), .CO(n35361), .S(n34915)
         );
  XNOR2_X1 U35416 ( .A(n34928), .B(n35361), .ZN(n35101) );
  XNOR2_X1 U35417 ( .A(n34929), .B(\fmem_data[6][7] ), .ZN(n35121) );
  INV_X1 U35418 ( .A(n34931), .ZN(n34935) );
  NAND2_X1 U35419 ( .A1(n34933), .A2(n34932), .ZN(n34934) );
  NAND2_X1 U35420 ( .A1(n34935), .A2(n34934), .ZN(n35068) );
  XNOR2_X1 U35421 ( .A(n35069), .B(n35068), .ZN(n34939) );
  FA_X1 U35422 ( .A(n34938), .B(n34937), .CI(n34936), .CO(n35067), .S(n34844)
         );
  XNOR2_X1 U35423 ( .A(n34939), .B(n35067), .ZN(n35100) );
  AOI21_X1 U35424 ( .B1(n34942), .B2(n34941), .A(n34940), .ZN(n34943) );
  AND2_X1 U35425 ( .A1(n34945), .A2(n34944), .ZN(n34946) );
  FA_X1 U35426 ( .A(n34950), .B(n34949), .CI(n34948), .CO(n35367), .S(n34914)
         );
  XNOR2_X1 U35427 ( .A(n35375), .B(n35374), .ZN(n34954) );
  FA_X1 U35428 ( .A(n34953), .B(n34952), .CI(n34951), .CO(n35373), .S(n34957)
         );
  XNOR2_X1 U35429 ( .A(n34954), .B(n35373), .ZN(n35386) );
  FA_X1 U35430 ( .A(n34957), .B(n34956), .CI(n34955), .CO(n35385), .S(n34895)
         );
  XNOR2_X1 U35431 ( .A(n35386), .B(n35385), .ZN(n34963) );
  OAI21_X1 U35432 ( .B1(n34960), .B2(n34959), .A(n34958), .ZN(n34962) );
  NAND2_X1 U35433 ( .A1(n34960), .A2(n34959), .ZN(n34961) );
  NAND2_X1 U35434 ( .A1(n34962), .A2(n34961), .ZN(n35384) );
  XNOR2_X1 U35435 ( .A(n34963), .B(n35384), .ZN(n35229) );
  OAI21_X1 U35436 ( .B1(n34965), .B2(n34966), .A(n34964), .ZN(n34968) );
  NAND2_X1 U35437 ( .A1(n34968), .A2(n34967), .ZN(n35477) );
  INV_X1 U35438 ( .A(n34969), .ZN(n34974) );
  NOR2_X1 U35439 ( .A1(n34971), .A2(n34970), .ZN(n34973) );
  OAI21_X1 U35440 ( .B1(n34974), .B2(n34973), .A(n34972), .ZN(n35298) );
  OAI21_X1 U35441 ( .B1(n34977), .B2(n34976), .A(n34975), .ZN(n34979) );
  NAND2_X1 U35442 ( .A1(n34979), .A2(n34978), .ZN(n35237) );
  INV_X1 U35443 ( .A(n34987), .ZN(n35267) );
  FA_X1 U35444 ( .A(n34994), .B(n34993), .CI(n34992), .CO(n35247), .S(n34975)
         );
  FA_X1 U35445 ( .A(n34997), .B(n34996), .CI(n34995), .CO(n35235), .S(n34998)
         );
  OAI21_X1 U35446 ( .B1(n34999), .B2(n35000), .A(n34998), .ZN(n35002) );
  NAND2_X1 U35447 ( .A1(n35000), .A2(n34999), .ZN(n35001) );
  NAND2_X1 U35448 ( .A1(n35002), .A2(n35001), .ZN(n35233) );
  FA_X1 U35449 ( .A(n35016), .B(n35015), .CI(n35014), .CO(n35278), .S(n34996)
         );
  INV_X1 U35450 ( .A(n35020), .ZN(n35262) );
  OAI21_X1 U35451 ( .B1(n35027), .B2(n35026), .A(n35025), .ZN(n35029) );
  NAND2_X1 U35452 ( .A1(n35027), .A2(n35026), .ZN(n35028) );
  NAND2_X1 U35453 ( .A1(n35029), .A2(n35028), .ZN(n35251) );
  INV_X1 U35454 ( .A(n35035), .ZN(n35282) );
  INV_X1 U35455 ( .A(n35042), .ZN(n35284) );
  FA_X1 U35456 ( .A(n35046), .B(n35045), .CI(n35044), .CO(n35263), .S(n34995)
         );
  FA_X1 U35457 ( .A(n35047), .B(n35048), .CI(n35049), .CO(n35304), .S(n32049)
         );
  FA_X1 U35458 ( .A(n35052), .B(n35051), .CI(n35050), .CO(n35303), .S(n34960)
         );
  XNOR2_X1 U35459 ( .A(n35304), .B(n35303), .ZN(n35056) );
  FA_X1 U35460 ( .A(n35055), .B(n35054), .CI(n35053), .CO(n35302), .S(n32050)
         );
  XNOR2_X1 U35461 ( .A(n35056), .B(n35302), .ZN(n35296) );
  OAI21_X1 U35462 ( .B1(n35059), .B2(n35058), .A(n35057), .ZN(n35061) );
  NAND2_X1 U35463 ( .A1(n35059), .A2(n35058), .ZN(n35060) );
  NAND2_X1 U35464 ( .A1(n35061), .A2(n35060), .ZN(n35390) );
  OAI21_X1 U35465 ( .B1(n35064), .B2(n35063), .A(n35062), .ZN(n35066) );
  NAND2_X1 U35466 ( .A1(n35064), .A2(n35063), .ZN(n35065) );
  NAND2_X1 U35467 ( .A1(n35066), .A2(n35065), .ZN(n35389) );
  XNOR2_X1 U35468 ( .A(n35072), .B(\fmem_data[22][7] ), .ZN(n35583) );
  XNOR2_X1 U35469 ( .A(n35073), .B(\fmem_data[22][7] ), .ZN(n35176) );
  XNOR2_X1 U35470 ( .A(n35074), .B(\fmem_data[17][7] ), .ZN(n35579) );
  OAI22_X1 U35471 ( .A1(n35707), .A2(n35709), .B1(n35077), .B2(n35708), .ZN(
        n35714) );
  FA_X1 U35472 ( .A(n35079), .B(n3496), .CI(n35078), .CO(n35732), .S(n35370)
         );
  FA_X1 U35473 ( .A(n35082), .B(n35081), .CI(n35080), .CO(n35152), .S(n35160)
         );
  AND2_X1 U35474 ( .A1(n35084), .A2(n35083), .ZN(n35085) );
  FA_X1 U35475 ( .A(n35093), .B(n35092), .CI(n35091), .CO(n35116), .S(n35080)
         );
  OAI21_X1 U35476 ( .B1(n35096), .B2(n35095), .A(n35094), .ZN(n35098) );
  NAND2_X1 U35477 ( .A1(n35098), .A2(n35097), .ZN(n35150) );
  FA_X1 U35478 ( .A(n35101), .B(n35100), .CI(n35099), .CO(n35766), .S(n35374)
         );
  XNOR2_X1 U35479 ( .A(n35104), .B(\fmem_data[13][7] ), .ZN(n35590) );
  XNOR2_X1 U35480 ( .A(n35106), .B(\fmem_data[26][7] ), .ZN(n35710) );
  OAI22_X1 U35481 ( .A1(n35711), .A2(n35107), .B1(n35710), .B2(n35712), .ZN(
        n35755) );
  XNOR2_X1 U35482 ( .A(n35108), .B(\fmem_data[18][7] ), .ZN(n35703) );
  OAI22_X1 U35483 ( .A1(n35703), .A2(n35705), .B1(n35109), .B2(n35704), .ZN(
        n35756) );
  XNOR2_X1 U35484 ( .A(n35755), .B(n35756), .ZN(n35717) );
  XNOR2_X1 U35485 ( .A(n35110), .B(\fmem_data[31][7] ), .ZN(n35257) );
  XNOR2_X1 U35486 ( .A(n35112), .B(\fmem_data[11][7] ), .ZN(n35239) );
  FA_X1 U35487 ( .A(n3879), .B(n35117), .CI(n35116), .CO(n35692), .S(n35151)
         );
  HA_X1 U35488 ( .A(n35119), .B(n35118), .CO(n35670), .S(n35333) );
  OAI22_X1 U35489 ( .A1(n35510), .A2(n35512), .B1(n35121), .B2(n35511), .ZN(
        n35669) );
  OAI22_X1 U35490 ( .A1(n35514), .A2(n35516), .B1(n35123), .B2(n35515), .ZN(
        n35668) );
  INV_X1 U35491 ( .A(n35133), .ZN(n35130) );
  NAND2_X1 U35492 ( .A1(n31823), .A2(n35130), .ZN(n35131) );
  NAND2_X1 U35493 ( .A1(n35132), .A2(n35131), .ZN(n35136) );
  NAND2_X1 U35494 ( .A1(n35136), .A2(n35135), .ZN(n35644) );
  FA_X1 U35495 ( .A(n35139), .B(n35138), .CI(n35137), .CO(n35693), .S(n35194)
         );
  XNOR2_X1 U35496 ( .A(n35140), .B(\fmem_data[7][7] ), .ZN(n35360) );
  FA_X1 U35497 ( .A(n35144), .B(n35143), .CI(n35142), .CO(n35168), .S(n35184)
         );
  XNOR2_X1 U35498 ( .A(n35145), .B(\fmem_data[27][7] ), .ZN(n35243) );
  OAI22_X1 U35499 ( .A1(n35146), .A2(n35641), .B1(n35243), .B2(n35642), .ZN(
        n35167) );
  FA_X1 U35500 ( .A(n35149), .B(n35148), .CI(n35147), .CO(n35192), .S(n35199)
         );
  FA_X1 U35501 ( .A(n35152), .B(n35151), .CI(n35150), .CO(n35767), .S(n35205)
         );
  OAI21_X1 U35502 ( .B1(n35155), .B2(n35154), .A(n35153), .ZN(n35157) );
  NAND2_X1 U35503 ( .A1(n35155), .A2(n35154), .ZN(n35156) );
  FA_X1 U35504 ( .A(n35160), .B(n35159), .CI(n35158), .CO(n35203), .S(n35211)
         );
  FA_X1 U35505 ( .A(n35163), .B(n35162), .CI(n35161), .CO(n35673), .S(n35172)
         );
  FA_X1 U35506 ( .A(n35166), .B(n35165), .CI(n35164), .CO(n35672), .S(n35171)
         );
  FA_X1 U35507 ( .A(n35169), .B(n35168), .CI(n35167), .CO(n35671), .S(n35193)
         );
  FA_X1 U35508 ( .A(n35170), .B(n35171), .CI(n35172), .CO(n35690), .S(n35191)
         );
  FA_X1 U35509 ( .A(n35175), .B(n35174), .CI(n35173), .CO(n35197), .S(n35155)
         );
  OAI22_X1 U35510 ( .A1(n35179), .A2(n35740), .B1(n35341), .B2(n35739), .ZN(
        n35393) );
  INV_X1 U35511 ( .A(n35183), .ZN(n35392) );
  OAI21_X1 U35512 ( .B1(n35185), .B2(n35186), .A(n35184), .ZN(n35188) );
  NAND2_X1 U35513 ( .A1(n35188), .A2(n35187), .ZN(n35195) );
  FA_X1 U35514 ( .A(n35191), .B(n35190), .CI(n35189), .CO(n35678), .S(n35426)
         );
  FA_X1 U35515 ( .A(n35194), .B(n35193), .CI(n35192), .CO(n35686), .S(n35208)
         );
  FA_X1 U35516 ( .A(n35197), .B(n35196), .CI(n35195), .CO(n35689), .S(n35207)
         );
  OAI21_X1 U35517 ( .B1(n35200), .B2(n35199), .A(n35198), .ZN(n35202) );
  NAND2_X1 U35518 ( .A1(n35200), .A2(n35199), .ZN(n35201) );
  NAND2_X1 U35519 ( .A1(n35202), .A2(n35201), .ZN(n35206) );
  FA_X1 U35520 ( .A(n35205), .B(n35204), .CI(n35203), .CO(n35683), .S(n35214)
         );
  FA_X1 U35521 ( .A(n35208), .B(n35207), .CI(n35206), .CO(n35677), .S(n35213)
         );
  FA_X1 U35522 ( .A(n35211), .B(n35210), .CI(n35209), .CO(n35212), .S(n35217)
         );
  FA_X1 U35523 ( .A(n35214), .B(n35213), .CI(n35212), .CO(n35680), .S(n35443)
         );
  FA_X1 U35524 ( .A(n35217), .B(n35216), .CI(n35215), .CO(n35442), .S(n35440)
         );
  OAI21_X1 U35525 ( .B1(n35219), .B2(n3419), .A(n35218), .ZN(n35222) );
  NAND2_X1 U35526 ( .A1(n3419), .A2(n35219), .ZN(n35221) );
  NAND2_X1 U35527 ( .A1(n35222), .A2(n35221), .ZN(n35446) );
  FA_X1 U35528 ( .A(n35225), .B(n35224), .CI(n35223), .CO(n35382), .S(n35445)
         );
  FA_X1 U35529 ( .A(n35228), .B(n35227), .CI(n35226), .CO(n35444), .S(n35451)
         );
  FA_X1 U35530 ( .A(n35231), .B(n35230), .CI(n35229), .CO(n35546), .S(n35478)
         );
  FA_X1 U35531 ( .A(n35232), .B(n35233), .CI(n35234), .CO(n35535), .S(n35297)
         );
  FA_X1 U35532 ( .A(n35237), .B(n35236), .CI(n35235), .CO(n35529), .S(n35234)
         );
  XNOR2_X1 U35533 ( .A(n35238), .B(\fmem_data[11][7] ), .ZN(n35632) );
  XNOR2_X1 U35534 ( .A(n35240), .B(\fmem_data[3][7] ), .ZN(n35636) );
  OAI22_X1 U35535 ( .A1(n35636), .A2(n35638), .B1(n35241), .B2(n35637), .ZN(
        n35501) );
  FA_X1 U35536 ( .A(n35246), .B(n35245), .CI(n35244), .CO(n35525), .S(n35353)
         );
  FA_X1 U35537 ( .A(n35249), .B(n35248), .CI(n35247), .CO(n35524), .S(n35236)
         );
  FA_X1 U35538 ( .A(n35252), .B(n35251), .CI(n35250), .CO(n35527), .S(n35232)
         );
  FA_X1 U35539 ( .A(n35255), .B(n35254), .CI(n35253), .CO(n35561), .S(n35308)
         );
  XNOR2_X1 U35540 ( .A(n3462), .B(\fmem_data[23][7] ), .ZN(n35650) );
  FA_X1 U35541 ( .A(n35262), .B(n35261), .CI(n35260), .CO(n35518), .S(n35277)
         );
  XNOR2_X1 U35542 ( .A(n35561), .B(n35562), .ZN(n35266) );
  FA_X1 U35543 ( .A(n35265), .B(n35264), .CI(n35263), .CO(n35563), .S(n35250)
         );
  XNOR2_X1 U35544 ( .A(n35266), .B(n35563), .ZN(n35532) );
  FA_X1 U35545 ( .A(n35269), .B(n35268), .CI(n35267), .CO(n35505), .S(n35249)
         );
  FA_X1 U35546 ( .A(n35279), .B(n35278), .CI(n35277), .CO(n35568), .S(n35252)
         );
  XNOR2_X1 U35547 ( .A(n35569), .B(n35568), .ZN(n35290) );
  XNOR2_X1 U35548 ( .A(n35280), .B(\fmem_data[1][7] ), .ZN(n35699) );
  OAI21_X1 U35549 ( .B1(n35284), .B2(n35283), .A(n35282), .ZN(n35286) );
  FA_X1 U35550 ( .A(n35289), .B(n35288), .CI(n35287), .CO(n35521), .S(n35254)
         );
  XNOR2_X1 U35551 ( .A(n35290), .B(n35567), .ZN(n35531) );
  OAI21_X1 U35552 ( .B1(n35292), .B2(n35293), .A(n35291), .ZN(n35295) );
  NAND2_X1 U35553 ( .A1(n35295), .A2(n35294), .ZN(n35530) );
  FA_X1 U35554 ( .A(n35297), .B(n35298), .CI(n35296), .CO(n35544), .S(n35391)
         );
  FA_X1 U35555 ( .A(n35301), .B(n35300), .CI(n35299), .CO(n35621), .S(n35429)
         );
  OAI21_X1 U35556 ( .B1(n35304), .B2(n35303), .A(n35302), .ZN(n35305) );
  NAND2_X1 U35557 ( .A1(n35306), .A2(n35305), .ZN(n35622) );
  XNOR2_X1 U35558 ( .A(n35621), .B(n35622), .ZN(n35351) );
  FA_X1 U35559 ( .A(n35307), .B(n35308), .CI(n35309), .CO(n35560), .S(n35301)
         );
  FA_X1 U35560 ( .A(n35312), .B(n35311), .CI(n35310), .CO(n35602), .S(n35291)
         );
  FA_X1 U35561 ( .A(n35315), .B(n35314), .CI(n35313), .CO(n35574), .S(n35255)
         );
  FA_X1 U35562 ( .A(n35320), .B(n35319), .CI(n35318), .CO(n35572), .S(n35312)
         );
  FA_X1 U35563 ( .A(n35323), .B(n35322), .CI(n35321), .CO(n35608), .S(n35408)
         );
  XNOR2_X1 U35564 ( .A(n35328), .B(\fmem_data[8][7] ), .ZN(n35728) );
  FA_X1 U35565 ( .A(n35332), .B(n35331), .CI(n35330), .CO(n35606), .S(n35346)
         );
  FA_X1 U35566 ( .A(n35335), .B(n35334), .CI(n35333), .CO(n35605), .S(n35409)
         );
  FA_X1 U35567 ( .A(n35344), .B(n35343), .CI(n35342), .CO(n35603), .S(n35345)
         );
  FA_X1 U35568 ( .A(n35347), .B(n35346), .CI(n35345), .CO(n35598), .S(n35419)
         );
  FA_X1 U35569 ( .A(n35350), .B(n35349), .CI(n35348), .CO(n35597), .S(n35417)
         );
  XNOR2_X1 U35570 ( .A(n35351), .B(n35623), .ZN(n35543) );
  FA_X1 U35571 ( .A(n35354), .B(n35353), .CI(n35352), .CO(n35771), .S(n35375)
         );
  XNOR2_X1 U35572 ( .A(n35355), .B(\fmem_data[10][7] ), .ZN(n35609) );
  XNOR2_X1 U35573 ( .A(n35359), .B(\fmem_data[7][7] ), .ZN(n35617) );
  FA_X1 U35574 ( .A(n35368), .B(n3714), .CI(n35367), .CO(n35763), .S(n35099)
         );
  XNOR2_X1 U35575 ( .A(n35771), .B(n35770), .ZN(n35372) );
  FA_X1 U35576 ( .A(n35371), .B(n35370), .CI(n35369), .CO(n35769), .S(n35380)
         );
  XNOR2_X1 U35577 ( .A(n35372), .B(n35769), .ZN(n35538) );
  FA_X1 U35578 ( .A(n35380), .B(n35379), .CI(n35378), .CO(n35536), .S(n35383)
         );
  FA_X1 U35579 ( .A(n35383), .B(n35382), .CI(n35381), .CO(n35541), .S(n35231)
         );
  FA_X1 U35580 ( .A(n35391), .B(n35390), .CI(n35389), .CO(n35549), .S(n35476)
         );
  FA_X1 U35581 ( .A(n35394), .B(n35393), .CI(n35392), .CO(n35631), .S(n35196)
         );
  XNOR2_X1 U35582 ( .A(n35397), .B(\fmem_data[16][7] ), .ZN(n35751) );
  XNOR2_X1 U35583 ( .A(n35399), .B(\fmem_data[28][7] ), .ZN(n35759) );
  OAI22_X1 U35584 ( .A1(n35759), .A2(n35761), .B1(n35400), .B2(n35760), .ZN(
        n35665) );
  OAI22_X1 U35585 ( .A1(n35496), .A2(n35498), .B1(n35406), .B2(n35497), .ZN(
        n35658) );
  FA_X1 U35586 ( .A(n35409), .B(n35408), .CI(n35407), .CO(n35648), .S(n35307)
         );
  OAI21_X1 U35587 ( .B1(n35412), .B2(n35411), .A(n35410), .ZN(n35414) );
  NAND2_X1 U35588 ( .A1(n35412), .A2(n35411), .ZN(n35413) );
  NAND2_X1 U35589 ( .A1(n35414), .A2(n35413), .ZN(n35647) );
  FA_X1 U35590 ( .A(n35417), .B(n35416), .CI(n35415), .CO(n35675), .S(n35423)
         );
  FA_X1 U35591 ( .A(n35420), .B(n35419), .CI(n35418), .CO(n35674), .S(n35422)
         );
  FA_X1 U35592 ( .A(n35422), .B(n35423), .CI(n35421), .CO(n35627), .S(n35431)
         );
  FA_X1 U35593 ( .A(n35426), .B(n35425), .CI(n35424), .CO(n35626), .S(n35430)
         );
  FA_X1 U35594 ( .A(n35429), .B(n35428), .CI(n35427), .CO(n35556), .S(n35435)
         );
  FA_X1 U35595 ( .A(n35432), .B(n35431), .CI(n35430), .CO(n35555), .S(n35433)
         );
  OAI21_X1 U35596 ( .B1(n35434), .B2(n35435), .A(n35433), .ZN(n35437) );
  NAND2_X1 U35597 ( .A1(n35435), .A2(n35434), .ZN(n35436) );
  NAND2_X1 U35598 ( .A1(n35437), .A2(n35436), .ZN(n35778) );
  XNOR2_X1 U35599 ( .A(n35779), .B(n35778), .ZN(n35453) );
  FA_X1 U35600 ( .A(n35440), .B(n35439), .CI(n35438), .CO(n35462), .S(n33406)
         );
  FA_X1 U35601 ( .A(n35443), .B(n35442), .CI(n35441), .CO(n35547), .S(n35461)
         );
  FA_X1 U35602 ( .A(n35446), .B(n35445), .CI(n35444), .CO(n35441), .S(n35465)
         );
  FA_X1 U35603 ( .A(n35447), .B(n35448), .CI(n35449), .CO(n35464), .S(n35468)
         );
  FA_X1 U35604 ( .A(n35452), .B(n35451), .CI(n35450), .CO(n35463), .S(n35470)
         );
  XNOR2_X1 U35605 ( .A(n35453), .B(n35777), .ZN(n35485) );
  INV_X1 U35606 ( .A(n35454), .ZN(n35459) );
  NOR2_X1 U35607 ( .A1(n3277), .A2(n35456), .ZN(n35458) );
  NAND2_X1 U35608 ( .A1(n35456), .A2(n3277), .ZN(n35457) );
  XNOR2_X1 U35609 ( .A(n35485), .B(n35484), .ZN(n35481) );
  FA_X1 U35610 ( .A(n35462), .B(n35461), .CI(n35460), .CO(n35777), .S(n36434)
         );
  FA_X1 U35611 ( .A(n35465), .B(n35464), .CI(n35463), .CO(n35460), .S(n36029)
         );
  FA_X1 U35612 ( .A(n35468), .B(n35467), .CI(n35466), .CO(n36028), .S(n36641)
         );
  OAI21_X1 U35613 ( .B1(n3355), .B2(n35470), .A(n35469), .ZN(n35473) );
  NAND2_X1 U35614 ( .A1(n3355), .A2(n35470), .ZN(n35472) );
  NAND2_X1 U35615 ( .A1(n35473), .A2(n35472), .ZN(n36030) );
  OAI21_X1 U35616 ( .B1(n36029), .B2(n36028), .A(n36030), .ZN(n35475) );
  NAND2_X1 U35617 ( .A1(n36029), .A2(n36028), .ZN(n35474) );
  NAND2_X1 U35618 ( .A1(n35475), .A2(n35474), .ZN(n36435) );
  FA_X1 U35619 ( .A(n35478), .B(n35477), .CI(n35476), .CO(n35554), .S(n36436)
         );
  OAI21_X1 U35620 ( .B1(n36434), .B2(n36435), .A(n36436), .ZN(n35480) );
  NAND2_X1 U35621 ( .A1(n36435), .A2(n36434), .ZN(n35479) );
  NAND2_X1 U35622 ( .A1(n35480), .A2(n35479), .ZN(n35483) );
  XNOR2_X1 U35623 ( .A(n35481), .B(n3422), .ZN(n36022) );
  INV_X1 U35624 ( .A(n37145), .ZN(n35785) );
  OR2_X1 U35625 ( .A1(n35485), .A2(n35484), .ZN(n35482) );
  NAND2_X1 U35626 ( .A1(n35483), .A2(n35482), .ZN(n35487) );
  NAND2_X1 U35627 ( .A1(n35485), .A2(n35484), .ZN(n35486) );
  NAND2_X1 U35628 ( .A1(n35487), .A2(n35486), .ZN(n36013) );
  FA_X1 U35629 ( .A(n35502), .B(n35501), .CI(n35500), .CO(n35817), .S(n35526)
         );
  FA_X1 U35630 ( .A(n35505), .B(n35504), .CI(n35503), .CO(n35816), .S(n35569)
         );
  FA_X1 U35631 ( .A(n35520), .B(n35519), .CI(n35518), .CO(n35814), .S(n35562)
         );
  FA_X1 U35632 ( .A(n35523), .B(n35522), .CI(n35521), .CO(n35813), .S(n35567)
         );
  FA_X1 U35633 ( .A(n35526), .B(n35525), .CI(n35524), .CO(n35828), .S(n35528)
         );
  FA_X1 U35634 ( .A(n35529), .B(n35528), .CI(n35527), .CO(n35790), .S(n35534)
         );
  FA_X1 U35635 ( .A(n35532), .B(n35531), .CI(n35530), .CO(n35789), .S(n35533)
         );
  FA_X1 U35636 ( .A(n35535), .B(n35534), .CI(n35533), .CO(n35909), .S(n35545)
         );
  FA_X1 U35637 ( .A(n35538), .B(n35537), .CI(n35536), .CO(n35910), .S(n35542)
         );
  FA_X1 U35638 ( .A(n35542), .B(n35541), .CI(n35540), .CO(n35949), .S(n35550)
         );
  FA_X1 U35639 ( .A(n35545), .B(n35544), .CI(n35543), .CO(n35948), .S(n35551)
         );
  FA_X1 U35640 ( .A(n35548), .B(n35547), .CI(n35546), .CO(n35971), .S(n35553)
         );
  FA_X1 U35641 ( .A(n35549), .B(n35550), .CI(n35551), .CO(n35970), .S(n35552)
         );
  XNOR2_X1 U35642 ( .A(n36013), .B(n36014), .ZN(n35784) );
  FA_X1 U35643 ( .A(n35554), .B(n35553), .CI(n35552), .CO(n35973), .S(n36023)
         );
  FA_X1 U35644 ( .A(n35557), .B(n35556), .CI(n35555), .CO(n35956), .S(n35779)
         );
  FA_X1 U35645 ( .A(n35560), .B(n35559), .CI(n35558), .CO(n35857), .S(n35623)
         );
  FA_X1 U35646 ( .A(n35574), .B(n35573), .CI(n35572), .CO(n35839), .S(n35601)
         );
  INV_X1 U35647 ( .A(n35578), .ZN(n35821) );
  INV_X1 U35648 ( .A(n35582), .ZN(n35820) );
  INV_X1 U35649 ( .A(n35586), .ZN(n35819) );
  FA_X1 U35650 ( .A(n35589), .B(n35588), .CI(n35587), .CO(n35827), .S(n35604)
         );
  INV_X1 U35651 ( .A(n35593), .ZN(n35826) );
  FA_X1 U35652 ( .A(n35596), .B(n35595), .CI(n35594), .CO(n35825), .S(n35607)
         );
  FA_X1 U35653 ( .A(n35599), .B(n35598), .CI(n35597), .CO(n35851), .S(n35558)
         );
  FA_X1 U35654 ( .A(n35602), .B(n35601), .CI(n35600), .CO(n35850), .S(n35559)
         );
  FA_X1 U35655 ( .A(n35605), .B(n35604), .CI(n35603), .CO(n35836), .S(n35599)
         );
  FA_X1 U35656 ( .A(n35608), .B(n35607), .CI(n35606), .CO(n35835), .S(n35600)
         );
  INV_X1 U35657 ( .A(n35612), .ZN(n35845) );
  INV_X1 U35658 ( .A(n35616), .ZN(n35844) );
  INV_X1 U35659 ( .A(n35620), .ZN(n35843) );
  FA_X1 U35660 ( .A(n35628), .B(n35627), .CI(n35626), .CO(n35786), .S(n35557)
         );
  FA_X1 U35661 ( .A(n35631), .B(n35630), .CI(n35629), .CO(n35884), .S(n35649)
         );
  INV_X1 U35662 ( .A(n35635), .ZN(n35842) );
  INV_X1 U35663 ( .A(n35639), .ZN(n35841) );
  INV_X1 U35664 ( .A(n35643), .ZN(n35840) );
  FA_X1 U35665 ( .A(n35646), .B(n35645), .CI(n35644), .CO(n35882), .S(n35687)
         );
  FA_X1 U35666 ( .A(n35649), .B(n35648), .CI(n35647), .CO(n35853), .S(n35676)
         );
  INV_X1 U35667 ( .A(n35653), .ZN(n35866) );
  INV_X1 U35668 ( .A(n35657), .ZN(n35865) );
  FA_X1 U35669 ( .A(n35660), .B(n35659), .CI(n35658), .CO(n35864), .S(n35629)
         );
  INV_X1 U35670 ( .A(n35664), .ZN(n35848) );
  FA_X1 U35671 ( .A(n35667), .B(n35666), .CI(n35665), .CO(n35847), .S(n35630)
         );
  FA_X1 U35672 ( .A(n35670), .B(n35669), .CI(n35668), .CO(n35846), .S(n35646)
         );
  FA_X1 U35673 ( .A(n35673), .B(n35672), .CI(n35671), .CO(n35879), .S(n35691)
         );
  FA_X1 U35674 ( .A(n35676), .B(n35675), .CI(n35674), .CO(n35859), .S(n35628)
         );
  FA_X1 U35675 ( .A(n35679), .B(n35678), .CI(n35677), .CO(n35858), .S(n35681)
         );
  FA_X1 U35676 ( .A(n35682), .B(n35681), .CI(n35680), .CO(n35946), .S(n35548)
         );
  FA_X1 U35677 ( .A(n35685), .B(n35684), .CI(n35683), .CO(n35905), .S(n35682)
         );
  FA_X1 U35678 ( .A(n35688), .B(n35687), .CI(n35686), .CO(n35893), .S(n35684)
         );
  FA_X1 U35679 ( .A(n35691), .B(n35690), .CI(n35689), .CO(n35892), .S(n35679)
         );
  FA_X1 U35680 ( .A(n35694), .B(n35693), .CI(n35692), .CO(n35797), .S(n35688)
         );
  INV_X1 U35681 ( .A(n35698), .ZN(n35863) );
  INV_X1 U35682 ( .A(n35702), .ZN(n35862) );
  INV_X1 U35683 ( .A(n35706), .ZN(n35868) );
  INV_X1 U35684 ( .A(n35713), .ZN(n35867) );
  FA_X1 U35685 ( .A(n35716), .B(n35715), .CI(n35714), .CO(n35803), .S(n35733)
         );
  FA_X1 U35686 ( .A(n35719), .B(n35718), .CI(n35717), .CO(n35802), .S(n35694)
         );
  AOI21_X1 U35687 ( .B1(n35722), .B2(n35721), .A(n35720), .ZN(n35723) );
  INV_X1 U35688 ( .A(n35723), .ZN(n35872) );
  INV_X1 U35689 ( .A(n35727), .ZN(n35871) );
  INV_X1 U35690 ( .A(n35731), .ZN(n35870) );
  FA_X1 U35691 ( .A(n35734), .B(n35733), .CI(n35732), .CO(n35794), .S(n35768)
         );
  FA_X1 U35692 ( .A(n35737), .B(n35736), .CI(n35735), .CO(n35800), .S(n35765)
         );
  INV_X1 U35693 ( .A(n35738), .ZN(n35742) );
  NAND2_X1 U35694 ( .A1(n35740), .A2(n35739), .ZN(n35741) );
  NAND2_X1 U35695 ( .A1(n35742), .A2(n35741), .ZN(n35809) );
  AOI21_X1 U35696 ( .B1(n35745), .B2(n35744), .A(n35743), .ZN(n35746) );
  INV_X1 U35697 ( .A(n35746), .ZN(n35808) );
  AOI21_X1 U35698 ( .B1(n35749), .B2(n35748), .A(n35747), .ZN(n35750) );
  INV_X1 U35699 ( .A(n35750), .ZN(n35807) );
  INV_X1 U35700 ( .A(n35754), .ZN(n35806) );
  INV_X1 U35701 ( .A(n35755), .ZN(n35758) );
  INV_X1 U35702 ( .A(n35756), .ZN(n35757) );
  NAND2_X1 U35703 ( .A1(n35758), .A2(n35757), .ZN(n35805) );
  INV_X1 U35704 ( .A(n35762), .ZN(n35804) );
  FA_X1 U35705 ( .A(n35765), .B(n35764), .CI(n35763), .CO(n35792), .S(n35770)
         );
  FA_X1 U35706 ( .A(n35768), .B(n35767), .CI(n35766), .CO(n35898), .S(n35685)
         );
  OAI21_X1 U35707 ( .B1(n35771), .B2(n35770), .A(n35769), .ZN(n35773) );
  NAND2_X1 U35708 ( .A1(n35771), .A2(n35770), .ZN(n35772) );
  NAND2_X1 U35709 ( .A1(n35773), .A2(n35772), .ZN(n35897) );
  INV_X1 U35710 ( .A(n35779), .ZN(n35775) );
  INV_X1 U35711 ( .A(n35778), .ZN(n35774) );
  NAND2_X1 U35712 ( .A1(n35775), .A2(n35774), .ZN(n35776) );
  NAND2_X1 U35713 ( .A1(n35777), .A2(n35776), .ZN(n35781) );
  NAND2_X1 U35714 ( .A1(n35781), .A2(n35780), .ZN(n35975) );
  XNOR2_X1 U35715 ( .A(n35974), .B(n35975), .ZN(n35782) );
  XNOR2_X1 U35716 ( .A(n35973), .B(n35782), .ZN(n36015) );
  INV_X1 U35717 ( .A(n36015), .ZN(n35783) );
  XNOR2_X1 U35718 ( .A(n35784), .B(n35783), .ZN(n37144) );
  NAND2_X1 U35719 ( .A1(n35785), .A2(n37144), .ZN(n37205) );
  INV_X1 U35720 ( .A(n37205), .ZN(n37232) );
  FA_X1 U35721 ( .A(n35788), .B(n35787), .CI(n35786), .CO(n35959), .S(n35955)
         );
  FA_X1 U35722 ( .A(n35791), .B(n35790), .CI(n35789), .CO(n35902), .S(n35911)
         );
  FA_X1 U35723 ( .A(n35794), .B(n35793), .CI(n35792), .CO(n35890), .S(n35899)
         );
  FA_X1 U35724 ( .A(n35797), .B(n35796), .CI(n35795), .CO(n35889), .S(n35891)
         );
  FA_X1 U35725 ( .A(n35800), .B(n35799), .CI(n35798), .CO(n35878), .S(n35793)
         );
  FA_X1 U35726 ( .A(n35803), .B(n35802), .CI(n35801), .CO(n35877), .S(n35795)
         );
  FA_X1 U35727 ( .A(n35806), .B(n35805), .CI(n35804), .CO(n35921), .S(n35798)
         );
  FA_X1 U35728 ( .A(n35809), .B(n35808), .CI(n35807), .CO(n35920), .S(n35799)
         );
  FA_X1 U35729 ( .A(n35812), .B(n35811), .CI(n35810), .CO(n35919), .S(n35818)
         );
  FA_X1 U35730 ( .A(n35815), .B(n35814), .CI(n35813), .CO(n35930), .S(n35829)
         );
  FA_X1 U35731 ( .A(n35818), .B(n35817), .CI(n35816), .CO(n35929), .S(n35830)
         );
  FA_X1 U35732 ( .A(n35821), .B(n35820), .CI(n35819), .CO(n35927), .S(n35838)
         );
  FA_X1 U35733 ( .A(n35824), .B(n35823), .CI(n35822), .CO(n35926), .S(n35815)
         );
  FA_X1 U35734 ( .A(n35827), .B(n35826), .CI(n35825), .CO(n35925), .S(n35837)
         );
  FA_X1 U35735 ( .A(n35830), .B(n35829), .CI(n35828), .CO(n35935), .S(n35791)
         );
  FA_X1 U35736 ( .A(n35833), .B(n35832), .CI(n35831), .CO(n35934), .S(n35856)
         );
  FA_X1 U35737 ( .A(n35836), .B(n35835), .CI(n35834), .CO(n35933), .S(n35849)
         );
  FA_X1 U35738 ( .A(n35839), .B(n35838), .CI(n35837), .CO(n35932), .S(n35831)
         );
  FA_X1 U35739 ( .A(n35842), .B(n35841), .CI(n35840), .CO(n35875), .S(n35883)
         );
  FA_X1 U35740 ( .A(n35845), .B(n35844), .CI(n35843), .CO(n35874), .S(n35834)
         );
  FA_X1 U35741 ( .A(n35848), .B(n35847), .CI(n35846), .CO(n35873), .S(n35880)
         );
  FA_X1 U35742 ( .A(n35851), .B(n35850), .CI(n35849), .CO(n35938), .S(n35855)
         );
  FA_X1 U35743 ( .A(n35854), .B(n35853), .CI(n35852), .CO(n35937), .S(n35860)
         );
  FA_X1 U35744 ( .A(n35857), .B(n35856), .CI(n35855), .CO(n35917), .S(n35788)
         );
  FA_X1 U35745 ( .A(n35860), .B(n35859), .CI(n35858), .CO(n35916), .S(n35947)
         );
  FA_X1 U35746 ( .A(n35863), .B(n35862), .CI(n35861), .CO(n35887), .S(n35796)
         );
  FA_X1 U35747 ( .A(n35866), .B(n35865), .CI(n35864), .CO(n35886), .S(n35881)
         );
  FA_X1 U35748 ( .A(n35868), .B(n35869), .CI(n35867), .CO(n35924), .S(n35861)
         );
  INV_X1 U35749 ( .A(n35869), .ZN(n35923) );
  FA_X1 U35750 ( .A(n35872), .B(n35871), .CI(n35870), .CO(n35922), .S(n35801)
         );
  FA_X1 U35751 ( .A(n35875), .B(n35874), .CI(n35873), .CO(n35988), .S(n35931)
         );
  FA_X1 U35752 ( .A(n35878), .B(n35877), .CI(n35876), .CO(n35987), .S(n35888)
         );
  FA_X1 U35753 ( .A(n35881), .B(n35880), .CI(n35879), .CO(n35896), .S(n35852)
         );
  FA_X1 U35754 ( .A(n35884), .B(n35883), .CI(n35882), .CO(n35895), .S(n35854)
         );
  FA_X1 U35755 ( .A(n35887), .B(n35886), .CI(n35885), .CO(n35989), .S(n35894)
         );
  FA_X1 U35756 ( .A(n35890), .B(n35889), .CI(n35888), .CO(n35993), .S(n35901)
         );
  FA_X1 U35757 ( .A(n35893), .B(n35892), .CI(n35891), .CO(n35908), .S(n35904)
         );
  FA_X1 U35758 ( .A(n35896), .B(n35895), .CI(n35894), .CO(n35994), .S(n35907)
         );
  FA_X1 U35759 ( .A(n35899), .B(n35898), .CI(n35897), .CO(n35906), .S(n35903)
         );
  FA_X1 U35760 ( .A(n35902), .B(n35901), .CI(n35900), .CO(n35999), .S(n35958)
         );
  FA_X1 U35761 ( .A(n35905), .B(n35904), .CI(n35903), .CO(n35941), .S(n35945)
         );
  FA_X1 U35762 ( .A(n35908), .B(n35907), .CI(n35906), .CO(n36000), .S(n35942)
         );
  OAI21_X1 U35763 ( .B1(n35911), .B2(n35910), .A(n35909), .ZN(n35913) );
  NAND2_X1 U35764 ( .A1(n35911), .A2(n35910), .ZN(n35912) );
  NAND2_X1 U35765 ( .A1(n35913), .A2(n35912), .ZN(n35943) );
  OAI21_X1 U35766 ( .B1(n35941), .B2(n35942), .A(n35943), .ZN(n35915) );
  NAND2_X1 U35767 ( .A1(n35942), .A2(n35941), .ZN(n35914) );
  NAND2_X1 U35768 ( .A1(n35915), .A2(n35914), .ZN(n36007) );
  FA_X1 U35769 ( .A(n35918), .B(n35917), .CI(n35916), .CO(n36005), .S(n35957)
         );
  FA_X1 U35770 ( .A(n35921), .B(n35920), .CI(n35919), .CO(n35986), .S(n35876)
         );
  FA_X1 U35771 ( .A(n35924), .B(n35923), .CI(n35922), .CO(n37172), .S(n35885)
         );
  INV_X1 U35772 ( .A(n37172), .ZN(n35985) );
  FA_X1 U35773 ( .A(n35927), .B(n35926), .CI(n35925), .CO(n35984), .S(n35928)
         );
  FA_X1 U35774 ( .A(n35930), .B(n35929), .CI(n35928), .CO(n35991), .S(n35936)
         );
  FA_X1 U35775 ( .A(n35933), .B(n35932), .CI(n35931), .CO(n35990), .S(n35939)
         );
  FA_X1 U35776 ( .A(n35936), .B(n35935), .CI(n35934), .CO(n35997), .S(n35900)
         );
  FA_X1 U35777 ( .A(n35939), .B(n35938), .CI(n35937), .CO(n35996), .S(n35918)
         );
  XNOR2_X1 U35778 ( .A(n36005), .B(n36004), .ZN(n35940) );
  XNOR2_X1 U35779 ( .A(n36007), .B(n35940), .ZN(n36009) );
  XNOR2_X1 U35780 ( .A(n35942), .B(n35941), .ZN(n35944) );
  XNOR2_X1 U35781 ( .A(n35944), .B(n35943), .ZN(n35961) );
  FA_X1 U35782 ( .A(n35947), .B(n35946), .CI(n35945), .CO(n35960), .S(n35954)
         );
  FA_X1 U35783 ( .A(n35950), .B(n35949), .CI(n35948), .CO(n35962), .S(n35972)
         );
  FA_X1 U35784 ( .A(n35956), .B(n35955), .CI(n35954), .CO(n35967), .S(n35974)
         );
  FA_X1 U35785 ( .A(n35959), .B(n35958), .CI(n35957), .CO(n36011), .S(n35966)
         );
  XNOR2_X1 U35786 ( .A(n35961), .B(n35960), .ZN(n35963) );
  XNOR2_X1 U35787 ( .A(n35963), .B(n35962), .ZN(n35968) );
  OAI21_X1 U35788 ( .B1(n35966), .B2(n35967), .A(n35968), .ZN(n35965) );
  NAND2_X1 U35789 ( .A1(n35967), .A2(n35966), .ZN(n35964) );
  NAND2_X1 U35790 ( .A1(n35965), .A2(n35964), .ZN(n35981) );
  XNOR2_X1 U35791 ( .A(n35967), .B(n35966), .ZN(n35969) );
  XNOR2_X1 U35792 ( .A(n35969), .B(n35968), .ZN(n36019) );
  FA_X1 U35793 ( .A(n35972), .B(n35971), .CI(n35970), .CO(n36018), .S(n36014)
         );
  INV_X1 U35794 ( .A(n35973), .ZN(n35978) );
  NOR2_X1 U35795 ( .A1(n35974), .A2(n35975), .ZN(n35977) );
  OAI21_X1 U35796 ( .B1(n35978), .B2(n35977), .A(n35976), .ZN(n36021) );
  OAI21_X1 U35797 ( .B1(n36019), .B2(n36018), .A(n36021), .ZN(n35980) );
  NAND2_X1 U35798 ( .A1(n36019), .A2(n36018), .ZN(n35979) );
  NAND2_X1 U35799 ( .A1(n35980), .A2(n35979), .ZN(n37149) );
  FA_X1 U35800 ( .A(n35983), .B(n35982), .CI(n35981), .CO(n37152), .S(n37150)
         );
  FA_X1 U35801 ( .A(n35986), .B(n35985), .CI(n35984), .CO(n37173), .S(n35992)
         );
  FA_X1 U35802 ( .A(n35989), .B(n35988), .CI(n35987), .CO(n37171), .S(n35995)
         );
  FA_X1 U35803 ( .A(n35992), .B(n35991), .CI(n35990), .CO(n37169), .S(n35998)
         );
  FA_X1 U35804 ( .A(n35995), .B(n35994), .CI(n35993), .CO(n37168), .S(n36001)
         );
  FA_X1 U35805 ( .A(n35998), .B(n35997), .CI(n35996), .CO(n37175), .S(n36004)
         );
  FA_X1 U35806 ( .A(n36001), .B(n36000), .CI(n35999), .CO(n37174), .S(n36010)
         );
  FA_X1 U35807 ( .A(n36011), .B(n36010), .CI(n36009), .CO(n37165), .S(n35983)
         );
  INV_X1 U35808 ( .A(n37228), .ZN(n36012) );
  OAI21_X1 U35809 ( .B1(n36014), .B2(n36015), .A(n36013), .ZN(n36017) );
  NAND2_X1 U35810 ( .A1(n36015), .A2(n36014), .ZN(n36016) );
  NAND2_X1 U35811 ( .A1(n36017), .A2(n36016), .ZN(n37147) );
  XNOR2_X1 U35812 ( .A(n36019), .B(n36018), .ZN(n36020) );
  XNOR2_X1 U35813 ( .A(n36020), .B(n36021), .ZN(n37148) );
  OR2_X2 U35814 ( .A1(n37147), .A2(n37148), .ZN(n37239) );
  NAND2_X1 U35815 ( .A1(n37154), .A2(n37239), .ZN(n37146) );
  NOR2_X1 U35816 ( .A1(n37232), .A2(n3370), .ZN(n37163) );
  FA_X1 U35817 ( .A(n36024), .B(n36023), .CI(n36022), .CO(n37145), .S(n37162)
         );
  FA_X1 U35818 ( .A(n36027), .B(n36026), .CI(n36025), .CO(n36439), .S(n36447)
         );
  XNOR2_X1 U35819 ( .A(n36029), .B(n36028), .ZN(n36031) );
  XNOR2_X1 U35820 ( .A(n36033), .B(n36032), .ZN(n36035) );
  XNOR2_X1 U35821 ( .A(n36035), .B(n36034), .ZN(n37123) );
  XNOR2_X1 U35822 ( .A(n36037), .B(n36036), .ZN(n36039) );
  XNOR2_X1 U35823 ( .A(n36039), .B(n36038), .ZN(n36757) );
  XNOR2_X1 U35824 ( .A(n36045), .B(n36044), .ZN(n36046) );
  XNOR2_X1 U35825 ( .A(n36047), .B(n36046), .ZN(n36765) );
  XNOR2_X1 U35826 ( .A(n36053), .B(n36052), .ZN(n36054) );
  XNOR2_X1 U35827 ( .A(n36055), .B(n36054), .ZN(n36814) );
  XNOR2_X1 U35828 ( .A(n36057), .B(n36056), .ZN(n36059) );
  XNOR2_X1 U35829 ( .A(n36059), .B(n36058), .ZN(n36502) );
  FA_X1 U35830 ( .A(n36062), .B(n36061), .CI(n36060), .CO(n34570), .S(n36501)
         );
  XNOR2_X1 U35831 ( .A(n36064), .B(n36063), .ZN(n36066) );
  XNOR2_X1 U35832 ( .A(n36066), .B(n36065), .ZN(n36500) );
  FA_X1 U35833 ( .A(n36069), .B(n36068), .CI(n36067), .CO(n34559), .S(n36494)
         );
  XNOR2_X1 U35834 ( .A(n36071), .B(n36070), .ZN(n36073) );
  XNOR2_X1 U35835 ( .A(n36073), .B(n36072), .ZN(n36493) );
  XNOR2_X1 U35836 ( .A(n36075), .B(n36074), .ZN(n36077) );
  XNOR2_X1 U35837 ( .A(n36077), .B(n36076), .ZN(n36768) );
  XNOR2_X1 U35838 ( .A(n36079), .B(n36078), .ZN(n36081) );
  XNOR2_X1 U35839 ( .A(n36081), .B(n36080), .ZN(n36767) );
  FA_X1 U35840 ( .A(n36084), .B(n36083), .CI(n36082), .CO(n36064), .S(n36547)
         );
  FA_X1 U35841 ( .A(n36087), .B(n36086), .CI(n36085), .CO(n34636), .S(n36599)
         );
  FA_X1 U35842 ( .A(n36090), .B(n36089), .CI(n36088), .CO(n34602), .S(n36598)
         );
  FA_X1 U35843 ( .A(n36093), .B(n36092), .CI(n36091), .CO(n34575), .S(n36597)
         );
  FA_X1 U35844 ( .A(n36096), .B(n36095), .CI(n36094), .CO(n36139), .S(n36577)
         );
  FA_X1 U35845 ( .A(n36099), .B(n36098), .CI(1'b0), .CO(n36137), .S(n36576) );
  FA_X1 U35846 ( .A(n36109), .B(n36108), .CI(n36107), .CO(n36127), .S(n36549)
         );
  NAND2_X1 U35847 ( .A1(n36114), .A2(n36113), .ZN(n36579) );
  OR2_X1 U35848 ( .A1(n36313), .A2(n3699), .ZN(n36115) );
  NAND2_X1 U35849 ( .A1(n36196), .A2(n36115), .ZN(n36578) );
  FA_X1 U35850 ( .A(n36118), .B(n36117), .CI(n36116), .CO(n36109), .S(n36573)
         );
  OAI22_X1 U35851 ( .A1(n36119), .A2(n3582), .B1(n36199), .B2(n36315), .ZN(
        n36586) );
  NAND2_X1 U35852 ( .A1(n36122), .A2(\fmem_data[7][1] ), .ZN(n36123) );
  NAND2_X1 U35853 ( .A1(n36218), .A2(n36123), .ZN(n36584) );
  FA_X1 U35854 ( .A(n36126), .B(n36125), .CI(n36124), .CO(n36072), .S(n36611)
         );
  FA_X1 U35855 ( .A(n36129), .B(n36128), .CI(n36127), .CO(n36124), .S(n36591)
         );
  FA_X1 U35856 ( .A(n36132), .B(n36131), .CI(n36130), .CO(n36164), .S(n36590)
         );
  FA_X1 U35857 ( .A(n36135), .B(n36134), .CI(n36133), .CO(n36175), .S(n36783)
         );
  XNOR2_X1 U35858 ( .A(n36137), .B(n36136), .ZN(n36138) );
  XNOR2_X1 U35859 ( .A(n36139), .B(n36138), .ZN(n36782) );
  FA_X1 U35860 ( .A(n36142), .B(n36141), .CI(n36140), .CO(n36192), .S(n36781)
         );
  OAI21_X1 U35861 ( .B1(n36612), .B2(n36611), .A(n36610), .ZN(n36144) );
  NAND2_X1 U35862 ( .A1(n36612), .A2(n36611), .ZN(n36143) );
  NAND2_X1 U35863 ( .A1(n36144), .A2(n36143), .ZN(n36766) );
  OAI21_X1 U35864 ( .B1(n36814), .B2(n36813), .A(n36815), .ZN(n36146) );
  NAND2_X1 U35865 ( .A1(n36814), .A2(n36813), .ZN(n36145) );
  NAND2_X1 U35866 ( .A1(n36146), .A2(n36145), .ZN(n36763) );
  OAI21_X1 U35867 ( .B1(n36757), .B2(n36755), .A(n36756), .ZN(n36148) );
  NAND2_X1 U35868 ( .A1(n36755), .A2(n36757), .ZN(n36147) );
  NAND2_X1 U35869 ( .A1(n36148), .A2(n36147), .ZN(n37122) );
  XNOR2_X1 U35870 ( .A(n36150), .B(n36149), .ZN(n36152) );
  XNOR2_X1 U35871 ( .A(n36152), .B(n36151), .ZN(n36752) );
  XNOR2_X1 U35872 ( .A(n36154), .B(n36153), .ZN(n36156) );
  XNOR2_X1 U35873 ( .A(n36156), .B(n36155), .ZN(n36759) );
  FA_X1 U35874 ( .A(n36159), .B(n36158), .CI(n36157), .CO(n36150), .S(n36762)
         );
  FA_X1 U35875 ( .A(n36162), .B(n36161), .CI(n36160), .CO(n36079), .S(n36807)
         );
  XNOR2_X1 U35876 ( .A(n36164), .B(n36163), .ZN(n36166) );
  XNOR2_X1 U35877 ( .A(n36166), .B(n36165), .ZN(n36806) );
  FA_X1 U35878 ( .A(n36169), .B(n36168), .CI(n36167), .CO(n36160), .S(n36773)
         );
  XNOR2_X1 U35879 ( .A(n36171), .B(n36170), .ZN(n36173) );
  XNOR2_X1 U35880 ( .A(n36173), .B(n36172), .ZN(n36775) );
  FA_X1 U35881 ( .A(n36182), .B(n36181), .CI(n36180), .CO(n36268), .S(n36769)
         );
  FA_X1 U35882 ( .A(n36185), .B(n36184), .CI(n36183), .CO(n36180), .S(n36810)
         );
  XNOR2_X1 U35883 ( .A(n36187), .B(n36186), .ZN(n36189) );
  FA_X1 U35884 ( .A(n36192), .B(n36191), .CI(n36190), .CO(n36188), .S(n36804)
         );
  FA_X1 U35885 ( .A(n36195), .B(n36194), .CI(n36193), .CO(n36174), .S(n36777)
         );
  OAI22_X1 U35886 ( .A1(n36197), .A2(n3577), .B1(n36196), .B2(n36313), .ZN(
        n36799) );
  NAND2_X1 U35887 ( .A1(n36199), .A2(n36198), .ZN(n36798) );
  INV_X1 U35888 ( .A(n36201), .ZN(n36202) );
  XNOR2_X1 U35889 ( .A(n36203), .B(n36202), .ZN(n36721) );
  XNOR2_X1 U35890 ( .A(n36205), .B(n36204), .ZN(n36207) );
  XNOR2_X1 U35891 ( .A(n36207), .B(n36206), .ZN(n36787) );
  OR2_X1 U35892 ( .A1(n36316), .A2(n3740), .ZN(n36208) );
  NAND2_X1 U35893 ( .A1(n36240), .A2(n36208), .ZN(n36796) );
  INV_X1 U35894 ( .A(n36314), .ZN(n36210) );
  OAI21_X1 U35895 ( .B1(n36789), .B2(n36787), .A(n36788), .ZN(n36213) );
  NAND2_X1 U35896 ( .A1(n36213), .A2(n36212), .ZN(n36778) );
  NOR2_X1 U35897 ( .A1(n36777), .A2(n36778), .ZN(n36232) );
  NAND2_X1 U35898 ( .A1(n36226), .A2(n36214), .ZN(n36691) );
  NAND2_X1 U35899 ( .A1(n36216), .A2(n36215), .ZN(n36690) );
  NAND2_X1 U35900 ( .A1(n36223), .A2(n36217), .ZN(n36689) );
  OAI22_X1 U35901 ( .A1(n36219), .A2(n3581), .B1(n36218), .B2(n36311), .ZN(
        n36793) );
  NAND2_X1 U35902 ( .A1(n36221), .A2(n36220), .ZN(n36792) );
  OR2_X1 U35903 ( .A1(n3116), .A2(n3735), .ZN(n36224) );
  NAND2_X1 U35904 ( .A1(n36241), .A2(n36224), .ZN(n36694) );
  INV_X1 U35905 ( .A(n36779), .ZN(n36231) );
  OAI21_X1 U35906 ( .B1(n36232), .B2(n36231), .A(n36230), .ZN(n36803) );
  FA_X1 U35907 ( .A(n36235), .B(n36234), .CI(n36233), .CO(n36190), .S(n36685)
         );
  FA_X1 U35908 ( .A(n36238), .B(n36237), .CI(n36236), .CO(n36193), .S(n36695)
         );
  OAI22_X1 U35909 ( .A1(n36316), .A2(n36240), .B1(n36239), .B2(n3482), .ZN(
        n36688) );
  OAI22_X1 U35910 ( .A1(n36242), .A2(n3662), .B1(n3116), .B2(n36241), .ZN(
        n36687) );
  OAI21_X1 U35911 ( .B1(n36695), .B2(n36696), .A(n36697), .ZN(n36251) );
  NAND2_X1 U35912 ( .A1(n36251), .A2(n36250), .ZN(n36684) );
  XOR2_X1 U35913 ( .A(n36254), .B(n36253), .Z(n36255) );
  XOR2_X1 U35914 ( .A(n36252), .B(n36255), .Z(n36701) );
  FA_X1 U35915 ( .A(n36258), .B(n36257), .CI(n36256), .CO(n36133), .S(n36700)
         );
  XNOR2_X1 U35916 ( .A(n36260), .B(n36259), .ZN(n36262) );
  XNOR2_X1 U35917 ( .A(n36262), .B(n36261), .ZN(n36699) );
  OAI21_X1 U35918 ( .B1(n36770), .B2(n36769), .A(n36771), .ZN(n36264) );
  NAND2_X1 U35919 ( .A1(n36264), .A2(n36263), .ZN(n36819) );
  FA_X1 U35920 ( .A(n36267), .B(n36266), .CI(n36265), .CO(n36154), .S(n36817)
         );
  FA_X1 U35921 ( .A(n36270), .B(n36269), .CI(n36268), .CO(n36155), .S(n36818)
         );
  OAI21_X1 U35922 ( .B1(n36819), .B2(n36817), .A(n36818), .ZN(n36272) );
  NAND2_X1 U35923 ( .A1(n36819), .A2(n36817), .ZN(n36271) );
  NAND2_X1 U35924 ( .A1(n36272), .A2(n36271), .ZN(n36760) );
  OAI21_X1 U35925 ( .B1(n36759), .B2(n36762), .A(n36760), .ZN(n36274) );
  NAND2_X1 U35926 ( .A1(n36759), .A2(n36762), .ZN(n36273) );
  NAND2_X1 U35927 ( .A1(n36274), .A2(n36273), .ZN(n36751) );
  FA_X1 U35928 ( .A(n36277), .B(n36276), .CI(n36275), .CO(n36381), .S(n36673)
         );
  FA_X1 U35929 ( .A(n36280), .B(n36279), .CI(n36278), .CO(n36276), .S(n36740)
         );
  FA_X1 U35930 ( .A(n36283), .B(n36282), .CI(n36281), .CO(n36376), .S(n36741)
         );
  XNOR2_X1 U35931 ( .A(n36285), .B(n36284), .ZN(n36287) );
  XNOR2_X1 U35932 ( .A(n36287), .B(n36286), .ZN(n36675) );
  XNOR2_X1 U35933 ( .A(n36289), .B(n36288), .ZN(n36291) );
  FA_X1 U35934 ( .A(n36294), .B(n36293), .CI(n36292), .CO(n36410), .S(n36703)
         );
  FA_X1 U35935 ( .A(n36303), .B(n36302), .CI(n36301), .CO(n36355), .S(n36715)
         );
  XNOR2_X1 U35936 ( .A(n36305), .B(n36304), .ZN(n36307) );
  FA_X1 U35937 ( .A(n36310), .B(n36309), .CI(n36308), .CO(n36348), .S(n36728)
         );
  AND2_X1 U35938 ( .A1(n36313), .A2(\fmem_data[11][0] ), .ZN(n36724) );
  AND2_X1 U35939 ( .A1(n36316), .A2(\fmem_data[27][0] ), .ZN(n36860) );
  OAI21_X1 U35940 ( .B1(n36728), .B2(n36727), .A(n36729), .ZN(n36318) );
  NAND2_X1 U35941 ( .A1(n36318), .A2(n36317), .ZN(n36709) );
  FA_X1 U35942 ( .A(n36321), .B(n36320), .CI(n36319), .CO(n36285), .S(n36679)
         );
  FA_X1 U35943 ( .A(n36324), .B(n36323), .CI(n36322), .CO(n36476), .S(n36851)
         );
  FA_X1 U35944 ( .A(n36327), .B(n36326), .CI(n36325), .CO(n36477), .S(n36850)
         );
  FA_X1 U35945 ( .A(n36330), .B(n36329), .CI(n36328), .CO(n36473), .S(n36852)
         );
  OAI21_X1 U35946 ( .B1(n36851), .B2(n36850), .A(n36852), .ZN(n36332) );
  NAND2_X1 U35947 ( .A1(n36851), .A2(n36850), .ZN(n36331) );
  NAND2_X1 U35948 ( .A1(n36332), .A2(n36331), .ZN(n36849) );
  XNOR2_X1 U35949 ( .A(n36334), .B(n36333), .ZN(n36336) );
  XNOR2_X1 U35950 ( .A(n36336), .B(n36335), .ZN(n36848) );
  AND2_X1 U35951 ( .A1(n36337), .A2(\fmem_data[19][0] ), .ZN(n36859) );
  FA_X1 U35952 ( .A(n36342), .B(n36341), .CI(n36340), .CO(n36475), .S(n36855)
         );
  XNOR2_X1 U35953 ( .A(n36344), .B(n36343), .ZN(n36346) );
  XNOR2_X1 U35954 ( .A(n36346), .B(n36345), .ZN(n36854) );
  FA_X1 U35955 ( .A(n36349), .B(n36348), .CI(n36347), .CO(n36408), .S(n36714)
         );
  XNOR2_X1 U35956 ( .A(n36353), .B(n36352), .ZN(n36713) );
  FA_X1 U35957 ( .A(n36356), .B(n36355), .CI(n36354), .CO(n36404), .S(n36712)
         );
  XNOR2_X1 U35958 ( .A(n36358), .B(n36357), .ZN(n36360) );
  XNOR2_X1 U35959 ( .A(n36360), .B(n36359), .ZN(n36705) );
  OAI21_X1 U35960 ( .B1(n36680), .B2(n36679), .A(n36681), .ZN(n36365) );
  NAND2_X1 U35961 ( .A1(n36680), .A2(n36679), .ZN(n36364) );
  NAND2_X1 U35962 ( .A1(n36365), .A2(n36364), .ZN(n36678) );
  FA_X1 U35963 ( .A(n36368), .B(n36367), .CI(n36366), .CO(n36278), .S(n36676)
         );
  OAI21_X1 U35964 ( .B1(n36675), .B2(n36678), .A(n36676), .ZN(n36370) );
  NAND2_X1 U35965 ( .A1(n36675), .A2(n36678), .ZN(n36369) );
  NAND2_X1 U35966 ( .A1(n36370), .A2(n36369), .ZN(n36743) );
  OAI21_X1 U35967 ( .B1(n36740), .B2(n36741), .A(n36743), .ZN(n36372) );
  NAND2_X1 U35968 ( .A1(n36740), .A2(n36741), .ZN(n36371) );
  NAND2_X1 U35969 ( .A1(n36372), .A2(n36371), .ZN(n36671) );
  XNOR2_X1 U35970 ( .A(n36374), .B(n36373), .ZN(n36375) );
  OAI21_X1 U35971 ( .B1(n36673), .B2(n36671), .A(n36672), .ZN(n36378) );
  NAND2_X1 U35972 ( .A1(n36673), .A2(n36671), .ZN(n36377) );
  NAND2_X1 U35973 ( .A1(n36378), .A2(n36377), .ZN(n36664) );
  XNOR2_X1 U35974 ( .A(n36380), .B(n36379), .ZN(n36382) );
  XNOR2_X1 U35975 ( .A(n36382), .B(n36381), .ZN(n36663) );
  XNOR2_X1 U35976 ( .A(n36384), .B(n36383), .ZN(n36386) );
  XNOR2_X1 U35977 ( .A(n36386), .B(n36385), .ZN(n36668) );
  XNOR2_X1 U35978 ( .A(n36388), .B(n36387), .ZN(n36390) );
  XNOR2_X1 U35979 ( .A(n36390), .B(n36389), .ZN(n36746) );
  XNOR2_X1 U35980 ( .A(n36392), .B(n36391), .ZN(n36394) );
  XNOR2_X1 U35981 ( .A(n36394), .B(n36393), .ZN(n36737) );
  FA_X1 U35982 ( .A(n36397), .B(n36396), .CI(n36395), .CO(n36420), .S(n36734)
         );
  XNOR2_X1 U35983 ( .A(n36399), .B(n36398), .ZN(n36401) );
  XNOR2_X1 U35984 ( .A(n36401), .B(n36400), .ZN(n36733) );
  XNOR2_X1 U35985 ( .A(n36403), .B(n36402), .ZN(n36405) );
  XNOR2_X1 U35986 ( .A(n36405), .B(n36404), .ZN(n36732) );
  FA_X1 U35987 ( .A(n36408), .B(n36407), .CI(n36406), .CO(n36414), .S(n36731)
         );
  XNOR2_X1 U35988 ( .A(n36410), .B(n36409), .ZN(n36412) );
  XNOR2_X1 U35989 ( .A(n36412), .B(n36411), .ZN(n36842) );
  XNOR2_X1 U35990 ( .A(n36414), .B(n36413), .ZN(n36416) );
  XNOR2_X1 U35991 ( .A(n36416), .B(n36415), .ZN(n36841) );
  OAI21_X1 U35992 ( .B1(n36737), .B2(n36734), .A(n36735), .ZN(n36418) );
  NAND2_X1 U35993 ( .A1(n36418), .A2(n36417), .ZN(n36745) );
  XNOR2_X1 U35994 ( .A(n36420), .B(n36419), .ZN(n36422) );
  XNOR2_X1 U35995 ( .A(n36422), .B(n36421), .ZN(n36744) );
  FA_X1 U35996 ( .A(n36425), .B(n36424), .CI(n36423), .CO(n36618), .S(n36669)
         );
  OAI21_X1 U35997 ( .B1(n36668), .B2(n36667), .A(n36669), .ZN(n36427) );
  NAND2_X1 U35998 ( .A1(n36668), .A2(n36667), .ZN(n36426) );
  NAND2_X1 U35999 ( .A1(n36427), .A2(n36426), .ZN(n36666) );
  OAI21_X1 U36000 ( .B1(n36664), .B2(n36663), .A(n36666), .ZN(n36429) );
  NAND2_X1 U36001 ( .A1(n36429), .A2(n36428), .ZN(n36753) );
  OAI21_X1 U36002 ( .B1(n36752), .B2(n36751), .A(n36753), .ZN(n36431) );
  NAND2_X1 U36003 ( .A1(n36751), .A2(n36752), .ZN(n36430) );
  NAND2_X1 U36004 ( .A1(n36431), .A2(n36430), .ZN(n37121) );
  OAI21_X1 U36005 ( .B1(n36447), .B2(n36446), .A(n36448), .ZN(n36433) );
  NAND2_X1 U36006 ( .A1(n36447), .A2(n36446), .ZN(n36432) );
  NAND2_X1 U36007 ( .A1(n36433), .A2(n36432), .ZN(n36656) );
  XNOR2_X1 U36008 ( .A(n36435), .B(n36434), .ZN(n36437) );
  XNOR2_X1 U36009 ( .A(n36437), .B(n36436), .ZN(n36655) );
  NAND2_X1 U36010 ( .A1(n3283), .A2(n36438), .ZN(n36443) );
  XNOR2_X1 U36011 ( .A(n36440), .B(n36439), .ZN(n36441) );
  XNOR2_X1 U36012 ( .A(n3122), .B(n36441), .ZN(n36657) );
  NAND2_X1 U36013 ( .A1(n36443), .A2(n36657), .ZN(n36445) );
  NAND2_X1 U36014 ( .A1(n36445), .A2(n36444), .ZN(n37161) );
  NOR2_X2 U36015 ( .A1(n37162), .A2(n37161), .ZN(n37254) );
  XNOR2_X1 U36016 ( .A(n36447), .B(n36446), .ZN(n36450) );
  XNOR2_X1 U36017 ( .A(n36450), .B(n36449), .ZN(n37130) );
  FA_X1 U36018 ( .A(n36453), .B(n36452), .CI(n36451), .CO(n36621), .S(n36831)
         );
  XNOR2_X1 U36019 ( .A(n36455), .B(n36454), .ZN(n36457) );
  XNOR2_X1 U36020 ( .A(n36457), .B(n36456), .ZN(n36834) );
  FA_X1 U36021 ( .A(n36460), .B(n36459), .CI(n36458), .CO(n36451), .S(n36833)
         );
  XNOR2_X1 U36022 ( .A(n36462), .B(n36461), .ZN(n36463) );
  XNOR2_X1 U36023 ( .A(n36464), .B(n36463), .ZN(n36837) );
  FA_X1 U36024 ( .A(n36467), .B(n36466), .CI(n36465), .CO(n36492), .S(n36840)
         );
  FA_X1 U36025 ( .A(n36470), .B(n36469), .CI(n36468), .CO(n36366), .S(n36839)
         );
  XNOR2_X1 U36026 ( .A(n36472), .B(n36471), .ZN(n36474) );
  XNOR2_X1 U36027 ( .A(n36474), .B(n36473), .ZN(n36868) );
  FA_X1 U36028 ( .A(n36477), .B(n36476), .CI(n36475), .CO(n36290), .S(n36867)
         );
  XNOR2_X1 U36029 ( .A(n36479), .B(n36478), .ZN(n36481) );
  XNOR2_X1 U36030 ( .A(n36481), .B(n36480), .ZN(n36866) );
  XNOR2_X1 U36031 ( .A(n36483), .B(n36482), .ZN(n36485) );
  XNOR2_X1 U36032 ( .A(n36485), .B(n36484), .ZN(n36845) );
  FA_X1 U36033 ( .A(n36488), .B(n36487), .CI(n36486), .CO(n36504), .S(n36844)
         );
  FA_X1 U36034 ( .A(n36495), .B(n36494), .CI(n36493), .CO(n36813), .S(n36879)
         );
  XNOR2_X1 U36035 ( .A(n36497), .B(n36496), .ZN(n36499) );
  XNOR2_X1 U36036 ( .A(n36499), .B(n36498), .ZN(n36876) );
  FA_X1 U36037 ( .A(n36502), .B(n36501), .CI(n36500), .CO(n36495), .S(n36874)
         );
  XNOR2_X1 U36038 ( .A(n36504), .B(n36503), .ZN(n36506) );
  FA_X1 U36039 ( .A(n36513), .B(n36512), .CI(n36511), .CO(n36607), .S(n36873)
         );
  FA_X1 U36040 ( .A(n36516), .B(n36515), .CI(n36514), .CO(n36508), .S(n36872)
         );
  FA_X1 U36041 ( .A(n36519), .B(n36518), .CI(n36517), .CO(n36555), .S(n36910)
         );
  FA_X1 U36042 ( .A(n36522), .B(n36521), .CI(n36520), .CO(n36518), .S(n36865)
         );
  AND2_X1 U36043 ( .A1(n3116), .A2(\fmem_data[23][0] ), .ZN(n36864) );
  FA_X1 U36044 ( .A(n36526), .B(n36525), .CI(n36524), .CO(n36532), .S(n36863)
         );
  FA_X1 U36045 ( .A(n36529), .B(n36528), .CI(n36527), .CO(n36554), .S(n36908)
         );
  FA_X1 U36046 ( .A(n36532), .B(n36531), .CI(n36530), .CO(n36480), .S(n36913)
         );
  FA_X1 U36047 ( .A(n36539), .B(n36538), .CI(n36537), .CO(n36540), .S(n36911)
         );
  FA_X1 U36048 ( .A(n36542), .B(n36541), .CI(n36540), .CO(n36513), .S(n36917)
         );
  OAI21_X1 U36049 ( .B1(n36876), .B2(n36874), .A(n36875), .ZN(n36544) );
  NAND2_X1 U36050 ( .A1(n36544), .A2(n36543), .ZN(n36878) );
  FA_X1 U36051 ( .A(n36547), .B(n36546), .CI(n36545), .CO(n36612), .S(n36947)
         );
  FA_X1 U36052 ( .A(n36550), .B(n36549), .CI(n36548), .CO(n36545), .S(n36924)
         );
  FA_X1 U36053 ( .A(n36553), .B(n36552), .CI(n36551), .CO(n36603), .S(n36922)
         );
  FA_X1 U36054 ( .A(n36556), .B(n36555), .CI(n36554), .CO(n36512), .S(n36921)
         );
  FA_X1 U36055 ( .A(n36559), .B(n36558), .CI(n36557), .CO(n36538), .S(n37071)
         );
  FA_X1 U36056 ( .A(n36562), .B(n36561), .CI(n36560), .CO(n36535), .S(n37070)
         );
  FA_X1 U36057 ( .A(n36565), .B(n36564), .CI(n36563), .CO(n36580), .S(n37069)
         );
  FA_X1 U36058 ( .A(n36568), .B(n36567), .CI(n36566), .CO(n36552), .S(n36915)
         );
  FA_X1 U36059 ( .A(n36571), .B(n36570), .CI(n36569), .CO(n36551), .S(n36914)
         );
  FA_X1 U36060 ( .A(n36574), .B(n36573), .CI(n36572), .CO(n36548), .S(n36960)
         );
  FA_X1 U36061 ( .A(n36577), .B(n36576), .CI(n36575), .CO(n36550), .S(n36959)
         );
  FA_X1 U36062 ( .A(n36580), .B(n36579), .CI(n36578), .CO(n36574), .S(n36954)
         );
  FA_X1 U36063 ( .A(n36583), .B(n36582), .CI(n36581), .CO(n36575), .S(n36953)
         );
  FA_X1 U36064 ( .A(n36586), .B(n36585), .CI(n36584), .CO(n36572), .S(n36952)
         );
  OAI21_X1 U36065 ( .B1(n36924), .B2(n36923), .A(n36925), .ZN(n36588) );
  NAND2_X1 U36066 ( .A1(n36588), .A2(n36587), .ZN(n36946) );
  FA_X1 U36067 ( .A(n36591), .B(n36590), .CI(n36589), .CO(n36610), .S(n36945)
         );
  OAI21_X1 U36068 ( .B1(n36947), .B2(n36946), .A(n36945), .ZN(n36593) );
  NAND2_X1 U36069 ( .A1(n36946), .A2(n36947), .ZN(n36592) );
  NAND2_X1 U36070 ( .A1(n36593), .A2(n36592), .ZN(n36898) );
  FA_X1 U36071 ( .A(n36596), .B(n36595), .CI(n36594), .CO(n36498), .S(n36901)
         );
  FA_X1 U36072 ( .A(n36599), .B(n36598), .CI(n36597), .CO(n36546), .S(n36907)
         );
  FA_X1 U36073 ( .A(n36602), .B(n36601), .CI(n36600), .CO(n36505), .S(n36906)
         );
  FA_X1 U36074 ( .A(n36605), .B(n36604), .CI(n36603), .CO(n36594), .S(n36905)
         );
  XNOR2_X1 U36075 ( .A(n36607), .B(n36606), .ZN(n36609) );
  XNOR2_X1 U36076 ( .A(n36609), .B(n36608), .ZN(n36899) );
  XNOR2_X1 U36077 ( .A(n36611), .B(n36610), .ZN(n36613) );
  OAI21_X1 U36078 ( .B1(n36879), .B2(n36878), .A(n36880), .ZN(n36615) );
  NAND2_X1 U36079 ( .A1(n36879), .A2(n36878), .ZN(n36614) );
  NAND2_X1 U36080 ( .A1(n36615), .A2(n36614), .ZN(n36829) );
  INV_X1 U36081 ( .A(n36750), .ZN(n36626) );
  XNOR2_X1 U36082 ( .A(n36621), .B(n36620), .ZN(n36623) );
  XNOR2_X1 U36083 ( .A(n36623), .B(n36622), .ZN(n36748) );
  NOR2_X1 U36084 ( .A1(n36747), .A2(n36748), .ZN(n36625) );
  NAND2_X1 U36085 ( .A1(n36747), .A2(n36748), .ZN(n36624) );
  OAI21_X1 U36086 ( .B1(n36626), .B2(n36625), .A(n36624), .ZN(n36660) );
  XNOR2_X1 U36087 ( .A(n36628), .B(n36627), .ZN(n36630) );
  XNOR2_X1 U36088 ( .A(n36630), .B(n36629), .ZN(n36659) );
  XNOR2_X1 U36089 ( .A(n36634), .B(n36633), .ZN(n36661) );
  OAI21_X1 U36090 ( .B1(n36660), .B2(n36659), .A(n36661), .ZN(n36636) );
  NAND2_X1 U36091 ( .A1(n36660), .A2(n36659), .ZN(n36635) );
  NAND2_X1 U36092 ( .A1(n36636), .A2(n36635), .ZN(n37115) );
  XNOR2_X1 U36093 ( .A(n36638), .B(n36637), .ZN(n36640) );
  XNOR2_X1 U36094 ( .A(n36640), .B(n36639), .ZN(n37114) );
  XNOR2_X1 U36095 ( .A(n36642), .B(n3284), .ZN(n36643) );
  XNOR2_X1 U36096 ( .A(n36644), .B(n36643), .ZN(n37116) );
  OAI21_X1 U36097 ( .B1(n37115), .B2(n37114), .A(n37116), .ZN(n36646) );
  NAND2_X1 U36098 ( .A1(n37115), .A2(n37114), .ZN(n36645) );
  NAND2_X1 U36099 ( .A1(n36646), .A2(n36645), .ZN(n37129) );
  INV_X1 U36100 ( .A(n37129), .ZN(n36651) );
  FA_X1 U36101 ( .A(n36649), .B(n36648), .CI(n36647), .CO(n36442), .S(n37128)
         );
  NAND2_X1 U36102 ( .A1(n36651), .A2(n36650), .ZN(n36652) );
  NAND2_X1 U36103 ( .A1(n37130), .A2(n36652), .ZN(n36654) );
  NAND2_X1 U36104 ( .A1(n37129), .A2(n37128), .ZN(n36653) );
  XNOR2_X1 U36105 ( .A(n36656), .B(n36655), .ZN(n36658) );
  XNOR2_X1 U36106 ( .A(n36658), .B(n36657), .ZN(n37159) );
  NOR2_X1 U36107 ( .A1(n37160), .A2(n37159), .ZN(n37187) );
  NOR2_X1 U36108 ( .A1(n37254), .A2(n37187), .ZN(n37206) );
  NAND2_X1 U36109 ( .A1(n37163), .A2(n37206), .ZN(n37158) );
  XNOR2_X1 U36110 ( .A(n36660), .B(n36659), .ZN(n36662) );
  XNOR2_X1 U36111 ( .A(n36668), .B(n36667), .ZN(n36670) );
  XNOR2_X1 U36112 ( .A(n36670), .B(n36669), .ZN(n36891) );
  XNOR2_X1 U36113 ( .A(n36676), .B(n36675), .ZN(n36677) );
  XNOR2_X1 U36114 ( .A(n36680), .B(n36679), .ZN(n36682) );
  XNOR2_X1 U36115 ( .A(n36682), .B(n36681), .ZN(n36989) );
  FA_X1 U36116 ( .A(n36685), .B(n36684), .CI(n36683), .CO(n36802), .S(n36970)
         );
  FA_X1 U36117 ( .A(n36688), .B(n36687), .CI(n36686), .CO(n36696), .S(n36957)
         );
  FA_X1 U36118 ( .A(n36691), .B(n36690), .CI(n36689), .CO(n36786), .S(n36956)
         );
  FA_X1 U36119 ( .A(n36694), .B(n36693), .CI(n36692), .CO(n36784), .S(n36955)
         );
  XNOR2_X1 U36120 ( .A(n36696), .B(n36695), .ZN(n36698) );
  XNOR2_X1 U36121 ( .A(n36698), .B(n36697), .ZN(n36975) );
  FA_X1 U36122 ( .A(n36701), .B(n36700), .CI(n36699), .CO(n36683), .S(n36974)
         );
  FA_X1 U36123 ( .A(n36704), .B(n36703), .CI(n36702), .CO(n36680), .S(n36968)
         );
  XNOR2_X1 U36124 ( .A(n36706), .B(n36705), .ZN(n36708) );
  XNOR2_X1 U36125 ( .A(n36708), .B(n36707), .ZN(n36983) );
  FA_X1 U36126 ( .A(n36711), .B(n36710), .CI(n36709), .CO(n36702), .S(n36973)
         );
  FA_X1 U36127 ( .A(n36714), .B(n36713), .CI(n36712), .CO(n36706), .S(n36972)
         );
  FA_X1 U36128 ( .A(n36717), .B(n36716), .CI(n36715), .CO(n36711), .S(n37013)
         );
  FA_X1 U36129 ( .A(n36720), .B(n36719), .CI(n36718), .CO(n36686), .S(n37068)
         );
  FA_X1 U36130 ( .A(n36723), .B(n36722), .CI(n36721), .CO(n36797), .S(n37067)
         );
  FA_X1 U36131 ( .A(n36726), .B(n36725), .CI(n36724), .CO(n36727), .S(n37066)
         );
  FA_X1 U36132 ( .A(n36733), .B(n36732), .CI(n36731), .CO(n36843), .S(n36981)
         );
  OAI21_X1 U36133 ( .B1(n36938), .B2(n36941), .A(n36939), .ZN(n36739) );
  NAND2_X1 U36134 ( .A1(n36739), .A2(n36738), .ZN(n36934) );
  FA_X1 U36135 ( .A(n36746), .B(n36745), .CI(n36744), .CO(n36667), .S(n36932)
         );
  XNOR2_X1 U36136 ( .A(n36748), .B(n36747), .ZN(n36749) );
  XNOR2_X1 U36137 ( .A(n36750), .B(n36749), .ZN(n36823) );
  XNOR2_X1 U36138 ( .A(n36752), .B(n36751), .ZN(n36754) );
  XNOR2_X1 U36139 ( .A(n36754), .B(n36753), .ZN(n37120) );
  XNOR2_X1 U36140 ( .A(n36756), .B(n36755), .ZN(n36758) );
  XNOR2_X1 U36141 ( .A(n36758), .B(n36757), .ZN(n37119) );
  XNOR2_X1 U36142 ( .A(n36760), .B(n36759), .ZN(n36761) );
  XNOR2_X1 U36143 ( .A(n36762), .B(n36761), .ZN(n36828) );
  FA_X1 U36144 ( .A(n36765), .B(n36764), .CI(n36763), .CO(n36756), .S(n36827)
         );
  FA_X1 U36145 ( .A(n36768), .B(n36767), .CI(n36766), .CO(n36815), .S(n36892)
         );
  XNOR2_X1 U36146 ( .A(n36770), .B(n36769), .ZN(n36772) );
  XNOR2_X1 U36147 ( .A(n36772), .B(n36771), .ZN(n36894) );
  XNOR2_X1 U36148 ( .A(n36774), .B(n36773), .ZN(n36776) );
  XNOR2_X1 U36149 ( .A(n36776), .B(n36775), .ZN(n36944) );
  XNOR2_X1 U36150 ( .A(n36778), .B(n36777), .ZN(n36780) );
  XNOR2_X1 U36151 ( .A(n36780), .B(n36779), .ZN(n36965) );
  FA_X1 U36152 ( .A(n36783), .B(n36782), .CI(n36781), .CO(n36589), .S(n36964)
         );
  FA_X1 U36153 ( .A(n36786), .B(n36785), .CI(n36784), .CO(n36779), .S(n36963)
         );
  XNOR2_X1 U36154 ( .A(n36788), .B(n36787), .ZN(n36790) );
  XNOR2_X1 U36155 ( .A(n36790), .B(n36789), .ZN(n36962) );
  FA_X1 U36156 ( .A(n36793), .B(n36792), .CI(n36791), .CO(n36785), .S(n36951)
         );
  FA_X1 U36157 ( .A(n36796), .B(n36795), .CI(n36794), .CO(n36788), .S(n36950)
         );
  FA_X1 U36158 ( .A(n36799), .B(n36798), .CI(n36797), .CO(n36789), .S(n36949)
         );
  OAI21_X1 U36159 ( .B1(n36965), .B2(n36964), .A(n36967), .ZN(n36801) );
  NAND2_X1 U36160 ( .A1(n36965), .A2(n36964), .ZN(n36800) );
  NAND2_X1 U36161 ( .A1(n36801), .A2(n36800), .ZN(n36943) );
  FA_X1 U36162 ( .A(n36804), .B(n36803), .CI(n36802), .CO(n36808), .S(n36942)
         );
  FA_X1 U36163 ( .A(n36807), .B(n36806), .CI(n36805), .CO(n36770), .S(n36930)
         );
  FA_X1 U36164 ( .A(n36810), .B(n36809), .CI(n36808), .CO(n36771), .S(n36929)
         );
  OAI21_X1 U36165 ( .B1(n36892), .B2(n36894), .A(n36893), .ZN(n36812) );
  NAND2_X1 U36166 ( .A1(n36892), .A2(n36894), .ZN(n36811) );
  NAND2_X1 U36167 ( .A1(n36812), .A2(n36811), .ZN(n36884) );
  XNOR2_X1 U36168 ( .A(n36818), .B(n36817), .ZN(n36820) );
  XNOR2_X1 U36169 ( .A(n36820), .B(n36819), .ZN(n36882) );
  OAI21_X1 U36170 ( .B1(n36884), .B2(n36883), .A(n36882), .ZN(n36821) );
  NAND2_X1 U36171 ( .A1(n36822), .A2(n36821), .ZN(n36826) );
  FA_X1 U36172 ( .A(n36825), .B(n36824), .CI(n36823), .CO(n37126), .S(n37104)
         );
  FA_X1 U36173 ( .A(n36828), .B(n36827), .CI(n36826), .CO(n37118), .S(n37103)
         );
  FA_X1 U36174 ( .A(n36831), .B(n36830), .CI(n36829), .CO(n36750), .S(n37036)
         );
  FA_X1 U36175 ( .A(n36834), .B(n36833), .CI(n36832), .CO(n36830), .S(n36937)
         );
  FA_X1 U36176 ( .A(n36837), .B(n36836), .CI(n36835), .CO(n36832), .S(n36998)
         );
  FA_X1 U36177 ( .A(n36840), .B(n36839), .CI(n36838), .CO(n36836), .S(n36992)
         );
  FA_X1 U36178 ( .A(n36843), .B(n36842), .CI(n36841), .CO(n36735), .S(n36991)
         );
  FA_X1 U36179 ( .A(n36846), .B(n36845), .CI(n36844), .CO(n36838), .S(n36986)
         );
  FA_X1 U36180 ( .A(n36849), .B(n36848), .CI(n36847), .CO(n36707), .S(n36977)
         );
  XNOR2_X1 U36181 ( .A(n36851), .B(n36850), .ZN(n36853) );
  XNOR2_X1 U36182 ( .A(n36853), .B(n36852), .ZN(n37010) );
  FA_X1 U36183 ( .A(n36856), .B(n36855), .CI(n36854), .CO(n36847), .S(n37009)
         );
  FA_X1 U36184 ( .A(n36859), .B(n36858), .CI(n36857), .CO(n36856), .S(n37074)
         );
  FA_X1 U36185 ( .A(n36862), .B(n36861), .CI(n36860), .CO(n36729), .S(n37073)
         );
  FA_X1 U36186 ( .A(n36865), .B(n36864), .CI(n36863), .CO(n36909), .S(n37072)
         );
  FA_X1 U36187 ( .A(n36868), .B(n36867), .CI(n36866), .CO(n36846), .S(n36978)
         );
  OAI21_X1 U36188 ( .B1(n36977), .B2(n36979), .A(n36978), .ZN(n36870) );
  NAND2_X1 U36189 ( .A1(n36870), .A2(n36869), .ZN(n36985) );
  FA_X1 U36190 ( .A(n36873), .B(n36872), .CI(n36871), .CO(n36902), .S(n36984)
         );
  XNOR2_X1 U36191 ( .A(n36875), .B(n36874), .ZN(n36877) );
  XNOR2_X1 U36192 ( .A(n36877), .B(n36876), .ZN(n36996) );
  XNOR2_X1 U36193 ( .A(n36879), .B(n36878), .ZN(n36881) );
  XNOR2_X1 U36194 ( .A(n36881), .B(n36880), .ZN(n36935) );
  XNOR2_X1 U36195 ( .A(n36883), .B(n36882), .ZN(n36885) );
  XNOR2_X1 U36196 ( .A(n36885), .B(n36884), .ZN(n37034) );
  NAND2_X1 U36197 ( .A1(n36888), .A2(n36887), .ZN(n37269) );
  NOR2_X1 U36198 ( .A1(n37270), .A2(n37269), .ZN(n37113) );
  FA_X1 U36199 ( .A(n36891), .B(n36890), .CI(n36889), .CO(n36824), .S(n37108)
         );
  FA_X1 U36200 ( .A(n36898), .B(n36897), .CI(n36896), .CO(n36880), .S(n36995)
         );
  FA_X1 U36201 ( .A(n36901), .B(n36900), .CI(n36899), .CO(n36897), .S(n37004)
         );
  FA_X1 U36202 ( .A(n36904), .B(n36903), .CI(n36902), .CO(n36875), .S(n37003)
         );
  FA_X1 U36203 ( .A(n36907), .B(n36906), .CI(n36905), .CO(n36900), .S(n37020)
         );
  FA_X1 U36204 ( .A(n36910), .B(n36909), .CI(n36908), .CO(n36919), .S(n37016)
         );
  FA_X1 U36205 ( .A(n36913), .B(n36912), .CI(n36911), .CO(n36918), .S(n37015)
         );
  FA_X1 U36206 ( .A(n36916), .B(n36915), .CI(n36914), .CO(n36920), .S(n37014)
         );
  FA_X1 U36207 ( .A(n36919), .B(n36918), .CI(n36917), .CO(n36871), .S(n37006)
         );
  FA_X1 U36208 ( .A(n36922), .B(n36921), .CI(n36920), .CO(n36923), .S(n37005)
         );
  XNOR2_X1 U36209 ( .A(n36924), .B(n36923), .ZN(n36926) );
  XNOR2_X1 U36210 ( .A(n36926), .B(n36925), .ZN(n37022) );
  OAI21_X1 U36211 ( .B1(n37020), .B2(n37021), .A(n37022), .ZN(n36928) );
  NAND2_X1 U36212 ( .A1(n37021), .A2(n37020), .ZN(n36927) );
  NAND2_X1 U36213 ( .A1(n36928), .A2(n36927), .ZN(n37002) );
  FA_X1 U36214 ( .A(n36931), .B(n36930), .CI(n36929), .CO(n36893), .S(n36993)
         );
  FA_X1 U36215 ( .A(n36934), .B(n36933), .CI(n36932), .CO(n36889), .S(n37041)
         );
  XNOR2_X1 U36216 ( .A(n37108), .B(n37107), .ZN(n37033) );
  FA_X1 U36217 ( .A(n36937), .B(n36936), .CI(n36935), .CO(n37035), .S(n37038)
         );
  FA_X1 U36218 ( .A(n36944), .B(n36943), .CI(n36942), .CO(n36931), .S(n37001)
         );
  XNOR2_X1 U36219 ( .A(n36946), .B(n36945), .ZN(n36948) );
  FA_X1 U36220 ( .A(n36951), .B(n36950), .CI(n36949), .CO(n36961), .S(n37065)
         );
  FA_X1 U36221 ( .A(n36954), .B(n36953), .CI(n36952), .CO(n36958), .S(n37064)
         );
  FA_X1 U36222 ( .A(n36957), .B(n36956), .CI(n36955), .CO(n36976), .S(n37063)
         );
  FA_X1 U36223 ( .A(n36960), .B(n36959), .CI(n36958), .CO(n36925), .S(n37018)
         );
  FA_X1 U36224 ( .A(n36963), .B(n36962), .CI(n36961), .CO(n36967), .S(n37017)
         );
  XNOR2_X1 U36225 ( .A(n36965), .B(n36964), .ZN(n36966) );
  FA_X1 U36226 ( .A(n36970), .B(n36969), .CI(n36968), .CO(n36988), .S(n37024)
         );
  FA_X1 U36227 ( .A(n36973), .B(n36972), .CI(n36971), .CO(n36982), .S(n37062)
         );
  FA_X1 U36228 ( .A(n36976), .B(n36975), .CI(n36974), .CO(n36969), .S(n37061)
         );
  FA_X1 U36229 ( .A(n36983), .B(n36982), .CI(n36981), .CO(n36987), .S(n37055)
         );
  FA_X1 U36230 ( .A(n36986), .B(n36985), .CI(n36984), .CO(n36990), .S(n37054)
         );
  FA_X1 U36231 ( .A(n36989), .B(n36988), .CI(n36987), .CO(n36941), .S(n37089)
         );
  FA_X1 U36232 ( .A(n36992), .B(n36991), .CI(n36990), .CO(n36997), .S(n37088)
         );
  FA_X1 U36233 ( .A(n36995), .B(n36994), .CI(n36993), .CO(n37042), .S(n37045)
         );
  FA_X1 U36234 ( .A(n36998), .B(n36997), .CI(n36996), .CO(n36936), .S(n37044)
         );
  FA_X1 U36235 ( .A(n37001), .B(n37000), .CI(n36999), .CO(n37049), .S(n37086)
         );
  FA_X1 U36236 ( .A(n37004), .B(n37003), .CI(n37002), .CO(n36994), .S(n37084)
         );
  FA_X1 U36237 ( .A(n37007), .B(n37006), .CI(n37005), .CO(n37021), .S(n37059)
         );
  FA_X1 U36238 ( .A(n37010), .B(n37009), .CI(n37008), .CO(n36979), .S(n37077)
         );
  FA_X1 U36239 ( .A(n37013), .B(n37012), .CI(n37011), .CO(n36971), .S(n37076)
         );
  FA_X1 U36240 ( .A(n37016), .B(n37015), .CI(n37014), .CO(n37007), .S(n37075)
         );
  FA_X1 U36241 ( .A(n37019), .B(n37018), .CI(n37017), .CO(n37026), .S(n37057)
         );
  FA_X1 U36242 ( .A(n37026), .B(n37025), .CI(n37024), .CO(n36999), .S(n37051)
         );
  OAI21_X1 U36243 ( .B1(n37086), .B2(n37084), .A(n37085), .ZN(n37028) );
  NAND2_X1 U36244 ( .A1(n37028), .A2(n37027), .ZN(n37046) );
  OAI21_X1 U36245 ( .B1(n37045), .B2(n37044), .A(n37046), .ZN(n37030) );
  NAND2_X1 U36246 ( .A1(n37045), .A2(n37044), .ZN(n37029) );
  NAND2_X1 U36247 ( .A1(n37030), .A2(n37029), .ZN(n37039) );
  OAI21_X1 U36248 ( .B1(n37038), .B2(n37037), .A(n37039), .ZN(n37032) );
  NAND2_X1 U36249 ( .A1(n37038), .A2(n37037), .ZN(n37031) );
  NAND2_X1 U36250 ( .A1(n37032), .A2(n37031), .ZN(n37106) );
  XNOR2_X1 U36251 ( .A(n37033), .B(n37106), .ZN(n37101) );
  FA_X1 U36252 ( .A(n37036), .B(n37035), .CI(n37034), .CO(n37102), .S(n37100)
         );
  NOR2_X1 U36253 ( .A1(n37101), .A2(n37100), .ZN(n37280) );
  XNOR2_X1 U36254 ( .A(n37038), .B(n37037), .ZN(n37040) );
  XNOR2_X1 U36255 ( .A(n37040), .B(n37039), .ZN(n37099) );
  FA_X1 U36256 ( .A(n37043), .B(n37042), .CI(n37041), .CO(n37107), .S(n37098)
         );
  XNOR2_X1 U36257 ( .A(n37045), .B(n37044), .ZN(n37047) );
  XNOR2_X1 U36258 ( .A(n37047), .B(n37046), .ZN(n37096) );
  FA_X1 U36259 ( .A(n37050), .B(n37049), .CI(n37048), .CO(n37037), .S(n37095)
         );
  NAND2_X1 U36260 ( .A1(n37096), .A2(n37095), .ZN(n37290) );
  FA_X1 U36261 ( .A(n37053), .B(n37052), .CI(n37051), .CO(n37085), .S(n37083)
         );
  FA_X1 U36262 ( .A(n37056), .B(n37055), .CI(n37054), .CO(n37090), .S(n37082)
         );
  FA_X1 U36263 ( .A(n37059), .B(n37058), .CI(n37057), .CO(n37053), .S(n37079)
         );
  FA_X1 U36264 ( .A(n37062), .B(n37061), .CI(n37060), .CO(n37056), .S(n37078)
         );
  FA_X1 U36265 ( .A(n37065), .B(n37064), .CI(n37063), .CO(n37019), .S(n37310)
         );
  FA_X1 U36266 ( .A(n37068), .B(n37067), .CI(n37066), .CO(n37012), .S(n37313)
         );
  FA_X1 U36267 ( .A(n37071), .B(n37070), .CI(n37069), .CO(n36916), .S(n37312)
         );
  FA_X1 U36268 ( .A(n37074), .B(n37073), .CI(n37072), .CO(n37008), .S(n37311)
         );
  FA_X1 U36269 ( .A(n37077), .B(n37076), .CI(n37075), .CO(n37058), .S(n37308)
         );
  INV_X1 U36270 ( .A(n37306), .ZN(n37080) );
  XNOR2_X1 U36271 ( .A(n37085), .B(n37084), .ZN(n37087) );
  XNOR2_X1 U36272 ( .A(n37087), .B(n37086), .ZN(n37092) );
  FA_X1 U36273 ( .A(n37090), .B(n37089), .CI(n37088), .CO(n37048), .S(n37091)
         );
  NAND2_X1 U36274 ( .A1(n37092), .A2(n37091), .ZN(n37294) );
  INV_X1 U36275 ( .A(n37294), .ZN(n37093) );
  AOI21_X1 U36276 ( .B1(n37296), .B2(n37295), .A(n37093), .ZN(n37094) );
  INV_X1 U36277 ( .A(n37094), .ZN(n37292) );
  NAND2_X1 U36278 ( .A1(n37292), .A2(n37291), .ZN(n37097) );
  NAND2_X1 U36279 ( .A1(n37290), .A2(n37097), .ZN(n37287) );
  AOI21_X1 U36280 ( .B1(n3708), .B2(n37287), .A(n37285), .ZN(n37284) );
  OAI21_X1 U36281 ( .B1(n37280), .B2(n37284), .A(n37281), .ZN(n37279) );
  XNOR2_X1 U36282 ( .A(n37103), .B(n37102), .ZN(n37105) );
  XNOR2_X1 U36283 ( .A(n37105), .B(n37104), .ZN(n37112) );
  AND2_X1 U36284 ( .A1(n37112), .A2(n37111), .ZN(n37275) );
  AOI21_X1 U36285 ( .B1(n37279), .B2(n37276), .A(n37275), .ZN(n37274) );
  OAI21_X1 U36286 ( .B1(n37113), .B2(n37274), .A(n37271), .ZN(n37258) );
  XNOR2_X1 U36287 ( .A(n37115), .B(n37114), .ZN(n37117) );
  XNOR2_X1 U36288 ( .A(n37117), .B(n37116), .ZN(n37133) );
  FA_X1 U36289 ( .A(n37120), .B(n37119), .CI(n37118), .CO(n37135), .S(n37125)
         );
  FA_X1 U36290 ( .A(n37123), .B(n37122), .CI(n37121), .CO(n36448), .S(n37134)
         );
  XNOR2_X1 U36291 ( .A(n37135), .B(n37134), .ZN(n37124) );
  XNOR2_X1 U36292 ( .A(n37133), .B(n37124), .ZN(n37139) );
  FA_X1 U36293 ( .A(n37127), .B(n37126), .CI(n37125), .CO(n37138), .S(n37270)
         );
  XNOR2_X1 U36294 ( .A(n37129), .B(n37128), .ZN(n37131) );
  XNOR2_X1 U36295 ( .A(n37131), .B(n37130), .ZN(n37140) );
  OR2_X1 U36296 ( .A1(n37135), .A2(n37134), .ZN(n37132) );
  NAND2_X1 U36297 ( .A1(n37133), .A2(n37132), .ZN(n37137) );
  NAND2_X1 U36298 ( .A1(n37135), .A2(n37134), .ZN(n37136) );
  NAND2_X1 U36299 ( .A1(n37137), .A2(n37136), .ZN(n37141) );
  NOR2_X1 U36300 ( .A1(n37264), .A2(n3435), .ZN(n37143) );
  NAND2_X1 U36301 ( .A1(n37139), .A2(n37138), .ZN(n37265) );
  NAND2_X1 U36302 ( .A1(n37140), .A2(n37141), .ZN(n37260) );
  OAI21_X1 U36303 ( .B1(n37259), .B2(n37265), .A(n37260), .ZN(n37142) );
  AOI21_X1 U36304 ( .B1(n37258), .B2(n37143), .A(n37142), .ZN(n37186) );
  OR2_X1 U36305 ( .A1(n37146), .A2(n37234), .ZN(n37156) );
  INV_X1 U36306 ( .A(n37238), .ZN(n37207) );
  AOI21_X1 U36307 ( .B1(n37154), .B2(n37207), .A(n37153), .ZN(n37155) );
  AND2_X1 U36308 ( .A1(n37156), .A2(n37155), .ZN(n37157) );
  OAI21_X1 U36309 ( .B1(n37158), .B2(n37186), .A(n37157), .ZN(n37244) );
  NAND2_X1 U36310 ( .A1(n37160), .A2(n37159), .ZN(n37250) );
  NAND2_X1 U36311 ( .A1(n37162), .A2(n37161), .ZN(n37255) );
  OAI21_X2 U36312 ( .B1(n37254), .B2(n37250), .A(n37255), .ZN(n37233) );
  NAND2_X1 U36313 ( .A1(n3273), .A2(n37233), .ZN(n37242) );
  INV_X1 U36314 ( .A(n37242), .ZN(n37164) );
  FA_X1 U36315 ( .A(n37167), .B(n37166), .CI(n37165), .CO(n37181), .S(n37151)
         );
  FA_X1 U36316 ( .A(n37170), .B(n37169), .CI(n37168), .CO(n37179), .S(n37176)
         );
  FA_X1 U36317 ( .A(n37173), .B(n37172), .CI(n37171), .CO(n37182), .S(n37170)
         );
  FA_X1 U36318 ( .A(n37176), .B(n37175), .CI(n37174), .CO(n37177), .S(n37167)
         );
  FA_X1 U36319 ( .A(n37179), .B(n37178), .CI(n37177), .CO(n37183), .S(n37180)
         );
  AOI21_X1 U36320 ( .B1(n37204), .B2(n37185), .A(n37184), .ZN(m_data_out_y[20]) );
  INV_X1 U36321 ( .A(n37186), .ZN(n37253) );
  XNOR2_X1 U36322 ( .A(n37253), .B(n37188), .ZN(m_data_out_y[12]) );
  NAND2_X1 U36323 ( .A1(n39051), .A2(n39001), .ZN(n37195) );
  INV_X1 U36324 ( .A(n37195), .ZN(n37189) );
  NAND2_X1 U36325 ( .A1(n37189), .A2(conv_pre_start), .ZN(n37314) );
  NAND2_X1 U36326 ( .A1(m_valid_y), .A2(m_ready_y), .ZN(n37194) );
  NAND4_X1 U36327 ( .A1(n37192), .A2(n37191), .A3(load_xaddr_val[6]), .A4(
        n37190), .ZN(n37196) );
  NOR3_X1 U36328 ( .A1(n37314), .A2(n37194), .A3(n37196), .ZN(n37193) );
  NOR2_X1 U36329 ( .A1(n37193), .A2(reset), .ZN(n37669) );
  INV_X1 U36330 ( .A(n37194), .ZN(n37197) );
  NOR2_X1 U36331 ( .A1(reset), .A2(n37195), .ZN(N229) );
  AND2_X1 U36332 ( .A1(conv_pre_start), .A2(N229), .ZN(
        \ctrl_conv_output_inst/N7 ) );
  NAND4_X1 U36333 ( .A1(n37197), .A2(\ctrl_conv_output_inst/N7 ), .A3(
        \ctrl_conv_output_inst/conv_start_reg ), .A4(n37196), .ZN(n38994) );
  NAND2_X1 U36334 ( .A1(n37669), .A2(n38994), .ZN(n38995) );
  OAI22_X1 U36335 ( .A1(n37199), .A2(n38995), .B1(n38994), .B2(n37198), .ZN(
        n37200) );
  INV_X1 U36336 ( .A(n37200), .ZN(n38996) );
  AOI21_X1 U36337 ( .B1(n37253), .B2(n37206), .A(n37233), .ZN(n37201) );
  XNOR2_X1 U36338 ( .A(n37201), .B(n4007), .ZN(m_data_out_y[14]) );
  XNOR2_X1 U36339 ( .A(n37204), .B(n37203), .ZN(m_data_out_y[18]) );
  NAND2_X1 U36340 ( .A1(n37205), .A2(n37239), .ZN(n37208) );
  INV_X1 U36341 ( .A(n37206), .ZN(n37231) );
  NOR2_X1 U36342 ( .A1(n37208), .A2(n37231), .ZN(n37213) );
  INV_X1 U36343 ( .A(n37234), .ZN(n37221) );
  AOI21_X1 U36344 ( .B1(n37239), .B2(n37221), .A(n37207), .ZN(n37211) );
  NAND2_X1 U36345 ( .A1(n37209), .A2(n37233), .ZN(n37210) );
  NAND2_X1 U36346 ( .A1(n37210), .A2(n37211), .ZN(n37212) );
  AOI21_X1 U36347 ( .B1(n37213), .B2(n37253), .A(n37212), .ZN(n37215) );
  XNOR2_X1 U36348 ( .A(n37215), .B(n37214), .ZN(m_data_out_y[16]) );
  INV_X1 U36349 ( .A(n37239), .ZN(n37217) );
  NOR2_X1 U36350 ( .A1(n37217), .A2(n37219), .ZN(n37222) );
  NAND2_X1 U36351 ( .A1(n37205), .A2(n37222), .ZN(n37225) );
  NOR2_X1 U36352 ( .A1(n37231), .A2(n37225), .ZN(n37227) );
  INV_X1 U36353 ( .A(n37233), .ZN(n37224) );
  OAI21_X1 U36354 ( .B1(n37225), .B2(n37224), .A(n37223), .ZN(n37226) );
  AOI21_X1 U36355 ( .B1(n37253), .B2(n37227), .A(n37226), .ZN(n37230) );
  XNOR2_X1 U36356 ( .A(n37230), .B(n4013), .ZN(m_data_out_y[17]) );
  NAND2_X1 U36357 ( .A1(n37233), .A2(n37205), .ZN(n37235) );
  NAND2_X1 U36358 ( .A1(n37235), .A2(n37234), .ZN(n37236) );
  AOI21_X1 U36359 ( .B1(n37237), .B2(n37253), .A(n37236), .ZN(n37240) );
  XNOR2_X1 U36360 ( .A(n37240), .B(n4000), .ZN(m_data_out_y[15]) );
  NAND2_X1 U36361 ( .A1(n37242), .A2(n37241), .ZN(n37245) );
  OAI21_X1 U36362 ( .B1(n37245), .B2(n37244), .A(n37243), .ZN(n37249) );
  XNOR2_X1 U36363 ( .A(n37249), .B(n4014), .ZN(m_data_out_y[19]) );
  AOI21_X1 U36364 ( .B1(n37253), .B2(n37252), .A(n37251), .ZN(n37257) );
  XNOR2_X1 U36365 ( .A(n37257), .B(n4011), .ZN(m_data_out_y[13]) );
  INV_X1 U36366 ( .A(n37258), .ZN(n37267) );
  INV_X1 U36367 ( .A(n3435), .ZN(n37261) );
  NAND2_X1 U36368 ( .A1(n37261), .A2(n37260), .ZN(n37262) );
  XNOR2_X1 U36369 ( .A(n37263), .B(n37262), .ZN(m_data_out_y[11]) );
  NAND2_X1 U36370 ( .A1(n37266), .A2(n37265), .ZN(n37268) );
  XOR2_X1 U36371 ( .A(n37268), .B(n37267), .Z(m_data_out_y[10]) );
  OR2_X1 U36372 ( .A1(n37270), .A2(n37269), .ZN(n37272) );
  NAND2_X1 U36373 ( .A1(n37272), .A2(n37271), .ZN(n37273) );
  XOR2_X1 U36374 ( .A(n37274), .B(n37273), .Z(m_data_out_y[9]) );
  NAND2_X1 U36375 ( .A1(n37277), .A2(n37276), .ZN(n37278) );
  XNOR2_X1 U36376 ( .A(n37279), .B(n37278), .ZN(m_data_out_y[8]) );
  INV_X1 U36377 ( .A(n37280), .ZN(n37282) );
  NAND2_X1 U36378 ( .A1(n37282), .A2(n37281), .ZN(n37283) );
  XOR2_X1 U36379 ( .A(n37284), .B(n37283), .Z(m_data_out_y[7]) );
  NAND2_X1 U36380 ( .A1(n3708), .A2(n37286), .ZN(n37289) );
  INV_X1 U36381 ( .A(n37287), .ZN(n37288) );
  XOR2_X1 U36382 ( .A(n37289), .B(n37288), .Z(m_data_out_y[6]) );
  NAND2_X1 U36383 ( .A1(n37291), .A2(n37290), .ZN(n37293) );
  XNOR2_X1 U36384 ( .A(n37293), .B(n37292), .ZN(m_data_out_y[5]) );
  NAND2_X1 U36385 ( .A1(n37295), .A2(n37294), .ZN(n37297) );
  XNOR2_X1 U36386 ( .A(n37297), .B(n37296), .ZN(m_data_out_y[4]) );
  INV_X1 U36387 ( .A(n37298), .ZN(n37300) );
  NAND2_X1 U36388 ( .A1(n37300), .A2(n37299), .ZN(n37302) );
  XOR2_X1 U36389 ( .A(n37302), .B(n37301), .Z(m_data_out_y[3]) );
  INV_X1 U36390 ( .A(n37303), .ZN(n37305) );
  NAND2_X1 U36391 ( .A1(n37305), .A2(n37304), .ZN(n37307) );
  XNOR2_X1 U36392 ( .A(n37307), .B(n37306), .ZN(m_data_out_y[2]) );
  FA_X1 U36393 ( .A(n37310), .B(n37309), .CI(n37308), .CO(n37306), .S(
        m_data_out_y[1]) );
  FA_X1 U36394 ( .A(n37313), .B(n37312), .CI(n37311), .CO(n37309), .S(
        m_data_out_y[0]) );
  INV_X1 U36395 ( .A(n37669), .ZN(n37661) );
  AOI221_X1 U36396 ( .B1(\ctrl_conv_output_inst/conv_start_reg ), .B2(n39050), 
        .C1(n37314), .C2(n39050), .A(n37661), .ZN(n3115) );
  OAI22_X1 U36397 ( .A1(n39040), .A2(n38995), .B1(n38994), .B2(n37315), .ZN(
        n3114) );
  NAND2_X1 U36398 ( .A1(s_ready_f), .A2(s_valid_f), .ZN(n37323) );
  INV_X1 U36399 ( .A(n37323), .ZN(n37320) );
  AND2_X1 U36400 ( .A1(n37320), .A2(fmem_addr[3]), .ZN(n37572) );
  NAND2_X1 U36401 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n37317) );
  NOR2_X1 U36402 ( .A1(n39000), .A2(n37317), .ZN(n37395) );
  NAND2_X1 U36403 ( .A1(n37572), .A2(n37395), .ZN(n37322) );
  INV_X1 U36404 ( .A(n37322), .ZN(n37478) );
  NAND2_X1 U36405 ( .A1(n37478), .A2(fmem_addr[4]), .ZN(n37659) );
  INV_X1 U36406 ( .A(n37659), .ZN(n37658) );
  OAI21_X1 U36407 ( .B1(n37658), .B2(n39001), .A(n37669), .ZN(n3113) );
  AOI221_X1 U36408 ( .B1(n37320), .B2(fmem_addr[0]), .C1(n37323), .C2(n39046), 
        .A(n37661), .ZN(n3112) );
  NOR2_X1 U36409 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n37364) );
  OAI221_X1 U36410 ( .B1(n37320), .B2(fmem_addr[1]), .C1(n37323), .C2(n37317), 
        .A(n37669), .ZN(n37316) );
  NOR2_X1 U36411 ( .A1(n37364), .A2(n37316), .ZN(n3111) );
  NOR2_X1 U36412 ( .A1(n37317), .A2(n37323), .ZN(n37319) );
  OAI21_X1 U36413 ( .B1(fmem_addr[2]), .B2(n37319), .A(n37669), .ZN(n37318) );
  AOI21_X1 U36414 ( .B1(fmem_addr[2]), .B2(n37319), .A(n37318), .ZN(n3110) );
  OAI221_X1 U36415 ( .B1(fmem_addr[3]), .B2(n37395), .C1(fmem_addr[3]), .C2(
        n37320), .A(n37669), .ZN(n37321) );
  NOR2_X1 U36416 ( .A1(n37478), .A2(n37321), .ZN(n3109) );
  AOI221_X1 U36417 ( .B1(n37478), .B2(fmem_addr[4]), .C1(n37322), .C2(n39045), 
        .A(n37661), .ZN(n3108) );
  NAND2_X1 U36418 ( .A1(n37364), .A2(n39000), .ZN(n37573) );
  NOR2_X1 U36419 ( .A1(fmem_addr[3]), .A2(n37323), .ZN(n37489) );
  NAND2_X1 U36420 ( .A1(n37489), .A2(n39045), .ZN(n37396) );
  NOR2_X1 U36421 ( .A1(n37573), .A2(n37396), .ZN(n37331) );
  INV_X1 U36422 ( .A(n37331), .ZN(n37332) );
  OAI22_X1 U36423 ( .A1(n37332), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[0][0] ), .B2(n37331), .ZN(n37324) );
  INV_X1 U36424 ( .A(n37324), .ZN(n3107) );
  OAI22_X1 U36425 ( .A1(n37332), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[0][1] ), .B2(n37331), .ZN(n37325) );
  INV_X1 U36426 ( .A(n37325), .ZN(n3106) );
  OAI22_X1 U36427 ( .A1(n37332), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[0][2] ), .B2(n37331), .ZN(n37326) );
  INV_X1 U36428 ( .A(n37326), .ZN(n3105) );
  OAI22_X1 U36429 ( .A1(n37332), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[0][3] ), .B2(n37331), .ZN(n37327) );
  INV_X1 U36430 ( .A(n37327), .ZN(n3104) );
  OAI22_X1 U36431 ( .A1(n37332), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[0][4] ), .B2(n37331), .ZN(n37328) );
  INV_X1 U36432 ( .A(n37328), .ZN(n3103) );
  OAI22_X1 U36433 ( .A1(n37332), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[0][5] ), .B2(n37331), .ZN(n37329) );
  INV_X1 U36434 ( .A(n37329), .ZN(n3102) );
  OAI22_X1 U36435 ( .A1(n37332), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[0][6] ), .B2(n37331), .ZN(n37330) );
  INV_X1 U36436 ( .A(n37330), .ZN(n3101) );
  OAI22_X1 U36437 ( .A1(n37332), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[0][7] ), .B2(n37331), .ZN(n37333) );
  INV_X1 U36438 ( .A(n37333), .ZN(n3100) );
  NAND3_X1 U36439 ( .A1(fmem_addr[0]), .A2(n39000), .A3(n39047), .ZN(n37584)
         );
  NOR2_X1 U36440 ( .A1(n37396), .A2(n37584), .ZN(n37341) );
  INV_X1 U36441 ( .A(n37341), .ZN(n37342) );
  OAI22_X1 U36442 ( .A1(n37342), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[1][0] ), .B2(n37341), .ZN(n37334) );
  INV_X1 U36443 ( .A(n37334), .ZN(n3099) );
  OAI22_X1 U36444 ( .A1(n37342), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[1][1] ), .B2(n37341), .ZN(n37335) );
  INV_X1 U36445 ( .A(n37335), .ZN(n3098) );
  OAI22_X1 U36446 ( .A1(n37342), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[1][2] ), .B2(n37341), .ZN(n37336) );
  INV_X1 U36447 ( .A(n37336), .ZN(n3097) );
  OAI22_X1 U36448 ( .A1(n37342), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[1][3] ), .B2(n37341), .ZN(n37337) );
  INV_X1 U36449 ( .A(n37337), .ZN(n3096) );
  OAI22_X1 U36450 ( .A1(n37342), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[1][4] ), .B2(n37341), .ZN(n37338) );
  INV_X1 U36451 ( .A(n37338), .ZN(n3095) );
  OAI22_X1 U36452 ( .A1(n37342), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[1][5] ), .B2(n37341), .ZN(n37339) );
  INV_X1 U36453 ( .A(n37339), .ZN(n3094) );
  OAI22_X1 U36454 ( .A1(n37342), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[1][6] ), .B2(n37341), .ZN(n37340) );
  INV_X1 U36455 ( .A(n37340), .ZN(n3093) );
  OAI22_X1 U36456 ( .A1(n37342), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[1][7] ), .B2(n37341), .ZN(n37343) );
  INV_X1 U36457 ( .A(n37343), .ZN(n3092) );
  NAND3_X1 U36458 ( .A1(fmem_addr[1]), .A2(n39000), .A3(n39046), .ZN(n37595)
         );
  NOR2_X1 U36459 ( .A1(n37396), .A2(n37595), .ZN(n37351) );
  INV_X1 U36460 ( .A(n37351), .ZN(n37352) );
  OAI22_X1 U36461 ( .A1(n37352), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[2][0] ), .B2(n37351), .ZN(n37344) );
  INV_X1 U36462 ( .A(n37344), .ZN(n3091) );
  OAI22_X1 U36463 ( .A1(n37352), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[2][1] ), .B2(n37351), .ZN(n37345) );
  INV_X1 U36464 ( .A(n37345), .ZN(n3090) );
  OAI22_X1 U36465 ( .A1(n37352), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[2][2] ), .B2(n37351), .ZN(n37346) );
  INV_X1 U36466 ( .A(n37346), .ZN(n3089) );
  OAI22_X1 U36467 ( .A1(n37352), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[2][3] ), .B2(n37351), .ZN(n37347) );
  INV_X1 U36468 ( .A(n37347), .ZN(n3088) );
  OAI22_X1 U36469 ( .A1(n37352), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[2][4] ), .B2(n37351), .ZN(n37348) );
  INV_X1 U36470 ( .A(n37348), .ZN(n3087) );
  OAI22_X1 U36471 ( .A1(n37352), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[2][5] ), .B2(n37351), .ZN(n37349) );
  INV_X1 U36472 ( .A(n37349), .ZN(n3086) );
  OAI22_X1 U36473 ( .A1(n37352), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[2][6] ), .B2(n37351), .ZN(n37350) );
  INV_X1 U36474 ( .A(n37350), .ZN(n3085) );
  OAI22_X1 U36475 ( .A1(n37352), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[2][7] ), .B2(n37351), .ZN(n37353) );
  INV_X1 U36476 ( .A(n37353), .ZN(n3084) );
  NAND3_X1 U36477 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .A3(n39000), .ZN(
        n37606) );
  NOR2_X1 U36478 ( .A1(n37606), .A2(n37396), .ZN(n37361) );
  INV_X1 U36479 ( .A(n37361), .ZN(n37362) );
  OAI22_X1 U36480 ( .A1(n37362), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[3][0] ), .B2(n37361), .ZN(n37354) );
  INV_X1 U36481 ( .A(n37354), .ZN(n3083) );
  OAI22_X1 U36482 ( .A1(n37362), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[3][1] ), .B2(n37361), .ZN(n37355) );
  INV_X1 U36483 ( .A(n37355), .ZN(n3082) );
  OAI22_X1 U36484 ( .A1(n37362), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[3][2] ), .B2(n37361), .ZN(n37356) );
  INV_X1 U36485 ( .A(n37356), .ZN(n3081) );
  OAI22_X1 U36486 ( .A1(n37362), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[3][3] ), .B2(n37361), .ZN(n37357) );
  INV_X1 U36487 ( .A(n37357), .ZN(n3080) );
  OAI22_X1 U36488 ( .A1(n37362), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[3][4] ), .B2(n37361), .ZN(n37358) );
  INV_X1 U36489 ( .A(n37358), .ZN(n3079) );
  OAI22_X1 U36490 ( .A1(n37362), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[3][5] ), .B2(n37361), .ZN(n37359) );
  INV_X1 U36491 ( .A(n37359), .ZN(n3078) );
  OAI22_X1 U36492 ( .A1(n37362), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[3][6] ), .B2(n37361), .ZN(n37360) );
  INV_X1 U36493 ( .A(n37360), .ZN(n3077) );
  OAI22_X1 U36494 ( .A1(n37362), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[3][7] ), .B2(n37361), .ZN(n37363) );
  INV_X1 U36495 ( .A(n37363), .ZN(n3076) );
  NAND2_X1 U36496 ( .A1(fmem_addr[2]), .A2(n37364), .ZN(n37617) );
  NOR2_X1 U36497 ( .A1(n37396), .A2(n37617), .ZN(n37372) );
  INV_X1 U36498 ( .A(n37372), .ZN(n37373) );
  OAI22_X1 U36499 ( .A1(n37373), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[4][0] ), .B2(n37372), .ZN(n37365) );
  INV_X1 U36500 ( .A(n37365), .ZN(n3075) );
  OAI22_X1 U36501 ( .A1(n37373), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[4][1] ), .B2(n37372), .ZN(n37366) );
  INV_X1 U36502 ( .A(n37366), .ZN(n3074) );
  OAI22_X1 U36503 ( .A1(n37373), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[4][2] ), .B2(n37372), .ZN(n37367) );
  INV_X1 U36504 ( .A(n37367), .ZN(n3073) );
  OAI22_X1 U36505 ( .A1(n37373), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[4][3] ), .B2(n37372), .ZN(n37368) );
  INV_X1 U36506 ( .A(n37368), .ZN(n3072) );
  OAI22_X1 U36507 ( .A1(n37373), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[4][4] ), .B2(n37372), .ZN(n37369) );
  INV_X1 U36508 ( .A(n37369), .ZN(n3071) );
  OAI22_X1 U36509 ( .A1(n37373), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[4][5] ), .B2(n37372), .ZN(n37370) );
  INV_X1 U36510 ( .A(n37370), .ZN(n3070) );
  OAI22_X1 U36511 ( .A1(n37373), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[4][6] ), .B2(n37372), .ZN(n37371) );
  INV_X1 U36512 ( .A(n37371), .ZN(n3069) );
  OAI22_X1 U36513 ( .A1(n37373), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[4][7] ), .B2(n37372), .ZN(n37374) );
  INV_X1 U36514 ( .A(n37374), .ZN(n3068) );
  NAND3_X1 U36515 ( .A1(fmem_addr[0]), .A2(fmem_addr[2]), .A3(n39047), .ZN(
        n37628) );
  NOR2_X1 U36516 ( .A1(n37396), .A2(n37628), .ZN(n37382) );
  INV_X1 U36517 ( .A(n37382), .ZN(n37383) );
  OAI22_X1 U36518 ( .A1(n37383), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[5][0] ), .B2(n37382), .ZN(n37375) );
  INV_X1 U36519 ( .A(n37375), .ZN(n3067) );
  OAI22_X1 U36520 ( .A1(n37383), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[5][1] ), .B2(n37382), .ZN(n37376) );
  INV_X1 U36521 ( .A(n37376), .ZN(n3066) );
  OAI22_X1 U36522 ( .A1(n37383), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[5][2] ), .B2(n37382), .ZN(n37377) );
  INV_X1 U36523 ( .A(n37377), .ZN(n3065) );
  OAI22_X1 U36524 ( .A1(n37383), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[5][3] ), .B2(n37382), .ZN(n37378) );
  INV_X1 U36525 ( .A(n37378), .ZN(n3064) );
  OAI22_X1 U36526 ( .A1(n37383), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[5][4] ), .B2(n37382), .ZN(n37379) );
  INV_X1 U36527 ( .A(n37379), .ZN(n3063) );
  OAI22_X1 U36528 ( .A1(n37383), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[5][5] ), .B2(n37382), .ZN(n37380) );
  INV_X1 U36529 ( .A(n37380), .ZN(n3062) );
  OAI22_X1 U36530 ( .A1(n37383), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[5][6] ), .B2(n37382), .ZN(n37381) );
  INV_X1 U36531 ( .A(n37381), .ZN(n3061) );
  OAI22_X1 U36532 ( .A1(n37383), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[5][7] ), .B2(n37382), .ZN(n37384) );
  INV_X1 U36533 ( .A(n37384), .ZN(n3060) );
  NAND3_X1 U36534 ( .A1(fmem_addr[2]), .A2(fmem_addr[1]), .A3(n39046), .ZN(
        n37640) );
  NOR2_X1 U36535 ( .A1(n37396), .A2(n37640), .ZN(n37392) );
  INV_X1 U36536 ( .A(n37392), .ZN(n37393) );
  OAI22_X1 U36537 ( .A1(n37393), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[6][0] ), .B2(n37392), .ZN(n37385) );
  INV_X1 U36538 ( .A(n37385), .ZN(n3059) );
  OAI22_X1 U36539 ( .A1(n37393), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[6][1] ), .B2(n37392), .ZN(n37386) );
  INV_X1 U36540 ( .A(n37386), .ZN(n3058) );
  OAI22_X1 U36541 ( .A1(n37393), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[6][2] ), .B2(n37392), .ZN(n37387) );
  INV_X1 U36542 ( .A(n37387), .ZN(n3057) );
  OAI22_X1 U36543 ( .A1(n37393), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[6][3] ), .B2(n37392), .ZN(n37388) );
  INV_X1 U36544 ( .A(n37388), .ZN(n3056) );
  OAI22_X1 U36545 ( .A1(n37393), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[6][4] ), .B2(n37392), .ZN(n37389) );
  INV_X1 U36546 ( .A(n37389), .ZN(n3055) );
  OAI22_X1 U36547 ( .A1(n37393), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[6][5] ), .B2(n37392), .ZN(n37390) );
  INV_X1 U36548 ( .A(n37390), .ZN(n3054) );
  OAI22_X1 U36549 ( .A1(n37393), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[6][6] ), .B2(n37392), .ZN(n37391) );
  INV_X1 U36550 ( .A(n37391), .ZN(n3053) );
  OAI22_X1 U36551 ( .A1(n37393), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[6][7] ), .B2(n37392), .ZN(n37394) );
  INV_X1 U36552 ( .A(n37394), .ZN(n3052) );
  INV_X1 U36553 ( .A(n37395), .ZN(n37561) );
  NOR2_X1 U36554 ( .A1(n37561), .A2(n37396), .ZN(n37404) );
  INV_X1 U36555 ( .A(n37404), .ZN(n37405) );
  OAI22_X1 U36556 ( .A1(n37405), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[7][0] ), .B2(n37404), .ZN(n37397) );
  INV_X1 U36557 ( .A(n37397), .ZN(n3051) );
  OAI22_X1 U36558 ( .A1(n37405), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[7][1] ), .B2(n37404), .ZN(n37398) );
  INV_X1 U36559 ( .A(n37398), .ZN(n3050) );
  OAI22_X1 U36560 ( .A1(n37405), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[7][2] ), .B2(n37404), .ZN(n37399) );
  INV_X1 U36561 ( .A(n37399), .ZN(n3049) );
  OAI22_X1 U36562 ( .A1(n37405), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[7][3] ), .B2(n37404), .ZN(n37400) );
  INV_X1 U36563 ( .A(n37400), .ZN(n3048) );
  OAI22_X1 U36564 ( .A1(n37405), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[7][4] ), .B2(n37404), .ZN(n37401) );
  INV_X1 U36565 ( .A(n37401), .ZN(n3047) );
  OAI22_X1 U36566 ( .A1(n37405), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[7][5] ), .B2(n37404), .ZN(n37402) );
  INV_X1 U36567 ( .A(n37402), .ZN(n3046) );
  OAI22_X1 U36568 ( .A1(n37405), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[7][6] ), .B2(n37404), .ZN(n37403) );
  INV_X1 U36569 ( .A(n37403), .ZN(n3045) );
  OAI22_X1 U36570 ( .A1(n37405), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[7][7] ), .B2(n37404), .ZN(n37406) );
  INV_X1 U36571 ( .A(n37406), .ZN(n3044) );
  NAND2_X1 U36572 ( .A1(n37572), .A2(n39045), .ZN(n37467) );
  NOR2_X1 U36573 ( .A1(n37573), .A2(n37467), .ZN(n37414) );
  INV_X1 U36574 ( .A(n37414), .ZN(n37415) );
  OAI22_X1 U36575 ( .A1(n37415), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[8][0] ), .B2(n37414), .ZN(n37407) );
  INV_X1 U36576 ( .A(n37407), .ZN(n3043) );
  OAI22_X1 U36577 ( .A1(n37415), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[8][1] ), .B2(n37414), .ZN(n37408) );
  INV_X1 U36578 ( .A(n37408), .ZN(n3042) );
  OAI22_X1 U36579 ( .A1(n37415), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[8][2] ), .B2(n37414), .ZN(n37409) );
  INV_X1 U36580 ( .A(n37409), .ZN(n3041) );
  OAI22_X1 U36581 ( .A1(n37415), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[8][3] ), .B2(n37414), .ZN(n37410) );
  INV_X1 U36582 ( .A(n37410), .ZN(n3040) );
  OAI22_X1 U36583 ( .A1(n37415), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[8][4] ), .B2(n37414), .ZN(n37411) );
  INV_X1 U36584 ( .A(n37411), .ZN(n3039) );
  OAI22_X1 U36585 ( .A1(n37415), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[8][5] ), .B2(n37414), .ZN(n37412) );
  INV_X1 U36586 ( .A(n37412), .ZN(n3038) );
  OAI22_X1 U36587 ( .A1(n37415), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[8][6] ), .B2(n37414), .ZN(n37413) );
  INV_X1 U36588 ( .A(n37413), .ZN(n3037) );
  OAI22_X1 U36589 ( .A1(n37415), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[8][7] ), .B2(n37414), .ZN(n37416) );
  INV_X1 U36590 ( .A(n37416), .ZN(n3036) );
  NOR2_X1 U36591 ( .A1(n37584), .A2(n37467), .ZN(n37424) );
  INV_X1 U36592 ( .A(n37424), .ZN(n37425) );
  OAI22_X1 U36593 ( .A1(n37425), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[9][0] ), .B2(n37424), .ZN(n37417) );
  INV_X1 U36594 ( .A(n37417), .ZN(n3035) );
  OAI22_X1 U36595 ( .A1(n37425), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[9][1] ), .B2(n37424), .ZN(n37418) );
  INV_X1 U36596 ( .A(n37418), .ZN(n3034) );
  OAI22_X1 U36597 ( .A1(n37425), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[9][2] ), .B2(n37424), .ZN(n37419) );
  INV_X1 U36598 ( .A(n37419), .ZN(n3033) );
  OAI22_X1 U36599 ( .A1(n37425), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[9][3] ), .B2(n37424), .ZN(n37420) );
  INV_X1 U36600 ( .A(n37420), .ZN(n3032) );
  OAI22_X1 U36601 ( .A1(n37425), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[9][4] ), .B2(n37424), .ZN(n37421) );
  INV_X1 U36602 ( .A(n37421), .ZN(n3031) );
  OAI22_X1 U36603 ( .A1(n37425), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[9][5] ), .B2(n37424), .ZN(n37422) );
  INV_X1 U36604 ( .A(n37422), .ZN(n3030) );
  OAI22_X1 U36605 ( .A1(n37425), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[9][6] ), .B2(n37424), .ZN(n37423) );
  INV_X1 U36606 ( .A(n37423), .ZN(n3029) );
  OAI22_X1 U36607 ( .A1(n37425), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[9][7] ), .B2(n37424), .ZN(n37426) );
  INV_X1 U36608 ( .A(n37426), .ZN(n3028) );
  NOR2_X1 U36609 ( .A1(n37595), .A2(n37467), .ZN(n37434) );
  INV_X1 U36610 ( .A(n37434), .ZN(n37435) );
  OAI22_X1 U36611 ( .A1(n37435), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[10][0] ), .B2(n37434), .ZN(n37427) );
  INV_X1 U36612 ( .A(n37427), .ZN(n3027) );
  OAI22_X1 U36613 ( .A1(n37435), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[10][1] ), .B2(n37434), .ZN(n37428) );
  INV_X1 U36614 ( .A(n37428), .ZN(n3026) );
  OAI22_X1 U36615 ( .A1(n37435), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[10][2] ), .B2(n37434), .ZN(n37429) );
  INV_X1 U36616 ( .A(n37429), .ZN(n3025) );
  OAI22_X1 U36617 ( .A1(n37435), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[10][3] ), .B2(n37434), .ZN(n37430) );
  INV_X1 U36618 ( .A(n37430), .ZN(n3024) );
  OAI22_X1 U36619 ( .A1(n37435), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[10][4] ), .B2(n37434), .ZN(n37431) );
  INV_X1 U36620 ( .A(n37431), .ZN(n3023) );
  OAI22_X1 U36621 ( .A1(n37435), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[10][5] ), .B2(n37434), .ZN(n37432) );
  INV_X1 U36622 ( .A(n37432), .ZN(n3022) );
  OAI22_X1 U36623 ( .A1(n37435), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[10][6] ), .B2(n37434), .ZN(n37433) );
  INV_X1 U36624 ( .A(n37433), .ZN(n3021) );
  OAI22_X1 U36625 ( .A1(n37435), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[10][7] ), .B2(n37434), .ZN(n37436) );
  INV_X1 U36626 ( .A(n37436), .ZN(n3020) );
  NOR2_X1 U36627 ( .A1(n37606), .A2(n37467), .ZN(n37444) );
  INV_X1 U36628 ( .A(n37444), .ZN(n37445) );
  OAI22_X1 U36629 ( .A1(n37445), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[11][0] ), .B2(n37444), .ZN(n37437) );
  INV_X1 U36630 ( .A(n37437), .ZN(n3019) );
  OAI22_X1 U36631 ( .A1(n37445), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[11][1] ), .B2(n37444), .ZN(n37438) );
  INV_X1 U36632 ( .A(n37438), .ZN(n3018) );
  OAI22_X1 U36633 ( .A1(n37445), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[11][2] ), .B2(n37444), .ZN(n37439) );
  INV_X1 U36634 ( .A(n37439), .ZN(n3017) );
  OAI22_X1 U36635 ( .A1(n37445), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[11][3] ), .B2(n37444), .ZN(n37440) );
  INV_X1 U36636 ( .A(n37440), .ZN(n3016) );
  OAI22_X1 U36637 ( .A1(n37445), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[11][4] ), .B2(n37444), .ZN(n37441) );
  INV_X1 U36638 ( .A(n37441), .ZN(n3015) );
  OAI22_X1 U36639 ( .A1(n37445), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[11][5] ), .B2(n37444), .ZN(n37442) );
  INV_X1 U36640 ( .A(n37442), .ZN(n3014) );
  OAI22_X1 U36641 ( .A1(n37445), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[11][6] ), .B2(n37444), .ZN(n37443) );
  INV_X1 U36642 ( .A(n37443), .ZN(n3013) );
  OAI22_X1 U36643 ( .A1(n37445), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[11][7] ), .B2(n37444), .ZN(n37446) );
  INV_X1 U36644 ( .A(n37446), .ZN(n3012) );
  NOR2_X1 U36645 ( .A1(n37617), .A2(n37467), .ZN(n37454) );
  INV_X1 U36646 ( .A(n37454), .ZN(n37455) );
  OAI22_X1 U36647 ( .A1(n37455), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[12][0] ), .B2(n37454), .ZN(n37447) );
  INV_X1 U36648 ( .A(n37447), .ZN(n3011) );
  OAI22_X1 U36649 ( .A1(n37455), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[12][1] ), .B2(n37454), .ZN(n37448) );
  INV_X1 U36650 ( .A(n37448), .ZN(n3010) );
  OAI22_X1 U36651 ( .A1(n37455), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[12][2] ), .B2(n37454), .ZN(n37449) );
  INV_X1 U36652 ( .A(n37449), .ZN(n3009) );
  OAI22_X1 U36653 ( .A1(n37455), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[12][3] ), .B2(n37454), .ZN(n37450) );
  INV_X1 U36654 ( .A(n37450), .ZN(n3008) );
  OAI22_X1 U36655 ( .A1(n37455), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[12][4] ), .B2(n37454), .ZN(n37451) );
  INV_X1 U36656 ( .A(n37451), .ZN(n3007) );
  OAI22_X1 U36657 ( .A1(n37455), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[12][5] ), .B2(n37454), .ZN(n37452) );
  INV_X1 U36658 ( .A(n37452), .ZN(n3006) );
  OAI22_X1 U36659 ( .A1(n37455), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[12][6] ), .B2(n37454), .ZN(n37453) );
  INV_X1 U36660 ( .A(n37453), .ZN(n3005) );
  OAI22_X1 U36661 ( .A1(n37455), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[12][7] ), .B2(n37454), .ZN(n37456) );
  INV_X1 U36662 ( .A(n37456), .ZN(n3004) );
  NOR2_X1 U36663 ( .A1(n37628), .A2(n37467), .ZN(n37464) );
  INV_X1 U36664 ( .A(n37464), .ZN(n37465) );
  OAI22_X1 U36665 ( .A1(n37465), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[13][0] ), .B2(n37464), .ZN(n37457) );
  INV_X1 U36666 ( .A(n37457), .ZN(n3003) );
  OAI22_X1 U36667 ( .A1(n37465), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[13][1] ), .B2(n37464), .ZN(n37458) );
  INV_X1 U36668 ( .A(n37458), .ZN(n3002) );
  OAI22_X1 U36669 ( .A1(n37465), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[13][2] ), .B2(n37464), .ZN(n37459) );
  INV_X1 U36670 ( .A(n37459), .ZN(n3001) );
  OAI22_X1 U36671 ( .A1(n37465), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[13][3] ), .B2(n37464), .ZN(n37460) );
  INV_X1 U36672 ( .A(n37460), .ZN(n3000) );
  OAI22_X1 U36673 ( .A1(n37465), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[13][4] ), .B2(n37464), .ZN(n37461) );
  INV_X1 U36674 ( .A(n37461), .ZN(n2999) );
  OAI22_X1 U36675 ( .A1(n37465), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[13][5] ), .B2(n37464), .ZN(n37462) );
  INV_X1 U36676 ( .A(n37462), .ZN(n2998) );
  OAI22_X1 U36677 ( .A1(n37465), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[13][6] ), .B2(n37464), .ZN(n37463) );
  INV_X1 U36678 ( .A(n37463), .ZN(n2997) );
  OAI22_X1 U36679 ( .A1(n37465), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[13][7] ), .B2(n37464), .ZN(n37466) );
  INV_X1 U36680 ( .A(n37466), .ZN(n2996) );
  NOR2_X1 U36681 ( .A1(n37640), .A2(n37467), .ZN(n37475) );
  INV_X1 U36682 ( .A(n37475), .ZN(n37476) );
  OAI22_X1 U36683 ( .A1(n37476), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[14][0] ), .B2(n37475), .ZN(n37468) );
  INV_X1 U36684 ( .A(n37468), .ZN(n2995) );
  OAI22_X1 U36685 ( .A1(n37476), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[14][1] ), .B2(n37475), .ZN(n37469) );
  INV_X1 U36686 ( .A(n37469), .ZN(n2994) );
  OAI22_X1 U36687 ( .A1(n37476), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[14][2] ), .B2(n37475), .ZN(n37470) );
  INV_X1 U36688 ( .A(n37470), .ZN(n2993) );
  OAI22_X1 U36689 ( .A1(n37476), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[14][3] ), .B2(n37475), .ZN(n37471) );
  INV_X1 U36690 ( .A(n37471), .ZN(n2992) );
  OAI22_X1 U36691 ( .A1(n37476), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[14][4] ), .B2(n37475), .ZN(n37472) );
  INV_X1 U36692 ( .A(n37472), .ZN(n2991) );
  OAI22_X1 U36693 ( .A1(n37476), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[14][5] ), .B2(n37475), .ZN(n37473) );
  INV_X1 U36694 ( .A(n37473), .ZN(n2990) );
  OAI22_X1 U36695 ( .A1(n37476), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[14][6] ), .B2(n37475), .ZN(n37474) );
  INV_X1 U36696 ( .A(n37474), .ZN(n2989) );
  OAI22_X1 U36697 ( .A1(n37476), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[14][7] ), .B2(n37475), .ZN(n37477) );
  INV_X1 U36698 ( .A(n37477), .ZN(n2988) );
  NAND2_X1 U36699 ( .A1(n39045), .A2(n37478), .ZN(n37487) );
  INV_X1 U36700 ( .A(n37487), .ZN(n37486) );
  OAI22_X1 U36701 ( .A1(n37487), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[15][0] ), .B2(n37486), .ZN(n37479) );
  INV_X1 U36702 ( .A(n37479), .ZN(n2987) );
  OAI22_X1 U36703 ( .A1(n37487), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[15][1] ), .B2(n37486), .ZN(n37480) );
  INV_X1 U36704 ( .A(n37480), .ZN(n2986) );
  OAI22_X1 U36705 ( .A1(n37487), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[15][2] ), .B2(n37486), .ZN(n37481) );
  INV_X1 U36706 ( .A(n37481), .ZN(n2985) );
  OAI22_X1 U36707 ( .A1(n37487), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[15][3] ), .B2(n37486), .ZN(n37482) );
  INV_X1 U36708 ( .A(n37482), .ZN(n2984) );
  OAI22_X1 U36709 ( .A1(n37487), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[15][4] ), .B2(n37486), .ZN(n37483) );
  INV_X1 U36710 ( .A(n37483), .ZN(n2983) );
  OAI22_X1 U36711 ( .A1(n37487), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[15][5] ), .B2(n37486), .ZN(n37484) );
  INV_X1 U36712 ( .A(n37484), .ZN(n2982) );
  OAI22_X1 U36713 ( .A1(n37487), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[15][6] ), .B2(n37486), .ZN(n37485) );
  INV_X1 U36714 ( .A(n37485), .ZN(n2981) );
  OAI22_X1 U36715 ( .A1(n37487), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[15][7] ), .B2(n37486), .ZN(n37488) );
  INV_X1 U36716 ( .A(n37488), .ZN(n2980) );
  NAND2_X1 U36717 ( .A1(fmem_addr[4]), .A2(n37489), .ZN(n37560) );
  NOR2_X1 U36718 ( .A1(n37573), .A2(n37560), .ZN(n37497) );
  INV_X1 U36719 ( .A(n37497), .ZN(n37498) );
  OAI22_X1 U36720 ( .A1(n37498), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[16][0] ), .B2(n37497), .ZN(n37490) );
  INV_X1 U36721 ( .A(n37490), .ZN(n2979) );
  OAI22_X1 U36722 ( .A1(n37498), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[16][1] ), .B2(n37497), .ZN(n37491) );
  INV_X1 U36723 ( .A(n37491), .ZN(n2978) );
  OAI22_X1 U36724 ( .A1(n37498), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[16][2] ), .B2(n37497), .ZN(n37492) );
  INV_X1 U36725 ( .A(n37492), .ZN(n2977) );
  OAI22_X1 U36726 ( .A1(n37498), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[16][3] ), .B2(n37497), .ZN(n37493) );
  INV_X1 U36727 ( .A(n37493), .ZN(n2976) );
  OAI22_X1 U36728 ( .A1(n37498), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[16][4] ), .B2(n37497), .ZN(n37494) );
  INV_X1 U36729 ( .A(n37494), .ZN(n2975) );
  OAI22_X1 U36730 ( .A1(n37498), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[16][5] ), .B2(n37497), .ZN(n37495) );
  INV_X1 U36731 ( .A(n37495), .ZN(n2974) );
  OAI22_X1 U36732 ( .A1(n37498), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[16][6] ), .B2(n37497), .ZN(n37496) );
  INV_X1 U36733 ( .A(n37496), .ZN(n2973) );
  OAI22_X1 U36734 ( .A1(n37498), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[16][7] ), .B2(n37497), .ZN(n37499) );
  INV_X1 U36735 ( .A(n37499), .ZN(n2972) );
  NOR2_X1 U36736 ( .A1(n37584), .A2(n37560), .ZN(n37507) );
  INV_X1 U36737 ( .A(n37507), .ZN(n37508) );
  OAI22_X1 U36738 ( .A1(n37508), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[17][0] ), .B2(n37507), .ZN(n37500) );
  INV_X1 U36739 ( .A(n37500), .ZN(n2971) );
  OAI22_X1 U36740 ( .A1(n37508), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[17][1] ), .B2(n37507), .ZN(n37501) );
  INV_X1 U36741 ( .A(n37501), .ZN(n2970) );
  OAI22_X1 U36742 ( .A1(n37508), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[17][2] ), .B2(n37507), .ZN(n37502) );
  INV_X1 U36743 ( .A(n37502), .ZN(n2969) );
  OAI22_X1 U36744 ( .A1(n37508), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[17][3] ), .B2(n37507), .ZN(n37503) );
  INV_X1 U36745 ( .A(n37503), .ZN(n2968) );
  OAI22_X1 U36746 ( .A1(n37508), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[17][4] ), .B2(n37507), .ZN(n37504) );
  INV_X1 U36747 ( .A(n37504), .ZN(n2967) );
  OAI22_X1 U36748 ( .A1(n37508), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[17][5] ), .B2(n37507), .ZN(n37505) );
  INV_X1 U36749 ( .A(n37505), .ZN(n2966) );
  OAI22_X1 U36750 ( .A1(n37508), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[17][6] ), .B2(n37507), .ZN(n37506) );
  INV_X1 U36751 ( .A(n37506), .ZN(n2965) );
  OAI22_X1 U36752 ( .A1(n37508), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[17][7] ), .B2(n37507), .ZN(n37509) );
  INV_X1 U36753 ( .A(n37509), .ZN(n2964) );
  NOR2_X1 U36754 ( .A1(n37595), .A2(n37560), .ZN(n37517) );
  INV_X1 U36755 ( .A(n37517), .ZN(n37518) );
  OAI22_X1 U36756 ( .A1(n37518), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[18][0] ), .B2(n37517), .ZN(n37510) );
  INV_X1 U36757 ( .A(n37510), .ZN(n2963) );
  OAI22_X1 U36758 ( .A1(n37518), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[18][1] ), .B2(n37517), .ZN(n37511) );
  INV_X1 U36759 ( .A(n37511), .ZN(n2962) );
  OAI22_X1 U36760 ( .A1(n37518), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[18][2] ), .B2(n37517), .ZN(n37512) );
  INV_X1 U36761 ( .A(n37512), .ZN(n2961) );
  OAI22_X1 U36762 ( .A1(n37518), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[18][3] ), .B2(n37517), .ZN(n37513) );
  INV_X1 U36763 ( .A(n37513), .ZN(n2960) );
  OAI22_X1 U36764 ( .A1(n37518), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[18][4] ), .B2(n37517), .ZN(n37514) );
  INV_X1 U36765 ( .A(n37514), .ZN(n2959) );
  OAI22_X1 U36766 ( .A1(n37518), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[18][5] ), .B2(n37517), .ZN(n37515) );
  INV_X1 U36767 ( .A(n37515), .ZN(n2958) );
  OAI22_X1 U36768 ( .A1(n37518), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[18][6] ), .B2(n37517), .ZN(n37516) );
  INV_X1 U36769 ( .A(n37516), .ZN(n2957) );
  OAI22_X1 U36770 ( .A1(n37518), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[18][7] ), .B2(n37517), .ZN(n37519) );
  INV_X1 U36771 ( .A(n37519), .ZN(n2956) );
  NOR2_X1 U36772 ( .A1(n37606), .A2(n37560), .ZN(n37527) );
  INV_X1 U36773 ( .A(n37527), .ZN(n37528) );
  OAI22_X1 U36774 ( .A1(n37528), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[19][0] ), .B2(n37527), .ZN(n37520) );
  INV_X1 U36775 ( .A(n37520), .ZN(n2955) );
  OAI22_X1 U36776 ( .A1(n37528), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[19][1] ), .B2(n37527), .ZN(n37521) );
  INV_X1 U36777 ( .A(n37521), .ZN(n2954) );
  OAI22_X1 U36778 ( .A1(n37528), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[19][2] ), .B2(n37527), .ZN(n37522) );
  INV_X1 U36779 ( .A(n37522), .ZN(n2953) );
  OAI22_X1 U36780 ( .A1(n37528), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[19][3] ), .B2(n37527), .ZN(n37523) );
  INV_X1 U36781 ( .A(n37523), .ZN(n2952) );
  OAI22_X1 U36782 ( .A1(n37528), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[19][4] ), .B2(n37527), .ZN(n37524) );
  INV_X1 U36783 ( .A(n37524), .ZN(n2951) );
  OAI22_X1 U36784 ( .A1(n37528), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[19][5] ), .B2(n37527), .ZN(n37525) );
  INV_X1 U36785 ( .A(n37525), .ZN(n2950) );
  OAI22_X1 U36786 ( .A1(n37528), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[19][6] ), .B2(n37527), .ZN(n37526) );
  INV_X1 U36787 ( .A(n37526), .ZN(n2949) );
  OAI22_X1 U36788 ( .A1(n37528), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[19][7] ), .B2(n37527), .ZN(n37529) );
  INV_X1 U36789 ( .A(n37529), .ZN(n2948) );
  NOR2_X1 U36790 ( .A1(n37617), .A2(n37560), .ZN(n37537) );
  INV_X1 U36791 ( .A(n37537), .ZN(n37538) );
  OAI22_X1 U36792 ( .A1(n37538), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[20][0] ), .B2(n37537), .ZN(n37530) );
  INV_X1 U36793 ( .A(n37530), .ZN(n2947) );
  OAI22_X1 U36794 ( .A1(n37538), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[20][1] ), .B2(n37537), .ZN(n37531) );
  INV_X1 U36795 ( .A(n37531), .ZN(n2946) );
  OAI22_X1 U36796 ( .A1(n37538), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[20][2] ), .B2(n37537), .ZN(n37532) );
  INV_X1 U36797 ( .A(n37532), .ZN(n2945) );
  OAI22_X1 U36798 ( .A1(n37538), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[20][3] ), .B2(n37537), .ZN(n37533) );
  INV_X1 U36799 ( .A(n37533), .ZN(n2944) );
  OAI22_X1 U36800 ( .A1(n37538), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[20][4] ), .B2(n37537), .ZN(n37534) );
  INV_X1 U36801 ( .A(n37534), .ZN(n2943) );
  OAI22_X1 U36802 ( .A1(n37538), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[20][5] ), .B2(n37537), .ZN(n37535) );
  INV_X1 U36803 ( .A(n37535), .ZN(n2942) );
  OAI22_X1 U36804 ( .A1(n37538), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[20][6] ), .B2(n37537), .ZN(n37536) );
  INV_X1 U36805 ( .A(n37536), .ZN(n2941) );
  OAI22_X1 U36806 ( .A1(n37538), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[20][7] ), .B2(n37537), .ZN(n37539) );
  INV_X1 U36807 ( .A(n37539), .ZN(n2940) );
  NOR2_X1 U36808 ( .A1(n37628), .A2(n37560), .ZN(n37547) );
  INV_X1 U36809 ( .A(n37547), .ZN(n37548) );
  OAI22_X1 U36810 ( .A1(n37548), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[21][0] ), .B2(n37547), .ZN(n37540) );
  INV_X1 U36811 ( .A(n37540), .ZN(n2939) );
  OAI22_X1 U36812 ( .A1(n37548), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[21][1] ), .B2(n37547), .ZN(n37541) );
  INV_X1 U36813 ( .A(n37541), .ZN(n2938) );
  OAI22_X1 U36814 ( .A1(n37548), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[21][2] ), .B2(n37547), .ZN(n37542) );
  INV_X1 U36815 ( .A(n37542), .ZN(n2937) );
  OAI22_X1 U36816 ( .A1(n37548), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[21][3] ), .B2(n37547), .ZN(n37543) );
  INV_X1 U36817 ( .A(n37543), .ZN(n2936) );
  OAI22_X1 U36818 ( .A1(n37548), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[21][4] ), .B2(n37547), .ZN(n37544) );
  INV_X1 U36819 ( .A(n37544), .ZN(n2935) );
  OAI22_X1 U36820 ( .A1(n37548), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[21][5] ), .B2(n37547), .ZN(n37545) );
  INV_X1 U36821 ( .A(n37545), .ZN(n2934) );
  OAI22_X1 U36822 ( .A1(n37548), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[21][6] ), .B2(n37547), .ZN(n37546) );
  INV_X1 U36823 ( .A(n37546), .ZN(n2933) );
  OAI22_X1 U36824 ( .A1(n37548), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[21][7] ), .B2(n37547), .ZN(n37549) );
  INV_X1 U36825 ( .A(n37549), .ZN(n2932) );
  NOR2_X1 U36826 ( .A1(n37640), .A2(n37560), .ZN(n37557) );
  INV_X1 U36827 ( .A(n37557), .ZN(n37558) );
  OAI22_X1 U36828 ( .A1(n37558), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[22][0] ), .B2(n37557), .ZN(n37550) );
  INV_X1 U36829 ( .A(n37550), .ZN(n2931) );
  OAI22_X1 U36830 ( .A1(n37558), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[22][1] ), .B2(n37557), .ZN(n37551) );
  INV_X1 U36831 ( .A(n37551), .ZN(n2930) );
  OAI22_X1 U36832 ( .A1(n37558), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[22][2] ), .B2(n37557), .ZN(n37552) );
  INV_X1 U36833 ( .A(n37552), .ZN(n2929) );
  OAI22_X1 U36834 ( .A1(n37558), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[22][3] ), .B2(n37557), .ZN(n37553) );
  INV_X1 U36835 ( .A(n37553), .ZN(n2928) );
  OAI22_X1 U36836 ( .A1(n37558), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[22][4] ), .B2(n37557), .ZN(n37554) );
  INV_X1 U36837 ( .A(n37554), .ZN(n2927) );
  OAI22_X1 U36838 ( .A1(n37558), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[22][5] ), .B2(n37557), .ZN(n37555) );
  INV_X1 U36839 ( .A(n37555), .ZN(n2926) );
  OAI22_X1 U36840 ( .A1(n37558), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[22][6] ), .B2(n37557), .ZN(n37556) );
  INV_X1 U36841 ( .A(n37556), .ZN(n2925) );
  OAI22_X1 U36842 ( .A1(n37558), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[22][7] ), .B2(n37557), .ZN(n37559) );
  INV_X1 U36843 ( .A(n37559), .ZN(n2924) );
  NOR2_X1 U36844 ( .A1(n37561), .A2(n37560), .ZN(n37569) );
  INV_X1 U36845 ( .A(n37569), .ZN(n37570) );
  OAI22_X1 U36846 ( .A1(n37570), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[23][0] ), .B2(n37569), .ZN(n37562) );
  INV_X1 U36847 ( .A(n37562), .ZN(n2923) );
  OAI22_X1 U36848 ( .A1(n37570), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[23][1] ), .B2(n37569), .ZN(n37563) );
  INV_X1 U36849 ( .A(n37563), .ZN(n2922) );
  OAI22_X1 U36850 ( .A1(n37570), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[23][2] ), .B2(n37569), .ZN(n37564) );
  INV_X1 U36851 ( .A(n37564), .ZN(n2921) );
  OAI22_X1 U36852 ( .A1(n37570), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[23][3] ), .B2(n37569), .ZN(n37565) );
  INV_X1 U36853 ( .A(n37565), .ZN(n2920) );
  OAI22_X1 U36854 ( .A1(n37570), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[23][4] ), .B2(n37569), .ZN(n37566) );
  INV_X1 U36855 ( .A(n37566), .ZN(n2919) );
  OAI22_X1 U36856 ( .A1(n37570), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[23][5] ), .B2(n37569), .ZN(n37567) );
  INV_X1 U36857 ( .A(n37567), .ZN(n2918) );
  OAI22_X1 U36858 ( .A1(n37570), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[23][6] ), .B2(n37569), .ZN(n37568) );
  INV_X1 U36859 ( .A(n37568), .ZN(n2917) );
  OAI22_X1 U36860 ( .A1(n37570), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[23][7] ), .B2(n37569), .ZN(n37571) );
  INV_X1 U36861 ( .A(n37571), .ZN(n2916) );
  NAND2_X1 U36862 ( .A1(n37572), .A2(fmem_addr[4]), .ZN(n37639) );
  NOR2_X1 U36863 ( .A1(n37573), .A2(n37639), .ZN(n37581) );
  INV_X1 U36864 ( .A(n37581), .ZN(n37582) );
  OAI22_X1 U36865 ( .A1(n37582), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[24][0] ), .B2(n37581), .ZN(n37574) );
  INV_X1 U36866 ( .A(n37574), .ZN(n2915) );
  OAI22_X1 U36867 ( .A1(n37582), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[24][1] ), .B2(n37581), .ZN(n37575) );
  INV_X1 U36868 ( .A(n37575), .ZN(n2914) );
  OAI22_X1 U36869 ( .A1(n37582), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[24][2] ), .B2(n37581), .ZN(n37576) );
  INV_X1 U36870 ( .A(n37576), .ZN(n2913) );
  OAI22_X1 U36871 ( .A1(n37582), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[24][3] ), .B2(n37581), .ZN(n37577) );
  INV_X1 U36872 ( .A(n37577), .ZN(n2912) );
  OAI22_X1 U36873 ( .A1(n37582), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[24][4] ), .B2(n37581), .ZN(n37578) );
  INV_X1 U36874 ( .A(n37578), .ZN(n2911) );
  OAI22_X1 U36875 ( .A1(n37582), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[24][5] ), .B2(n37581), .ZN(n37579) );
  INV_X1 U36876 ( .A(n37579), .ZN(n2910) );
  OAI22_X1 U36877 ( .A1(n37582), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[24][6] ), .B2(n37581), .ZN(n37580) );
  INV_X1 U36878 ( .A(n37580), .ZN(n2909) );
  OAI22_X1 U36879 ( .A1(n37582), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[24][7] ), .B2(n37581), .ZN(n37583) );
  INV_X1 U36880 ( .A(n37583), .ZN(n2908) );
  NOR2_X1 U36881 ( .A1(n37584), .A2(n37639), .ZN(n37592) );
  INV_X1 U36882 ( .A(n37592), .ZN(n37593) );
  OAI22_X1 U36883 ( .A1(n37593), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[25][0] ), .B2(n37592), .ZN(n37585) );
  INV_X1 U36884 ( .A(n37585), .ZN(n2907) );
  OAI22_X1 U36885 ( .A1(n37593), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[25][1] ), .B2(n37592), .ZN(n37586) );
  INV_X1 U36886 ( .A(n37586), .ZN(n2906) );
  OAI22_X1 U36887 ( .A1(n37593), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[25][2] ), .B2(n37592), .ZN(n37587) );
  INV_X1 U36888 ( .A(n37587), .ZN(n2905) );
  OAI22_X1 U36889 ( .A1(n37593), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[25][3] ), .B2(n37592), .ZN(n37588) );
  INV_X1 U36890 ( .A(n37588), .ZN(n2904) );
  OAI22_X1 U36891 ( .A1(n37593), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[25][4] ), .B2(n37592), .ZN(n37589) );
  INV_X1 U36892 ( .A(n37589), .ZN(n2903) );
  OAI22_X1 U36893 ( .A1(n37593), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[25][5] ), .B2(n37592), .ZN(n37590) );
  INV_X1 U36894 ( .A(n37590), .ZN(n2902) );
  OAI22_X1 U36895 ( .A1(n37593), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[25][6] ), .B2(n37592), .ZN(n37591) );
  INV_X1 U36896 ( .A(n37591), .ZN(n2901) );
  OAI22_X1 U36897 ( .A1(n37593), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[25][7] ), .B2(n37592), .ZN(n37594) );
  INV_X1 U36898 ( .A(n37594), .ZN(n2900) );
  NOR2_X1 U36899 ( .A1(n37595), .A2(n37639), .ZN(n37603) );
  INV_X1 U36900 ( .A(n37603), .ZN(n37604) );
  OAI22_X1 U36901 ( .A1(n37604), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[26][0] ), .B2(n37603), .ZN(n37596) );
  INV_X1 U36902 ( .A(n37596), .ZN(n2899) );
  OAI22_X1 U36903 ( .A1(n37604), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[26][1] ), .B2(n37603), .ZN(n37597) );
  INV_X1 U36904 ( .A(n37597), .ZN(n2898) );
  OAI22_X1 U36905 ( .A1(n37604), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[26][2] ), .B2(n37603), .ZN(n37598) );
  INV_X1 U36906 ( .A(n37598), .ZN(n2897) );
  OAI22_X1 U36907 ( .A1(n37604), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[26][3] ), .B2(n37603), .ZN(n37599) );
  INV_X1 U36908 ( .A(n37599), .ZN(n2896) );
  OAI22_X1 U36909 ( .A1(n37604), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[26][4] ), .B2(n37603), .ZN(n37600) );
  INV_X1 U36910 ( .A(n37600), .ZN(n2895) );
  OAI22_X1 U36911 ( .A1(n37604), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[26][5] ), .B2(n37603), .ZN(n37601) );
  INV_X1 U36912 ( .A(n37601), .ZN(n2894) );
  OAI22_X1 U36913 ( .A1(n37604), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[26][6] ), .B2(n37603), .ZN(n37602) );
  INV_X1 U36914 ( .A(n37602), .ZN(n2893) );
  OAI22_X1 U36915 ( .A1(n37604), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[26][7] ), .B2(n37603), .ZN(n37605) );
  INV_X1 U36916 ( .A(n37605), .ZN(n2892) );
  NOR2_X1 U36917 ( .A1(n37606), .A2(n37639), .ZN(n37614) );
  INV_X1 U36918 ( .A(n37614), .ZN(n37615) );
  OAI22_X1 U36919 ( .A1(n37615), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[27][0] ), .B2(n37614), .ZN(n37607) );
  INV_X1 U36920 ( .A(n37607), .ZN(n2891) );
  OAI22_X1 U36921 ( .A1(n37615), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[27][1] ), .B2(n37614), .ZN(n37608) );
  INV_X1 U36922 ( .A(n37608), .ZN(n2890) );
  OAI22_X1 U36923 ( .A1(n37615), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[27][2] ), .B2(n37614), .ZN(n37609) );
  INV_X1 U36924 ( .A(n37609), .ZN(n2889) );
  OAI22_X1 U36925 ( .A1(n37615), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[27][3] ), .B2(n37614), .ZN(n37610) );
  INV_X1 U36926 ( .A(n37610), .ZN(n2888) );
  OAI22_X1 U36927 ( .A1(n37615), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[27][4] ), .B2(n37614), .ZN(n37611) );
  INV_X1 U36928 ( .A(n37611), .ZN(n2887) );
  OAI22_X1 U36929 ( .A1(n37615), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[27][5] ), .B2(n37614), .ZN(n37612) );
  INV_X1 U36930 ( .A(n37612), .ZN(n2886) );
  OAI22_X1 U36931 ( .A1(n37615), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[27][6] ), .B2(n37614), .ZN(n37613) );
  INV_X1 U36932 ( .A(n37613), .ZN(n2885) );
  OAI22_X1 U36933 ( .A1(n37615), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[27][7] ), .B2(n37614), .ZN(n37616) );
  INV_X1 U36934 ( .A(n37616), .ZN(n2884) );
  NOR2_X1 U36935 ( .A1(n37617), .A2(n37639), .ZN(n37625) );
  INV_X1 U36936 ( .A(n37625), .ZN(n37626) );
  OAI22_X1 U36937 ( .A1(n37626), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[28][0] ), .B2(n37625), .ZN(n37618) );
  INV_X1 U36938 ( .A(n37618), .ZN(n2883) );
  OAI22_X1 U36939 ( .A1(n37626), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[28][1] ), .B2(n37625), .ZN(n37619) );
  INV_X1 U36940 ( .A(n37619), .ZN(n2882) );
  OAI22_X1 U36941 ( .A1(n37626), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[28][2] ), .B2(n37625), .ZN(n37620) );
  INV_X1 U36942 ( .A(n37620), .ZN(n2881) );
  OAI22_X1 U36943 ( .A1(n37626), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[28][3] ), .B2(n37625), .ZN(n37621) );
  INV_X1 U36944 ( .A(n37621), .ZN(n2880) );
  OAI22_X1 U36945 ( .A1(n37626), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[28][4] ), .B2(n37625), .ZN(n37622) );
  INV_X1 U36946 ( .A(n37622), .ZN(n2879) );
  OAI22_X1 U36947 ( .A1(n37626), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[28][5] ), .B2(n37625), .ZN(n37623) );
  INV_X1 U36948 ( .A(n37623), .ZN(n2878) );
  OAI22_X1 U36949 ( .A1(n37626), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[28][6] ), .B2(n37625), .ZN(n37624) );
  INV_X1 U36950 ( .A(n37624), .ZN(n2877) );
  OAI22_X1 U36951 ( .A1(n37626), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[28][7] ), .B2(n37625), .ZN(n37627) );
  INV_X1 U36952 ( .A(n37627), .ZN(n2876) );
  NOR2_X1 U36953 ( .A1(n37628), .A2(n37639), .ZN(n37636) );
  INV_X1 U36954 ( .A(n37636), .ZN(n37637) );
  OAI22_X1 U36955 ( .A1(n37637), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[29][0] ), .B2(n37636), .ZN(n37629) );
  INV_X1 U36956 ( .A(n37629), .ZN(n2875) );
  OAI22_X1 U36957 ( .A1(n37637), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[29][1] ), .B2(n37636), .ZN(n37630) );
  INV_X1 U36958 ( .A(n37630), .ZN(n2874) );
  OAI22_X1 U36959 ( .A1(n37637), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[29][2] ), .B2(n37636), .ZN(n37631) );
  INV_X1 U36960 ( .A(n37631), .ZN(n2873) );
  OAI22_X1 U36961 ( .A1(n37637), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[29][3] ), .B2(n37636), .ZN(n37632) );
  INV_X1 U36962 ( .A(n37632), .ZN(n2872) );
  OAI22_X1 U36963 ( .A1(n37637), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[29][4] ), .B2(n37636), .ZN(n37633) );
  INV_X1 U36964 ( .A(n37633), .ZN(n2871) );
  OAI22_X1 U36965 ( .A1(n37637), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[29][5] ), .B2(n37636), .ZN(n37634) );
  INV_X1 U36966 ( .A(n37634), .ZN(n2870) );
  OAI22_X1 U36967 ( .A1(n37637), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[29][6] ), .B2(n37636), .ZN(n37635) );
  INV_X1 U36968 ( .A(n37635), .ZN(n2869) );
  OAI22_X1 U36969 ( .A1(n37637), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[29][7] ), .B2(n37636), .ZN(n37638) );
  INV_X1 U36970 ( .A(n37638), .ZN(n2868) );
  NOR2_X1 U36971 ( .A1(n37640), .A2(n37639), .ZN(n37648) );
  INV_X1 U36972 ( .A(n37648), .ZN(n37649) );
  OAI22_X1 U36973 ( .A1(n37649), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[30][0] ), .B2(n37648), .ZN(n37641) );
  INV_X1 U36974 ( .A(n37641), .ZN(n2867) );
  OAI22_X1 U36975 ( .A1(n37649), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[30][1] ), .B2(n37648), .ZN(n37642) );
  INV_X1 U36976 ( .A(n37642), .ZN(n2866) );
  OAI22_X1 U36977 ( .A1(n37649), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[30][2] ), .B2(n37648), .ZN(n37643) );
  INV_X1 U36978 ( .A(n37643), .ZN(n2865) );
  OAI22_X1 U36979 ( .A1(n37649), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[30][3] ), .B2(n37648), .ZN(n37644) );
  INV_X1 U36980 ( .A(n37644), .ZN(n2864) );
  OAI22_X1 U36981 ( .A1(n37649), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[30][4] ), .B2(n37648), .ZN(n37645) );
  INV_X1 U36982 ( .A(n37645), .ZN(n2863) );
  OAI22_X1 U36983 ( .A1(n37649), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[30][5] ), .B2(n37648), .ZN(n37646) );
  INV_X1 U36984 ( .A(n37646), .ZN(n2862) );
  OAI22_X1 U36985 ( .A1(n37649), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[30][6] ), .B2(n37648), .ZN(n37647) );
  INV_X1 U36986 ( .A(n37647), .ZN(n2861) );
  OAI22_X1 U36987 ( .A1(n37649), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[30][7] ), .B2(n37648), .ZN(n37650) );
  INV_X1 U36988 ( .A(n37650), .ZN(n2860) );
  OAI22_X1 U36989 ( .A1(n37659), .A2(s_data_in_f[0]), .B1(
        \fmem_inst/mem[31][0] ), .B2(n37658), .ZN(n37651) );
  INV_X1 U36990 ( .A(n37651), .ZN(n2859) );
  OAI22_X1 U36991 ( .A1(n37659), .A2(s_data_in_f[1]), .B1(
        \fmem_inst/mem[31][1] ), .B2(n37658), .ZN(n37652) );
  INV_X1 U36992 ( .A(n37652), .ZN(n2858) );
  OAI22_X1 U36993 ( .A1(n37659), .A2(s_data_in_f[2]), .B1(
        \fmem_inst/mem[31][2] ), .B2(n37658), .ZN(n37653) );
  INV_X1 U36994 ( .A(n37653), .ZN(n2857) );
  OAI22_X1 U36995 ( .A1(n37659), .A2(s_data_in_f[3]), .B1(
        \fmem_inst/mem[31][3] ), .B2(n37658), .ZN(n37654) );
  INV_X1 U36996 ( .A(n37654), .ZN(n2856) );
  OAI22_X1 U36997 ( .A1(n37659), .A2(s_data_in_f[4]), .B1(
        \fmem_inst/mem[31][4] ), .B2(n37658), .ZN(n37655) );
  INV_X1 U36998 ( .A(n37655), .ZN(n2855) );
  OAI22_X1 U36999 ( .A1(n37659), .A2(s_data_in_f[5]), .B1(
        \fmem_inst/mem[31][5] ), .B2(n37658), .ZN(n37656) );
  INV_X1 U37000 ( .A(n37656), .ZN(n2854) );
  OAI22_X1 U37001 ( .A1(n37659), .A2(s_data_in_f[6]), .B1(
        \fmem_inst/mem[31][6] ), .B2(n37658), .ZN(n37657) );
  INV_X1 U37002 ( .A(n37657), .ZN(n2853) );
  OAI22_X1 U37003 ( .A1(n37659), .A2(s_data_in_f[7]), .B1(
        \fmem_inst/mem[31][7] ), .B2(n37658), .ZN(n37660) );
  INV_X1 U37004 ( .A(n37660), .ZN(n2852) );
  NAND2_X1 U37005 ( .A1(xmem_addr[0]), .A2(xmem_addr[1]), .ZN(n37705) );
  NOR2_X1 U37006 ( .A1(n37705), .A2(n38999), .ZN(n37664) );
  INV_X1 U37007 ( .A(n37664), .ZN(n37663) );
  NOR2_X1 U37008 ( .A1(n39044), .A2(n37663), .ZN(n37666) );
  INV_X1 U37009 ( .A(n37666), .ZN(n38803) );
  NAND2_X1 U37010 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n37674) );
  NOR2_X1 U37011 ( .A1(n37674), .A2(n39042), .ZN(n38489) );
  NAND3_X1 U37012 ( .A1(xmem_addr[6]), .A2(xmem_addr[5]), .A3(n38489), .ZN(
        n38969) );
  NOR2_X1 U37013 ( .A1(n38803), .A2(n38969), .ZN(n38987) );
  OAI21_X1 U37014 ( .B1(n38987), .B2(n39051), .A(n37669), .ZN(n2851) );
  NAND2_X1 U37015 ( .A1(n37669), .A2(n37674), .ZN(n37668) );
  OR2_X1 U37016 ( .A1(n37661), .A2(n37674), .ZN(n37672) );
  AOI22_X1 U37017 ( .A1(xmem_addr[0]), .A2(n37668), .B1(n37672), .B2(n39048), 
        .ZN(n2850) );
  NOR2_X1 U37018 ( .A1(xmem_addr[0]), .A2(n39049), .ZN(n37823) );
  NOR2_X1 U37019 ( .A1(xmem_addr[1]), .A2(n39048), .ZN(n37811) );
  NOR2_X1 U37020 ( .A1(n37823), .A2(n37811), .ZN(n37662) );
  OAI22_X1 U37021 ( .A1(n37662), .A2(n37672), .B1(n37668), .B2(n39049), .ZN(
        n2849) );
  OAI21_X1 U37022 ( .B1(n37674), .B2(n37663), .A(n37669), .ZN(n37665) );
  AOI221_X1 U37023 ( .B1(n37705), .B2(n38999), .C1(n37672), .C2(n38999), .A(
        n37665), .ZN(n2848) );
  NAND2_X1 U37024 ( .A1(n37664), .A2(n39044), .ZN(n38891) );
  OAI22_X1 U37025 ( .A1(n37665), .A2(n39044), .B1(n37672), .B2(n38891), .ZN(
        n2847) );
  NAND2_X1 U37026 ( .A1(n37666), .A2(xmem_addr[4]), .ZN(n37671) );
  OAI21_X1 U37027 ( .B1(n37666), .B2(xmem_addr[4]), .A(n37671), .ZN(n37667) );
  OAI22_X1 U37028 ( .A1(n37668), .A2(n39042), .B1(n37672), .B2(n37667), .ZN(
        n2846) );
  OR3_X1 U37029 ( .A1(n37674), .A2(n37671), .A3(n38998), .ZN(n37670) );
  NAND2_X1 U37030 ( .A1(n37670), .A2(n37669), .ZN(n37673) );
  AOI221_X1 U37031 ( .B1(n37672), .B2(n38998), .C1(n37671), .C2(n38998), .A(
        n37673), .ZN(n2845) );
  NAND3_X1 U37032 ( .A1(n39043), .A2(xmem_addr[5]), .A3(n38489), .ZN(n38307)
         );
  NOR2_X1 U37033 ( .A1(n38803), .A2(n38307), .ZN(n38325) );
  INV_X1 U37034 ( .A(n38325), .ZN(n38326) );
  OAI22_X1 U37035 ( .A1(n37673), .A2(n39043), .B1(n37672), .B2(n38326), .ZN(
        n2844) );
  NOR2_X1 U37036 ( .A1(xmem_addr[0]), .A2(xmem_addr[1]), .ZN(n37800) );
  NOR2_X1 U37037 ( .A1(xmem_addr[3]), .A2(xmem_addr[2]), .ZN(n37706) );
  NAND2_X1 U37038 ( .A1(n37800), .A2(n37706), .ZN(n38814) );
  NOR2_X1 U37039 ( .A1(xmem_addr[4]), .A2(n37674), .ZN(n38651) );
  NAND3_X1 U37040 ( .A1(n38651), .A2(n39043), .A3(n38998), .ZN(n37834) );
  NOR2_X1 U37041 ( .A1(n38814), .A2(n37834), .ZN(n37682) );
  INV_X1 U37042 ( .A(n37682), .ZN(n37683) );
  OAI22_X1 U37043 ( .A1(n37683), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[0][0] ), .B2(n37682), .ZN(n37675) );
  INV_X1 U37044 ( .A(n37675), .ZN(n2843) );
  OAI22_X1 U37045 ( .A1(n37683), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[0][1] ), .B2(n37682), .ZN(n37676) );
  INV_X1 U37046 ( .A(n37676), .ZN(n2842) );
  OAI22_X1 U37047 ( .A1(n37683), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[0][2] ), .B2(n37682), .ZN(n37677) );
  INV_X1 U37048 ( .A(n37677), .ZN(n2841) );
  OAI22_X1 U37049 ( .A1(n37683), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[0][3] ), .B2(n37682), .ZN(n37678) );
  INV_X1 U37050 ( .A(n37678), .ZN(n2840) );
  OAI22_X1 U37051 ( .A1(n37683), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[0][4] ), .B2(n37682), .ZN(n37679) );
  INV_X1 U37052 ( .A(n37679), .ZN(n2839) );
  OAI22_X1 U37053 ( .A1(n37683), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[0][5] ), .B2(n37682), .ZN(n37680) );
  INV_X1 U37054 ( .A(n37680), .ZN(n2838) );
  OAI22_X1 U37055 ( .A1(n37683), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[0][6] ), .B2(n37682), .ZN(n37681) );
  INV_X1 U37056 ( .A(n37681), .ZN(n2837) );
  OAI22_X1 U37057 ( .A1(n37683), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[0][7] ), .B2(n37682), .ZN(n37684) );
  INV_X1 U37058 ( .A(n37684), .ZN(n2836) );
  NAND2_X1 U37059 ( .A1(n37811), .A2(n37706), .ZN(n38825) );
  NOR2_X1 U37060 ( .A1(n37834), .A2(n38825), .ZN(n37692) );
  INV_X1 U37061 ( .A(n37692), .ZN(n37693) );
  OAI22_X1 U37062 ( .A1(n37693), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[1][0] ), .B2(n37692), .ZN(n37685) );
  INV_X1 U37063 ( .A(n37685), .ZN(n2835) );
  OAI22_X1 U37064 ( .A1(n37693), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[1][1] ), .B2(n37692), .ZN(n37686) );
  INV_X1 U37065 ( .A(n37686), .ZN(n2834) );
  OAI22_X1 U37066 ( .A1(n37693), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[1][2] ), .B2(n37692), .ZN(n37687) );
  INV_X1 U37067 ( .A(n37687), .ZN(n2833) );
  OAI22_X1 U37068 ( .A1(n37693), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[1][3] ), .B2(n37692), .ZN(n37688) );
  INV_X1 U37069 ( .A(n37688), .ZN(n2832) );
  OAI22_X1 U37070 ( .A1(n37693), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[1][4] ), .B2(n37692), .ZN(n37689) );
  INV_X1 U37071 ( .A(n37689), .ZN(n2831) );
  OAI22_X1 U37072 ( .A1(n37693), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[1][5] ), .B2(n37692), .ZN(n37690) );
  INV_X1 U37073 ( .A(n37690), .ZN(n2830) );
  OAI22_X1 U37074 ( .A1(n37693), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[1][6] ), .B2(n37692), .ZN(n37691) );
  INV_X1 U37075 ( .A(n37691), .ZN(n2829) );
  OAI22_X1 U37076 ( .A1(n37693), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[1][7] ), .B2(n37692), .ZN(n37694) );
  INV_X1 U37077 ( .A(n37694), .ZN(n2828) );
  NAND2_X1 U37078 ( .A1(n37823), .A2(n37706), .ZN(n38836) );
  NOR2_X1 U37079 ( .A1(n37834), .A2(n38836), .ZN(n37702) );
  INV_X1 U37080 ( .A(n37702), .ZN(n37703) );
  OAI22_X1 U37081 ( .A1(n37703), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[2][0] ), .B2(n37702), .ZN(n37695) );
  INV_X1 U37082 ( .A(n37695), .ZN(n2827) );
  OAI22_X1 U37083 ( .A1(n37703), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[2][1] ), .B2(n37702), .ZN(n37696) );
  INV_X1 U37084 ( .A(n37696), .ZN(n2826) );
  OAI22_X1 U37085 ( .A1(n37703), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[2][2] ), .B2(n37702), .ZN(n37697) );
  INV_X1 U37086 ( .A(n37697), .ZN(n2825) );
  OAI22_X1 U37087 ( .A1(n37703), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[2][3] ), .B2(n37702), .ZN(n37698) );
  INV_X1 U37088 ( .A(n37698), .ZN(n2824) );
  OAI22_X1 U37089 ( .A1(n37703), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[2][4] ), .B2(n37702), .ZN(n37699) );
  INV_X1 U37090 ( .A(n37699), .ZN(n2823) );
  OAI22_X1 U37091 ( .A1(n37703), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[2][5] ), .B2(n37702), .ZN(n37700) );
  INV_X1 U37092 ( .A(n37700), .ZN(n2822) );
  OAI22_X1 U37093 ( .A1(n37703), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[2][6] ), .B2(n37702), .ZN(n37701) );
  INV_X1 U37094 ( .A(n37701), .ZN(n2821) );
  OAI22_X1 U37095 ( .A1(n37703), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[2][7] ), .B2(n37702), .ZN(n37704) );
  INV_X1 U37096 ( .A(n37704), .ZN(n2820) );
  INV_X1 U37097 ( .A(n37705), .ZN(n37789) );
  NAND2_X1 U37098 ( .A1(n37789), .A2(n37706), .ZN(n38847) );
  NOR2_X1 U37099 ( .A1(n37834), .A2(n38847), .ZN(n37714) );
  INV_X1 U37100 ( .A(n37714), .ZN(n37715) );
  OAI22_X1 U37101 ( .A1(n37715), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[3][0] ), .B2(n37714), .ZN(n37707) );
  INV_X1 U37102 ( .A(n37707), .ZN(n2819) );
  OAI22_X1 U37103 ( .A1(n37715), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[3][1] ), .B2(n37714), .ZN(n37708) );
  INV_X1 U37104 ( .A(n37708), .ZN(n2818) );
  OAI22_X1 U37105 ( .A1(n37715), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[3][2] ), .B2(n37714), .ZN(n37709) );
  INV_X1 U37106 ( .A(n37709), .ZN(n2817) );
  OAI22_X1 U37107 ( .A1(n37715), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[3][3] ), .B2(n37714), .ZN(n37710) );
  INV_X1 U37108 ( .A(n37710), .ZN(n2816) );
  OAI22_X1 U37109 ( .A1(n37715), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[3][4] ), .B2(n37714), .ZN(n37711) );
  INV_X1 U37110 ( .A(n37711), .ZN(n2815) );
  OAI22_X1 U37111 ( .A1(n37715), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[3][5] ), .B2(n37714), .ZN(n37712) );
  INV_X1 U37112 ( .A(n37712), .ZN(n2814) );
  OAI22_X1 U37113 ( .A1(n37715), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[3][6] ), .B2(n37714), .ZN(n37713) );
  INV_X1 U37114 ( .A(n37713), .ZN(n2813) );
  OAI22_X1 U37115 ( .A1(n37715), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[3][7] ), .B2(n37714), .ZN(n37716) );
  INV_X1 U37116 ( .A(n37716), .ZN(n2812) );
  NOR2_X1 U37117 ( .A1(xmem_addr[3]), .A2(n38999), .ZN(n37737) );
  NAND2_X1 U37118 ( .A1(n37800), .A2(n37737), .ZN(n38858) );
  NOR2_X1 U37119 ( .A1(n37834), .A2(n38858), .ZN(n37724) );
  INV_X1 U37120 ( .A(n37724), .ZN(n37725) );
  OAI22_X1 U37121 ( .A1(n37725), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[4][0] ), .B2(n37724), .ZN(n37717) );
  INV_X1 U37122 ( .A(n37717), .ZN(n2811) );
  OAI22_X1 U37123 ( .A1(n37725), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[4][1] ), .B2(n37724), .ZN(n37718) );
  INV_X1 U37124 ( .A(n37718), .ZN(n2810) );
  OAI22_X1 U37125 ( .A1(n37725), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[4][2] ), .B2(n37724), .ZN(n37719) );
  INV_X1 U37126 ( .A(n37719), .ZN(n2809) );
  OAI22_X1 U37127 ( .A1(n37725), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[4][3] ), .B2(n37724), .ZN(n37720) );
  INV_X1 U37128 ( .A(n37720), .ZN(n2808) );
  OAI22_X1 U37129 ( .A1(n37725), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[4][4] ), .B2(n37724), .ZN(n37721) );
  INV_X1 U37130 ( .A(n37721), .ZN(n2807) );
  OAI22_X1 U37131 ( .A1(n37725), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[4][5] ), .B2(n37724), .ZN(n37722) );
  INV_X1 U37132 ( .A(n37722), .ZN(n2806) );
  OAI22_X1 U37133 ( .A1(n37725), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[4][6] ), .B2(n37724), .ZN(n37723) );
  INV_X1 U37134 ( .A(n37723), .ZN(n2805) );
  OAI22_X1 U37135 ( .A1(n37725), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[4][7] ), .B2(n37724), .ZN(n37726) );
  INV_X1 U37136 ( .A(n37726), .ZN(n2804) );
  NAND2_X1 U37137 ( .A1(n37811), .A2(n37737), .ZN(n38869) );
  NOR2_X1 U37138 ( .A1(n37834), .A2(n38869), .ZN(n37734) );
  INV_X1 U37139 ( .A(n37734), .ZN(n37735) );
  OAI22_X1 U37140 ( .A1(n37735), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[5][0] ), .B2(n37734), .ZN(n37727) );
  INV_X1 U37141 ( .A(n37727), .ZN(n2803) );
  OAI22_X1 U37142 ( .A1(n37735), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[5][1] ), .B2(n37734), .ZN(n37728) );
  INV_X1 U37143 ( .A(n37728), .ZN(n2802) );
  OAI22_X1 U37144 ( .A1(n37735), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[5][2] ), .B2(n37734), .ZN(n37729) );
  INV_X1 U37145 ( .A(n37729), .ZN(n2801) );
  OAI22_X1 U37146 ( .A1(n37735), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[5][3] ), .B2(n37734), .ZN(n37730) );
  INV_X1 U37147 ( .A(n37730), .ZN(n2800) );
  OAI22_X1 U37148 ( .A1(n37735), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[5][4] ), .B2(n37734), .ZN(n37731) );
  INV_X1 U37149 ( .A(n37731), .ZN(n2799) );
  OAI22_X1 U37150 ( .A1(n37735), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[5][5] ), .B2(n37734), .ZN(n37732) );
  INV_X1 U37151 ( .A(n37732), .ZN(n2798) );
  OAI22_X1 U37152 ( .A1(n37735), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[5][6] ), .B2(n37734), .ZN(n37733) );
  INV_X1 U37153 ( .A(n37733), .ZN(n2797) );
  OAI22_X1 U37154 ( .A1(n37735), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[5][7] ), .B2(n37734), .ZN(n37736) );
  INV_X1 U37155 ( .A(n37736), .ZN(n2796) );
  NAND2_X1 U37156 ( .A1(n37823), .A2(n37737), .ZN(n38880) );
  NOR2_X1 U37157 ( .A1(n37834), .A2(n38880), .ZN(n37745) );
  INV_X1 U37158 ( .A(n37745), .ZN(n37746) );
  OAI22_X1 U37159 ( .A1(n37746), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[6][0] ), .B2(n37745), .ZN(n37738) );
  INV_X1 U37160 ( .A(n37738), .ZN(n2795) );
  OAI22_X1 U37161 ( .A1(n37746), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[6][1] ), .B2(n37745), .ZN(n37739) );
  INV_X1 U37162 ( .A(n37739), .ZN(n2794) );
  OAI22_X1 U37163 ( .A1(n37746), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[6][2] ), .B2(n37745), .ZN(n37740) );
  INV_X1 U37164 ( .A(n37740), .ZN(n2793) );
  OAI22_X1 U37165 ( .A1(n37746), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[6][3] ), .B2(n37745), .ZN(n37741) );
  INV_X1 U37166 ( .A(n37741), .ZN(n2792) );
  OAI22_X1 U37167 ( .A1(n37746), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[6][4] ), .B2(n37745), .ZN(n37742) );
  INV_X1 U37168 ( .A(n37742), .ZN(n2791) );
  OAI22_X1 U37169 ( .A1(n37746), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[6][5] ), .B2(n37745), .ZN(n37743) );
  INV_X1 U37170 ( .A(n37743), .ZN(n2790) );
  OAI22_X1 U37171 ( .A1(n37746), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[6][6] ), .B2(n37745), .ZN(n37744) );
  INV_X1 U37172 ( .A(n37744), .ZN(n2789) );
  OAI22_X1 U37173 ( .A1(n37746), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[6][7] ), .B2(n37745), .ZN(n37747) );
  INV_X1 U37174 ( .A(n37747), .ZN(n2788) );
  NOR2_X1 U37175 ( .A1(n38891), .A2(n37834), .ZN(n37755) );
  INV_X1 U37176 ( .A(n37755), .ZN(n37756) );
  OAI22_X1 U37177 ( .A1(n37756), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[7][0] ), .B2(n37755), .ZN(n37748) );
  INV_X1 U37178 ( .A(n37748), .ZN(n2787) );
  OAI22_X1 U37179 ( .A1(n37756), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[7][1] ), .B2(n37755), .ZN(n37749) );
  INV_X1 U37180 ( .A(n37749), .ZN(n2786) );
  OAI22_X1 U37181 ( .A1(n37756), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[7][2] ), .B2(n37755), .ZN(n37750) );
  INV_X1 U37182 ( .A(n37750), .ZN(n2785) );
  OAI22_X1 U37183 ( .A1(n37756), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[7][3] ), .B2(n37755), .ZN(n37751) );
  INV_X1 U37184 ( .A(n37751), .ZN(n2784) );
  OAI22_X1 U37185 ( .A1(n37756), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[7][4] ), .B2(n37755), .ZN(n37752) );
  INV_X1 U37186 ( .A(n37752), .ZN(n2783) );
  OAI22_X1 U37187 ( .A1(n37756), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[7][5] ), .B2(n37755), .ZN(n37753) );
  INV_X1 U37188 ( .A(n37753), .ZN(n2782) );
  OAI22_X1 U37189 ( .A1(n37756), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[7][6] ), .B2(n37755), .ZN(n37754) );
  INV_X1 U37190 ( .A(n37754), .ZN(n2781) );
  OAI22_X1 U37191 ( .A1(n37756), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[7][7] ), .B2(n37755), .ZN(n37757) );
  INV_X1 U37192 ( .A(n37757), .ZN(n2780) );
  NOR2_X1 U37193 ( .A1(xmem_addr[2]), .A2(n39044), .ZN(n37788) );
  NAND2_X1 U37194 ( .A1(n37800), .A2(n37788), .ZN(n38902) );
  NOR2_X1 U37195 ( .A1(n37834), .A2(n38902), .ZN(n37765) );
  INV_X1 U37196 ( .A(n37765), .ZN(n37766) );
  OAI22_X1 U37197 ( .A1(n37766), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[8][0] ), .B2(n37765), .ZN(n37758) );
  INV_X1 U37198 ( .A(n37758), .ZN(n2779) );
  OAI22_X1 U37199 ( .A1(n37766), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[8][1] ), .B2(n37765), .ZN(n37759) );
  INV_X1 U37200 ( .A(n37759), .ZN(n2778) );
  OAI22_X1 U37201 ( .A1(n37766), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[8][2] ), .B2(n37765), .ZN(n37760) );
  INV_X1 U37202 ( .A(n37760), .ZN(n2777) );
  OAI22_X1 U37203 ( .A1(n37766), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[8][3] ), .B2(n37765), .ZN(n37761) );
  INV_X1 U37204 ( .A(n37761), .ZN(n2776) );
  OAI22_X1 U37205 ( .A1(n37766), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[8][4] ), .B2(n37765), .ZN(n37762) );
  INV_X1 U37206 ( .A(n37762), .ZN(n2775) );
  OAI22_X1 U37207 ( .A1(n37766), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[8][5] ), .B2(n37765), .ZN(n37763) );
  INV_X1 U37208 ( .A(n37763), .ZN(n2774) );
  OAI22_X1 U37209 ( .A1(n37766), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[8][6] ), .B2(n37765), .ZN(n37764) );
  INV_X1 U37210 ( .A(n37764), .ZN(n2773) );
  OAI22_X1 U37211 ( .A1(n37766), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[8][7] ), .B2(n37765), .ZN(n37767) );
  INV_X1 U37212 ( .A(n37767), .ZN(n2772) );
  NAND2_X1 U37213 ( .A1(n37811), .A2(n37788), .ZN(n38913) );
  NOR2_X1 U37214 ( .A1(n37834), .A2(n38913), .ZN(n37775) );
  INV_X1 U37215 ( .A(n37775), .ZN(n37776) );
  OAI22_X1 U37216 ( .A1(n37776), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[9][0] ), .B2(n37775), .ZN(n37768) );
  INV_X1 U37217 ( .A(n37768), .ZN(n2771) );
  OAI22_X1 U37218 ( .A1(n37776), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[9][1] ), .B2(n37775), .ZN(n37769) );
  INV_X1 U37219 ( .A(n37769), .ZN(n2770) );
  OAI22_X1 U37220 ( .A1(n37776), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[9][2] ), .B2(n37775), .ZN(n37770) );
  INV_X1 U37221 ( .A(n37770), .ZN(n2769) );
  OAI22_X1 U37222 ( .A1(n37776), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[9][3] ), .B2(n37775), .ZN(n37771) );
  INV_X1 U37223 ( .A(n37771), .ZN(n2768) );
  OAI22_X1 U37224 ( .A1(n37776), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[9][4] ), .B2(n37775), .ZN(n37772) );
  INV_X1 U37225 ( .A(n37772), .ZN(n2767) );
  OAI22_X1 U37226 ( .A1(n37776), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[9][5] ), .B2(n37775), .ZN(n37773) );
  INV_X1 U37227 ( .A(n37773), .ZN(n2766) );
  OAI22_X1 U37228 ( .A1(n37776), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[9][6] ), .B2(n37775), .ZN(n37774) );
  INV_X1 U37229 ( .A(n37774), .ZN(n2765) );
  OAI22_X1 U37230 ( .A1(n37776), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[9][7] ), .B2(n37775), .ZN(n37777) );
  INV_X1 U37231 ( .A(n37777), .ZN(n2764) );
  NAND2_X1 U37232 ( .A1(n37823), .A2(n37788), .ZN(n38924) );
  NOR2_X1 U37233 ( .A1(n37834), .A2(n38924), .ZN(n37785) );
  INV_X1 U37234 ( .A(n37785), .ZN(n37786) );
  OAI22_X1 U37235 ( .A1(n37786), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[10][0] ), .B2(n37785), .ZN(n37778) );
  INV_X1 U37236 ( .A(n37778), .ZN(n2763) );
  OAI22_X1 U37237 ( .A1(n37786), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[10][1] ), .B2(n37785), .ZN(n37779) );
  INV_X1 U37238 ( .A(n37779), .ZN(n2762) );
  OAI22_X1 U37239 ( .A1(n37786), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[10][2] ), .B2(n37785), .ZN(n37780) );
  INV_X1 U37240 ( .A(n37780), .ZN(n2761) );
  OAI22_X1 U37241 ( .A1(n37786), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[10][3] ), .B2(n37785), .ZN(n37781) );
  INV_X1 U37242 ( .A(n37781), .ZN(n2760) );
  OAI22_X1 U37243 ( .A1(n37786), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[10][4] ), .B2(n37785), .ZN(n37782) );
  INV_X1 U37244 ( .A(n37782), .ZN(n2759) );
  OAI22_X1 U37245 ( .A1(n37786), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[10][5] ), .B2(n37785), .ZN(n37783) );
  INV_X1 U37246 ( .A(n37783), .ZN(n2758) );
  OAI22_X1 U37247 ( .A1(n37786), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[10][6] ), .B2(n37785), .ZN(n37784) );
  INV_X1 U37248 ( .A(n37784), .ZN(n2757) );
  OAI22_X1 U37249 ( .A1(n37786), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[10][7] ), .B2(n37785), .ZN(n37787) );
  INV_X1 U37250 ( .A(n37787), .ZN(n2756) );
  NAND2_X1 U37251 ( .A1(n37789), .A2(n37788), .ZN(n38935) );
  NOR2_X1 U37252 ( .A1(n37834), .A2(n38935), .ZN(n37797) );
  INV_X1 U37253 ( .A(n37797), .ZN(n37798) );
  OAI22_X1 U37254 ( .A1(n37798), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[11][0] ), .B2(n37797), .ZN(n37790) );
  INV_X1 U37255 ( .A(n37790), .ZN(n2755) );
  OAI22_X1 U37256 ( .A1(n37798), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[11][1] ), .B2(n37797), .ZN(n37791) );
  INV_X1 U37257 ( .A(n37791), .ZN(n2754) );
  OAI22_X1 U37258 ( .A1(n37798), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[11][2] ), .B2(n37797), .ZN(n37792) );
  INV_X1 U37259 ( .A(n37792), .ZN(n2753) );
  OAI22_X1 U37260 ( .A1(n37798), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[11][3] ), .B2(n37797), .ZN(n37793) );
  INV_X1 U37261 ( .A(n37793), .ZN(n2752) );
  OAI22_X1 U37262 ( .A1(n37798), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[11][4] ), .B2(n37797), .ZN(n37794) );
  INV_X1 U37263 ( .A(n37794), .ZN(n2751) );
  OAI22_X1 U37264 ( .A1(n37798), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[11][5] ), .B2(n37797), .ZN(n37795) );
  INV_X1 U37265 ( .A(n37795), .ZN(n2750) );
  OAI22_X1 U37266 ( .A1(n37798), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[11][6] ), .B2(n37797), .ZN(n37796) );
  INV_X1 U37267 ( .A(n37796), .ZN(n2749) );
  OAI22_X1 U37268 ( .A1(n37798), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[11][7] ), .B2(n37797), .ZN(n37799) );
  INV_X1 U37269 ( .A(n37799), .ZN(n2748) );
  NOR2_X1 U37270 ( .A1(n39044), .A2(n38999), .ZN(n37822) );
  NAND2_X1 U37271 ( .A1(n37800), .A2(n37822), .ZN(n38946) );
  NOR2_X1 U37272 ( .A1(n37834), .A2(n38946), .ZN(n37808) );
  INV_X1 U37273 ( .A(n37808), .ZN(n37809) );
  OAI22_X1 U37274 ( .A1(n37809), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[12][0] ), .B2(n37808), .ZN(n37801) );
  INV_X1 U37275 ( .A(n37801), .ZN(n2747) );
  OAI22_X1 U37276 ( .A1(n37809), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[12][1] ), .B2(n37808), .ZN(n37802) );
  INV_X1 U37277 ( .A(n37802), .ZN(n2746) );
  OAI22_X1 U37278 ( .A1(n37809), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[12][2] ), .B2(n37808), .ZN(n37803) );
  INV_X1 U37279 ( .A(n37803), .ZN(n2745) );
  OAI22_X1 U37280 ( .A1(n37809), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[12][3] ), .B2(n37808), .ZN(n37804) );
  INV_X1 U37281 ( .A(n37804), .ZN(n2744) );
  OAI22_X1 U37282 ( .A1(n37809), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[12][4] ), .B2(n37808), .ZN(n37805) );
  INV_X1 U37283 ( .A(n37805), .ZN(n2743) );
  OAI22_X1 U37284 ( .A1(n37809), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[12][5] ), .B2(n37808), .ZN(n37806) );
  INV_X1 U37285 ( .A(n37806), .ZN(n2742) );
  OAI22_X1 U37286 ( .A1(n37809), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[12][6] ), .B2(n37808), .ZN(n37807) );
  INV_X1 U37287 ( .A(n37807), .ZN(n2741) );
  OAI22_X1 U37288 ( .A1(n37809), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[12][7] ), .B2(n37808), .ZN(n37810) );
  INV_X1 U37289 ( .A(n37810), .ZN(n2740) );
  NAND2_X1 U37290 ( .A1(n37811), .A2(n37822), .ZN(n38957) );
  NOR2_X1 U37291 ( .A1(n37834), .A2(n38957), .ZN(n37819) );
  INV_X1 U37292 ( .A(n37819), .ZN(n37820) );
  OAI22_X1 U37293 ( .A1(n37820), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[13][0] ), .B2(n37819), .ZN(n37812) );
  INV_X1 U37294 ( .A(n37812), .ZN(n2739) );
  OAI22_X1 U37295 ( .A1(n37820), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[13][1] ), .B2(n37819), .ZN(n37813) );
  INV_X1 U37296 ( .A(n37813), .ZN(n2738) );
  OAI22_X1 U37297 ( .A1(n37820), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[13][2] ), .B2(n37819), .ZN(n37814) );
  INV_X1 U37298 ( .A(n37814), .ZN(n2737) );
  OAI22_X1 U37299 ( .A1(n37820), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[13][3] ), .B2(n37819), .ZN(n37815) );
  INV_X1 U37300 ( .A(n37815), .ZN(n2736) );
  OAI22_X1 U37301 ( .A1(n37820), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[13][4] ), .B2(n37819), .ZN(n37816) );
  INV_X1 U37302 ( .A(n37816), .ZN(n2735) );
  OAI22_X1 U37303 ( .A1(n37820), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[13][5] ), .B2(n37819), .ZN(n37817) );
  INV_X1 U37304 ( .A(n37817), .ZN(n2734) );
  OAI22_X1 U37305 ( .A1(n37820), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[13][6] ), .B2(n37819), .ZN(n37818) );
  INV_X1 U37306 ( .A(n37818), .ZN(n2733) );
  OAI22_X1 U37307 ( .A1(n37820), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[13][7] ), .B2(n37819), .ZN(n37821) );
  INV_X1 U37308 ( .A(n37821), .ZN(n2732) );
  NAND2_X1 U37309 ( .A1(n37823), .A2(n37822), .ZN(n38968) );
  NOR2_X1 U37310 ( .A1(n37834), .A2(n38968), .ZN(n37831) );
  INV_X1 U37311 ( .A(n37831), .ZN(n37832) );
  OAI22_X1 U37312 ( .A1(n37832), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[14][0] ), .B2(n37831), .ZN(n37824) );
  INV_X1 U37313 ( .A(n37824), .ZN(n2731) );
  OAI22_X1 U37314 ( .A1(n37832), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[14][1] ), .B2(n37831), .ZN(n37825) );
  INV_X1 U37315 ( .A(n37825), .ZN(n2730) );
  OAI22_X1 U37316 ( .A1(n37832), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[14][2] ), .B2(n37831), .ZN(n37826) );
  INV_X1 U37317 ( .A(n37826), .ZN(n2729) );
  OAI22_X1 U37318 ( .A1(n37832), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[14][3] ), .B2(n37831), .ZN(n37827) );
  INV_X1 U37319 ( .A(n37827), .ZN(n2728) );
  OAI22_X1 U37320 ( .A1(n37832), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[14][4] ), .B2(n37831), .ZN(n37828) );
  INV_X1 U37321 ( .A(n37828), .ZN(n2727) );
  OAI22_X1 U37322 ( .A1(n37832), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[14][5] ), .B2(n37831), .ZN(n37829) );
  INV_X1 U37323 ( .A(n37829), .ZN(n2726) );
  OAI22_X1 U37324 ( .A1(n37832), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[14][6] ), .B2(n37831), .ZN(n37830) );
  INV_X1 U37325 ( .A(n37830), .ZN(n2725) );
  OAI22_X1 U37326 ( .A1(n37832), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[14][7] ), .B2(n37831), .ZN(n37833) );
  INV_X1 U37327 ( .A(n37833), .ZN(n2724) );
  NOR2_X1 U37328 ( .A1(n38803), .A2(n37834), .ZN(n37842) );
  INV_X1 U37329 ( .A(n37842), .ZN(n37843) );
  OAI22_X1 U37330 ( .A1(n37843), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[15][0] ), .B2(n37842), .ZN(n37835) );
  INV_X1 U37331 ( .A(n37835), .ZN(n2723) );
  OAI22_X1 U37332 ( .A1(n37843), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[15][1] ), .B2(n37842), .ZN(n37836) );
  INV_X1 U37333 ( .A(n37836), .ZN(n2722) );
  OAI22_X1 U37334 ( .A1(n37843), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[15][2] ), .B2(n37842), .ZN(n37837) );
  INV_X1 U37335 ( .A(n37837), .ZN(n2721) );
  OAI22_X1 U37336 ( .A1(n37843), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[15][3] ), .B2(n37842), .ZN(n37838) );
  INV_X1 U37337 ( .A(n37838), .ZN(n2720) );
  OAI22_X1 U37338 ( .A1(n37843), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[15][4] ), .B2(n37842), .ZN(n37839) );
  INV_X1 U37339 ( .A(n37839), .ZN(n2719) );
  OAI22_X1 U37340 ( .A1(n37843), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[15][5] ), .B2(n37842), .ZN(n37840) );
  INV_X1 U37341 ( .A(n37840), .ZN(n2718) );
  OAI22_X1 U37342 ( .A1(n37843), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[15][6] ), .B2(n37842), .ZN(n37841) );
  INV_X1 U37343 ( .A(n37841), .ZN(n2717) );
  OAI22_X1 U37344 ( .A1(n37843), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[15][7] ), .B2(n37842), .ZN(n37844) );
  INV_X1 U37345 ( .A(n37844), .ZN(n2716) );
  NAND3_X1 U37346 ( .A1(n38489), .A2(n39043), .A3(n38998), .ZN(n37995) );
  NOR2_X1 U37347 ( .A1(n38814), .A2(n37995), .ZN(n37852) );
  INV_X1 U37348 ( .A(n37852), .ZN(n37853) );
  OAI22_X1 U37349 ( .A1(n37853), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[16][0] ), .B2(n37852), .ZN(n37845) );
  INV_X1 U37350 ( .A(n37845), .ZN(n2715) );
  OAI22_X1 U37351 ( .A1(n37853), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[16][1] ), .B2(n37852), .ZN(n37846) );
  INV_X1 U37352 ( .A(n37846), .ZN(n2714) );
  OAI22_X1 U37353 ( .A1(n37853), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[16][2] ), .B2(n37852), .ZN(n37847) );
  INV_X1 U37354 ( .A(n37847), .ZN(n2713) );
  OAI22_X1 U37355 ( .A1(n37853), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[16][3] ), .B2(n37852), .ZN(n37848) );
  INV_X1 U37356 ( .A(n37848), .ZN(n2712) );
  OAI22_X1 U37357 ( .A1(n37853), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[16][4] ), .B2(n37852), .ZN(n37849) );
  INV_X1 U37358 ( .A(n37849), .ZN(n2711) );
  OAI22_X1 U37359 ( .A1(n37853), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[16][5] ), .B2(n37852), .ZN(n37850) );
  INV_X1 U37360 ( .A(n37850), .ZN(n2710) );
  OAI22_X1 U37361 ( .A1(n37853), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[16][6] ), .B2(n37852), .ZN(n37851) );
  INV_X1 U37362 ( .A(n37851), .ZN(n2709) );
  OAI22_X1 U37363 ( .A1(n37853), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[16][7] ), .B2(n37852), .ZN(n37854) );
  INV_X1 U37364 ( .A(n37854), .ZN(n2708) );
  NOR2_X1 U37365 ( .A1(n38825), .A2(n37995), .ZN(n37862) );
  INV_X1 U37366 ( .A(n37862), .ZN(n37863) );
  OAI22_X1 U37367 ( .A1(n37863), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[17][0] ), .B2(n37862), .ZN(n37855) );
  INV_X1 U37368 ( .A(n37855), .ZN(n2707) );
  OAI22_X1 U37369 ( .A1(n37863), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[17][1] ), .B2(n37862), .ZN(n37856) );
  INV_X1 U37370 ( .A(n37856), .ZN(n2706) );
  OAI22_X1 U37371 ( .A1(n37863), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[17][2] ), .B2(n37862), .ZN(n37857) );
  INV_X1 U37372 ( .A(n37857), .ZN(n2705) );
  OAI22_X1 U37373 ( .A1(n37863), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[17][3] ), .B2(n37862), .ZN(n37858) );
  INV_X1 U37374 ( .A(n37858), .ZN(n2704) );
  OAI22_X1 U37375 ( .A1(n37863), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[17][4] ), .B2(n37862), .ZN(n37859) );
  INV_X1 U37376 ( .A(n37859), .ZN(n2703) );
  OAI22_X1 U37377 ( .A1(n37863), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[17][5] ), .B2(n37862), .ZN(n37860) );
  INV_X1 U37378 ( .A(n37860), .ZN(n2702) );
  OAI22_X1 U37379 ( .A1(n37863), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[17][6] ), .B2(n37862), .ZN(n37861) );
  INV_X1 U37380 ( .A(n37861), .ZN(n2701) );
  OAI22_X1 U37381 ( .A1(n37863), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[17][7] ), .B2(n37862), .ZN(n37864) );
  INV_X1 U37382 ( .A(n37864), .ZN(n2700) );
  NOR2_X1 U37383 ( .A1(n38836), .A2(n37995), .ZN(n37872) );
  INV_X1 U37384 ( .A(n37872), .ZN(n37873) );
  OAI22_X1 U37385 ( .A1(n37873), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[18][0] ), .B2(n37872), .ZN(n37865) );
  INV_X1 U37386 ( .A(n37865), .ZN(n2699) );
  OAI22_X1 U37387 ( .A1(n37873), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[18][1] ), .B2(n37872), .ZN(n37866) );
  INV_X1 U37388 ( .A(n37866), .ZN(n2698) );
  OAI22_X1 U37389 ( .A1(n37873), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[18][2] ), .B2(n37872), .ZN(n37867) );
  INV_X1 U37390 ( .A(n37867), .ZN(n2697) );
  OAI22_X1 U37391 ( .A1(n37873), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[18][3] ), .B2(n37872), .ZN(n37868) );
  INV_X1 U37392 ( .A(n37868), .ZN(n2696) );
  OAI22_X1 U37393 ( .A1(n37873), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[18][4] ), .B2(n37872), .ZN(n37869) );
  INV_X1 U37394 ( .A(n37869), .ZN(n2695) );
  OAI22_X1 U37395 ( .A1(n37873), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[18][5] ), .B2(n37872), .ZN(n37870) );
  INV_X1 U37396 ( .A(n37870), .ZN(n2694) );
  OAI22_X1 U37397 ( .A1(n37873), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[18][6] ), .B2(n37872), .ZN(n37871) );
  INV_X1 U37398 ( .A(n37871), .ZN(n2693) );
  OAI22_X1 U37399 ( .A1(n37873), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[18][7] ), .B2(n37872), .ZN(n37874) );
  INV_X1 U37400 ( .A(n37874), .ZN(n2692) );
  NOR2_X1 U37401 ( .A1(n38847), .A2(n37995), .ZN(n37882) );
  INV_X1 U37402 ( .A(n37882), .ZN(n37883) );
  OAI22_X1 U37403 ( .A1(n37883), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[19][0] ), .B2(n37882), .ZN(n37875) );
  INV_X1 U37404 ( .A(n37875), .ZN(n2691) );
  OAI22_X1 U37405 ( .A1(n37883), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[19][1] ), .B2(n37882), .ZN(n37876) );
  INV_X1 U37406 ( .A(n37876), .ZN(n2690) );
  OAI22_X1 U37407 ( .A1(n37883), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[19][2] ), .B2(n37882), .ZN(n37877) );
  INV_X1 U37408 ( .A(n37877), .ZN(n2689) );
  OAI22_X1 U37409 ( .A1(n37883), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[19][3] ), .B2(n37882), .ZN(n37878) );
  INV_X1 U37410 ( .A(n37878), .ZN(n2688) );
  OAI22_X1 U37411 ( .A1(n37883), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[19][4] ), .B2(n37882), .ZN(n37879) );
  INV_X1 U37412 ( .A(n37879), .ZN(n2687) );
  OAI22_X1 U37413 ( .A1(n37883), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[19][5] ), .B2(n37882), .ZN(n37880) );
  INV_X1 U37414 ( .A(n37880), .ZN(n2686) );
  OAI22_X1 U37415 ( .A1(n37883), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[19][6] ), .B2(n37882), .ZN(n37881) );
  INV_X1 U37416 ( .A(n37881), .ZN(n2685) );
  OAI22_X1 U37417 ( .A1(n37883), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[19][7] ), .B2(n37882), .ZN(n37884) );
  INV_X1 U37418 ( .A(n37884), .ZN(n2684) );
  NOR2_X1 U37419 ( .A1(n38858), .A2(n37995), .ZN(n37892) );
  INV_X1 U37420 ( .A(n37892), .ZN(n37893) );
  OAI22_X1 U37421 ( .A1(n37893), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[20][0] ), .B2(n37892), .ZN(n37885) );
  INV_X1 U37422 ( .A(n37885), .ZN(n2683) );
  OAI22_X1 U37423 ( .A1(n37893), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[20][1] ), .B2(n37892), .ZN(n37886) );
  INV_X1 U37424 ( .A(n37886), .ZN(n2682) );
  OAI22_X1 U37425 ( .A1(n37893), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[20][2] ), .B2(n37892), .ZN(n37887) );
  INV_X1 U37426 ( .A(n37887), .ZN(n2681) );
  OAI22_X1 U37427 ( .A1(n37893), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[20][3] ), .B2(n37892), .ZN(n37888) );
  INV_X1 U37428 ( .A(n37888), .ZN(n2680) );
  OAI22_X1 U37429 ( .A1(n37893), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[20][4] ), .B2(n37892), .ZN(n37889) );
  INV_X1 U37430 ( .A(n37889), .ZN(n2679) );
  OAI22_X1 U37431 ( .A1(n37893), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[20][5] ), .B2(n37892), .ZN(n37890) );
  INV_X1 U37432 ( .A(n37890), .ZN(n2678) );
  OAI22_X1 U37433 ( .A1(n37893), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[20][6] ), .B2(n37892), .ZN(n37891) );
  INV_X1 U37434 ( .A(n37891), .ZN(n2677) );
  OAI22_X1 U37435 ( .A1(n37893), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[20][7] ), .B2(n37892), .ZN(n37894) );
  INV_X1 U37436 ( .A(n37894), .ZN(n2676) );
  NOR2_X1 U37437 ( .A1(n38869), .A2(n37995), .ZN(n37902) );
  INV_X1 U37438 ( .A(n37902), .ZN(n37903) );
  OAI22_X1 U37439 ( .A1(n37903), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[21][0] ), .B2(n37902), .ZN(n37895) );
  INV_X1 U37440 ( .A(n37895), .ZN(n2675) );
  OAI22_X1 U37441 ( .A1(n37903), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[21][1] ), .B2(n37902), .ZN(n37896) );
  INV_X1 U37442 ( .A(n37896), .ZN(n2674) );
  OAI22_X1 U37443 ( .A1(n37903), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[21][2] ), .B2(n37902), .ZN(n37897) );
  INV_X1 U37444 ( .A(n37897), .ZN(n2673) );
  OAI22_X1 U37445 ( .A1(n37903), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[21][3] ), .B2(n37902), .ZN(n37898) );
  INV_X1 U37446 ( .A(n37898), .ZN(n2672) );
  OAI22_X1 U37447 ( .A1(n37903), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[21][4] ), .B2(n37902), .ZN(n37899) );
  INV_X1 U37448 ( .A(n37899), .ZN(n2671) );
  OAI22_X1 U37449 ( .A1(n37903), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[21][5] ), .B2(n37902), .ZN(n37900) );
  INV_X1 U37450 ( .A(n37900), .ZN(n2670) );
  OAI22_X1 U37451 ( .A1(n37903), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[21][6] ), .B2(n37902), .ZN(n37901) );
  INV_X1 U37452 ( .A(n37901), .ZN(n2669) );
  OAI22_X1 U37453 ( .A1(n37903), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[21][7] ), .B2(n37902), .ZN(n37904) );
  INV_X1 U37454 ( .A(n37904), .ZN(n2668) );
  NOR2_X1 U37455 ( .A1(n38880), .A2(n37995), .ZN(n37912) );
  INV_X1 U37456 ( .A(n37912), .ZN(n37913) );
  OAI22_X1 U37457 ( .A1(n37913), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[22][0] ), .B2(n37912), .ZN(n37905) );
  INV_X1 U37458 ( .A(n37905), .ZN(n2667) );
  OAI22_X1 U37459 ( .A1(n37913), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[22][1] ), .B2(n37912), .ZN(n37906) );
  INV_X1 U37460 ( .A(n37906), .ZN(n2666) );
  OAI22_X1 U37461 ( .A1(n37913), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[22][2] ), .B2(n37912), .ZN(n37907) );
  INV_X1 U37462 ( .A(n37907), .ZN(n2665) );
  OAI22_X1 U37463 ( .A1(n37913), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[22][3] ), .B2(n37912), .ZN(n37908) );
  INV_X1 U37464 ( .A(n37908), .ZN(n2664) );
  OAI22_X1 U37465 ( .A1(n37913), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[22][4] ), .B2(n37912), .ZN(n37909) );
  INV_X1 U37466 ( .A(n37909), .ZN(n2663) );
  OAI22_X1 U37467 ( .A1(n37913), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[22][5] ), .B2(n37912), .ZN(n37910) );
  INV_X1 U37468 ( .A(n37910), .ZN(n2662) );
  OAI22_X1 U37469 ( .A1(n37913), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[22][6] ), .B2(n37912), .ZN(n37911) );
  INV_X1 U37470 ( .A(n37911), .ZN(n2661) );
  OAI22_X1 U37471 ( .A1(n37913), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[22][7] ), .B2(n37912), .ZN(n37914) );
  INV_X1 U37472 ( .A(n37914), .ZN(n2660) );
  NOR2_X1 U37473 ( .A1(n38891), .A2(n37995), .ZN(n37922) );
  INV_X1 U37474 ( .A(n37922), .ZN(n37923) );
  OAI22_X1 U37475 ( .A1(n37923), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[23][0] ), .B2(n37922), .ZN(n37915) );
  INV_X1 U37476 ( .A(n37915), .ZN(n2659) );
  OAI22_X1 U37477 ( .A1(n37923), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[23][1] ), .B2(n37922), .ZN(n37916) );
  INV_X1 U37478 ( .A(n37916), .ZN(n2658) );
  OAI22_X1 U37479 ( .A1(n37923), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[23][2] ), .B2(n37922), .ZN(n37917) );
  INV_X1 U37480 ( .A(n37917), .ZN(n2657) );
  OAI22_X1 U37481 ( .A1(n37923), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[23][3] ), .B2(n37922), .ZN(n37918) );
  INV_X1 U37482 ( .A(n37918), .ZN(n2656) );
  OAI22_X1 U37483 ( .A1(n37923), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[23][4] ), .B2(n37922), .ZN(n37919) );
  INV_X1 U37484 ( .A(n37919), .ZN(n2655) );
  OAI22_X1 U37485 ( .A1(n37923), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[23][5] ), .B2(n37922), .ZN(n37920) );
  INV_X1 U37486 ( .A(n37920), .ZN(n2654) );
  OAI22_X1 U37487 ( .A1(n37923), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[23][6] ), .B2(n37922), .ZN(n37921) );
  INV_X1 U37488 ( .A(n37921), .ZN(n2653) );
  OAI22_X1 U37489 ( .A1(n37923), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[23][7] ), .B2(n37922), .ZN(n37924) );
  INV_X1 U37490 ( .A(n37924), .ZN(n2652) );
  NOR2_X1 U37491 ( .A1(n38902), .A2(n37995), .ZN(n37932) );
  INV_X1 U37492 ( .A(n37932), .ZN(n37933) );
  OAI22_X1 U37493 ( .A1(n37933), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[24][0] ), .B2(n37932), .ZN(n37925) );
  INV_X1 U37494 ( .A(n37925), .ZN(n2651) );
  OAI22_X1 U37495 ( .A1(n37933), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[24][1] ), .B2(n37932), .ZN(n37926) );
  INV_X1 U37496 ( .A(n37926), .ZN(n2650) );
  OAI22_X1 U37497 ( .A1(n37933), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[24][2] ), .B2(n37932), .ZN(n37927) );
  INV_X1 U37498 ( .A(n37927), .ZN(n2649) );
  OAI22_X1 U37499 ( .A1(n37933), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[24][3] ), .B2(n37932), .ZN(n37928) );
  INV_X1 U37500 ( .A(n37928), .ZN(n2648) );
  OAI22_X1 U37501 ( .A1(n37933), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[24][4] ), .B2(n37932), .ZN(n37929) );
  INV_X1 U37502 ( .A(n37929), .ZN(n2647) );
  OAI22_X1 U37503 ( .A1(n37933), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[24][5] ), .B2(n37932), .ZN(n37930) );
  INV_X1 U37504 ( .A(n37930), .ZN(n2646) );
  OAI22_X1 U37505 ( .A1(n37933), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[24][6] ), .B2(n37932), .ZN(n37931) );
  INV_X1 U37506 ( .A(n37931), .ZN(n2645) );
  OAI22_X1 U37507 ( .A1(n37933), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[24][7] ), .B2(n37932), .ZN(n37934) );
  INV_X1 U37508 ( .A(n37934), .ZN(n2644) );
  NOR2_X1 U37509 ( .A1(n38913), .A2(n37995), .ZN(n37942) );
  INV_X1 U37510 ( .A(n37942), .ZN(n37943) );
  OAI22_X1 U37511 ( .A1(n37943), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[25][0] ), .B2(n37942), .ZN(n37935) );
  INV_X1 U37512 ( .A(n37935), .ZN(n2643) );
  OAI22_X1 U37513 ( .A1(n37943), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[25][1] ), .B2(n37942), .ZN(n37936) );
  INV_X1 U37514 ( .A(n37936), .ZN(n2642) );
  OAI22_X1 U37515 ( .A1(n37943), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[25][2] ), .B2(n37942), .ZN(n37937) );
  INV_X1 U37516 ( .A(n37937), .ZN(n2641) );
  OAI22_X1 U37517 ( .A1(n37943), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[25][3] ), .B2(n37942), .ZN(n37938) );
  INV_X1 U37518 ( .A(n37938), .ZN(n2640) );
  OAI22_X1 U37519 ( .A1(n37943), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[25][4] ), .B2(n37942), .ZN(n37939) );
  INV_X1 U37520 ( .A(n37939), .ZN(n2639) );
  OAI22_X1 U37521 ( .A1(n37943), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[25][5] ), .B2(n37942), .ZN(n37940) );
  INV_X1 U37522 ( .A(n37940), .ZN(n2638) );
  OAI22_X1 U37523 ( .A1(n37943), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[25][6] ), .B2(n37942), .ZN(n37941) );
  INV_X1 U37524 ( .A(n37941), .ZN(n2637) );
  OAI22_X1 U37525 ( .A1(n37943), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[25][7] ), .B2(n37942), .ZN(n37944) );
  INV_X1 U37526 ( .A(n37944), .ZN(n2636) );
  NOR2_X1 U37527 ( .A1(n38924), .A2(n37995), .ZN(n37952) );
  INV_X1 U37528 ( .A(n37952), .ZN(n37953) );
  OAI22_X1 U37529 ( .A1(n37953), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[26][0] ), .B2(n37952), .ZN(n37945) );
  INV_X1 U37530 ( .A(n37945), .ZN(n2635) );
  OAI22_X1 U37531 ( .A1(n37953), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[26][1] ), .B2(n37952), .ZN(n37946) );
  INV_X1 U37532 ( .A(n37946), .ZN(n2634) );
  OAI22_X1 U37533 ( .A1(n37953), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[26][2] ), .B2(n37952), .ZN(n37947) );
  INV_X1 U37534 ( .A(n37947), .ZN(n2633) );
  OAI22_X1 U37535 ( .A1(n37953), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[26][3] ), .B2(n37952), .ZN(n37948) );
  INV_X1 U37536 ( .A(n37948), .ZN(n2632) );
  OAI22_X1 U37537 ( .A1(n37953), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[26][4] ), .B2(n37952), .ZN(n37949) );
  INV_X1 U37538 ( .A(n37949), .ZN(n2631) );
  OAI22_X1 U37539 ( .A1(n37953), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[26][5] ), .B2(n37952), .ZN(n37950) );
  INV_X1 U37540 ( .A(n37950), .ZN(n2630) );
  OAI22_X1 U37541 ( .A1(n37953), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[26][6] ), .B2(n37952), .ZN(n37951) );
  INV_X1 U37542 ( .A(n37951), .ZN(n2629) );
  OAI22_X1 U37543 ( .A1(n37953), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[26][7] ), .B2(n37952), .ZN(n37954) );
  INV_X1 U37544 ( .A(n37954), .ZN(n2628) );
  NOR2_X1 U37545 ( .A1(n38935), .A2(n37995), .ZN(n37962) );
  INV_X1 U37546 ( .A(n37962), .ZN(n37963) );
  OAI22_X1 U37547 ( .A1(n37963), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[27][0] ), .B2(n37962), .ZN(n37955) );
  INV_X1 U37548 ( .A(n37955), .ZN(n2627) );
  OAI22_X1 U37549 ( .A1(n37963), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[27][1] ), .B2(n37962), .ZN(n37956) );
  INV_X1 U37550 ( .A(n37956), .ZN(n2626) );
  OAI22_X1 U37551 ( .A1(n37963), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[27][2] ), .B2(n37962), .ZN(n37957) );
  INV_X1 U37552 ( .A(n37957), .ZN(n2625) );
  OAI22_X1 U37553 ( .A1(n37963), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[27][3] ), .B2(n37962), .ZN(n37958) );
  INV_X1 U37554 ( .A(n37958), .ZN(n2624) );
  OAI22_X1 U37555 ( .A1(n37963), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[27][4] ), .B2(n37962), .ZN(n37959) );
  INV_X1 U37556 ( .A(n37959), .ZN(n2623) );
  OAI22_X1 U37557 ( .A1(n37963), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[27][5] ), .B2(n37962), .ZN(n37960) );
  INV_X1 U37558 ( .A(n37960), .ZN(n2622) );
  OAI22_X1 U37559 ( .A1(n37963), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[27][6] ), .B2(n37962), .ZN(n37961) );
  INV_X1 U37560 ( .A(n37961), .ZN(n2621) );
  OAI22_X1 U37561 ( .A1(n37963), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[27][7] ), .B2(n37962), .ZN(n37964) );
  INV_X1 U37562 ( .A(n37964), .ZN(n2620) );
  NOR2_X1 U37563 ( .A1(n38946), .A2(n37995), .ZN(n37972) );
  INV_X1 U37564 ( .A(n37972), .ZN(n37973) );
  OAI22_X1 U37565 ( .A1(n37973), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[28][0] ), .B2(n37972), .ZN(n37965) );
  INV_X1 U37566 ( .A(n37965), .ZN(n2619) );
  OAI22_X1 U37567 ( .A1(n37973), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[28][1] ), .B2(n37972), .ZN(n37966) );
  INV_X1 U37568 ( .A(n37966), .ZN(n2618) );
  OAI22_X1 U37569 ( .A1(n37973), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[28][2] ), .B2(n37972), .ZN(n37967) );
  INV_X1 U37570 ( .A(n37967), .ZN(n2617) );
  OAI22_X1 U37571 ( .A1(n37973), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[28][3] ), .B2(n37972), .ZN(n37968) );
  INV_X1 U37572 ( .A(n37968), .ZN(n2616) );
  OAI22_X1 U37573 ( .A1(n37973), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[28][4] ), .B2(n37972), .ZN(n37969) );
  INV_X1 U37574 ( .A(n37969), .ZN(n2615) );
  OAI22_X1 U37575 ( .A1(n37973), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[28][5] ), .B2(n37972), .ZN(n37970) );
  INV_X1 U37576 ( .A(n37970), .ZN(n2614) );
  OAI22_X1 U37577 ( .A1(n37973), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[28][6] ), .B2(n37972), .ZN(n37971) );
  INV_X1 U37578 ( .A(n37971), .ZN(n2613) );
  OAI22_X1 U37579 ( .A1(n37973), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[28][7] ), .B2(n37972), .ZN(n37974) );
  INV_X1 U37580 ( .A(n37974), .ZN(n2612) );
  NOR2_X1 U37581 ( .A1(n38957), .A2(n37995), .ZN(n37982) );
  INV_X1 U37582 ( .A(n37982), .ZN(n37983) );
  OAI22_X1 U37583 ( .A1(n37983), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[29][0] ), .B2(n37982), .ZN(n37975) );
  INV_X1 U37584 ( .A(n37975), .ZN(n2611) );
  OAI22_X1 U37585 ( .A1(n37983), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[29][1] ), .B2(n37982), .ZN(n37976) );
  INV_X1 U37586 ( .A(n37976), .ZN(n2610) );
  OAI22_X1 U37587 ( .A1(n37983), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[29][2] ), .B2(n37982), .ZN(n37977) );
  INV_X1 U37588 ( .A(n37977), .ZN(n2609) );
  OAI22_X1 U37589 ( .A1(n37983), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[29][3] ), .B2(n37982), .ZN(n37978) );
  INV_X1 U37590 ( .A(n37978), .ZN(n2608) );
  OAI22_X1 U37591 ( .A1(n37983), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[29][4] ), .B2(n37982), .ZN(n37979) );
  INV_X1 U37592 ( .A(n37979), .ZN(n2607) );
  OAI22_X1 U37593 ( .A1(n37983), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[29][5] ), .B2(n37982), .ZN(n37980) );
  INV_X1 U37594 ( .A(n37980), .ZN(n2606) );
  OAI22_X1 U37595 ( .A1(n37983), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[29][6] ), .B2(n37982), .ZN(n37981) );
  INV_X1 U37596 ( .A(n37981), .ZN(n2605) );
  OAI22_X1 U37597 ( .A1(n37983), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[29][7] ), .B2(n37982), .ZN(n37984) );
  INV_X1 U37598 ( .A(n37984), .ZN(n2604) );
  NOR2_X1 U37599 ( .A1(n38968), .A2(n37995), .ZN(n37992) );
  INV_X1 U37600 ( .A(n37992), .ZN(n37993) );
  OAI22_X1 U37601 ( .A1(n37993), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[30][0] ), .B2(n37992), .ZN(n37985) );
  INV_X1 U37602 ( .A(n37985), .ZN(n2603) );
  OAI22_X1 U37603 ( .A1(n37993), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[30][1] ), .B2(n37992), .ZN(n37986) );
  INV_X1 U37604 ( .A(n37986), .ZN(n2602) );
  OAI22_X1 U37605 ( .A1(n37993), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[30][2] ), .B2(n37992), .ZN(n37987) );
  INV_X1 U37606 ( .A(n37987), .ZN(n2601) );
  OAI22_X1 U37607 ( .A1(n37993), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[30][3] ), .B2(n37992), .ZN(n37988) );
  INV_X1 U37608 ( .A(n37988), .ZN(n2600) );
  OAI22_X1 U37609 ( .A1(n37993), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[30][4] ), .B2(n37992), .ZN(n37989) );
  INV_X1 U37610 ( .A(n37989), .ZN(n2599) );
  OAI22_X1 U37611 ( .A1(n37993), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[30][5] ), .B2(n37992), .ZN(n37990) );
  INV_X1 U37612 ( .A(n37990), .ZN(n2598) );
  OAI22_X1 U37613 ( .A1(n37993), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[30][6] ), .B2(n37992), .ZN(n37991) );
  INV_X1 U37614 ( .A(n37991), .ZN(n2597) );
  OAI22_X1 U37615 ( .A1(n37993), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[30][7] ), .B2(n37992), .ZN(n37994) );
  INV_X1 U37616 ( .A(n37994), .ZN(n2596) );
  NOR2_X1 U37617 ( .A1(n38803), .A2(n37995), .ZN(n38003) );
  INV_X1 U37618 ( .A(n38003), .ZN(n38004) );
  OAI22_X1 U37619 ( .A1(n38004), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[31][0] ), .B2(n38003), .ZN(n37996) );
  INV_X1 U37620 ( .A(n37996), .ZN(n2595) );
  OAI22_X1 U37621 ( .A1(n38004), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[31][1] ), .B2(n38003), .ZN(n37997) );
  INV_X1 U37622 ( .A(n37997), .ZN(n2594) );
  OAI22_X1 U37623 ( .A1(n38004), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[31][2] ), .B2(n38003), .ZN(n37998) );
  INV_X1 U37624 ( .A(n37998), .ZN(n2593) );
  OAI22_X1 U37625 ( .A1(n38004), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[31][3] ), .B2(n38003), .ZN(n37999) );
  INV_X1 U37626 ( .A(n37999), .ZN(n2592) );
  OAI22_X1 U37627 ( .A1(n38004), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[31][4] ), .B2(n38003), .ZN(n38000) );
  INV_X1 U37628 ( .A(n38000), .ZN(n2591) );
  OAI22_X1 U37629 ( .A1(n38004), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[31][5] ), .B2(n38003), .ZN(n38001) );
  INV_X1 U37630 ( .A(n38001), .ZN(n2590) );
  OAI22_X1 U37631 ( .A1(n38004), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[31][6] ), .B2(n38003), .ZN(n38002) );
  INV_X1 U37632 ( .A(n38002), .ZN(n2589) );
  OAI22_X1 U37633 ( .A1(n38004), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[31][7] ), .B2(n38003), .ZN(n38005) );
  INV_X1 U37634 ( .A(n38005), .ZN(n2588) );
  NAND3_X1 U37635 ( .A1(xmem_addr[5]), .A2(n38651), .A3(n39043), .ZN(n38156)
         );
  NOR2_X1 U37636 ( .A1(n38814), .A2(n38156), .ZN(n38013) );
  INV_X1 U37637 ( .A(n38013), .ZN(n38014) );
  OAI22_X1 U37638 ( .A1(n38014), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[32][0] ), .B2(n38013), .ZN(n38006) );
  INV_X1 U37639 ( .A(n38006), .ZN(n2587) );
  OAI22_X1 U37640 ( .A1(n38014), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[32][1] ), .B2(n38013), .ZN(n38007) );
  INV_X1 U37641 ( .A(n38007), .ZN(n2586) );
  OAI22_X1 U37642 ( .A1(n38014), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[32][2] ), .B2(n38013), .ZN(n38008) );
  INV_X1 U37643 ( .A(n38008), .ZN(n2585) );
  OAI22_X1 U37644 ( .A1(n38014), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[32][3] ), .B2(n38013), .ZN(n38009) );
  INV_X1 U37645 ( .A(n38009), .ZN(n2584) );
  OAI22_X1 U37646 ( .A1(n38014), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[32][4] ), .B2(n38013), .ZN(n38010) );
  INV_X1 U37647 ( .A(n38010), .ZN(n2583) );
  OAI22_X1 U37648 ( .A1(n38014), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[32][5] ), .B2(n38013), .ZN(n38011) );
  INV_X1 U37649 ( .A(n38011), .ZN(n2582) );
  OAI22_X1 U37650 ( .A1(n38014), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[32][6] ), .B2(n38013), .ZN(n38012) );
  INV_X1 U37651 ( .A(n38012), .ZN(n2581) );
  OAI22_X1 U37652 ( .A1(n38014), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[32][7] ), .B2(n38013), .ZN(n38015) );
  INV_X1 U37653 ( .A(n38015), .ZN(n2580) );
  NOR2_X1 U37654 ( .A1(n38825), .A2(n38156), .ZN(n38023) );
  INV_X1 U37655 ( .A(n38023), .ZN(n38024) );
  OAI22_X1 U37656 ( .A1(n38024), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[33][0] ), .B2(n38023), .ZN(n38016) );
  INV_X1 U37657 ( .A(n38016), .ZN(n2579) );
  OAI22_X1 U37658 ( .A1(n38024), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[33][1] ), .B2(n38023), .ZN(n38017) );
  INV_X1 U37659 ( .A(n38017), .ZN(n2578) );
  OAI22_X1 U37660 ( .A1(n38024), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[33][2] ), .B2(n38023), .ZN(n38018) );
  INV_X1 U37661 ( .A(n38018), .ZN(n2577) );
  OAI22_X1 U37662 ( .A1(n38024), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[33][3] ), .B2(n38023), .ZN(n38019) );
  INV_X1 U37663 ( .A(n38019), .ZN(n2576) );
  OAI22_X1 U37664 ( .A1(n38024), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[33][4] ), .B2(n38023), .ZN(n38020) );
  INV_X1 U37665 ( .A(n38020), .ZN(n2575) );
  OAI22_X1 U37666 ( .A1(n38024), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[33][5] ), .B2(n38023), .ZN(n38021) );
  INV_X1 U37667 ( .A(n38021), .ZN(n2574) );
  OAI22_X1 U37668 ( .A1(n38024), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[33][6] ), .B2(n38023), .ZN(n38022) );
  INV_X1 U37669 ( .A(n38022), .ZN(n2573) );
  OAI22_X1 U37670 ( .A1(n38024), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[33][7] ), .B2(n38023), .ZN(n38025) );
  INV_X1 U37671 ( .A(n38025), .ZN(n2572) );
  NOR2_X1 U37672 ( .A1(n38836), .A2(n38156), .ZN(n38033) );
  INV_X1 U37673 ( .A(n38033), .ZN(n38034) );
  OAI22_X1 U37674 ( .A1(n38034), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[34][0] ), .B2(n38033), .ZN(n38026) );
  INV_X1 U37675 ( .A(n38026), .ZN(n2571) );
  OAI22_X1 U37676 ( .A1(n38034), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[34][1] ), .B2(n38033), .ZN(n38027) );
  INV_X1 U37677 ( .A(n38027), .ZN(n2570) );
  OAI22_X1 U37678 ( .A1(n38034), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[34][2] ), .B2(n38033), .ZN(n38028) );
  INV_X1 U37679 ( .A(n38028), .ZN(n2569) );
  OAI22_X1 U37680 ( .A1(n38034), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[34][3] ), .B2(n38033), .ZN(n38029) );
  INV_X1 U37681 ( .A(n38029), .ZN(n2568) );
  OAI22_X1 U37682 ( .A1(n38034), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[34][4] ), .B2(n38033), .ZN(n38030) );
  INV_X1 U37683 ( .A(n38030), .ZN(n2567) );
  OAI22_X1 U37684 ( .A1(n38034), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[34][5] ), .B2(n38033), .ZN(n38031) );
  INV_X1 U37685 ( .A(n38031), .ZN(n2566) );
  OAI22_X1 U37686 ( .A1(n38034), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[34][6] ), .B2(n38033), .ZN(n38032) );
  INV_X1 U37687 ( .A(n38032), .ZN(n2565) );
  OAI22_X1 U37688 ( .A1(n38034), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[34][7] ), .B2(n38033), .ZN(n38035) );
  INV_X1 U37689 ( .A(n38035), .ZN(n2564) );
  NOR2_X1 U37690 ( .A1(n38847), .A2(n38156), .ZN(n38043) );
  INV_X1 U37691 ( .A(n38043), .ZN(n38044) );
  OAI22_X1 U37692 ( .A1(n38044), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[35][0] ), .B2(n38043), .ZN(n38036) );
  INV_X1 U37693 ( .A(n38036), .ZN(n2563) );
  OAI22_X1 U37694 ( .A1(n38044), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[35][1] ), .B2(n38043), .ZN(n38037) );
  INV_X1 U37695 ( .A(n38037), .ZN(n2562) );
  OAI22_X1 U37696 ( .A1(n38044), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[35][2] ), .B2(n38043), .ZN(n38038) );
  INV_X1 U37697 ( .A(n38038), .ZN(n2561) );
  OAI22_X1 U37698 ( .A1(n38044), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[35][3] ), .B2(n38043), .ZN(n38039) );
  INV_X1 U37699 ( .A(n38039), .ZN(n2560) );
  OAI22_X1 U37700 ( .A1(n38044), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[35][4] ), .B2(n38043), .ZN(n38040) );
  INV_X1 U37701 ( .A(n38040), .ZN(n2559) );
  OAI22_X1 U37702 ( .A1(n38044), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[35][5] ), .B2(n38043), .ZN(n38041) );
  INV_X1 U37703 ( .A(n38041), .ZN(n2558) );
  OAI22_X1 U37704 ( .A1(n38044), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[35][6] ), .B2(n38043), .ZN(n38042) );
  INV_X1 U37705 ( .A(n38042), .ZN(n2557) );
  OAI22_X1 U37706 ( .A1(n38044), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[35][7] ), .B2(n38043), .ZN(n38045) );
  INV_X1 U37707 ( .A(n38045), .ZN(n2556) );
  NOR2_X1 U37708 ( .A1(n38858), .A2(n38156), .ZN(n38053) );
  INV_X1 U37709 ( .A(n38053), .ZN(n38054) );
  OAI22_X1 U37710 ( .A1(n38054), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[36][0] ), .B2(n38053), .ZN(n38046) );
  INV_X1 U37711 ( .A(n38046), .ZN(n2555) );
  OAI22_X1 U37712 ( .A1(n38054), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[36][1] ), .B2(n38053), .ZN(n38047) );
  INV_X1 U37713 ( .A(n38047), .ZN(n2554) );
  OAI22_X1 U37714 ( .A1(n38054), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[36][2] ), .B2(n38053), .ZN(n38048) );
  INV_X1 U37715 ( .A(n38048), .ZN(n2553) );
  OAI22_X1 U37716 ( .A1(n38054), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[36][3] ), .B2(n38053), .ZN(n38049) );
  INV_X1 U37717 ( .A(n38049), .ZN(n2552) );
  OAI22_X1 U37718 ( .A1(n38054), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[36][4] ), .B2(n38053), .ZN(n38050) );
  INV_X1 U37719 ( .A(n38050), .ZN(n2551) );
  OAI22_X1 U37720 ( .A1(n38054), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[36][5] ), .B2(n38053), .ZN(n38051) );
  INV_X1 U37721 ( .A(n38051), .ZN(n2550) );
  OAI22_X1 U37722 ( .A1(n38054), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[36][6] ), .B2(n38053), .ZN(n38052) );
  INV_X1 U37723 ( .A(n38052), .ZN(n2549) );
  OAI22_X1 U37724 ( .A1(n38054), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[36][7] ), .B2(n38053), .ZN(n38055) );
  INV_X1 U37725 ( .A(n38055), .ZN(n2548) );
  NOR2_X1 U37726 ( .A1(n38869), .A2(n38156), .ZN(n38063) );
  INV_X1 U37727 ( .A(n38063), .ZN(n38064) );
  OAI22_X1 U37728 ( .A1(n38064), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[37][0] ), .B2(n38063), .ZN(n38056) );
  INV_X1 U37729 ( .A(n38056), .ZN(n2547) );
  OAI22_X1 U37730 ( .A1(n38064), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[37][1] ), .B2(n38063), .ZN(n38057) );
  INV_X1 U37731 ( .A(n38057), .ZN(n2546) );
  OAI22_X1 U37732 ( .A1(n38064), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[37][2] ), .B2(n38063), .ZN(n38058) );
  INV_X1 U37733 ( .A(n38058), .ZN(n2545) );
  OAI22_X1 U37734 ( .A1(n38064), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[37][3] ), .B2(n38063), .ZN(n38059) );
  INV_X1 U37735 ( .A(n38059), .ZN(n2544) );
  OAI22_X1 U37736 ( .A1(n38064), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[37][4] ), .B2(n38063), .ZN(n38060) );
  INV_X1 U37737 ( .A(n38060), .ZN(n2543) );
  OAI22_X1 U37738 ( .A1(n38064), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[37][5] ), .B2(n38063), .ZN(n38061) );
  INV_X1 U37739 ( .A(n38061), .ZN(n2542) );
  OAI22_X1 U37740 ( .A1(n38064), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[37][6] ), .B2(n38063), .ZN(n38062) );
  INV_X1 U37741 ( .A(n38062), .ZN(n2541) );
  OAI22_X1 U37742 ( .A1(n38064), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[37][7] ), .B2(n38063), .ZN(n38065) );
  INV_X1 U37743 ( .A(n38065), .ZN(n2540) );
  NOR2_X1 U37744 ( .A1(n38880), .A2(n38156), .ZN(n38073) );
  INV_X1 U37745 ( .A(n38073), .ZN(n38074) );
  OAI22_X1 U37746 ( .A1(n38074), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[38][0] ), .B2(n38073), .ZN(n38066) );
  INV_X1 U37747 ( .A(n38066), .ZN(n2539) );
  OAI22_X1 U37748 ( .A1(n38074), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[38][1] ), .B2(n38073), .ZN(n38067) );
  INV_X1 U37749 ( .A(n38067), .ZN(n2538) );
  OAI22_X1 U37750 ( .A1(n38074), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[38][2] ), .B2(n38073), .ZN(n38068) );
  INV_X1 U37751 ( .A(n38068), .ZN(n2537) );
  OAI22_X1 U37752 ( .A1(n38074), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[38][3] ), .B2(n38073), .ZN(n38069) );
  INV_X1 U37753 ( .A(n38069), .ZN(n2536) );
  OAI22_X1 U37754 ( .A1(n38074), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[38][4] ), .B2(n38073), .ZN(n38070) );
  INV_X1 U37755 ( .A(n38070), .ZN(n2535) );
  OAI22_X1 U37756 ( .A1(n38074), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[38][5] ), .B2(n38073), .ZN(n38071) );
  INV_X1 U37757 ( .A(n38071), .ZN(n2534) );
  OAI22_X1 U37758 ( .A1(n38074), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[38][6] ), .B2(n38073), .ZN(n38072) );
  INV_X1 U37759 ( .A(n38072), .ZN(n2533) );
  OAI22_X1 U37760 ( .A1(n38074), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[38][7] ), .B2(n38073), .ZN(n38075) );
  INV_X1 U37761 ( .A(n38075), .ZN(n2532) );
  NOR2_X1 U37762 ( .A1(n38891), .A2(n38156), .ZN(n38083) );
  INV_X1 U37763 ( .A(n38083), .ZN(n38084) );
  OAI22_X1 U37764 ( .A1(n38084), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[39][0] ), .B2(n38083), .ZN(n38076) );
  INV_X1 U37765 ( .A(n38076), .ZN(n2531) );
  OAI22_X1 U37766 ( .A1(n38084), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[39][1] ), .B2(n38083), .ZN(n38077) );
  INV_X1 U37767 ( .A(n38077), .ZN(n2530) );
  OAI22_X1 U37768 ( .A1(n38084), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[39][2] ), .B2(n38083), .ZN(n38078) );
  INV_X1 U37769 ( .A(n38078), .ZN(n2529) );
  OAI22_X1 U37770 ( .A1(n38084), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[39][3] ), .B2(n38083), .ZN(n38079) );
  INV_X1 U37771 ( .A(n38079), .ZN(n2528) );
  OAI22_X1 U37772 ( .A1(n38084), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[39][4] ), .B2(n38083), .ZN(n38080) );
  INV_X1 U37773 ( .A(n38080), .ZN(n2527) );
  OAI22_X1 U37774 ( .A1(n38084), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[39][5] ), .B2(n38083), .ZN(n38081) );
  INV_X1 U37775 ( .A(n38081), .ZN(n2526) );
  OAI22_X1 U37776 ( .A1(n38084), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[39][6] ), .B2(n38083), .ZN(n38082) );
  INV_X1 U37777 ( .A(n38082), .ZN(n2525) );
  OAI22_X1 U37778 ( .A1(n38084), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[39][7] ), .B2(n38083), .ZN(n38085) );
  INV_X1 U37779 ( .A(n38085), .ZN(n2524) );
  NOR2_X1 U37780 ( .A1(n38902), .A2(n38156), .ZN(n38093) );
  INV_X1 U37781 ( .A(n38093), .ZN(n38094) );
  OAI22_X1 U37782 ( .A1(n38094), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[40][0] ), .B2(n38093), .ZN(n38086) );
  INV_X1 U37783 ( .A(n38086), .ZN(n2523) );
  OAI22_X1 U37784 ( .A1(n38094), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[40][1] ), .B2(n38093), .ZN(n38087) );
  INV_X1 U37785 ( .A(n38087), .ZN(n2522) );
  OAI22_X1 U37786 ( .A1(n38094), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[40][2] ), .B2(n38093), .ZN(n38088) );
  INV_X1 U37787 ( .A(n38088), .ZN(n2521) );
  OAI22_X1 U37788 ( .A1(n38094), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[40][3] ), .B2(n38093), .ZN(n38089) );
  INV_X1 U37789 ( .A(n38089), .ZN(n2520) );
  OAI22_X1 U37790 ( .A1(n38094), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[40][4] ), .B2(n38093), .ZN(n38090) );
  INV_X1 U37791 ( .A(n38090), .ZN(n2519) );
  OAI22_X1 U37792 ( .A1(n38094), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[40][5] ), .B2(n38093), .ZN(n38091) );
  INV_X1 U37793 ( .A(n38091), .ZN(n2518) );
  OAI22_X1 U37794 ( .A1(n38094), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[40][6] ), .B2(n38093), .ZN(n38092) );
  INV_X1 U37795 ( .A(n38092), .ZN(n2517) );
  OAI22_X1 U37796 ( .A1(n38094), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[40][7] ), .B2(n38093), .ZN(n38095) );
  INV_X1 U37797 ( .A(n38095), .ZN(n2516) );
  NOR2_X1 U37798 ( .A1(n38913), .A2(n38156), .ZN(n38103) );
  INV_X1 U37799 ( .A(n38103), .ZN(n38104) );
  OAI22_X1 U37800 ( .A1(n38104), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[41][0] ), .B2(n38103), .ZN(n38096) );
  INV_X1 U37801 ( .A(n38096), .ZN(n2515) );
  OAI22_X1 U37802 ( .A1(n38104), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[41][1] ), .B2(n38103), .ZN(n38097) );
  INV_X1 U37803 ( .A(n38097), .ZN(n2514) );
  OAI22_X1 U37804 ( .A1(n38104), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[41][2] ), .B2(n38103), .ZN(n38098) );
  INV_X1 U37805 ( .A(n38098), .ZN(n2513) );
  OAI22_X1 U37806 ( .A1(n38104), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[41][3] ), .B2(n38103), .ZN(n38099) );
  INV_X1 U37807 ( .A(n38099), .ZN(n2512) );
  OAI22_X1 U37808 ( .A1(n38104), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[41][4] ), .B2(n38103), .ZN(n38100) );
  INV_X1 U37809 ( .A(n38100), .ZN(n2511) );
  OAI22_X1 U37810 ( .A1(n38104), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[41][5] ), .B2(n38103), .ZN(n38101) );
  INV_X1 U37811 ( .A(n38101), .ZN(n2510) );
  OAI22_X1 U37812 ( .A1(n38104), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[41][6] ), .B2(n38103), .ZN(n38102) );
  INV_X1 U37813 ( .A(n38102), .ZN(n2509) );
  OAI22_X1 U37814 ( .A1(n38104), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[41][7] ), .B2(n38103), .ZN(n38105) );
  INV_X1 U37815 ( .A(n38105), .ZN(n2508) );
  NOR2_X1 U37816 ( .A1(n38924), .A2(n38156), .ZN(n38113) );
  INV_X1 U37817 ( .A(n38113), .ZN(n38114) );
  OAI22_X1 U37818 ( .A1(n38114), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[42][0] ), .B2(n38113), .ZN(n38106) );
  INV_X1 U37819 ( .A(n38106), .ZN(n2507) );
  OAI22_X1 U37820 ( .A1(n38114), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[42][1] ), .B2(n38113), .ZN(n38107) );
  INV_X1 U37821 ( .A(n38107), .ZN(n2506) );
  OAI22_X1 U37822 ( .A1(n38114), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[42][2] ), .B2(n38113), .ZN(n38108) );
  INV_X1 U37823 ( .A(n38108), .ZN(n2505) );
  OAI22_X1 U37824 ( .A1(n38114), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[42][3] ), .B2(n38113), .ZN(n38109) );
  INV_X1 U37825 ( .A(n38109), .ZN(n2504) );
  OAI22_X1 U37826 ( .A1(n38114), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[42][4] ), .B2(n38113), .ZN(n38110) );
  INV_X1 U37827 ( .A(n38110), .ZN(n2503) );
  OAI22_X1 U37828 ( .A1(n38114), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[42][5] ), .B2(n38113), .ZN(n38111) );
  INV_X1 U37829 ( .A(n38111), .ZN(n2502) );
  OAI22_X1 U37830 ( .A1(n38114), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[42][6] ), .B2(n38113), .ZN(n38112) );
  INV_X1 U37831 ( .A(n38112), .ZN(n2501) );
  OAI22_X1 U37832 ( .A1(n38114), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[42][7] ), .B2(n38113), .ZN(n38115) );
  INV_X1 U37833 ( .A(n38115), .ZN(n2500) );
  NOR2_X1 U37834 ( .A1(n38935), .A2(n38156), .ZN(n38123) );
  INV_X1 U37835 ( .A(n38123), .ZN(n38124) );
  OAI22_X1 U37836 ( .A1(n38124), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[43][0] ), .B2(n38123), .ZN(n38116) );
  INV_X1 U37837 ( .A(n38116), .ZN(n2499) );
  OAI22_X1 U37838 ( .A1(n38124), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[43][1] ), .B2(n38123), .ZN(n38117) );
  INV_X1 U37839 ( .A(n38117), .ZN(n2498) );
  OAI22_X1 U37840 ( .A1(n38124), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[43][2] ), .B2(n38123), .ZN(n38118) );
  INV_X1 U37841 ( .A(n38118), .ZN(n2497) );
  OAI22_X1 U37842 ( .A1(n38124), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[43][3] ), .B2(n38123), .ZN(n38119) );
  INV_X1 U37843 ( .A(n38119), .ZN(n2496) );
  OAI22_X1 U37844 ( .A1(n38124), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[43][4] ), .B2(n38123), .ZN(n38120) );
  INV_X1 U37845 ( .A(n38120), .ZN(n2495) );
  OAI22_X1 U37846 ( .A1(n38124), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[43][5] ), .B2(n38123), .ZN(n38121) );
  INV_X1 U37847 ( .A(n38121), .ZN(n2494) );
  OAI22_X1 U37848 ( .A1(n38124), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[43][6] ), .B2(n38123), .ZN(n38122) );
  INV_X1 U37849 ( .A(n38122), .ZN(n2493) );
  OAI22_X1 U37850 ( .A1(n38124), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[43][7] ), .B2(n38123), .ZN(n38125) );
  INV_X1 U37851 ( .A(n38125), .ZN(n2492) );
  NOR2_X1 U37852 ( .A1(n38946), .A2(n38156), .ZN(n38133) );
  INV_X1 U37853 ( .A(n38133), .ZN(n38134) );
  OAI22_X1 U37854 ( .A1(n38134), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[44][0] ), .B2(n38133), .ZN(n38126) );
  INV_X1 U37855 ( .A(n38126), .ZN(n2491) );
  OAI22_X1 U37856 ( .A1(n38134), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[44][1] ), .B2(n38133), .ZN(n38127) );
  INV_X1 U37857 ( .A(n38127), .ZN(n2490) );
  OAI22_X1 U37858 ( .A1(n38134), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[44][2] ), .B2(n38133), .ZN(n38128) );
  INV_X1 U37859 ( .A(n38128), .ZN(n2489) );
  OAI22_X1 U37860 ( .A1(n38134), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[44][3] ), .B2(n38133), .ZN(n38129) );
  INV_X1 U37861 ( .A(n38129), .ZN(n2488) );
  OAI22_X1 U37862 ( .A1(n38134), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[44][4] ), .B2(n38133), .ZN(n38130) );
  INV_X1 U37863 ( .A(n38130), .ZN(n2487) );
  OAI22_X1 U37864 ( .A1(n38134), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[44][5] ), .B2(n38133), .ZN(n38131) );
  INV_X1 U37865 ( .A(n38131), .ZN(n2486) );
  OAI22_X1 U37866 ( .A1(n38134), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[44][6] ), .B2(n38133), .ZN(n38132) );
  INV_X1 U37867 ( .A(n38132), .ZN(n2485) );
  OAI22_X1 U37868 ( .A1(n38134), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[44][7] ), .B2(n38133), .ZN(n38135) );
  INV_X1 U37869 ( .A(n38135), .ZN(n2484) );
  NOR2_X1 U37870 ( .A1(n38957), .A2(n38156), .ZN(n38143) );
  INV_X1 U37871 ( .A(n38143), .ZN(n38144) );
  OAI22_X1 U37872 ( .A1(n38144), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[45][0] ), .B2(n38143), .ZN(n38136) );
  INV_X1 U37873 ( .A(n38136), .ZN(n2483) );
  OAI22_X1 U37874 ( .A1(n38144), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[45][1] ), .B2(n38143), .ZN(n38137) );
  INV_X1 U37875 ( .A(n38137), .ZN(n2482) );
  OAI22_X1 U37876 ( .A1(n38144), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[45][2] ), .B2(n38143), .ZN(n38138) );
  INV_X1 U37877 ( .A(n38138), .ZN(n2481) );
  OAI22_X1 U37878 ( .A1(n38144), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[45][3] ), .B2(n38143), .ZN(n38139) );
  INV_X1 U37879 ( .A(n38139), .ZN(n2480) );
  OAI22_X1 U37880 ( .A1(n38144), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[45][4] ), .B2(n38143), .ZN(n38140) );
  INV_X1 U37881 ( .A(n38140), .ZN(n2479) );
  OAI22_X1 U37882 ( .A1(n38144), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[45][5] ), .B2(n38143), .ZN(n38141) );
  INV_X1 U37883 ( .A(n38141), .ZN(n2478) );
  OAI22_X1 U37884 ( .A1(n38144), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[45][6] ), .B2(n38143), .ZN(n38142) );
  INV_X1 U37885 ( .A(n38142), .ZN(n2477) );
  OAI22_X1 U37886 ( .A1(n38144), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[45][7] ), .B2(n38143), .ZN(n38145) );
  INV_X1 U37887 ( .A(n38145), .ZN(n2476) );
  NOR2_X1 U37888 ( .A1(n38968), .A2(n38156), .ZN(n38153) );
  INV_X1 U37889 ( .A(n38153), .ZN(n38154) );
  OAI22_X1 U37890 ( .A1(n38154), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[46][0] ), .B2(n38153), .ZN(n38146) );
  INV_X1 U37891 ( .A(n38146), .ZN(n2475) );
  OAI22_X1 U37892 ( .A1(n38154), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[46][1] ), .B2(n38153), .ZN(n38147) );
  INV_X1 U37893 ( .A(n38147), .ZN(n2474) );
  OAI22_X1 U37894 ( .A1(n38154), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[46][2] ), .B2(n38153), .ZN(n38148) );
  INV_X1 U37895 ( .A(n38148), .ZN(n2473) );
  OAI22_X1 U37896 ( .A1(n38154), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[46][3] ), .B2(n38153), .ZN(n38149) );
  INV_X1 U37897 ( .A(n38149), .ZN(n2472) );
  OAI22_X1 U37898 ( .A1(n38154), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[46][4] ), .B2(n38153), .ZN(n38150) );
  INV_X1 U37899 ( .A(n38150), .ZN(n2471) );
  OAI22_X1 U37900 ( .A1(n38154), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[46][5] ), .B2(n38153), .ZN(n38151) );
  INV_X1 U37901 ( .A(n38151), .ZN(n2470) );
  OAI22_X1 U37902 ( .A1(n38154), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[46][6] ), .B2(n38153), .ZN(n38152) );
  INV_X1 U37903 ( .A(n38152), .ZN(n2469) );
  OAI22_X1 U37904 ( .A1(n38154), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[46][7] ), .B2(n38153), .ZN(n38155) );
  INV_X1 U37905 ( .A(n38155), .ZN(n2468) );
  NOR2_X1 U37906 ( .A1(n38803), .A2(n38156), .ZN(n38164) );
  INV_X1 U37907 ( .A(n38164), .ZN(n38165) );
  OAI22_X1 U37908 ( .A1(n38165), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[47][0] ), .B2(n38164), .ZN(n38157) );
  INV_X1 U37909 ( .A(n38157), .ZN(n2467) );
  OAI22_X1 U37910 ( .A1(n38165), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[47][1] ), .B2(n38164), .ZN(n38158) );
  INV_X1 U37911 ( .A(n38158), .ZN(n2466) );
  OAI22_X1 U37912 ( .A1(n38165), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[47][2] ), .B2(n38164), .ZN(n38159) );
  INV_X1 U37913 ( .A(n38159), .ZN(n2465) );
  OAI22_X1 U37914 ( .A1(n38165), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[47][3] ), .B2(n38164), .ZN(n38160) );
  INV_X1 U37915 ( .A(n38160), .ZN(n2464) );
  OAI22_X1 U37916 ( .A1(n38165), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[47][4] ), .B2(n38164), .ZN(n38161) );
  INV_X1 U37917 ( .A(n38161), .ZN(n2463) );
  OAI22_X1 U37918 ( .A1(n38165), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[47][5] ), .B2(n38164), .ZN(n38162) );
  INV_X1 U37919 ( .A(n38162), .ZN(n2462) );
  OAI22_X1 U37920 ( .A1(n38165), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[47][6] ), .B2(n38164), .ZN(n38163) );
  INV_X1 U37921 ( .A(n38163), .ZN(n2461) );
  OAI22_X1 U37922 ( .A1(n38165), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[47][7] ), .B2(n38164), .ZN(n38166) );
  INV_X1 U37923 ( .A(n38166), .ZN(n2460) );
  NOR2_X1 U37924 ( .A1(n38307), .A2(n38814), .ZN(n38174) );
  INV_X1 U37925 ( .A(n38174), .ZN(n38175) );
  OAI22_X1 U37926 ( .A1(n38175), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[48][0] ), .B2(n38174), .ZN(n38167) );
  INV_X1 U37927 ( .A(n38167), .ZN(n2459) );
  OAI22_X1 U37928 ( .A1(n38175), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[48][1] ), .B2(n38174), .ZN(n38168) );
  INV_X1 U37929 ( .A(n38168), .ZN(n2458) );
  OAI22_X1 U37930 ( .A1(n38175), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[48][2] ), .B2(n38174), .ZN(n38169) );
  INV_X1 U37931 ( .A(n38169), .ZN(n2457) );
  OAI22_X1 U37932 ( .A1(n38175), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[48][3] ), .B2(n38174), .ZN(n38170) );
  INV_X1 U37933 ( .A(n38170), .ZN(n2456) );
  OAI22_X1 U37934 ( .A1(n38175), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[48][4] ), .B2(n38174), .ZN(n38171) );
  INV_X1 U37935 ( .A(n38171), .ZN(n2455) );
  OAI22_X1 U37936 ( .A1(n38175), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[48][5] ), .B2(n38174), .ZN(n38172) );
  INV_X1 U37937 ( .A(n38172), .ZN(n2454) );
  OAI22_X1 U37938 ( .A1(n38175), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[48][6] ), .B2(n38174), .ZN(n38173) );
  INV_X1 U37939 ( .A(n38173), .ZN(n2453) );
  OAI22_X1 U37940 ( .A1(n38175), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[48][7] ), .B2(n38174), .ZN(n38176) );
  INV_X1 U37941 ( .A(n38176), .ZN(n2452) );
  NOR2_X1 U37942 ( .A1(n38307), .A2(n38825), .ZN(n38184) );
  INV_X1 U37943 ( .A(n38184), .ZN(n38185) );
  OAI22_X1 U37944 ( .A1(n38185), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[49][0] ), .B2(n38184), .ZN(n38177) );
  INV_X1 U37945 ( .A(n38177), .ZN(n2451) );
  OAI22_X1 U37946 ( .A1(n38185), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[49][1] ), .B2(n38184), .ZN(n38178) );
  INV_X1 U37947 ( .A(n38178), .ZN(n2450) );
  OAI22_X1 U37948 ( .A1(n38185), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[49][2] ), .B2(n38184), .ZN(n38179) );
  INV_X1 U37949 ( .A(n38179), .ZN(n2449) );
  OAI22_X1 U37950 ( .A1(n38185), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[49][3] ), .B2(n38184), .ZN(n38180) );
  INV_X1 U37951 ( .A(n38180), .ZN(n2448) );
  OAI22_X1 U37952 ( .A1(n38185), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[49][4] ), .B2(n38184), .ZN(n38181) );
  INV_X1 U37953 ( .A(n38181), .ZN(n2447) );
  OAI22_X1 U37954 ( .A1(n38185), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[49][5] ), .B2(n38184), .ZN(n38182) );
  INV_X1 U37955 ( .A(n38182), .ZN(n2446) );
  OAI22_X1 U37956 ( .A1(n38185), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[49][6] ), .B2(n38184), .ZN(n38183) );
  INV_X1 U37957 ( .A(n38183), .ZN(n2445) );
  OAI22_X1 U37958 ( .A1(n38185), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[49][7] ), .B2(n38184), .ZN(n38186) );
  INV_X1 U37959 ( .A(n38186), .ZN(n2444) );
  NOR2_X1 U37960 ( .A1(n38307), .A2(n38836), .ZN(n38194) );
  INV_X1 U37961 ( .A(n38194), .ZN(n38195) );
  OAI22_X1 U37962 ( .A1(n38195), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[50][0] ), .B2(n38194), .ZN(n38187) );
  INV_X1 U37963 ( .A(n38187), .ZN(n2443) );
  OAI22_X1 U37964 ( .A1(n38195), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[50][1] ), .B2(n38194), .ZN(n38188) );
  INV_X1 U37965 ( .A(n38188), .ZN(n2442) );
  OAI22_X1 U37966 ( .A1(n38195), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[50][2] ), .B2(n38194), .ZN(n38189) );
  INV_X1 U37967 ( .A(n38189), .ZN(n2441) );
  OAI22_X1 U37968 ( .A1(n38195), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[50][3] ), .B2(n38194), .ZN(n38190) );
  INV_X1 U37969 ( .A(n38190), .ZN(n2440) );
  OAI22_X1 U37970 ( .A1(n38195), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[50][4] ), .B2(n38194), .ZN(n38191) );
  INV_X1 U37971 ( .A(n38191), .ZN(n2439) );
  OAI22_X1 U37972 ( .A1(n38195), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[50][5] ), .B2(n38194), .ZN(n38192) );
  INV_X1 U37973 ( .A(n38192), .ZN(n2438) );
  OAI22_X1 U37974 ( .A1(n38195), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[50][6] ), .B2(n38194), .ZN(n38193) );
  INV_X1 U37975 ( .A(n38193), .ZN(n2437) );
  OAI22_X1 U37976 ( .A1(n38195), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[50][7] ), .B2(n38194), .ZN(n38196) );
  INV_X1 U37977 ( .A(n38196), .ZN(n2436) );
  NOR2_X1 U37978 ( .A1(n38307), .A2(n38847), .ZN(n38204) );
  INV_X1 U37979 ( .A(n38204), .ZN(n38205) );
  OAI22_X1 U37980 ( .A1(n38205), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[51][0] ), .B2(n38204), .ZN(n38197) );
  INV_X1 U37981 ( .A(n38197), .ZN(n2435) );
  OAI22_X1 U37982 ( .A1(n38205), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[51][1] ), .B2(n38204), .ZN(n38198) );
  INV_X1 U37983 ( .A(n38198), .ZN(n2434) );
  OAI22_X1 U37984 ( .A1(n38205), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[51][2] ), .B2(n38204), .ZN(n38199) );
  INV_X1 U37985 ( .A(n38199), .ZN(n2433) );
  OAI22_X1 U37986 ( .A1(n38205), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[51][3] ), .B2(n38204), .ZN(n38200) );
  INV_X1 U37987 ( .A(n38200), .ZN(n2432) );
  OAI22_X1 U37988 ( .A1(n38205), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[51][4] ), .B2(n38204), .ZN(n38201) );
  INV_X1 U37989 ( .A(n38201), .ZN(n2431) );
  OAI22_X1 U37990 ( .A1(n38205), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[51][5] ), .B2(n38204), .ZN(n38202) );
  INV_X1 U37991 ( .A(n38202), .ZN(n2430) );
  OAI22_X1 U37992 ( .A1(n38205), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[51][6] ), .B2(n38204), .ZN(n38203) );
  INV_X1 U37993 ( .A(n38203), .ZN(n2429) );
  OAI22_X1 U37994 ( .A1(n38205), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[51][7] ), .B2(n38204), .ZN(n38206) );
  INV_X1 U37995 ( .A(n38206), .ZN(n2428) );
  NOR2_X1 U37996 ( .A1(n38307), .A2(n38858), .ZN(n38214) );
  INV_X1 U37997 ( .A(n38214), .ZN(n38215) );
  OAI22_X1 U37998 ( .A1(n38215), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[52][0] ), .B2(n38214), .ZN(n38207) );
  INV_X1 U37999 ( .A(n38207), .ZN(n2427) );
  OAI22_X1 U38000 ( .A1(n38215), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[52][1] ), .B2(n38214), .ZN(n38208) );
  INV_X1 U38001 ( .A(n38208), .ZN(n2426) );
  OAI22_X1 U38002 ( .A1(n38215), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[52][2] ), .B2(n38214), .ZN(n38209) );
  INV_X1 U38003 ( .A(n38209), .ZN(n2425) );
  OAI22_X1 U38004 ( .A1(n38215), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[52][3] ), .B2(n38214), .ZN(n38210) );
  INV_X1 U38005 ( .A(n38210), .ZN(n2424) );
  OAI22_X1 U38006 ( .A1(n38215), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[52][4] ), .B2(n38214), .ZN(n38211) );
  INV_X1 U38007 ( .A(n38211), .ZN(n2423) );
  OAI22_X1 U38008 ( .A1(n38215), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[52][5] ), .B2(n38214), .ZN(n38212) );
  INV_X1 U38009 ( .A(n38212), .ZN(n2422) );
  OAI22_X1 U38010 ( .A1(n38215), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[52][6] ), .B2(n38214), .ZN(n38213) );
  INV_X1 U38011 ( .A(n38213), .ZN(n2421) );
  OAI22_X1 U38012 ( .A1(n38215), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[52][7] ), .B2(n38214), .ZN(n38216) );
  INV_X1 U38013 ( .A(n38216), .ZN(n2420) );
  NOR2_X1 U38014 ( .A1(n38307), .A2(n38869), .ZN(n38224) );
  INV_X1 U38015 ( .A(n38224), .ZN(n38225) );
  OAI22_X1 U38016 ( .A1(n38225), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[53][0] ), .B2(n38224), .ZN(n38217) );
  INV_X1 U38017 ( .A(n38217), .ZN(n2419) );
  OAI22_X1 U38018 ( .A1(n38225), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[53][1] ), .B2(n38224), .ZN(n38218) );
  INV_X1 U38019 ( .A(n38218), .ZN(n2418) );
  OAI22_X1 U38020 ( .A1(n38225), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[53][2] ), .B2(n38224), .ZN(n38219) );
  INV_X1 U38021 ( .A(n38219), .ZN(n2417) );
  OAI22_X1 U38022 ( .A1(n38225), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[53][3] ), .B2(n38224), .ZN(n38220) );
  INV_X1 U38023 ( .A(n38220), .ZN(n2416) );
  OAI22_X1 U38024 ( .A1(n38225), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[53][4] ), .B2(n38224), .ZN(n38221) );
  INV_X1 U38025 ( .A(n38221), .ZN(n2415) );
  OAI22_X1 U38026 ( .A1(n38225), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[53][5] ), .B2(n38224), .ZN(n38222) );
  INV_X1 U38027 ( .A(n38222), .ZN(n2414) );
  OAI22_X1 U38028 ( .A1(n38225), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[53][6] ), .B2(n38224), .ZN(n38223) );
  INV_X1 U38029 ( .A(n38223), .ZN(n2413) );
  OAI22_X1 U38030 ( .A1(n38225), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[53][7] ), .B2(n38224), .ZN(n38226) );
  INV_X1 U38031 ( .A(n38226), .ZN(n2412) );
  NOR2_X1 U38032 ( .A1(n38307), .A2(n38880), .ZN(n38234) );
  INV_X1 U38033 ( .A(n38234), .ZN(n38235) );
  OAI22_X1 U38034 ( .A1(n38235), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[54][0] ), .B2(n38234), .ZN(n38227) );
  INV_X1 U38035 ( .A(n38227), .ZN(n2411) );
  OAI22_X1 U38036 ( .A1(n38235), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[54][1] ), .B2(n38234), .ZN(n38228) );
  INV_X1 U38037 ( .A(n38228), .ZN(n2410) );
  OAI22_X1 U38038 ( .A1(n38235), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[54][2] ), .B2(n38234), .ZN(n38229) );
  INV_X1 U38039 ( .A(n38229), .ZN(n2409) );
  OAI22_X1 U38040 ( .A1(n38235), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[54][3] ), .B2(n38234), .ZN(n38230) );
  INV_X1 U38041 ( .A(n38230), .ZN(n2408) );
  OAI22_X1 U38042 ( .A1(n38235), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[54][4] ), .B2(n38234), .ZN(n38231) );
  INV_X1 U38043 ( .A(n38231), .ZN(n2407) );
  OAI22_X1 U38044 ( .A1(n38235), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[54][5] ), .B2(n38234), .ZN(n38232) );
  INV_X1 U38045 ( .A(n38232), .ZN(n2406) );
  OAI22_X1 U38046 ( .A1(n38235), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[54][6] ), .B2(n38234), .ZN(n38233) );
  INV_X1 U38047 ( .A(n38233), .ZN(n2405) );
  OAI22_X1 U38048 ( .A1(n38235), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[54][7] ), .B2(n38234), .ZN(n38236) );
  INV_X1 U38049 ( .A(n38236), .ZN(n2404) );
  NOR2_X1 U38050 ( .A1(n38891), .A2(n38307), .ZN(n38244) );
  INV_X1 U38051 ( .A(n38244), .ZN(n38245) );
  OAI22_X1 U38052 ( .A1(n38245), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[55][0] ), .B2(n38244), .ZN(n38237) );
  INV_X1 U38053 ( .A(n38237), .ZN(n2403) );
  OAI22_X1 U38054 ( .A1(n38245), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[55][1] ), .B2(n38244), .ZN(n38238) );
  INV_X1 U38055 ( .A(n38238), .ZN(n2402) );
  OAI22_X1 U38056 ( .A1(n38245), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[55][2] ), .B2(n38244), .ZN(n38239) );
  INV_X1 U38057 ( .A(n38239), .ZN(n2401) );
  OAI22_X1 U38058 ( .A1(n38245), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[55][3] ), .B2(n38244), .ZN(n38240) );
  INV_X1 U38059 ( .A(n38240), .ZN(n2400) );
  OAI22_X1 U38060 ( .A1(n38245), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[55][4] ), .B2(n38244), .ZN(n38241) );
  INV_X1 U38061 ( .A(n38241), .ZN(n2399) );
  OAI22_X1 U38062 ( .A1(n38245), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[55][5] ), .B2(n38244), .ZN(n38242) );
  INV_X1 U38063 ( .A(n38242), .ZN(n2398) );
  OAI22_X1 U38064 ( .A1(n38245), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[55][6] ), .B2(n38244), .ZN(n38243) );
  INV_X1 U38065 ( .A(n38243), .ZN(n2397) );
  OAI22_X1 U38066 ( .A1(n38245), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[55][7] ), .B2(n38244), .ZN(n38246) );
  INV_X1 U38067 ( .A(n38246), .ZN(n2396) );
  NOR2_X1 U38068 ( .A1(n38307), .A2(n38902), .ZN(n38254) );
  INV_X1 U38069 ( .A(n38254), .ZN(n38255) );
  OAI22_X1 U38070 ( .A1(n38255), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[56][0] ), .B2(n38254), .ZN(n38247) );
  INV_X1 U38071 ( .A(n38247), .ZN(n2395) );
  OAI22_X1 U38072 ( .A1(n38255), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[56][1] ), .B2(n38254), .ZN(n38248) );
  INV_X1 U38073 ( .A(n38248), .ZN(n2394) );
  OAI22_X1 U38074 ( .A1(n38255), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[56][2] ), .B2(n38254), .ZN(n38249) );
  INV_X1 U38075 ( .A(n38249), .ZN(n2393) );
  OAI22_X1 U38076 ( .A1(n38255), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[56][3] ), .B2(n38254), .ZN(n38250) );
  INV_X1 U38077 ( .A(n38250), .ZN(n2392) );
  OAI22_X1 U38078 ( .A1(n38255), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[56][4] ), .B2(n38254), .ZN(n38251) );
  INV_X1 U38079 ( .A(n38251), .ZN(n2391) );
  OAI22_X1 U38080 ( .A1(n38255), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[56][5] ), .B2(n38254), .ZN(n38252) );
  INV_X1 U38081 ( .A(n38252), .ZN(n2390) );
  OAI22_X1 U38082 ( .A1(n38255), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[56][6] ), .B2(n38254), .ZN(n38253) );
  INV_X1 U38083 ( .A(n38253), .ZN(n2389) );
  OAI22_X1 U38084 ( .A1(n38255), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[56][7] ), .B2(n38254), .ZN(n38256) );
  INV_X1 U38085 ( .A(n38256), .ZN(n2388) );
  NOR2_X1 U38086 ( .A1(n38307), .A2(n38913), .ZN(n38264) );
  INV_X1 U38087 ( .A(n38264), .ZN(n38265) );
  OAI22_X1 U38088 ( .A1(n38265), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[57][0] ), .B2(n38264), .ZN(n38257) );
  INV_X1 U38089 ( .A(n38257), .ZN(n2387) );
  OAI22_X1 U38090 ( .A1(n38265), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[57][1] ), .B2(n38264), .ZN(n38258) );
  INV_X1 U38091 ( .A(n38258), .ZN(n2386) );
  OAI22_X1 U38092 ( .A1(n38265), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[57][2] ), .B2(n38264), .ZN(n38259) );
  INV_X1 U38093 ( .A(n38259), .ZN(n2385) );
  OAI22_X1 U38094 ( .A1(n38265), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[57][3] ), .B2(n38264), .ZN(n38260) );
  INV_X1 U38095 ( .A(n38260), .ZN(n2384) );
  OAI22_X1 U38096 ( .A1(n38265), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[57][4] ), .B2(n38264), .ZN(n38261) );
  INV_X1 U38097 ( .A(n38261), .ZN(n2383) );
  OAI22_X1 U38098 ( .A1(n38265), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[57][5] ), .B2(n38264), .ZN(n38262) );
  INV_X1 U38099 ( .A(n38262), .ZN(n2382) );
  OAI22_X1 U38100 ( .A1(n38265), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[57][6] ), .B2(n38264), .ZN(n38263) );
  INV_X1 U38101 ( .A(n38263), .ZN(n2381) );
  OAI22_X1 U38102 ( .A1(n38265), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[57][7] ), .B2(n38264), .ZN(n38266) );
  INV_X1 U38103 ( .A(n38266), .ZN(n2380) );
  NOR2_X1 U38104 ( .A1(n38307), .A2(n38924), .ZN(n38274) );
  INV_X1 U38105 ( .A(n38274), .ZN(n38275) );
  OAI22_X1 U38106 ( .A1(n38275), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[58][0] ), .B2(n38274), .ZN(n38267) );
  INV_X1 U38107 ( .A(n38267), .ZN(n2379) );
  OAI22_X1 U38108 ( .A1(n38275), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[58][1] ), .B2(n38274), .ZN(n38268) );
  INV_X1 U38109 ( .A(n38268), .ZN(n2378) );
  OAI22_X1 U38110 ( .A1(n38275), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[58][2] ), .B2(n38274), .ZN(n38269) );
  INV_X1 U38111 ( .A(n38269), .ZN(n2377) );
  OAI22_X1 U38112 ( .A1(n38275), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[58][3] ), .B2(n38274), .ZN(n38270) );
  INV_X1 U38113 ( .A(n38270), .ZN(n2376) );
  OAI22_X1 U38114 ( .A1(n38275), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[58][4] ), .B2(n38274), .ZN(n38271) );
  INV_X1 U38115 ( .A(n38271), .ZN(n2375) );
  OAI22_X1 U38116 ( .A1(n38275), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[58][5] ), .B2(n38274), .ZN(n38272) );
  INV_X1 U38117 ( .A(n38272), .ZN(n2374) );
  OAI22_X1 U38118 ( .A1(n38275), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[58][6] ), .B2(n38274), .ZN(n38273) );
  INV_X1 U38119 ( .A(n38273), .ZN(n2373) );
  OAI22_X1 U38120 ( .A1(n38275), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[58][7] ), .B2(n38274), .ZN(n38276) );
  INV_X1 U38121 ( .A(n38276), .ZN(n2372) );
  NOR2_X1 U38122 ( .A1(n38307), .A2(n38935), .ZN(n38284) );
  INV_X1 U38123 ( .A(n38284), .ZN(n38285) );
  OAI22_X1 U38124 ( .A1(n38285), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[59][0] ), .B2(n38284), .ZN(n38277) );
  INV_X1 U38125 ( .A(n38277), .ZN(n2371) );
  OAI22_X1 U38126 ( .A1(n38285), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[59][1] ), .B2(n38284), .ZN(n38278) );
  INV_X1 U38127 ( .A(n38278), .ZN(n2370) );
  OAI22_X1 U38128 ( .A1(n38285), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[59][2] ), .B2(n38284), .ZN(n38279) );
  INV_X1 U38129 ( .A(n38279), .ZN(n2369) );
  OAI22_X1 U38130 ( .A1(n38285), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[59][3] ), .B2(n38284), .ZN(n38280) );
  INV_X1 U38131 ( .A(n38280), .ZN(n2368) );
  OAI22_X1 U38132 ( .A1(n38285), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[59][4] ), .B2(n38284), .ZN(n38281) );
  INV_X1 U38133 ( .A(n38281), .ZN(n2367) );
  OAI22_X1 U38134 ( .A1(n38285), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[59][5] ), .B2(n38284), .ZN(n38282) );
  INV_X1 U38135 ( .A(n38282), .ZN(n2366) );
  OAI22_X1 U38136 ( .A1(n38285), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[59][6] ), .B2(n38284), .ZN(n38283) );
  INV_X1 U38137 ( .A(n38283), .ZN(n2365) );
  OAI22_X1 U38138 ( .A1(n38285), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[59][7] ), .B2(n38284), .ZN(n38286) );
  INV_X1 U38139 ( .A(n38286), .ZN(n2364) );
  NOR2_X1 U38140 ( .A1(n38307), .A2(n38946), .ZN(n38294) );
  INV_X1 U38141 ( .A(n38294), .ZN(n38295) );
  OAI22_X1 U38142 ( .A1(n38295), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[60][0] ), .B2(n38294), .ZN(n38287) );
  INV_X1 U38143 ( .A(n38287), .ZN(n2363) );
  OAI22_X1 U38144 ( .A1(n38295), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[60][1] ), .B2(n38294), .ZN(n38288) );
  INV_X1 U38145 ( .A(n38288), .ZN(n2362) );
  OAI22_X1 U38146 ( .A1(n38295), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[60][2] ), .B2(n38294), .ZN(n38289) );
  INV_X1 U38147 ( .A(n38289), .ZN(n2361) );
  OAI22_X1 U38148 ( .A1(n38295), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[60][3] ), .B2(n38294), .ZN(n38290) );
  INV_X1 U38149 ( .A(n38290), .ZN(n2360) );
  OAI22_X1 U38150 ( .A1(n38295), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[60][4] ), .B2(n38294), .ZN(n38291) );
  INV_X1 U38151 ( .A(n38291), .ZN(n2359) );
  OAI22_X1 U38152 ( .A1(n38295), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[60][5] ), .B2(n38294), .ZN(n38292) );
  INV_X1 U38153 ( .A(n38292), .ZN(n2358) );
  OAI22_X1 U38154 ( .A1(n38295), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[60][6] ), .B2(n38294), .ZN(n38293) );
  INV_X1 U38155 ( .A(n38293), .ZN(n2357) );
  OAI22_X1 U38156 ( .A1(n38295), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[60][7] ), .B2(n38294), .ZN(n38296) );
  INV_X1 U38157 ( .A(n38296), .ZN(n2356) );
  NOR2_X1 U38158 ( .A1(n38307), .A2(n38957), .ZN(n38304) );
  INV_X1 U38159 ( .A(n38304), .ZN(n38305) );
  OAI22_X1 U38160 ( .A1(n38305), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[61][0] ), .B2(n38304), .ZN(n38297) );
  INV_X1 U38161 ( .A(n38297), .ZN(n2355) );
  OAI22_X1 U38162 ( .A1(n38305), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[61][1] ), .B2(n38304), .ZN(n38298) );
  INV_X1 U38163 ( .A(n38298), .ZN(n2354) );
  OAI22_X1 U38164 ( .A1(n38305), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[61][2] ), .B2(n38304), .ZN(n38299) );
  INV_X1 U38165 ( .A(n38299), .ZN(n2353) );
  OAI22_X1 U38166 ( .A1(n38305), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[61][3] ), .B2(n38304), .ZN(n38300) );
  INV_X1 U38167 ( .A(n38300), .ZN(n2352) );
  OAI22_X1 U38168 ( .A1(n38305), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[61][4] ), .B2(n38304), .ZN(n38301) );
  INV_X1 U38169 ( .A(n38301), .ZN(n2351) );
  OAI22_X1 U38170 ( .A1(n38305), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[61][5] ), .B2(n38304), .ZN(n38302) );
  INV_X1 U38171 ( .A(n38302), .ZN(n2350) );
  OAI22_X1 U38172 ( .A1(n38305), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[61][6] ), .B2(n38304), .ZN(n38303) );
  INV_X1 U38173 ( .A(n38303), .ZN(n2349) );
  OAI22_X1 U38174 ( .A1(n38305), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[61][7] ), .B2(n38304), .ZN(n38306) );
  INV_X1 U38175 ( .A(n38306), .ZN(n2348) );
  NOR2_X1 U38176 ( .A1(n38307), .A2(n38968), .ZN(n38315) );
  INV_X1 U38177 ( .A(n38315), .ZN(n38316) );
  OAI22_X1 U38178 ( .A1(n38316), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[62][0] ), .B2(n38315), .ZN(n38308) );
  INV_X1 U38179 ( .A(n38308), .ZN(n2347) );
  OAI22_X1 U38180 ( .A1(n38316), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[62][1] ), .B2(n38315), .ZN(n38309) );
  INV_X1 U38181 ( .A(n38309), .ZN(n2346) );
  OAI22_X1 U38182 ( .A1(n38316), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[62][2] ), .B2(n38315), .ZN(n38310) );
  INV_X1 U38183 ( .A(n38310), .ZN(n2345) );
  OAI22_X1 U38184 ( .A1(n38316), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[62][3] ), .B2(n38315), .ZN(n38311) );
  INV_X1 U38185 ( .A(n38311), .ZN(n2344) );
  OAI22_X1 U38186 ( .A1(n38316), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[62][4] ), .B2(n38315), .ZN(n38312) );
  INV_X1 U38187 ( .A(n38312), .ZN(n2343) );
  OAI22_X1 U38188 ( .A1(n38316), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[62][5] ), .B2(n38315), .ZN(n38313) );
  INV_X1 U38189 ( .A(n38313), .ZN(n2342) );
  OAI22_X1 U38190 ( .A1(n38316), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[62][6] ), .B2(n38315), .ZN(n38314) );
  INV_X1 U38191 ( .A(n38314), .ZN(n2341) );
  OAI22_X1 U38192 ( .A1(n38316), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[62][7] ), .B2(n38315), .ZN(n38317) );
  INV_X1 U38193 ( .A(n38317), .ZN(n2340) );
  OAI22_X1 U38194 ( .A1(n38326), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[63][0] ), .B2(n38325), .ZN(n38318) );
  INV_X1 U38195 ( .A(n38318), .ZN(n2339) );
  OAI22_X1 U38196 ( .A1(n38326), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[63][1] ), .B2(n38325), .ZN(n38319) );
  INV_X1 U38197 ( .A(n38319), .ZN(n2338) );
  OAI22_X1 U38198 ( .A1(n38326), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[63][2] ), .B2(n38325), .ZN(n38320) );
  INV_X1 U38199 ( .A(n38320), .ZN(n2337) );
  OAI22_X1 U38200 ( .A1(n38326), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[63][3] ), .B2(n38325), .ZN(n38321) );
  INV_X1 U38201 ( .A(n38321), .ZN(n2336) );
  OAI22_X1 U38202 ( .A1(n38326), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[63][4] ), .B2(n38325), .ZN(n38322) );
  INV_X1 U38203 ( .A(n38322), .ZN(n2335) );
  OAI22_X1 U38204 ( .A1(n38326), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[63][5] ), .B2(n38325), .ZN(n38323) );
  INV_X1 U38205 ( .A(n38323), .ZN(n2334) );
  OAI22_X1 U38206 ( .A1(n38326), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[63][6] ), .B2(n38325), .ZN(n38324) );
  INV_X1 U38207 ( .A(n38324), .ZN(n2333) );
  OAI22_X1 U38208 ( .A1(n38326), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[63][7] ), .B2(n38325), .ZN(n38327) );
  INV_X1 U38209 ( .A(n38327), .ZN(n2332) );
  NAND3_X1 U38210 ( .A1(xmem_addr[6]), .A2(n38651), .A3(n38998), .ZN(n38478)
         );
  NOR2_X1 U38211 ( .A1(n38814), .A2(n38478), .ZN(n38335) );
  INV_X1 U38212 ( .A(n38335), .ZN(n38336) );
  OAI22_X1 U38213 ( .A1(n38336), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[64][0] ), .B2(n38335), .ZN(n38328) );
  INV_X1 U38214 ( .A(n38328), .ZN(n2331) );
  OAI22_X1 U38215 ( .A1(n38336), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[64][1] ), .B2(n38335), .ZN(n38329) );
  INV_X1 U38216 ( .A(n38329), .ZN(n2330) );
  OAI22_X1 U38217 ( .A1(n38336), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[64][2] ), .B2(n38335), .ZN(n38330) );
  INV_X1 U38218 ( .A(n38330), .ZN(n2329) );
  OAI22_X1 U38219 ( .A1(n38336), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[64][3] ), .B2(n38335), .ZN(n38331) );
  INV_X1 U38220 ( .A(n38331), .ZN(n2328) );
  OAI22_X1 U38221 ( .A1(n38336), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[64][4] ), .B2(n38335), .ZN(n38332) );
  INV_X1 U38222 ( .A(n38332), .ZN(n2327) );
  OAI22_X1 U38223 ( .A1(n38336), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[64][5] ), .B2(n38335), .ZN(n38333) );
  INV_X1 U38224 ( .A(n38333), .ZN(n2326) );
  OAI22_X1 U38225 ( .A1(n38336), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[64][6] ), .B2(n38335), .ZN(n38334) );
  INV_X1 U38226 ( .A(n38334), .ZN(n2325) );
  OAI22_X1 U38227 ( .A1(n38336), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[64][7] ), .B2(n38335), .ZN(n38337) );
  INV_X1 U38228 ( .A(n38337), .ZN(n2324) );
  NOR2_X1 U38229 ( .A1(n38825), .A2(n38478), .ZN(n38345) );
  INV_X1 U38230 ( .A(n38345), .ZN(n38346) );
  OAI22_X1 U38231 ( .A1(n38346), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[65][0] ), .B2(n38345), .ZN(n38338) );
  INV_X1 U38232 ( .A(n38338), .ZN(n2323) );
  OAI22_X1 U38233 ( .A1(n38346), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[65][1] ), .B2(n38345), .ZN(n38339) );
  INV_X1 U38234 ( .A(n38339), .ZN(n2322) );
  OAI22_X1 U38235 ( .A1(n38346), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[65][2] ), .B2(n38345), .ZN(n38340) );
  INV_X1 U38236 ( .A(n38340), .ZN(n2321) );
  OAI22_X1 U38237 ( .A1(n38346), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[65][3] ), .B2(n38345), .ZN(n38341) );
  INV_X1 U38238 ( .A(n38341), .ZN(n2320) );
  OAI22_X1 U38239 ( .A1(n38346), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[65][4] ), .B2(n38345), .ZN(n38342) );
  INV_X1 U38240 ( .A(n38342), .ZN(n2319) );
  OAI22_X1 U38241 ( .A1(n38346), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[65][5] ), .B2(n38345), .ZN(n38343) );
  INV_X1 U38242 ( .A(n38343), .ZN(n2318) );
  OAI22_X1 U38243 ( .A1(n38346), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[65][6] ), .B2(n38345), .ZN(n38344) );
  INV_X1 U38244 ( .A(n38344), .ZN(n2317) );
  OAI22_X1 U38245 ( .A1(n38346), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[65][7] ), .B2(n38345), .ZN(n38347) );
  INV_X1 U38246 ( .A(n38347), .ZN(n2316) );
  NOR2_X1 U38247 ( .A1(n38836), .A2(n38478), .ZN(n38355) );
  INV_X1 U38248 ( .A(n38355), .ZN(n38356) );
  OAI22_X1 U38249 ( .A1(n38356), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[66][0] ), .B2(n38355), .ZN(n38348) );
  INV_X1 U38250 ( .A(n38348), .ZN(n2315) );
  OAI22_X1 U38251 ( .A1(n38356), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[66][1] ), .B2(n38355), .ZN(n38349) );
  INV_X1 U38252 ( .A(n38349), .ZN(n2314) );
  OAI22_X1 U38253 ( .A1(n38356), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[66][2] ), .B2(n38355), .ZN(n38350) );
  INV_X1 U38254 ( .A(n38350), .ZN(n2313) );
  OAI22_X1 U38255 ( .A1(n38356), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[66][3] ), .B2(n38355), .ZN(n38351) );
  INV_X1 U38256 ( .A(n38351), .ZN(n2312) );
  OAI22_X1 U38257 ( .A1(n38356), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[66][4] ), .B2(n38355), .ZN(n38352) );
  INV_X1 U38258 ( .A(n38352), .ZN(n2311) );
  OAI22_X1 U38259 ( .A1(n38356), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[66][5] ), .B2(n38355), .ZN(n38353) );
  INV_X1 U38260 ( .A(n38353), .ZN(n2310) );
  OAI22_X1 U38261 ( .A1(n38356), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[66][6] ), .B2(n38355), .ZN(n38354) );
  INV_X1 U38262 ( .A(n38354), .ZN(n2309) );
  OAI22_X1 U38263 ( .A1(n38356), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[66][7] ), .B2(n38355), .ZN(n38357) );
  INV_X1 U38264 ( .A(n38357), .ZN(n2308) );
  NOR2_X1 U38265 ( .A1(n38847), .A2(n38478), .ZN(n38365) );
  INV_X1 U38266 ( .A(n38365), .ZN(n38366) );
  OAI22_X1 U38267 ( .A1(n38366), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[67][0] ), .B2(n38365), .ZN(n38358) );
  INV_X1 U38268 ( .A(n38358), .ZN(n2307) );
  OAI22_X1 U38269 ( .A1(n38366), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[67][1] ), .B2(n38365), .ZN(n38359) );
  INV_X1 U38270 ( .A(n38359), .ZN(n2306) );
  OAI22_X1 U38271 ( .A1(n38366), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[67][2] ), .B2(n38365), .ZN(n38360) );
  INV_X1 U38272 ( .A(n38360), .ZN(n2305) );
  OAI22_X1 U38273 ( .A1(n38366), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[67][3] ), .B2(n38365), .ZN(n38361) );
  INV_X1 U38274 ( .A(n38361), .ZN(n2304) );
  OAI22_X1 U38275 ( .A1(n38366), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[67][4] ), .B2(n38365), .ZN(n38362) );
  INV_X1 U38276 ( .A(n38362), .ZN(n2303) );
  OAI22_X1 U38277 ( .A1(n38366), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[67][5] ), .B2(n38365), .ZN(n38363) );
  INV_X1 U38278 ( .A(n38363), .ZN(n2302) );
  OAI22_X1 U38279 ( .A1(n38366), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[67][6] ), .B2(n38365), .ZN(n38364) );
  INV_X1 U38280 ( .A(n38364), .ZN(n2301) );
  OAI22_X1 U38281 ( .A1(n38366), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[67][7] ), .B2(n38365), .ZN(n38367) );
  INV_X1 U38282 ( .A(n38367), .ZN(n2300) );
  NOR2_X1 U38283 ( .A1(n38858), .A2(n38478), .ZN(n38375) );
  INV_X1 U38284 ( .A(n38375), .ZN(n38376) );
  OAI22_X1 U38285 ( .A1(n38376), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[68][0] ), .B2(n38375), .ZN(n38368) );
  INV_X1 U38286 ( .A(n38368), .ZN(n2299) );
  OAI22_X1 U38287 ( .A1(n38376), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[68][1] ), .B2(n38375), .ZN(n38369) );
  INV_X1 U38288 ( .A(n38369), .ZN(n2298) );
  OAI22_X1 U38289 ( .A1(n38376), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[68][2] ), .B2(n38375), .ZN(n38370) );
  INV_X1 U38290 ( .A(n38370), .ZN(n2297) );
  OAI22_X1 U38291 ( .A1(n38376), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[68][3] ), .B2(n38375), .ZN(n38371) );
  INV_X1 U38292 ( .A(n38371), .ZN(n2296) );
  OAI22_X1 U38293 ( .A1(n38376), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[68][4] ), .B2(n38375), .ZN(n38372) );
  INV_X1 U38294 ( .A(n38372), .ZN(n2295) );
  OAI22_X1 U38295 ( .A1(n38376), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[68][5] ), .B2(n38375), .ZN(n38373) );
  INV_X1 U38296 ( .A(n38373), .ZN(n2294) );
  OAI22_X1 U38297 ( .A1(n38376), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[68][6] ), .B2(n38375), .ZN(n38374) );
  INV_X1 U38298 ( .A(n38374), .ZN(n2293) );
  OAI22_X1 U38299 ( .A1(n38376), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[68][7] ), .B2(n38375), .ZN(n38377) );
  INV_X1 U38300 ( .A(n38377), .ZN(n2292) );
  NOR2_X1 U38301 ( .A1(n38869), .A2(n38478), .ZN(n38385) );
  INV_X1 U38302 ( .A(n38385), .ZN(n38386) );
  OAI22_X1 U38303 ( .A1(n38386), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[69][0] ), .B2(n38385), .ZN(n38378) );
  INV_X1 U38304 ( .A(n38378), .ZN(n2291) );
  OAI22_X1 U38305 ( .A1(n38386), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[69][1] ), .B2(n38385), .ZN(n38379) );
  INV_X1 U38306 ( .A(n38379), .ZN(n2290) );
  OAI22_X1 U38307 ( .A1(n38386), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[69][2] ), .B2(n38385), .ZN(n38380) );
  INV_X1 U38308 ( .A(n38380), .ZN(n2289) );
  OAI22_X1 U38309 ( .A1(n38386), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[69][3] ), .B2(n38385), .ZN(n38381) );
  INV_X1 U38310 ( .A(n38381), .ZN(n2288) );
  OAI22_X1 U38311 ( .A1(n38386), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[69][4] ), .B2(n38385), .ZN(n38382) );
  INV_X1 U38312 ( .A(n38382), .ZN(n2287) );
  OAI22_X1 U38313 ( .A1(n38386), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[69][5] ), .B2(n38385), .ZN(n38383) );
  INV_X1 U38314 ( .A(n38383), .ZN(n2286) );
  OAI22_X1 U38315 ( .A1(n38386), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[69][6] ), .B2(n38385), .ZN(n38384) );
  INV_X1 U38316 ( .A(n38384), .ZN(n2285) );
  OAI22_X1 U38317 ( .A1(n38386), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[69][7] ), .B2(n38385), .ZN(n38387) );
  INV_X1 U38318 ( .A(n38387), .ZN(n2284) );
  NOR2_X1 U38319 ( .A1(n38880), .A2(n38478), .ZN(n38395) );
  INV_X1 U38320 ( .A(n38395), .ZN(n38396) );
  OAI22_X1 U38321 ( .A1(n38396), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[70][0] ), .B2(n38395), .ZN(n38388) );
  INV_X1 U38322 ( .A(n38388), .ZN(n2283) );
  OAI22_X1 U38323 ( .A1(n38396), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[70][1] ), .B2(n38395), .ZN(n38389) );
  INV_X1 U38324 ( .A(n38389), .ZN(n2282) );
  OAI22_X1 U38325 ( .A1(n38396), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[70][2] ), .B2(n38395), .ZN(n38390) );
  INV_X1 U38326 ( .A(n38390), .ZN(n2281) );
  OAI22_X1 U38327 ( .A1(n38396), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[70][3] ), .B2(n38395), .ZN(n38391) );
  INV_X1 U38328 ( .A(n38391), .ZN(n2280) );
  OAI22_X1 U38329 ( .A1(n38396), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[70][4] ), .B2(n38395), .ZN(n38392) );
  INV_X1 U38330 ( .A(n38392), .ZN(n2279) );
  OAI22_X1 U38331 ( .A1(n38396), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[70][5] ), .B2(n38395), .ZN(n38393) );
  INV_X1 U38332 ( .A(n38393), .ZN(n2278) );
  OAI22_X1 U38333 ( .A1(n38396), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[70][6] ), .B2(n38395), .ZN(n38394) );
  INV_X1 U38334 ( .A(n38394), .ZN(n2277) );
  OAI22_X1 U38335 ( .A1(n38396), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[70][7] ), .B2(n38395), .ZN(n38397) );
  INV_X1 U38336 ( .A(n38397), .ZN(n2276) );
  NOR2_X1 U38337 ( .A1(n38891), .A2(n38478), .ZN(n38405) );
  INV_X1 U38338 ( .A(n38405), .ZN(n38406) );
  OAI22_X1 U38339 ( .A1(n38406), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[71][0] ), .B2(n38405), .ZN(n38398) );
  INV_X1 U38340 ( .A(n38398), .ZN(n2275) );
  OAI22_X1 U38341 ( .A1(n38406), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[71][1] ), .B2(n38405), .ZN(n38399) );
  INV_X1 U38342 ( .A(n38399), .ZN(n2274) );
  OAI22_X1 U38343 ( .A1(n38406), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[71][2] ), .B2(n38405), .ZN(n38400) );
  INV_X1 U38344 ( .A(n38400), .ZN(n2273) );
  OAI22_X1 U38345 ( .A1(n38406), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[71][3] ), .B2(n38405), .ZN(n38401) );
  INV_X1 U38346 ( .A(n38401), .ZN(n2272) );
  OAI22_X1 U38347 ( .A1(n38406), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[71][4] ), .B2(n38405), .ZN(n38402) );
  INV_X1 U38348 ( .A(n38402), .ZN(n2271) );
  OAI22_X1 U38349 ( .A1(n38406), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[71][5] ), .B2(n38405), .ZN(n38403) );
  INV_X1 U38350 ( .A(n38403), .ZN(n2270) );
  OAI22_X1 U38351 ( .A1(n38406), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[71][6] ), .B2(n38405), .ZN(n38404) );
  INV_X1 U38352 ( .A(n38404), .ZN(n2269) );
  OAI22_X1 U38353 ( .A1(n38406), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[71][7] ), .B2(n38405), .ZN(n38407) );
  INV_X1 U38354 ( .A(n38407), .ZN(n2268) );
  NOR2_X1 U38355 ( .A1(n38902), .A2(n38478), .ZN(n38415) );
  INV_X1 U38356 ( .A(n38415), .ZN(n38416) );
  OAI22_X1 U38357 ( .A1(n38416), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[72][0] ), .B2(n38415), .ZN(n38408) );
  INV_X1 U38358 ( .A(n38408), .ZN(n2267) );
  OAI22_X1 U38359 ( .A1(n38416), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[72][1] ), .B2(n38415), .ZN(n38409) );
  INV_X1 U38360 ( .A(n38409), .ZN(n2266) );
  OAI22_X1 U38361 ( .A1(n38416), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[72][2] ), .B2(n38415), .ZN(n38410) );
  INV_X1 U38362 ( .A(n38410), .ZN(n2265) );
  OAI22_X1 U38363 ( .A1(n38416), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[72][3] ), .B2(n38415), .ZN(n38411) );
  INV_X1 U38364 ( .A(n38411), .ZN(n2264) );
  OAI22_X1 U38365 ( .A1(n38416), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[72][4] ), .B2(n38415), .ZN(n38412) );
  INV_X1 U38366 ( .A(n38412), .ZN(n2263) );
  OAI22_X1 U38367 ( .A1(n38416), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[72][5] ), .B2(n38415), .ZN(n38413) );
  INV_X1 U38368 ( .A(n38413), .ZN(n2262) );
  OAI22_X1 U38369 ( .A1(n38416), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[72][6] ), .B2(n38415), .ZN(n38414) );
  INV_X1 U38370 ( .A(n38414), .ZN(n2261) );
  OAI22_X1 U38371 ( .A1(n38416), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[72][7] ), .B2(n38415), .ZN(n38417) );
  INV_X1 U38372 ( .A(n38417), .ZN(n2260) );
  NOR2_X1 U38373 ( .A1(n38913), .A2(n38478), .ZN(n38425) );
  INV_X1 U38374 ( .A(n38425), .ZN(n38426) );
  OAI22_X1 U38375 ( .A1(n38426), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[73][0] ), .B2(n38425), .ZN(n38418) );
  INV_X1 U38376 ( .A(n38418), .ZN(n2259) );
  OAI22_X1 U38377 ( .A1(n38426), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[73][1] ), .B2(n38425), .ZN(n38419) );
  INV_X1 U38378 ( .A(n38419), .ZN(n2258) );
  OAI22_X1 U38379 ( .A1(n38426), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[73][2] ), .B2(n38425), .ZN(n38420) );
  INV_X1 U38380 ( .A(n38420), .ZN(n2257) );
  OAI22_X1 U38381 ( .A1(n38426), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[73][3] ), .B2(n38425), .ZN(n38421) );
  INV_X1 U38382 ( .A(n38421), .ZN(n2256) );
  OAI22_X1 U38383 ( .A1(n38426), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[73][4] ), .B2(n38425), .ZN(n38422) );
  INV_X1 U38384 ( .A(n38422), .ZN(n2255) );
  OAI22_X1 U38385 ( .A1(n38426), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[73][5] ), .B2(n38425), .ZN(n38423) );
  INV_X1 U38386 ( .A(n38423), .ZN(n2254) );
  OAI22_X1 U38387 ( .A1(n38426), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[73][6] ), .B2(n38425), .ZN(n38424) );
  INV_X1 U38388 ( .A(n38424), .ZN(n2253) );
  OAI22_X1 U38389 ( .A1(n38426), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[73][7] ), .B2(n38425), .ZN(n38427) );
  INV_X1 U38390 ( .A(n38427), .ZN(n2252) );
  NOR2_X1 U38391 ( .A1(n38924), .A2(n38478), .ZN(n38435) );
  INV_X1 U38392 ( .A(n38435), .ZN(n38436) );
  OAI22_X1 U38393 ( .A1(n38436), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[74][0] ), .B2(n38435), .ZN(n38428) );
  INV_X1 U38394 ( .A(n38428), .ZN(n2251) );
  OAI22_X1 U38395 ( .A1(n38436), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[74][1] ), .B2(n38435), .ZN(n38429) );
  INV_X1 U38396 ( .A(n38429), .ZN(n2250) );
  OAI22_X1 U38397 ( .A1(n38436), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[74][2] ), .B2(n38435), .ZN(n38430) );
  INV_X1 U38398 ( .A(n38430), .ZN(n2249) );
  OAI22_X1 U38399 ( .A1(n38436), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[74][3] ), .B2(n38435), .ZN(n38431) );
  INV_X1 U38400 ( .A(n38431), .ZN(n2248) );
  OAI22_X1 U38401 ( .A1(n38436), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[74][4] ), .B2(n38435), .ZN(n38432) );
  INV_X1 U38402 ( .A(n38432), .ZN(n2247) );
  OAI22_X1 U38403 ( .A1(n38436), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[74][5] ), .B2(n38435), .ZN(n38433) );
  INV_X1 U38404 ( .A(n38433), .ZN(n2246) );
  OAI22_X1 U38405 ( .A1(n38436), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[74][6] ), .B2(n38435), .ZN(n38434) );
  INV_X1 U38406 ( .A(n38434), .ZN(n2245) );
  OAI22_X1 U38407 ( .A1(n38436), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[74][7] ), .B2(n38435), .ZN(n38437) );
  INV_X1 U38408 ( .A(n38437), .ZN(n2244) );
  NOR2_X1 U38409 ( .A1(n38935), .A2(n38478), .ZN(n38445) );
  INV_X1 U38410 ( .A(n38445), .ZN(n38446) );
  OAI22_X1 U38411 ( .A1(n38446), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[75][0] ), .B2(n38445), .ZN(n38438) );
  INV_X1 U38412 ( .A(n38438), .ZN(n2243) );
  OAI22_X1 U38413 ( .A1(n38446), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[75][1] ), .B2(n38445), .ZN(n38439) );
  INV_X1 U38414 ( .A(n38439), .ZN(n2242) );
  OAI22_X1 U38415 ( .A1(n38446), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[75][2] ), .B2(n38445), .ZN(n38440) );
  INV_X1 U38416 ( .A(n38440), .ZN(n2241) );
  OAI22_X1 U38417 ( .A1(n38446), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[75][3] ), .B2(n38445), .ZN(n38441) );
  INV_X1 U38418 ( .A(n38441), .ZN(n2240) );
  OAI22_X1 U38419 ( .A1(n38446), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[75][4] ), .B2(n38445), .ZN(n38442) );
  INV_X1 U38420 ( .A(n38442), .ZN(n2239) );
  OAI22_X1 U38421 ( .A1(n38446), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[75][5] ), .B2(n38445), .ZN(n38443) );
  INV_X1 U38422 ( .A(n38443), .ZN(n2238) );
  OAI22_X1 U38423 ( .A1(n38446), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[75][6] ), .B2(n38445), .ZN(n38444) );
  INV_X1 U38424 ( .A(n38444), .ZN(n2237) );
  OAI22_X1 U38425 ( .A1(n38446), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[75][7] ), .B2(n38445), .ZN(n38447) );
  INV_X1 U38426 ( .A(n38447), .ZN(n2236) );
  NOR2_X1 U38427 ( .A1(n38946), .A2(n38478), .ZN(n38455) );
  INV_X1 U38428 ( .A(n38455), .ZN(n38456) );
  OAI22_X1 U38429 ( .A1(n38456), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[76][0] ), .B2(n38455), .ZN(n38448) );
  INV_X1 U38430 ( .A(n38448), .ZN(n2235) );
  OAI22_X1 U38431 ( .A1(n38456), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[76][1] ), .B2(n38455), .ZN(n38449) );
  INV_X1 U38432 ( .A(n38449), .ZN(n2234) );
  OAI22_X1 U38433 ( .A1(n38456), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[76][2] ), .B2(n38455), .ZN(n38450) );
  INV_X1 U38434 ( .A(n38450), .ZN(n2233) );
  OAI22_X1 U38435 ( .A1(n38456), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[76][3] ), .B2(n38455), .ZN(n38451) );
  INV_X1 U38436 ( .A(n38451), .ZN(n2232) );
  OAI22_X1 U38437 ( .A1(n38456), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[76][4] ), .B2(n38455), .ZN(n38452) );
  INV_X1 U38438 ( .A(n38452), .ZN(n2231) );
  OAI22_X1 U38439 ( .A1(n38456), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[76][5] ), .B2(n38455), .ZN(n38453) );
  INV_X1 U38440 ( .A(n38453), .ZN(n2230) );
  OAI22_X1 U38441 ( .A1(n38456), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[76][6] ), .B2(n38455), .ZN(n38454) );
  INV_X1 U38442 ( .A(n38454), .ZN(n2229) );
  OAI22_X1 U38443 ( .A1(n38456), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[76][7] ), .B2(n38455), .ZN(n38457) );
  INV_X1 U38444 ( .A(n38457), .ZN(n2228) );
  NOR2_X1 U38445 ( .A1(n38957), .A2(n38478), .ZN(n38465) );
  INV_X1 U38446 ( .A(n38465), .ZN(n38466) );
  OAI22_X1 U38447 ( .A1(n38466), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[77][0] ), .B2(n38465), .ZN(n38458) );
  INV_X1 U38448 ( .A(n38458), .ZN(n2227) );
  OAI22_X1 U38449 ( .A1(n38466), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[77][1] ), .B2(n38465), .ZN(n38459) );
  INV_X1 U38450 ( .A(n38459), .ZN(n2226) );
  OAI22_X1 U38451 ( .A1(n38466), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[77][2] ), .B2(n38465), .ZN(n38460) );
  INV_X1 U38452 ( .A(n38460), .ZN(n2225) );
  OAI22_X1 U38453 ( .A1(n38466), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[77][3] ), .B2(n38465), .ZN(n38461) );
  INV_X1 U38454 ( .A(n38461), .ZN(n2224) );
  OAI22_X1 U38455 ( .A1(n38466), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[77][4] ), .B2(n38465), .ZN(n38462) );
  INV_X1 U38456 ( .A(n38462), .ZN(n2223) );
  OAI22_X1 U38457 ( .A1(n38466), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[77][5] ), .B2(n38465), .ZN(n38463) );
  INV_X1 U38458 ( .A(n38463), .ZN(n2222) );
  OAI22_X1 U38459 ( .A1(n38466), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[77][6] ), .B2(n38465), .ZN(n38464) );
  INV_X1 U38460 ( .A(n38464), .ZN(n2221) );
  OAI22_X1 U38461 ( .A1(n38466), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[77][7] ), .B2(n38465), .ZN(n38467) );
  INV_X1 U38462 ( .A(n38467), .ZN(n2220) );
  NOR2_X1 U38463 ( .A1(n38968), .A2(n38478), .ZN(n38475) );
  INV_X1 U38464 ( .A(n38475), .ZN(n38476) );
  OAI22_X1 U38465 ( .A1(n38476), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[78][0] ), .B2(n38475), .ZN(n38468) );
  INV_X1 U38466 ( .A(n38468), .ZN(n2219) );
  OAI22_X1 U38467 ( .A1(n38476), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[78][1] ), .B2(n38475), .ZN(n38469) );
  INV_X1 U38468 ( .A(n38469), .ZN(n2218) );
  OAI22_X1 U38469 ( .A1(n38476), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[78][2] ), .B2(n38475), .ZN(n38470) );
  INV_X1 U38470 ( .A(n38470), .ZN(n2217) );
  OAI22_X1 U38471 ( .A1(n38476), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[78][3] ), .B2(n38475), .ZN(n38471) );
  INV_X1 U38472 ( .A(n38471), .ZN(n2216) );
  OAI22_X1 U38473 ( .A1(n38476), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[78][4] ), .B2(n38475), .ZN(n38472) );
  INV_X1 U38474 ( .A(n38472), .ZN(n2215) );
  OAI22_X1 U38475 ( .A1(n38476), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[78][5] ), .B2(n38475), .ZN(n38473) );
  INV_X1 U38476 ( .A(n38473), .ZN(n2214) );
  OAI22_X1 U38477 ( .A1(n38476), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[78][6] ), .B2(n38475), .ZN(n38474) );
  INV_X1 U38478 ( .A(n38474), .ZN(n2213) );
  OAI22_X1 U38479 ( .A1(n38476), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[78][7] ), .B2(n38475), .ZN(n38477) );
  INV_X1 U38480 ( .A(n38477), .ZN(n2212) );
  NOR2_X1 U38481 ( .A1(n38803), .A2(n38478), .ZN(n38486) );
  INV_X1 U38482 ( .A(n38486), .ZN(n38487) );
  OAI22_X1 U38483 ( .A1(n38487), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[79][0] ), .B2(n38486), .ZN(n38479) );
  INV_X1 U38484 ( .A(n38479), .ZN(n2211) );
  OAI22_X1 U38485 ( .A1(n38487), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[79][1] ), .B2(n38486), .ZN(n38480) );
  INV_X1 U38486 ( .A(n38480), .ZN(n2210) );
  OAI22_X1 U38487 ( .A1(n38487), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[79][2] ), .B2(n38486), .ZN(n38481) );
  INV_X1 U38488 ( .A(n38481), .ZN(n2209) );
  OAI22_X1 U38489 ( .A1(n38487), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[79][3] ), .B2(n38486), .ZN(n38482) );
  INV_X1 U38490 ( .A(n38482), .ZN(n2208) );
  OAI22_X1 U38491 ( .A1(n38487), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[79][4] ), .B2(n38486), .ZN(n38483) );
  INV_X1 U38492 ( .A(n38483), .ZN(n2207) );
  OAI22_X1 U38493 ( .A1(n38487), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[79][5] ), .B2(n38486), .ZN(n38484) );
  INV_X1 U38494 ( .A(n38484), .ZN(n2206) );
  OAI22_X1 U38495 ( .A1(n38487), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[79][6] ), .B2(n38486), .ZN(n38485) );
  INV_X1 U38496 ( .A(n38485), .ZN(n2205) );
  OAI22_X1 U38497 ( .A1(n38487), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[79][7] ), .B2(n38486), .ZN(n38488) );
  INV_X1 U38498 ( .A(n38488), .ZN(n2204) );
  NAND3_X1 U38499 ( .A1(xmem_addr[6]), .A2(n38489), .A3(n38998), .ZN(n38640)
         );
  NOR2_X1 U38500 ( .A1(n38814), .A2(n38640), .ZN(n38497) );
  INV_X1 U38501 ( .A(n38497), .ZN(n38498) );
  OAI22_X1 U38502 ( .A1(n38498), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[80][0] ), .B2(n38497), .ZN(n38490) );
  INV_X1 U38503 ( .A(n38490), .ZN(n2203) );
  OAI22_X1 U38504 ( .A1(n38498), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[80][1] ), .B2(n38497), .ZN(n38491) );
  INV_X1 U38505 ( .A(n38491), .ZN(n2202) );
  OAI22_X1 U38506 ( .A1(n38498), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[80][2] ), .B2(n38497), .ZN(n38492) );
  INV_X1 U38507 ( .A(n38492), .ZN(n2201) );
  OAI22_X1 U38508 ( .A1(n38498), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[80][3] ), .B2(n38497), .ZN(n38493) );
  INV_X1 U38509 ( .A(n38493), .ZN(n2200) );
  OAI22_X1 U38510 ( .A1(n38498), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[80][4] ), .B2(n38497), .ZN(n38494) );
  INV_X1 U38511 ( .A(n38494), .ZN(n2199) );
  OAI22_X1 U38512 ( .A1(n38498), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[80][5] ), .B2(n38497), .ZN(n38495) );
  INV_X1 U38513 ( .A(n38495), .ZN(n2198) );
  OAI22_X1 U38514 ( .A1(n38498), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[80][6] ), .B2(n38497), .ZN(n38496) );
  INV_X1 U38515 ( .A(n38496), .ZN(n2197) );
  OAI22_X1 U38516 ( .A1(n38498), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[80][7] ), .B2(n38497), .ZN(n38499) );
  INV_X1 U38517 ( .A(n38499), .ZN(n2196) );
  NOR2_X1 U38518 ( .A1(n38825), .A2(n38640), .ZN(n38507) );
  INV_X1 U38519 ( .A(n38507), .ZN(n38508) );
  OAI22_X1 U38520 ( .A1(n38508), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[81][0] ), .B2(n38507), .ZN(n38500) );
  INV_X1 U38521 ( .A(n38500), .ZN(n2195) );
  OAI22_X1 U38522 ( .A1(n38508), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[81][1] ), .B2(n38507), .ZN(n38501) );
  INV_X1 U38523 ( .A(n38501), .ZN(n2194) );
  OAI22_X1 U38524 ( .A1(n38508), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[81][2] ), .B2(n38507), .ZN(n38502) );
  INV_X1 U38525 ( .A(n38502), .ZN(n2193) );
  OAI22_X1 U38526 ( .A1(n38508), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[81][3] ), .B2(n38507), .ZN(n38503) );
  INV_X1 U38527 ( .A(n38503), .ZN(n2192) );
  OAI22_X1 U38528 ( .A1(n38508), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[81][4] ), .B2(n38507), .ZN(n38504) );
  INV_X1 U38529 ( .A(n38504), .ZN(n2191) );
  OAI22_X1 U38530 ( .A1(n38508), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[81][5] ), .B2(n38507), .ZN(n38505) );
  INV_X1 U38531 ( .A(n38505), .ZN(n2190) );
  OAI22_X1 U38532 ( .A1(n38508), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[81][6] ), .B2(n38507), .ZN(n38506) );
  INV_X1 U38533 ( .A(n38506), .ZN(n2189) );
  OAI22_X1 U38534 ( .A1(n38508), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[81][7] ), .B2(n38507), .ZN(n38509) );
  INV_X1 U38535 ( .A(n38509), .ZN(n2188) );
  NOR2_X1 U38536 ( .A1(n38836), .A2(n38640), .ZN(n38517) );
  INV_X1 U38537 ( .A(n38517), .ZN(n38518) );
  OAI22_X1 U38538 ( .A1(n38518), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[82][0] ), .B2(n38517), .ZN(n38510) );
  INV_X1 U38539 ( .A(n38510), .ZN(n2187) );
  OAI22_X1 U38540 ( .A1(n38518), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[82][1] ), .B2(n38517), .ZN(n38511) );
  INV_X1 U38541 ( .A(n38511), .ZN(n2186) );
  OAI22_X1 U38542 ( .A1(n38518), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[82][2] ), .B2(n38517), .ZN(n38512) );
  INV_X1 U38543 ( .A(n38512), .ZN(n2185) );
  OAI22_X1 U38544 ( .A1(n38518), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[82][3] ), .B2(n38517), .ZN(n38513) );
  INV_X1 U38545 ( .A(n38513), .ZN(n2184) );
  OAI22_X1 U38546 ( .A1(n38518), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[82][4] ), .B2(n38517), .ZN(n38514) );
  INV_X1 U38547 ( .A(n38514), .ZN(n2183) );
  OAI22_X1 U38548 ( .A1(n38518), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[82][5] ), .B2(n38517), .ZN(n38515) );
  INV_X1 U38549 ( .A(n38515), .ZN(n2182) );
  OAI22_X1 U38550 ( .A1(n38518), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[82][6] ), .B2(n38517), .ZN(n38516) );
  INV_X1 U38551 ( .A(n38516), .ZN(n2181) );
  OAI22_X1 U38552 ( .A1(n38518), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[82][7] ), .B2(n38517), .ZN(n38519) );
  INV_X1 U38553 ( .A(n38519), .ZN(n2180) );
  NOR2_X1 U38554 ( .A1(n38847), .A2(n38640), .ZN(n38527) );
  INV_X1 U38555 ( .A(n38527), .ZN(n38528) );
  OAI22_X1 U38556 ( .A1(n38528), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[83][0] ), .B2(n38527), .ZN(n38520) );
  INV_X1 U38557 ( .A(n38520), .ZN(n2179) );
  OAI22_X1 U38558 ( .A1(n38528), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[83][1] ), .B2(n38527), .ZN(n38521) );
  INV_X1 U38559 ( .A(n38521), .ZN(n2178) );
  OAI22_X1 U38560 ( .A1(n38528), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[83][2] ), .B2(n38527), .ZN(n38522) );
  INV_X1 U38561 ( .A(n38522), .ZN(n2177) );
  OAI22_X1 U38562 ( .A1(n38528), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[83][3] ), .B2(n38527), .ZN(n38523) );
  INV_X1 U38563 ( .A(n38523), .ZN(n2176) );
  OAI22_X1 U38564 ( .A1(n38528), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[83][4] ), .B2(n38527), .ZN(n38524) );
  INV_X1 U38565 ( .A(n38524), .ZN(n2175) );
  OAI22_X1 U38566 ( .A1(n38528), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[83][5] ), .B2(n38527), .ZN(n38525) );
  INV_X1 U38567 ( .A(n38525), .ZN(n2174) );
  OAI22_X1 U38568 ( .A1(n38528), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[83][6] ), .B2(n38527), .ZN(n38526) );
  INV_X1 U38569 ( .A(n38526), .ZN(n2173) );
  OAI22_X1 U38570 ( .A1(n38528), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[83][7] ), .B2(n38527), .ZN(n38529) );
  INV_X1 U38571 ( .A(n38529), .ZN(n2172) );
  NOR2_X1 U38572 ( .A1(n38858), .A2(n38640), .ZN(n38537) );
  INV_X1 U38573 ( .A(n38537), .ZN(n38538) );
  OAI22_X1 U38574 ( .A1(n38538), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[84][0] ), .B2(n38537), .ZN(n38530) );
  INV_X1 U38575 ( .A(n38530), .ZN(n2171) );
  OAI22_X1 U38576 ( .A1(n38538), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[84][1] ), .B2(n38537), .ZN(n38531) );
  INV_X1 U38577 ( .A(n38531), .ZN(n2170) );
  OAI22_X1 U38578 ( .A1(n38538), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[84][2] ), .B2(n38537), .ZN(n38532) );
  INV_X1 U38579 ( .A(n38532), .ZN(n2169) );
  OAI22_X1 U38580 ( .A1(n38538), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[84][3] ), .B2(n38537), .ZN(n38533) );
  INV_X1 U38581 ( .A(n38533), .ZN(n2168) );
  OAI22_X1 U38582 ( .A1(n38538), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[84][4] ), .B2(n38537), .ZN(n38534) );
  INV_X1 U38583 ( .A(n38534), .ZN(n2167) );
  OAI22_X1 U38584 ( .A1(n38538), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[84][5] ), .B2(n38537), .ZN(n38535) );
  INV_X1 U38585 ( .A(n38535), .ZN(n2166) );
  OAI22_X1 U38586 ( .A1(n38538), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[84][6] ), .B2(n38537), .ZN(n38536) );
  INV_X1 U38587 ( .A(n38536), .ZN(n2165) );
  OAI22_X1 U38588 ( .A1(n38538), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[84][7] ), .B2(n38537), .ZN(n38539) );
  INV_X1 U38589 ( .A(n38539), .ZN(n2164) );
  NOR2_X1 U38590 ( .A1(n38869), .A2(n38640), .ZN(n38547) );
  INV_X1 U38591 ( .A(n38547), .ZN(n38548) );
  OAI22_X1 U38592 ( .A1(n38548), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[85][0] ), .B2(n38547), .ZN(n38540) );
  INV_X1 U38593 ( .A(n38540), .ZN(n2163) );
  OAI22_X1 U38594 ( .A1(n38548), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[85][1] ), .B2(n38547), .ZN(n38541) );
  INV_X1 U38595 ( .A(n38541), .ZN(n2162) );
  OAI22_X1 U38596 ( .A1(n38548), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[85][2] ), .B2(n38547), .ZN(n38542) );
  INV_X1 U38597 ( .A(n38542), .ZN(n2161) );
  OAI22_X1 U38598 ( .A1(n38548), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[85][3] ), .B2(n38547), .ZN(n38543) );
  INV_X1 U38599 ( .A(n38543), .ZN(n2160) );
  OAI22_X1 U38600 ( .A1(n38548), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[85][4] ), .B2(n38547), .ZN(n38544) );
  INV_X1 U38601 ( .A(n38544), .ZN(n2159) );
  OAI22_X1 U38602 ( .A1(n38548), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[85][5] ), .B2(n38547), .ZN(n38545) );
  INV_X1 U38603 ( .A(n38545), .ZN(n2158) );
  OAI22_X1 U38604 ( .A1(n38548), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[85][6] ), .B2(n38547), .ZN(n38546) );
  INV_X1 U38605 ( .A(n38546), .ZN(n2157) );
  OAI22_X1 U38606 ( .A1(n38548), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[85][7] ), .B2(n38547), .ZN(n38549) );
  INV_X1 U38607 ( .A(n38549), .ZN(n2156) );
  NOR2_X1 U38608 ( .A1(n38880), .A2(n38640), .ZN(n38557) );
  INV_X1 U38609 ( .A(n38557), .ZN(n38558) );
  OAI22_X1 U38610 ( .A1(n38558), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[86][0] ), .B2(n38557), .ZN(n38550) );
  INV_X1 U38611 ( .A(n38550), .ZN(n2155) );
  OAI22_X1 U38612 ( .A1(n38558), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[86][1] ), .B2(n38557), .ZN(n38551) );
  INV_X1 U38613 ( .A(n38551), .ZN(n2154) );
  OAI22_X1 U38614 ( .A1(n38558), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[86][2] ), .B2(n38557), .ZN(n38552) );
  INV_X1 U38615 ( .A(n38552), .ZN(n2153) );
  OAI22_X1 U38616 ( .A1(n38558), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[86][3] ), .B2(n38557), .ZN(n38553) );
  INV_X1 U38617 ( .A(n38553), .ZN(n2152) );
  OAI22_X1 U38618 ( .A1(n38558), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[86][4] ), .B2(n38557), .ZN(n38554) );
  INV_X1 U38619 ( .A(n38554), .ZN(n2151) );
  OAI22_X1 U38620 ( .A1(n38558), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[86][5] ), .B2(n38557), .ZN(n38555) );
  INV_X1 U38621 ( .A(n38555), .ZN(n2150) );
  OAI22_X1 U38622 ( .A1(n38558), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[86][6] ), .B2(n38557), .ZN(n38556) );
  INV_X1 U38623 ( .A(n38556), .ZN(n2149) );
  OAI22_X1 U38624 ( .A1(n38558), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[86][7] ), .B2(n38557), .ZN(n38559) );
  INV_X1 U38625 ( .A(n38559), .ZN(n2148) );
  NOR2_X1 U38626 ( .A1(n38891), .A2(n38640), .ZN(n38567) );
  INV_X1 U38627 ( .A(n38567), .ZN(n38568) );
  OAI22_X1 U38628 ( .A1(n38568), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[87][0] ), .B2(n38567), .ZN(n38560) );
  INV_X1 U38629 ( .A(n38560), .ZN(n2147) );
  OAI22_X1 U38630 ( .A1(n38568), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[87][1] ), .B2(n38567), .ZN(n38561) );
  INV_X1 U38631 ( .A(n38561), .ZN(n2146) );
  OAI22_X1 U38632 ( .A1(n38568), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[87][2] ), .B2(n38567), .ZN(n38562) );
  INV_X1 U38633 ( .A(n38562), .ZN(n2145) );
  OAI22_X1 U38634 ( .A1(n38568), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[87][3] ), .B2(n38567), .ZN(n38563) );
  INV_X1 U38635 ( .A(n38563), .ZN(n2144) );
  OAI22_X1 U38636 ( .A1(n38568), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[87][4] ), .B2(n38567), .ZN(n38564) );
  INV_X1 U38637 ( .A(n38564), .ZN(n2143) );
  OAI22_X1 U38638 ( .A1(n38568), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[87][5] ), .B2(n38567), .ZN(n38565) );
  INV_X1 U38639 ( .A(n38565), .ZN(n2142) );
  OAI22_X1 U38640 ( .A1(n38568), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[87][6] ), .B2(n38567), .ZN(n38566) );
  INV_X1 U38641 ( .A(n38566), .ZN(n2141) );
  OAI22_X1 U38642 ( .A1(n38568), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[87][7] ), .B2(n38567), .ZN(n38569) );
  INV_X1 U38643 ( .A(n38569), .ZN(n2140) );
  NOR2_X1 U38644 ( .A1(n38902), .A2(n38640), .ZN(n38577) );
  INV_X1 U38645 ( .A(n38577), .ZN(n38578) );
  OAI22_X1 U38646 ( .A1(n38578), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[88][0] ), .B2(n38577), .ZN(n38570) );
  INV_X1 U38647 ( .A(n38570), .ZN(n2139) );
  OAI22_X1 U38648 ( .A1(n38578), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[88][1] ), .B2(n38577), .ZN(n38571) );
  INV_X1 U38649 ( .A(n38571), .ZN(n2138) );
  OAI22_X1 U38650 ( .A1(n38578), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[88][2] ), .B2(n38577), .ZN(n38572) );
  INV_X1 U38651 ( .A(n38572), .ZN(n2137) );
  OAI22_X1 U38652 ( .A1(n38578), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[88][3] ), .B2(n38577), .ZN(n38573) );
  INV_X1 U38653 ( .A(n38573), .ZN(n2136) );
  OAI22_X1 U38654 ( .A1(n38578), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[88][4] ), .B2(n38577), .ZN(n38574) );
  INV_X1 U38655 ( .A(n38574), .ZN(n2135) );
  OAI22_X1 U38656 ( .A1(n38578), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[88][5] ), .B2(n38577), .ZN(n38575) );
  INV_X1 U38657 ( .A(n38575), .ZN(n2134) );
  OAI22_X1 U38658 ( .A1(n38578), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[88][6] ), .B2(n38577), .ZN(n38576) );
  INV_X1 U38659 ( .A(n38576), .ZN(n2133) );
  OAI22_X1 U38660 ( .A1(n38578), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[88][7] ), .B2(n38577), .ZN(n38579) );
  INV_X1 U38661 ( .A(n38579), .ZN(n2132) );
  NOR2_X1 U38662 ( .A1(n38913), .A2(n38640), .ZN(n38587) );
  INV_X1 U38663 ( .A(n38587), .ZN(n38588) );
  OAI22_X1 U38664 ( .A1(n38588), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[89][0] ), .B2(n38587), .ZN(n38580) );
  INV_X1 U38665 ( .A(n38580), .ZN(n2131) );
  OAI22_X1 U38666 ( .A1(n38588), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[89][1] ), .B2(n38587), .ZN(n38581) );
  INV_X1 U38667 ( .A(n38581), .ZN(n2130) );
  OAI22_X1 U38668 ( .A1(n38588), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[89][2] ), .B2(n38587), .ZN(n38582) );
  INV_X1 U38669 ( .A(n38582), .ZN(n2129) );
  OAI22_X1 U38670 ( .A1(n38588), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[89][3] ), .B2(n38587), .ZN(n38583) );
  INV_X1 U38671 ( .A(n38583), .ZN(n2128) );
  OAI22_X1 U38672 ( .A1(n38588), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[89][4] ), .B2(n38587), .ZN(n38584) );
  INV_X1 U38673 ( .A(n38584), .ZN(n2127) );
  OAI22_X1 U38674 ( .A1(n38588), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[89][5] ), .B2(n38587), .ZN(n38585) );
  INV_X1 U38675 ( .A(n38585), .ZN(n2126) );
  OAI22_X1 U38676 ( .A1(n38588), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[89][6] ), .B2(n38587), .ZN(n38586) );
  INV_X1 U38677 ( .A(n38586), .ZN(n2125) );
  OAI22_X1 U38678 ( .A1(n38588), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[89][7] ), .B2(n38587), .ZN(n38589) );
  INV_X1 U38679 ( .A(n38589), .ZN(n2124) );
  NOR2_X1 U38680 ( .A1(n38924), .A2(n38640), .ZN(n38597) );
  INV_X1 U38681 ( .A(n38597), .ZN(n38598) );
  OAI22_X1 U38682 ( .A1(n38598), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[90][0] ), .B2(n38597), .ZN(n38590) );
  INV_X1 U38683 ( .A(n38590), .ZN(n2123) );
  OAI22_X1 U38684 ( .A1(n38598), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[90][1] ), .B2(n38597), .ZN(n38591) );
  INV_X1 U38685 ( .A(n38591), .ZN(n2122) );
  OAI22_X1 U38686 ( .A1(n38598), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[90][2] ), .B2(n38597), .ZN(n38592) );
  INV_X1 U38687 ( .A(n38592), .ZN(n2121) );
  OAI22_X1 U38688 ( .A1(n38598), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[90][3] ), .B2(n38597), .ZN(n38593) );
  INV_X1 U38689 ( .A(n38593), .ZN(n2120) );
  OAI22_X1 U38690 ( .A1(n38598), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[90][4] ), .B2(n38597), .ZN(n38594) );
  INV_X1 U38691 ( .A(n38594), .ZN(n2119) );
  OAI22_X1 U38692 ( .A1(n38598), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[90][5] ), .B2(n38597), .ZN(n38595) );
  INV_X1 U38693 ( .A(n38595), .ZN(n2118) );
  OAI22_X1 U38694 ( .A1(n38598), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[90][6] ), .B2(n38597), .ZN(n38596) );
  INV_X1 U38695 ( .A(n38596), .ZN(n2117) );
  OAI22_X1 U38696 ( .A1(n38598), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[90][7] ), .B2(n38597), .ZN(n38599) );
  INV_X1 U38697 ( .A(n38599), .ZN(n2116) );
  NOR2_X1 U38698 ( .A1(n38935), .A2(n38640), .ZN(n38607) );
  INV_X1 U38699 ( .A(n38607), .ZN(n38608) );
  OAI22_X1 U38700 ( .A1(n38608), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[91][0] ), .B2(n38607), .ZN(n38600) );
  INV_X1 U38701 ( .A(n38600), .ZN(n2115) );
  OAI22_X1 U38702 ( .A1(n38608), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[91][1] ), .B2(n38607), .ZN(n38601) );
  INV_X1 U38703 ( .A(n38601), .ZN(n2114) );
  OAI22_X1 U38704 ( .A1(n38608), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[91][2] ), .B2(n38607), .ZN(n38602) );
  INV_X1 U38705 ( .A(n38602), .ZN(n2113) );
  OAI22_X1 U38706 ( .A1(n38608), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[91][3] ), .B2(n38607), .ZN(n38603) );
  INV_X1 U38707 ( .A(n38603), .ZN(n2112) );
  OAI22_X1 U38708 ( .A1(n38608), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[91][4] ), .B2(n38607), .ZN(n38604) );
  INV_X1 U38709 ( .A(n38604), .ZN(n2111) );
  OAI22_X1 U38710 ( .A1(n38608), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[91][5] ), .B2(n38607), .ZN(n38605) );
  INV_X1 U38711 ( .A(n38605), .ZN(n2110) );
  OAI22_X1 U38712 ( .A1(n38608), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[91][6] ), .B2(n38607), .ZN(n38606) );
  INV_X1 U38713 ( .A(n38606), .ZN(n2109) );
  OAI22_X1 U38714 ( .A1(n38608), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[91][7] ), .B2(n38607), .ZN(n38609) );
  INV_X1 U38715 ( .A(n38609), .ZN(n2108) );
  NOR2_X1 U38716 ( .A1(n38946), .A2(n38640), .ZN(n38617) );
  INV_X1 U38717 ( .A(n38617), .ZN(n38618) );
  OAI22_X1 U38718 ( .A1(n38618), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[92][0] ), .B2(n38617), .ZN(n38610) );
  INV_X1 U38719 ( .A(n38610), .ZN(n2107) );
  OAI22_X1 U38720 ( .A1(n38618), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[92][1] ), .B2(n38617), .ZN(n38611) );
  INV_X1 U38721 ( .A(n38611), .ZN(n2106) );
  OAI22_X1 U38722 ( .A1(n38618), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[92][2] ), .B2(n38617), .ZN(n38612) );
  INV_X1 U38723 ( .A(n38612), .ZN(n2105) );
  OAI22_X1 U38724 ( .A1(n38618), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[92][3] ), .B2(n38617), .ZN(n38613) );
  INV_X1 U38725 ( .A(n38613), .ZN(n2104) );
  OAI22_X1 U38726 ( .A1(n38618), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[92][4] ), .B2(n38617), .ZN(n38614) );
  INV_X1 U38727 ( .A(n38614), .ZN(n2103) );
  OAI22_X1 U38728 ( .A1(n38618), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[92][5] ), .B2(n38617), .ZN(n38615) );
  INV_X1 U38729 ( .A(n38615), .ZN(n2102) );
  OAI22_X1 U38730 ( .A1(n38618), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[92][6] ), .B2(n38617), .ZN(n38616) );
  INV_X1 U38731 ( .A(n38616), .ZN(n2101) );
  OAI22_X1 U38732 ( .A1(n38618), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[92][7] ), .B2(n38617), .ZN(n38619) );
  INV_X1 U38733 ( .A(n38619), .ZN(n2100) );
  NOR2_X1 U38734 ( .A1(n38957), .A2(n38640), .ZN(n38627) );
  INV_X1 U38735 ( .A(n38627), .ZN(n38628) );
  OAI22_X1 U38736 ( .A1(n38628), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[93][0] ), .B2(n38627), .ZN(n38620) );
  INV_X1 U38737 ( .A(n38620), .ZN(n2099) );
  OAI22_X1 U38738 ( .A1(n38628), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[93][1] ), .B2(n38627), .ZN(n38621) );
  INV_X1 U38739 ( .A(n38621), .ZN(n2098) );
  OAI22_X1 U38740 ( .A1(n38628), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[93][2] ), .B2(n38627), .ZN(n38622) );
  INV_X1 U38741 ( .A(n38622), .ZN(n2097) );
  OAI22_X1 U38742 ( .A1(n38628), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[93][3] ), .B2(n38627), .ZN(n38623) );
  INV_X1 U38743 ( .A(n38623), .ZN(n2096) );
  OAI22_X1 U38744 ( .A1(n38628), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[93][4] ), .B2(n38627), .ZN(n38624) );
  INV_X1 U38745 ( .A(n38624), .ZN(n2095) );
  OAI22_X1 U38746 ( .A1(n38628), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[93][5] ), .B2(n38627), .ZN(n38625) );
  INV_X1 U38747 ( .A(n38625), .ZN(n2094) );
  OAI22_X1 U38748 ( .A1(n38628), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[93][6] ), .B2(n38627), .ZN(n38626) );
  INV_X1 U38749 ( .A(n38626), .ZN(n2093) );
  OAI22_X1 U38750 ( .A1(n38628), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[93][7] ), .B2(n38627), .ZN(n38629) );
  INV_X1 U38751 ( .A(n38629), .ZN(n2092) );
  NOR2_X1 U38752 ( .A1(n38968), .A2(n38640), .ZN(n38637) );
  INV_X1 U38753 ( .A(n38637), .ZN(n38638) );
  OAI22_X1 U38754 ( .A1(n38638), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[94][0] ), .B2(n38637), .ZN(n38630) );
  INV_X1 U38755 ( .A(n38630), .ZN(n2091) );
  OAI22_X1 U38756 ( .A1(n38638), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[94][1] ), .B2(n38637), .ZN(n38631) );
  INV_X1 U38757 ( .A(n38631), .ZN(n2090) );
  OAI22_X1 U38758 ( .A1(n38638), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[94][2] ), .B2(n38637), .ZN(n38632) );
  INV_X1 U38759 ( .A(n38632), .ZN(n2089) );
  OAI22_X1 U38760 ( .A1(n38638), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[94][3] ), .B2(n38637), .ZN(n38633) );
  INV_X1 U38761 ( .A(n38633), .ZN(n2088) );
  OAI22_X1 U38762 ( .A1(n38638), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[94][4] ), .B2(n38637), .ZN(n38634) );
  INV_X1 U38763 ( .A(n38634), .ZN(n2087) );
  OAI22_X1 U38764 ( .A1(n38638), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[94][5] ), .B2(n38637), .ZN(n38635) );
  INV_X1 U38765 ( .A(n38635), .ZN(n2086) );
  OAI22_X1 U38766 ( .A1(n38638), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[94][6] ), .B2(n38637), .ZN(n38636) );
  INV_X1 U38767 ( .A(n38636), .ZN(n2085) );
  OAI22_X1 U38768 ( .A1(n38638), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[94][7] ), .B2(n38637), .ZN(n38639) );
  INV_X1 U38769 ( .A(n38639), .ZN(n2084) );
  NOR2_X1 U38770 ( .A1(n38803), .A2(n38640), .ZN(n38648) );
  INV_X1 U38771 ( .A(n38648), .ZN(n38649) );
  OAI22_X1 U38772 ( .A1(n38649), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[95][0] ), .B2(n38648), .ZN(n38641) );
  INV_X1 U38773 ( .A(n38641), .ZN(n2083) );
  OAI22_X1 U38774 ( .A1(n38649), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[95][1] ), .B2(n38648), .ZN(n38642) );
  INV_X1 U38775 ( .A(n38642), .ZN(n2082) );
  OAI22_X1 U38776 ( .A1(n38649), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[95][2] ), .B2(n38648), .ZN(n38643) );
  INV_X1 U38777 ( .A(n38643), .ZN(n2081) );
  OAI22_X1 U38778 ( .A1(n38649), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[95][3] ), .B2(n38648), .ZN(n38644) );
  INV_X1 U38779 ( .A(n38644), .ZN(n2080) );
  OAI22_X1 U38780 ( .A1(n38649), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[95][4] ), .B2(n38648), .ZN(n38645) );
  INV_X1 U38781 ( .A(n38645), .ZN(n2079) );
  OAI22_X1 U38782 ( .A1(n38649), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[95][5] ), .B2(n38648), .ZN(n38646) );
  INV_X1 U38783 ( .A(n38646), .ZN(n2078) );
  OAI22_X1 U38784 ( .A1(n38649), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[95][6] ), .B2(n38648), .ZN(n38647) );
  INV_X1 U38785 ( .A(n38647), .ZN(n2077) );
  OAI22_X1 U38786 ( .A1(n38649), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[95][7] ), .B2(n38648), .ZN(n38650) );
  INV_X1 U38787 ( .A(n38650), .ZN(n2076) );
  NAND3_X1 U38788 ( .A1(xmem_addr[6]), .A2(xmem_addr[5]), .A3(n38651), .ZN(
        n38802) );
  NOR2_X1 U38789 ( .A1(n38814), .A2(n38802), .ZN(n38659) );
  INV_X1 U38790 ( .A(n38659), .ZN(n38660) );
  OAI22_X1 U38791 ( .A1(n38660), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[96][0] ), .B2(n38659), .ZN(n38652) );
  INV_X1 U38792 ( .A(n38652), .ZN(n2075) );
  OAI22_X1 U38793 ( .A1(n38660), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[96][1] ), .B2(n38659), .ZN(n38653) );
  INV_X1 U38794 ( .A(n38653), .ZN(n2074) );
  OAI22_X1 U38795 ( .A1(n38660), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[96][2] ), .B2(n38659), .ZN(n38654) );
  INV_X1 U38796 ( .A(n38654), .ZN(n2073) );
  OAI22_X1 U38797 ( .A1(n38660), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[96][3] ), .B2(n38659), .ZN(n38655) );
  INV_X1 U38798 ( .A(n38655), .ZN(n2072) );
  OAI22_X1 U38799 ( .A1(n38660), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[96][4] ), .B2(n38659), .ZN(n38656) );
  INV_X1 U38800 ( .A(n38656), .ZN(n2071) );
  OAI22_X1 U38801 ( .A1(n38660), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[96][5] ), .B2(n38659), .ZN(n38657) );
  INV_X1 U38802 ( .A(n38657), .ZN(n2070) );
  OAI22_X1 U38803 ( .A1(n38660), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[96][6] ), .B2(n38659), .ZN(n38658) );
  INV_X1 U38804 ( .A(n38658), .ZN(n2069) );
  OAI22_X1 U38805 ( .A1(n38660), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[96][7] ), .B2(n38659), .ZN(n38661) );
  INV_X1 U38806 ( .A(n38661), .ZN(n2068) );
  NOR2_X1 U38807 ( .A1(n38825), .A2(n38802), .ZN(n38669) );
  INV_X1 U38808 ( .A(n38669), .ZN(n38670) );
  OAI22_X1 U38809 ( .A1(n38670), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[97][0] ), .B2(n38669), .ZN(n38662) );
  INV_X1 U38810 ( .A(n38662), .ZN(n2067) );
  OAI22_X1 U38811 ( .A1(n38670), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[97][1] ), .B2(n38669), .ZN(n38663) );
  INV_X1 U38812 ( .A(n38663), .ZN(n2066) );
  OAI22_X1 U38813 ( .A1(n38670), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[97][2] ), .B2(n38669), .ZN(n38664) );
  INV_X1 U38814 ( .A(n38664), .ZN(n2065) );
  OAI22_X1 U38815 ( .A1(n38670), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[97][3] ), .B2(n38669), .ZN(n38665) );
  INV_X1 U38816 ( .A(n38665), .ZN(n2064) );
  OAI22_X1 U38817 ( .A1(n38670), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[97][4] ), .B2(n38669), .ZN(n38666) );
  INV_X1 U38818 ( .A(n38666), .ZN(n2063) );
  OAI22_X1 U38819 ( .A1(n38670), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[97][5] ), .B2(n38669), .ZN(n38667) );
  INV_X1 U38820 ( .A(n38667), .ZN(n2062) );
  OAI22_X1 U38821 ( .A1(n38670), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[97][6] ), .B2(n38669), .ZN(n38668) );
  INV_X1 U38822 ( .A(n38668), .ZN(n2061) );
  OAI22_X1 U38823 ( .A1(n38670), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[97][7] ), .B2(n38669), .ZN(n38671) );
  INV_X1 U38824 ( .A(n38671), .ZN(n2060) );
  NOR2_X1 U38825 ( .A1(n38836), .A2(n38802), .ZN(n38679) );
  INV_X1 U38826 ( .A(n38679), .ZN(n38680) );
  OAI22_X1 U38827 ( .A1(n38680), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[98][0] ), .B2(n38679), .ZN(n38672) );
  INV_X1 U38828 ( .A(n38672), .ZN(n2059) );
  OAI22_X1 U38829 ( .A1(n38680), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[98][1] ), .B2(n38679), .ZN(n38673) );
  INV_X1 U38830 ( .A(n38673), .ZN(n2058) );
  OAI22_X1 U38831 ( .A1(n38680), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[98][2] ), .B2(n38679), .ZN(n38674) );
  INV_X1 U38832 ( .A(n38674), .ZN(n2057) );
  OAI22_X1 U38833 ( .A1(n38680), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[98][3] ), .B2(n38679), .ZN(n38675) );
  INV_X1 U38834 ( .A(n38675), .ZN(n2056) );
  OAI22_X1 U38835 ( .A1(n38680), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[98][4] ), .B2(n38679), .ZN(n38676) );
  INV_X1 U38836 ( .A(n38676), .ZN(n2055) );
  OAI22_X1 U38837 ( .A1(n38680), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[98][5] ), .B2(n38679), .ZN(n38677) );
  INV_X1 U38838 ( .A(n38677), .ZN(n2054) );
  OAI22_X1 U38839 ( .A1(n38680), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[98][6] ), .B2(n38679), .ZN(n38678) );
  INV_X1 U38840 ( .A(n38678), .ZN(n2053) );
  OAI22_X1 U38841 ( .A1(n38680), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[98][7] ), .B2(n38679), .ZN(n38681) );
  INV_X1 U38842 ( .A(n38681), .ZN(n2052) );
  NOR2_X1 U38843 ( .A1(n38847), .A2(n38802), .ZN(n38689) );
  INV_X1 U38844 ( .A(n38689), .ZN(n38690) );
  OAI22_X1 U38845 ( .A1(n38690), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[99][0] ), .B2(n38689), .ZN(n38682) );
  INV_X1 U38846 ( .A(n38682), .ZN(n2051) );
  OAI22_X1 U38847 ( .A1(n38690), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[99][1] ), .B2(n38689), .ZN(n38683) );
  INV_X1 U38848 ( .A(n38683), .ZN(n2050) );
  OAI22_X1 U38849 ( .A1(n38690), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[99][2] ), .B2(n38689), .ZN(n38684) );
  INV_X1 U38850 ( .A(n38684), .ZN(n2049) );
  OAI22_X1 U38851 ( .A1(n38690), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[99][3] ), .B2(n38689), .ZN(n38685) );
  INV_X1 U38852 ( .A(n38685), .ZN(n2048) );
  OAI22_X1 U38853 ( .A1(n38690), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[99][4] ), .B2(n38689), .ZN(n38686) );
  INV_X1 U38854 ( .A(n38686), .ZN(n2047) );
  OAI22_X1 U38855 ( .A1(n38690), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[99][5] ), .B2(n38689), .ZN(n38687) );
  INV_X1 U38856 ( .A(n38687), .ZN(n2046) );
  OAI22_X1 U38857 ( .A1(n38690), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[99][6] ), .B2(n38689), .ZN(n38688) );
  INV_X1 U38858 ( .A(n38688), .ZN(n2045) );
  OAI22_X1 U38859 ( .A1(n38690), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[99][7] ), .B2(n38689), .ZN(n38691) );
  INV_X1 U38860 ( .A(n38691), .ZN(n2044) );
  NOR2_X1 U38861 ( .A1(n38858), .A2(n38802), .ZN(n38699) );
  INV_X1 U38862 ( .A(n38699), .ZN(n38700) );
  OAI22_X1 U38863 ( .A1(n38700), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[100][0] ), .B2(n38699), .ZN(n38692) );
  INV_X1 U38864 ( .A(n38692), .ZN(n2043) );
  OAI22_X1 U38865 ( .A1(n38700), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[100][1] ), .B2(n38699), .ZN(n38693) );
  INV_X1 U38866 ( .A(n38693), .ZN(n2042) );
  OAI22_X1 U38867 ( .A1(n38700), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[100][2] ), .B2(n38699), .ZN(n38694) );
  INV_X1 U38868 ( .A(n38694), .ZN(n2041) );
  OAI22_X1 U38869 ( .A1(n38700), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[100][3] ), .B2(n38699), .ZN(n38695) );
  INV_X1 U38870 ( .A(n38695), .ZN(n2040) );
  OAI22_X1 U38871 ( .A1(n38700), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[100][4] ), .B2(n38699), .ZN(n38696) );
  INV_X1 U38872 ( .A(n38696), .ZN(n2039) );
  OAI22_X1 U38873 ( .A1(n38700), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[100][5] ), .B2(n38699), .ZN(n38697) );
  INV_X1 U38874 ( .A(n38697), .ZN(n2038) );
  OAI22_X1 U38875 ( .A1(n38700), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[100][6] ), .B2(n38699), .ZN(n38698) );
  INV_X1 U38876 ( .A(n38698), .ZN(n2037) );
  OAI22_X1 U38877 ( .A1(n38700), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[100][7] ), .B2(n38699), .ZN(n38701) );
  INV_X1 U38878 ( .A(n38701), .ZN(n2036) );
  NOR2_X1 U38879 ( .A1(n38869), .A2(n38802), .ZN(n38709) );
  INV_X1 U38880 ( .A(n38709), .ZN(n38710) );
  OAI22_X1 U38881 ( .A1(n38710), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[101][0] ), .B2(n38709), .ZN(n38702) );
  INV_X1 U38882 ( .A(n38702), .ZN(n2035) );
  OAI22_X1 U38883 ( .A1(n38710), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[101][1] ), .B2(n38709), .ZN(n38703) );
  INV_X1 U38884 ( .A(n38703), .ZN(n2034) );
  OAI22_X1 U38885 ( .A1(n38710), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[101][2] ), .B2(n38709), .ZN(n38704) );
  INV_X1 U38886 ( .A(n38704), .ZN(n2033) );
  OAI22_X1 U38887 ( .A1(n38710), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[101][3] ), .B2(n38709), .ZN(n38705) );
  INV_X1 U38888 ( .A(n38705), .ZN(n2032) );
  OAI22_X1 U38889 ( .A1(n38710), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[101][4] ), .B2(n38709), .ZN(n38706) );
  INV_X1 U38890 ( .A(n38706), .ZN(n2031) );
  OAI22_X1 U38891 ( .A1(n38710), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[101][5] ), .B2(n38709), .ZN(n38707) );
  INV_X1 U38892 ( .A(n38707), .ZN(n2030) );
  OAI22_X1 U38893 ( .A1(n38710), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[101][6] ), .B2(n38709), .ZN(n38708) );
  INV_X1 U38894 ( .A(n38708), .ZN(n2029) );
  OAI22_X1 U38895 ( .A1(n38710), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[101][7] ), .B2(n38709), .ZN(n38711) );
  INV_X1 U38896 ( .A(n38711), .ZN(n2028) );
  NOR2_X1 U38897 ( .A1(n38880), .A2(n38802), .ZN(n38719) );
  INV_X1 U38898 ( .A(n38719), .ZN(n38720) );
  OAI22_X1 U38899 ( .A1(n38720), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[102][0] ), .B2(n38719), .ZN(n38712) );
  INV_X1 U38900 ( .A(n38712), .ZN(n2027) );
  OAI22_X1 U38901 ( .A1(n38720), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[102][1] ), .B2(n38719), .ZN(n38713) );
  INV_X1 U38902 ( .A(n38713), .ZN(n2026) );
  OAI22_X1 U38903 ( .A1(n38720), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[102][2] ), .B2(n38719), .ZN(n38714) );
  INV_X1 U38904 ( .A(n38714), .ZN(n2025) );
  OAI22_X1 U38905 ( .A1(n38720), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[102][3] ), .B2(n38719), .ZN(n38715) );
  INV_X1 U38906 ( .A(n38715), .ZN(n2024) );
  OAI22_X1 U38907 ( .A1(n38720), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[102][4] ), .B2(n38719), .ZN(n38716) );
  INV_X1 U38908 ( .A(n38716), .ZN(n2023) );
  OAI22_X1 U38909 ( .A1(n38720), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[102][5] ), .B2(n38719), .ZN(n38717) );
  INV_X1 U38910 ( .A(n38717), .ZN(n2022) );
  OAI22_X1 U38911 ( .A1(n38720), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[102][6] ), .B2(n38719), .ZN(n38718) );
  INV_X1 U38912 ( .A(n38718), .ZN(n2021) );
  OAI22_X1 U38913 ( .A1(n38720), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[102][7] ), .B2(n38719), .ZN(n38721) );
  INV_X1 U38914 ( .A(n38721), .ZN(n2020) );
  NOR2_X1 U38915 ( .A1(n38891), .A2(n38802), .ZN(n38729) );
  INV_X1 U38916 ( .A(n38729), .ZN(n38730) );
  OAI22_X1 U38917 ( .A1(n38730), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[103][0] ), .B2(n38729), .ZN(n38722) );
  INV_X1 U38918 ( .A(n38722), .ZN(n2019) );
  OAI22_X1 U38919 ( .A1(n38730), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[103][1] ), .B2(n38729), .ZN(n38723) );
  INV_X1 U38920 ( .A(n38723), .ZN(n2018) );
  OAI22_X1 U38921 ( .A1(n38730), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[103][2] ), .B2(n38729), .ZN(n38724) );
  INV_X1 U38922 ( .A(n38724), .ZN(n2017) );
  OAI22_X1 U38923 ( .A1(n38730), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[103][3] ), .B2(n38729), .ZN(n38725) );
  INV_X1 U38924 ( .A(n38725), .ZN(n2016) );
  OAI22_X1 U38925 ( .A1(n38730), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[103][4] ), .B2(n38729), .ZN(n38726) );
  INV_X1 U38926 ( .A(n38726), .ZN(n2015) );
  OAI22_X1 U38927 ( .A1(n38730), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[103][5] ), .B2(n38729), .ZN(n38727) );
  INV_X1 U38928 ( .A(n38727), .ZN(n2014) );
  OAI22_X1 U38929 ( .A1(n38730), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[103][6] ), .B2(n38729), .ZN(n38728) );
  INV_X1 U38930 ( .A(n38728), .ZN(n2013) );
  OAI22_X1 U38931 ( .A1(n38730), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[103][7] ), .B2(n38729), .ZN(n38731) );
  INV_X1 U38932 ( .A(n38731), .ZN(n2012) );
  NOR2_X1 U38933 ( .A1(n38902), .A2(n38802), .ZN(n38739) );
  INV_X1 U38934 ( .A(n38739), .ZN(n38740) );
  OAI22_X1 U38935 ( .A1(n38740), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[104][0] ), .B2(n38739), .ZN(n38732) );
  INV_X1 U38936 ( .A(n38732), .ZN(n2011) );
  OAI22_X1 U38937 ( .A1(n38740), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[104][1] ), .B2(n38739), .ZN(n38733) );
  INV_X1 U38938 ( .A(n38733), .ZN(n2010) );
  OAI22_X1 U38939 ( .A1(n38740), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[104][2] ), .B2(n38739), .ZN(n38734) );
  INV_X1 U38940 ( .A(n38734), .ZN(n2009) );
  OAI22_X1 U38941 ( .A1(n38740), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[104][3] ), .B2(n38739), .ZN(n38735) );
  INV_X1 U38942 ( .A(n38735), .ZN(n2008) );
  OAI22_X1 U38943 ( .A1(n38740), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[104][4] ), .B2(n38739), .ZN(n38736) );
  INV_X1 U38944 ( .A(n38736), .ZN(n2007) );
  OAI22_X1 U38945 ( .A1(n38740), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[104][5] ), .B2(n38739), .ZN(n38737) );
  INV_X1 U38946 ( .A(n38737), .ZN(n2006) );
  OAI22_X1 U38947 ( .A1(n38740), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[104][6] ), .B2(n38739), .ZN(n38738) );
  INV_X1 U38948 ( .A(n38738), .ZN(n2005) );
  OAI22_X1 U38949 ( .A1(n38740), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[104][7] ), .B2(n38739), .ZN(n38741) );
  INV_X1 U38950 ( .A(n38741), .ZN(n2004) );
  NOR2_X1 U38951 ( .A1(n38913), .A2(n38802), .ZN(n38749) );
  INV_X1 U38952 ( .A(n38749), .ZN(n38750) );
  OAI22_X1 U38953 ( .A1(n38750), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[105][0] ), .B2(n38749), .ZN(n38742) );
  INV_X1 U38954 ( .A(n38742), .ZN(n2003) );
  OAI22_X1 U38955 ( .A1(n38750), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[105][1] ), .B2(n38749), .ZN(n38743) );
  INV_X1 U38956 ( .A(n38743), .ZN(n2002) );
  OAI22_X1 U38957 ( .A1(n38750), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[105][2] ), .B2(n38749), .ZN(n38744) );
  INV_X1 U38958 ( .A(n38744), .ZN(n2001) );
  OAI22_X1 U38959 ( .A1(n38750), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[105][3] ), .B2(n38749), .ZN(n38745) );
  INV_X1 U38960 ( .A(n38745), .ZN(n2000) );
  OAI22_X1 U38961 ( .A1(n38750), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[105][4] ), .B2(n38749), .ZN(n38746) );
  INV_X1 U38962 ( .A(n38746), .ZN(n1999) );
  OAI22_X1 U38963 ( .A1(n38750), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[105][5] ), .B2(n38749), .ZN(n38747) );
  INV_X1 U38964 ( .A(n38747), .ZN(n1998) );
  OAI22_X1 U38965 ( .A1(n38750), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[105][6] ), .B2(n38749), .ZN(n38748) );
  INV_X1 U38966 ( .A(n38748), .ZN(n1997) );
  OAI22_X1 U38967 ( .A1(n38750), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[105][7] ), .B2(n38749), .ZN(n38751) );
  INV_X1 U38968 ( .A(n38751), .ZN(n1996) );
  NOR2_X1 U38969 ( .A1(n38924), .A2(n38802), .ZN(n38759) );
  INV_X1 U38970 ( .A(n38759), .ZN(n38760) );
  OAI22_X1 U38971 ( .A1(n38760), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[106][0] ), .B2(n38759), .ZN(n38752) );
  INV_X1 U38972 ( .A(n38752), .ZN(n1995) );
  OAI22_X1 U38973 ( .A1(n38760), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[106][1] ), .B2(n38759), .ZN(n38753) );
  INV_X1 U38974 ( .A(n38753), .ZN(n1994) );
  OAI22_X1 U38975 ( .A1(n38760), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[106][2] ), .B2(n38759), .ZN(n38754) );
  INV_X1 U38976 ( .A(n38754), .ZN(n1993) );
  OAI22_X1 U38977 ( .A1(n38760), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[106][3] ), .B2(n38759), .ZN(n38755) );
  INV_X1 U38978 ( .A(n38755), .ZN(n1992) );
  OAI22_X1 U38979 ( .A1(n38760), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[106][4] ), .B2(n38759), .ZN(n38756) );
  INV_X1 U38980 ( .A(n38756), .ZN(n1991) );
  OAI22_X1 U38981 ( .A1(n38760), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[106][5] ), .B2(n38759), .ZN(n38757) );
  INV_X1 U38982 ( .A(n38757), .ZN(n1990) );
  OAI22_X1 U38983 ( .A1(n38760), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[106][6] ), .B2(n38759), .ZN(n38758) );
  INV_X1 U38984 ( .A(n38758), .ZN(n1989) );
  OAI22_X1 U38985 ( .A1(n38760), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[106][7] ), .B2(n38759), .ZN(n38761) );
  INV_X1 U38986 ( .A(n38761), .ZN(n1988) );
  NOR2_X1 U38987 ( .A1(n38935), .A2(n38802), .ZN(n38769) );
  INV_X1 U38988 ( .A(n38769), .ZN(n38770) );
  OAI22_X1 U38989 ( .A1(n38770), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[107][0] ), .B2(n38769), .ZN(n38762) );
  INV_X1 U38990 ( .A(n38762), .ZN(n1987) );
  OAI22_X1 U38991 ( .A1(n38770), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[107][1] ), .B2(n38769), .ZN(n38763) );
  INV_X1 U38992 ( .A(n38763), .ZN(n1986) );
  OAI22_X1 U38993 ( .A1(n38770), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[107][2] ), .B2(n38769), .ZN(n38764) );
  INV_X1 U38994 ( .A(n38764), .ZN(n1985) );
  OAI22_X1 U38995 ( .A1(n38770), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[107][3] ), .B2(n38769), .ZN(n38765) );
  INV_X1 U38996 ( .A(n38765), .ZN(n1984) );
  OAI22_X1 U38997 ( .A1(n38770), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[107][4] ), .B2(n38769), .ZN(n38766) );
  INV_X1 U38998 ( .A(n38766), .ZN(n1983) );
  OAI22_X1 U38999 ( .A1(n38770), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[107][5] ), .B2(n38769), .ZN(n38767) );
  INV_X1 U39000 ( .A(n38767), .ZN(n1982) );
  OAI22_X1 U39001 ( .A1(n38770), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[107][6] ), .B2(n38769), .ZN(n38768) );
  INV_X1 U39002 ( .A(n38768), .ZN(n1981) );
  OAI22_X1 U39003 ( .A1(n38770), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[107][7] ), .B2(n38769), .ZN(n38771) );
  INV_X1 U39004 ( .A(n38771), .ZN(n1980) );
  NOR2_X1 U39005 ( .A1(n38946), .A2(n38802), .ZN(n38779) );
  INV_X1 U39006 ( .A(n38779), .ZN(n38780) );
  OAI22_X1 U39007 ( .A1(n38780), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[108][0] ), .B2(n38779), .ZN(n38772) );
  INV_X1 U39008 ( .A(n38772), .ZN(n1979) );
  OAI22_X1 U39009 ( .A1(n38780), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[108][1] ), .B2(n38779), .ZN(n38773) );
  INV_X1 U39010 ( .A(n38773), .ZN(n1978) );
  OAI22_X1 U39011 ( .A1(n38780), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[108][2] ), .B2(n38779), .ZN(n38774) );
  INV_X1 U39012 ( .A(n38774), .ZN(n1977) );
  OAI22_X1 U39013 ( .A1(n38780), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[108][3] ), .B2(n38779), .ZN(n38775) );
  INV_X1 U39014 ( .A(n38775), .ZN(n1976) );
  OAI22_X1 U39015 ( .A1(n38780), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[108][4] ), .B2(n38779), .ZN(n38776) );
  INV_X1 U39016 ( .A(n38776), .ZN(n1975) );
  OAI22_X1 U39017 ( .A1(n38780), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[108][5] ), .B2(n38779), .ZN(n38777) );
  INV_X1 U39018 ( .A(n38777), .ZN(n1974) );
  OAI22_X1 U39019 ( .A1(n38780), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[108][6] ), .B2(n38779), .ZN(n38778) );
  INV_X1 U39020 ( .A(n38778), .ZN(n1973) );
  OAI22_X1 U39021 ( .A1(n38780), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[108][7] ), .B2(n38779), .ZN(n38781) );
  INV_X1 U39022 ( .A(n38781), .ZN(n1972) );
  NOR2_X1 U39023 ( .A1(n38957), .A2(n38802), .ZN(n38789) );
  INV_X1 U39024 ( .A(n38789), .ZN(n38790) );
  OAI22_X1 U39025 ( .A1(n38790), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[109][0] ), .B2(n38789), .ZN(n38782) );
  INV_X1 U39026 ( .A(n38782), .ZN(n1971) );
  OAI22_X1 U39027 ( .A1(n38790), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[109][1] ), .B2(n38789), .ZN(n38783) );
  INV_X1 U39028 ( .A(n38783), .ZN(n1970) );
  OAI22_X1 U39029 ( .A1(n38790), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[109][2] ), .B2(n38789), .ZN(n38784) );
  INV_X1 U39030 ( .A(n38784), .ZN(n1969) );
  OAI22_X1 U39031 ( .A1(n38790), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[109][3] ), .B2(n38789), .ZN(n38785) );
  INV_X1 U39032 ( .A(n38785), .ZN(n1968) );
  OAI22_X1 U39033 ( .A1(n38790), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[109][4] ), .B2(n38789), .ZN(n38786) );
  INV_X1 U39034 ( .A(n38786), .ZN(n1967) );
  OAI22_X1 U39035 ( .A1(n38790), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[109][5] ), .B2(n38789), .ZN(n38787) );
  INV_X1 U39036 ( .A(n38787), .ZN(n1966) );
  OAI22_X1 U39037 ( .A1(n38790), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[109][6] ), .B2(n38789), .ZN(n38788) );
  INV_X1 U39038 ( .A(n38788), .ZN(n1965) );
  OAI22_X1 U39039 ( .A1(n38790), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[109][7] ), .B2(n38789), .ZN(n38791) );
  INV_X1 U39040 ( .A(n38791), .ZN(n1964) );
  NOR2_X1 U39041 ( .A1(n38968), .A2(n38802), .ZN(n38799) );
  INV_X1 U39042 ( .A(n38799), .ZN(n38800) );
  OAI22_X1 U39043 ( .A1(n38800), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[110][0] ), .B2(n38799), .ZN(n38792) );
  INV_X1 U39044 ( .A(n38792), .ZN(n1963) );
  OAI22_X1 U39045 ( .A1(n38800), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[110][1] ), .B2(n38799), .ZN(n38793) );
  INV_X1 U39046 ( .A(n38793), .ZN(n1962) );
  OAI22_X1 U39047 ( .A1(n38800), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[110][2] ), .B2(n38799), .ZN(n38794) );
  INV_X1 U39048 ( .A(n38794), .ZN(n1961) );
  OAI22_X1 U39049 ( .A1(n38800), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[110][3] ), .B2(n38799), .ZN(n38795) );
  INV_X1 U39050 ( .A(n38795), .ZN(n1960) );
  OAI22_X1 U39051 ( .A1(n38800), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[110][4] ), .B2(n38799), .ZN(n38796) );
  INV_X1 U39052 ( .A(n38796), .ZN(n1959) );
  OAI22_X1 U39053 ( .A1(n38800), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[110][5] ), .B2(n38799), .ZN(n38797) );
  INV_X1 U39054 ( .A(n38797), .ZN(n1958) );
  OAI22_X1 U39055 ( .A1(n38800), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[110][6] ), .B2(n38799), .ZN(n38798) );
  INV_X1 U39056 ( .A(n38798), .ZN(n1957) );
  OAI22_X1 U39057 ( .A1(n38800), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[110][7] ), .B2(n38799), .ZN(n38801) );
  INV_X1 U39058 ( .A(n38801), .ZN(n1956) );
  NOR2_X1 U39059 ( .A1(n38803), .A2(n38802), .ZN(n38811) );
  INV_X1 U39060 ( .A(n38811), .ZN(n38812) );
  OAI22_X1 U39061 ( .A1(n38812), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[111][0] ), .B2(n38811), .ZN(n38804) );
  INV_X1 U39062 ( .A(n38804), .ZN(n1955) );
  OAI22_X1 U39063 ( .A1(n38812), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[111][1] ), .B2(n38811), .ZN(n38805) );
  INV_X1 U39064 ( .A(n38805), .ZN(n1954) );
  OAI22_X1 U39065 ( .A1(n38812), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[111][2] ), .B2(n38811), .ZN(n38806) );
  INV_X1 U39066 ( .A(n38806), .ZN(n1953) );
  OAI22_X1 U39067 ( .A1(n38812), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[111][3] ), .B2(n38811), .ZN(n38807) );
  INV_X1 U39068 ( .A(n38807), .ZN(n1952) );
  OAI22_X1 U39069 ( .A1(n38812), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[111][4] ), .B2(n38811), .ZN(n38808) );
  INV_X1 U39070 ( .A(n38808), .ZN(n1951) );
  OAI22_X1 U39071 ( .A1(n38812), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[111][5] ), .B2(n38811), .ZN(n38809) );
  INV_X1 U39072 ( .A(n38809), .ZN(n1950) );
  OAI22_X1 U39073 ( .A1(n38812), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[111][6] ), .B2(n38811), .ZN(n38810) );
  INV_X1 U39074 ( .A(n38810), .ZN(n1949) );
  OAI22_X1 U39075 ( .A1(n38812), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[111][7] ), .B2(n38811), .ZN(n38813) );
  INV_X1 U39076 ( .A(n38813), .ZN(n1948) );
  NOR2_X1 U39077 ( .A1(n38969), .A2(n38814), .ZN(n38822) );
  INV_X1 U39078 ( .A(n38822), .ZN(n38823) );
  OAI22_X1 U39079 ( .A1(n38823), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[112][0] ), .B2(n38822), .ZN(n38815) );
  INV_X1 U39080 ( .A(n38815), .ZN(n1947) );
  OAI22_X1 U39081 ( .A1(n38823), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[112][1] ), .B2(n38822), .ZN(n38816) );
  INV_X1 U39082 ( .A(n38816), .ZN(n1946) );
  OAI22_X1 U39083 ( .A1(n38823), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[112][2] ), .B2(n38822), .ZN(n38817) );
  INV_X1 U39084 ( .A(n38817), .ZN(n1945) );
  OAI22_X1 U39085 ( .A1(n38823), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[112][3] ), .B2(n38822), .ZN(n38818) );
  INV_X1 U39086 ( .A(n38818), .ZN(n1944) );
  OAI22_X1 U39087 ( .A1(n38823), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[112][4] ), .B2(n38822), .ZN(n38819) );
  INV_X1 U39088 ( .A(n38819), .ZN(n1943) );
  OAI22_X1 U39089 ( .A1(n38823), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[112][5] ), .B2(n38822), .ZN(n38820) );
  INV_X1 U39090 ( .A(n38820), .ZN(n1942) );
  OAI22_X1 U39091 ( .A1(n38823), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[112][6] ), .B2(n38822), .ZN(n38821) );
  INV_X1 U39092 ( .A(n38821), .ZN(n1941) );
  OAI22_X1 U39093 ( .A1(n38823), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[112][7] ), .B2(n38822), .ZN(n38824) );
  INV_X1 U39094 ( .A(n38824), .ZN(n1940) );
  NOR2_X1 U39095 ( .A1(n38969), .A2(n38825), .ZN(n38833) );
  INV_X1 U39096 ( .A(n38833), .ZN(n38834) );
  OAI22_X1 U39097 ( .A1(n38834), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[113][0] ), .B2(n38833), .ZN(n38826) );
  INV_X1 U39098 ( .A(n38826), .ZN(n1939) );
  OAI22_X1 U39099 ( .A1(n38834), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[113][1] ), .B2(n38833), .ZN(n38827) );
  INV_X1 U39100 ( .A(n38827), .ZN(n1938) );
  OAI22_X1 U39101 ( .A1(n38834), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[113][2] ), .B2(n38833), .ZN(n38828) );
  INV_X1 U39102 ( .A(n38828), .ZN(n1937) );
  OAI22_X1 U39103 ( .A1(n38834), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[113][3] ), .B2(n38833), .ZN(n38829) );
  INV_X1 U39104 ( .A(n38829), .ZN(n1936) );
  OAI22_X1 U39105 ( .A1(n38834), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[113][4] ), .B2(n38833), .ZN(n38830) );
  INV_X1 U39106 ( .A(n38830), .ZN(n1935) );
  OAI22_X1 U39107 ( .A1(n38834), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[113][5] ), .B2(n38833), .ZN(n38831) );
  INV_X1 U39108 ( .A(n38831), .ZN(n1934) );
  OAI22_X1 U39109 ( .A1(n38834), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[113][6] ), .B2(n38833), .ZN(n38832) );
  INV_X1 U39110 ( .A(n38832), .ZN(n1933) );
  OAI22_X1 U39111 ( .A1(n38834), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[113][7] ), .B2(n38833), .ZN(n38835) );
  INV_X1 U39112 ( .A(n38835), .ZN(n1932) );
  NOR2_X1 U39113 ( .A1(n38969), .A2(n38836), .ZN(n38844) );
  INV_X1 U39114 ( .A(n38844), .ZN(n38845) );
  OAI22_X1 U39115 ( .A1(n38845), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[114][0] ), .B2(n38844), .ZN(n38837) );
  INV_X1 U39116 ( .A(n38837), .ZN(n1931) );
  OAI22_X1 U39117 ( .A1(n38845), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[114][1] ), .B2(n38844), .ZN(n38838) );
  INV_X1 U39118 ( .A(n38838), .ZN(n1930) );
  OAI22_X1 U39119 ( .A1(n38845), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[114][2] ), .B2(n38844), .ZN(n38839) );
  INV_X1 U39120 ( .A(n38839), .ZN(n1929) );
  OAI22_X1 U39121 ( .A1(n38845), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[114][3] ), .B2(n38844), .ZN(n38840) );
  INV_X1 U39122 ( .A(n38840), .ZN(n1928) );
  OAI22_X1 U39123 ( .A1(n38845), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[114][4] ), .B2(n38844), .ZN(n38841) );
  INV_X1 U39124 ( .A(n38841), .ZN(n1927) );
  OAI22_X1 U39125 ( .A1(n38845), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[114][5] ), .B2(n38844), .ZN(n38842) );
  INV_X1 U39126 ( .A(n38842), .ZN(n1926) );
  OAI22_X1 U39127 ( .A1(n38845), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[114][6] ), .B2(n38844), .ZN(n38843) );
  INV_X1 U39128 ( .A(n38843), .ZN(n1925) );
  OAI22_X1 U39129 ( .A1(n38845), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[114][7] ), .B2(n38844), .ZN(n38846) );
  INV_X1 U39130 ( .A(n38846), .ZN(n1924) );
  NOR2_X1 U39131 ( .A1(n38969), .A2(n38847), .ZN(n38855) );
  INV_X1 U39132 ( .A(n38855), .ZN(n38856) );
  OAI22_X1 U39133 ( .A1(n38856), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[115][0] ), .B2(n38855), .ZN(n38848) );
  INV_X1 U39134 ( .A(n38848), .ZN(n1923) );
  OAI22_X1 U39135 ( .A1(n38856), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[115][1] ), .B2(n38855), .ZN(n38849) );
  INV_X1 U39136 ( .A(n38849), .ZN(n1922) );
  OAI22_X1 U39137 ( .A1(n38856), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[115][2] ), .B2(n38855), .ZN(n38850) );
  INV_X1 U39138 ( .A(n38850), .ZN(n1921) );
  OAI22_X1 U39139 ( .A1(n38856), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[115][3] ), .B2(n38855), .ZN(n38851) );
  INV_X1 U39140 ( .A(n38851), .ZN(n1920) );
  OAI22_X1 U39141 ( .A1(n38856), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[115][4] ), .B2(n38855), .ZN(n38852) );
  INV_X1 U39142 ( .A(n38852), .ZN(n1919) );
  OAI22_X1 U39143 ( .A1(n38856), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[115][5] ), .B2(n38855), .ZN(n38853) );
  INV_X1 U39144 ( .A(n38853), .ZN(n1918) );
  OAI22_X1 U39145 ( .A1(n38856), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[115][6] ), .B2(n38855), .ZN(n38854) );
  INV_X1 U39146 ( .A(n38854), .ZN(n1917) );
  OAI22_X1 U39147 ( .A1(n38856), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[115][7] ), .B2(n38855), .ZN(n38857) );
  INV_X1 U39148 ( .A(n38857), .ZN(n1916) );
  NOR2_X1 U39149 ( .A1(n38969), .A2(n38858), .ZN(n38866) );
  INV_X1 U39150 ( .A(n38866), .ZN(n38867) );
  OAI22_X1 U39151 ( .A1(n38867), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[116][0] ), .B2(n38866), .ZN(n38859) );
  INV_X1 U39152 ( .A(n38859), .ZN(n1915) );
  OAI22_X1 U39153 ( .A1(n38867), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[116][1] ), .B2(n38866), .ZN(n38860) );
  INV_X1 U39154 ( .A(n38860), .ZN(n1914) );
  OAI22_X1 U39155 ( .A1(n38867), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[116][2] ), .B2(n38866), .ZN(n38861) );
  INV_X1 U39156 ( .A(n38861), .ZN(n1913) );
  OAI22_X1 U39157 ( .A1(n38867), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[116][3] ), .B2(n38866), .ZN(n38862) );
  INV_X1 U39158 ( .A(n38862), .ZN(n1912) );
  OAI22_X1 U39159 ( .A1(n38867), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[116][4] ), .B2(n38866), .ZN(n38863) );
  INV_X1 U39160 ( .A(n38863), .ZN(n1911) );
  OAI22_X1 U39161 ( .A1(n38867), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[116][5] ), .B2(n38866), .ZN(n38864) );
  INV_X1 U39162 ( .A(n38864), .ZN(n1910) );
  OAI22_X1 U39163 ( .A1(n38867), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[116][6] ), .B2(n38866), .ZN(n38865) );
  INV_X1 U39164 ( .A(n38865), .ZN(n1909) );
  OAI22_X1 U39165 ( .A1(n38867), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[116][7] ), .B2(n38866), .ZN(n38868) );
  INV_X1 U39166 ( .A(n38868), .ZN(n1908) );
  NOR2_X1 U39167 ( .A1(n38969), .A2(n38869), .ZN(n38877) );
  INV_X1 U39168 ( .A(n38877), .ZN(n38878) );
  OAI22_X1 U39169 ( .A1(n38878), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[117][0] ), .B2(n38877), .ZN(n38870) );
  INV_X1 U39170 ( .A(n38870), .ZN(n1907) );
  OAI22_X1 U39171 ( .A1(n38878), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[117][1] ), .B2(n38877), .ZN(n38871) );
  INV_X1 U39172 ( .A(n38871), .ZN(n1906) );
  OAI22_X1 U39173 ( .A1(n38878), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[117][2] ), .B2(n38877), .ZN(n38872) );
  INV_X1 U39174 ( .A(n38872), .ZN(n1905) );
  OAI22_X1 U39175 ( .A1(n38878), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[117][3] ), .B2(n38877), .ZN(n38873) );
  INV_X1 U39176 ( .A(n38873), .ZN(n1904) );
  OAI22_X1 U39177 ( .A1(n38878), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[117][4] ), .B2(n38877), .ZN(n38874) );
  INV_X1 U39178 ( .A(n38874), .ZN(n1903) );
  OAI22_X1 U39179 ( .A1(n38878), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[117][5] ), .B2(n38877), .ZN(n38875) );
  INV_X1 U39180 ( .A(n38875), .ZN(n1902) );
  OAI22_X1 U39181 ( .A1(n38878), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[117][6] ), .B2(n38877), .ZN(n38876) );
  INV_X1 U39182 ( .A(n38876), .ZN(n1901) );
  OAI22_X1 U39183 ( .A1(n38878), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[117][7] ), .B2(n38877), .ZN(n38879) );
  INV_X1 U39184 ( .A(n38879), .ZN(n1900) );
  NOR2_X1 U39185 ( .A1(n38969), .A2(n38880), .ZN(n38888) );
  INV_X1 U39186 ( .A(n38888), .ZN(n38889) );
  OAI22_X1 U39187 ( .A1(n38889), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[118][0] ), .B2(n38888), .ZN(n38881) );
  INV_X1 U39188 ( .A(n38881), .ZN(n1899) );
  OAI22_X1 U39189 ( .A1(n38889), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[118][1] ), .B2(n38888), .ZN(n38882) );
  INV_X1 U39190 ( .A(n38882), .ZN(n1898) );
  OAI22_X1 U39191 ( .A1(n38889), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[118][2] ), .B2(n38888), .ZN(n38883) );
  INV_X1 U39192 ( .A(n38883), .ZN(n1897) );
  OAI22_X1 U39193 ( .A1(n38889), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[118][3] ), .B2(n38888), .ZN(n38884) );
  INV_X1 U39194 ( .A(n38884), .ZN(n1896) );
  OAI22_X1 U39195 ( .A1(n38889), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[118][4] ), .B2(n38888), .ZN(n38885) );
  INV_X1 U39196 ( .A(n38885), .ZN(n1895) );
  OAI22_X1 U39197 ( .A1(n38889), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[118][5] ), .B2(n38888), .ZN(n38886) );
  INV_X1 U39198 ( .A(n38886), .ZN(n1894) );
  OAI22_X1 U39199 ( .A1(n38889), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[118][6] ), .B2(n38888), .ZN(n38887) );
  INV_X1 U39200 ( .A(n38887), .ZN(n1893) );
  OAI22_X1 U39201 ( .A1(n38889), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[118][7] ), .B2(n38888), .ZN(n38890) );
  INV_X1 U39202 ( .A(n38890), .ZN(n1892) );
  NOR2_X1 U39203 ( .A1(n38891), .A2(n38969), .ZN(n38899) );
  INV_X1 U39204 ( .A(n38899), .ZN(n38900) );
  OAI22_X1 U39205 ( .A1(n38900), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[119][0] ), .B2(n38899), .ZN(n38892) );
  INV_X1 U39206 ( .A(n38892), .ZN(n1891) );
  OAI22_X1 U39207 ( .A1(n38900), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[119][1] ), .B2(n38899), .ZN(n38893) );
  INV_X1 U39208 ( .A(n38893), .ZN(n1890) );
  OAI22_X1 U39209 ( .A1(n38900), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[119][2] ), .B2(n38899), .ZN(n38894) );
  INV_X1 U39210 ( .A(n38894), .ZN(n1889) );
  OAI22_X1 U39211 ( .A1(n38900), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[119][3] ), .B2(n38899), .ZN(n38895) );
  INV_X1 U39212 ( .A(n38895), .ZN(n1888) );
  OAI22_X1 U39213 ( .A1(n38900), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[119][4] ), .B2(n38899), .ZN(n38896) );
  INV_X1 U39214 ( .A(n38896), .ZN(n1887) );
  OAI22_X1 U39215 ( .A1(n38900), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[119][5] ), .B2(n38899), .ZN(n38897) );
  INV_X1 U39216 ( .A(n38897), .ZN(n1886) );
  OAI22_X1 U39217 ( .A1(n38900), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[119][6] ), .B2(n38899), .ZN(n38898) );
  INV_X1 U39218 ( .A(n38898), .ZN(n1885) );
  OAI22_X1 U39219 ( .A1(n38900), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[119][7] ), .B2(n38899), .ZN(n38901) );
  INV_X1 U39220 ( .A(n38901), .ZN(n1884) );
  NOR2_X1 U39221 ( .A1(n38969), .A2(n38902), .ZN(n38910) );
  INV_X1 U39222 ( .A(n38910), .ZN(n38911) );
  OAI22_X1 U39223 ( .A1(n38911), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[120][0] ), .B2(n38910), .ZN(n38903) );
  INV_X1 U39224 ( .A(n38903), .ZN(n1883) );
  OAI22_X1 U39225 ( .A1(n38911), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[120][1] ), .B2(n38910), .ZN(n38904) );
  INV_X1 U39226 ( .A(n38904), .ZN(n1882) );
  OAI22_X1 U39227 ( .A1(n38911), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[120][2] ), .B2(n38910), .ZN(n38905) );
  INV_X1 U39228 ( .A(n38905), .ZN(n1881) );
  OAI22_X1 U39229 ( .A1(n38911), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[120][3] ), .B2(n38910), .ZN(n38906) );
  INV_X1 U39230 ( .A(n38906), .ZN(n1880) );
  OAI22_X1 U39231 ( .A1(n38911), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[120][4] ), .B2(n38910), .ZN(n38907) );
  INV_X1 U39232 ( .A(n38907), .ZN(n1879) );
  OAI22_X1 U39233 ( .A1(n38911), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[120][5] ), .B2(n38910), .ZN(n38908) );
  INV_X1 U39234 ( .A(n38908), .ZN(n1878) );
  OAI22_X1 U39235 ( .A1(n38911), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[120][6] ), .B2(n38910), .ZN(n38909) );
  INV_X1 U39236 ( .A(n38909), .ZN(n1877) );
  OAI22_X1 U39237 ( .A1(n38911), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[120][7] ), .B2(n38910), .ZN(n38912) );
  INV_X1 U39238 ( .A(n38912), .ZN(n1876) );
  NOR2_X1 U39239 ( .A1(n38969), .A2(n38913), .ZN(n38921) );
  INV_X1 U39240 ( .A(n38921), .ZN(n38922) );
  OAI22_X1 U39241 ( .A1(n38922), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[121][0] ), .B2(n38921), .ZN(n38914) );
  INV_X1 U39242 ( .A(n38914), .ZN(n1875) );
  OAI22_X1 U39243 ( .A1(n38922), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[121][1] ), .B2(n38921), .ZN(n38915) );
  INV_X1 U39244 ( .A(n38915), .ZN(n1874) );
  OAI22_X1 U39245 ( .A1(n38922), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[121][2] ), .B2(n38921), .ZN(n38916) );
  INV_X1 U39246 ( .A(n38916), .ZN(n1873) );
  OAI22_X1 U39247 ( .A1(n38922), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[121][3] ), .B2(n38921), .ZN(n38917) );
  INV_X1 U39248 ( .A(n38917), .ZN(n1872) );
  OAI22_X1 U39249 ( .A1(n38922), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[121][4] ), .B2(n38921), .ZN(n38918) );
  INV_X1 U39250 ( .A(n38918), .ZN(n1871) );
  OAI22_X1 U39251 ( .A1(n38922), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[121][5] ), .B2(n38921), .ZN(n38919) );
  INV_X1 U39252 ( .A(n38919), .ZN(n1870) );
  OAI22_X1 U39253 ( .A1(n38922), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[121][6] ), .B2(n38921), .ZN(n38920) );
  INV_X1 U39254 ( .A(n38920), .ZN(n1869) );
  OAI22_X1 U39255 ( .A1(n38922), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[121][7] ), .B2(n38921), .ZN(n38923) );
  INV_X1 U39256 ( .A(n38923), .ZN(n1868) );
  NOR2_X1 U39257 ( .A1(n38969), .A2(n38924), .ZN(n38932) );
  INV_X1 U39258 ( .A(n38932), .ZN(n38933) );
  OAI22_X1 U39259 ( .A1(n38933), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[122][0] ), .B2(n38932), .ZN(n38925) );
  INV_X1 U39260 ( .A(n38925), .ZN(n1867) );
  OAI22_X1 U39261 ( .A1(n38933), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[122][1] ), .B2(n38932), .ZN(n38926) );
  INV_X1 U39262 ( .A(n38926), .ZN(n1866) );
  OAI22_X1 U39263 ( .A1(n38933), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[122][2] ), .B2(n38932), .ZN(n38927) );
  INV_X1 U39264 ( .A(n38927), .ZN(n1865) );
  OAI22_X1 U39265 ( .A1(n38933), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[122][3] ), .B2(n38932), .ZN(n38928) );
  INV_X1 U39266 ( .A(n38928), .ZN(n1864) );
  OAI22_X1 U39267 ( .A1(n38933), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[122][4] ), .B2(n38932), .ZN(n38929) );
  INV_X1 U39268 ( .A(n38929), .ZN(n1863) );
  OAI22_X1 U39269 ( .A1(n38933), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[122][5] ), .B2(n38932), .ZN(n38930) );
  INV_X1 U39270 ( .A(n38930), .ZN(n1862) );
  OAI22_X1 U39271 ( .A1(n38933), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[122][6] ), .B2(n38932), .ZN(n38931) );
  INV_X1 U39272 ( .A(n38931), .ZN(n1861) );
  OAI22_X1 U39273 ( .A1(n38933), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[122][7] ), .B2(n38932), .ZN(n38934) );
  INV_X1 U39274 ( .A(n38934), .ZN(n1860) );
  NOR2_X1 U39275 ( .A1(n38969), .A2(n38935), .ZN(n38943) );
  INV_X1 U39276 ( .A(n38943), .ZN(n38944) );
  OAI22_X1 U39277 ( .A1(n38944), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[123][0] ), .B2(n38943), .ZN(n38936) );
  INV_X1 U39278 ( .A(n38936), .ZN(n1859) );
  OAI22_X1 U39279 ( .A1(n38944), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[123][1] ), .B2(n38943), .ZN(n38937) );
  INV_X1 U39280 ( .A(n38937), .ZN(n1858) );
  OAI22_X1 U39281 ( .A1(n38944), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[123][2] ), .B2(n38943), .ZN(n38938) );
  INV_X1 U39282 ( .A(n38938), .ZN(n1857) );
  OAI22_X1 U39283 ( .A1(n38944), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[123][3] ), .B2(n38943), .ZN(n38939) );
  INV_X1 U39284 ( .A(n38939), .ZN(n1856) );
  OAI22_X1 U39285 ( .A1(n38944), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[123][4] ), .B2(n38943), .ZN(n38940) );
  INV_X1 U39286 ( .A(n38940), .ZN(n1855) );
  OAI22_X1 U39287 ( .A1(n38944), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[123][5] ), .B2(n38943), .ZN(n38941) );
  INV_X1 U39288 ( .A(n38941), .ZN(n1854) );
  OAI22_X1 U39289 ( .A1(n38944), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[123][6] ), .B2(n38943), .ZN(n38942) );
  INV_X1 U39290 ( .A(n38942), .ZN(n1853) );
  OAI22_X1 U39291 ( .A1(n38944), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[123][7] ), .B2(n38943), .ZN(n38945) );
  INV_X1 U39292 ( .A(n38945), .ZN(n1852) );
  NOR2_X1 U39293 ( .A1(n38969), .A2(n38946), .ZN(n38954) );
  INV_X1 U39294 ( .A(n38954), .ZN(n38955) );
  OAI22_X1 U39295 ( .A1(n38955), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[124][0] ), .B2(n38954), .ZN(n38947) );
  INV_X1 U39296 ( .A(n38947), .ZN(n1851) );
  OAI22_X1 U39297 ( .A1(n38955), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[124][1] ), .B2(n38954), .ZN(n38948) );
  INV_X1 U39298 ( .A(n38948), .ZN(n1850) );
  OAI22_X1 U39299 ( .A1(n38955), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[124][2] ), .B2(n38954), .ZN(n38949) );
  INV_X1 U39300 ( .A(n38949), .ZN(n1849) );
  OAI22_X1 U39301 ( .A1(n38955), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[124][3] ), .B2(n38954), .ZN(n38950) );
  INV_X1 U39302 ( .A(n38950), .ZN(n1848) );
  OAI22_X1 U39303 ( .A1(n38955), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[124][4] ), .B2(n38954), .ZN(n38951) );
  INV_X1 U39304 ( .A(n38951), .ZN(n1847) );
  OAI22_X1 U39305 ( .A1(n38955), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[124][5] ), .B2(n38954), .ZN(n38952) );
  INV_X1 U39306 ( .A(n38952), .ZN(n1846) );
  OAI22_X1 U39307 ( .A1(n38955), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[124][6] ), .B2(n38954), .ZN(n38953) );
  INV_X1 U39308 ( .A(n38953), .ZN(n1845) );
  OAI22_X1 U39309 ( .A1(n38955), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[124][7] ), .B2(n38954), .ZN(n38956) );
  INV_X1 U39310 ( .A(n38956), .ZN(n1844) );
  NOR2_X1 U39311 ( .A1(n38969), .A2(n38957), .ZN(n38965) );
  INV_X1 U39312 ( .A(n38965), .ZN(n38966) );
  OAI22_X1 U39313 ( .A1(n38966), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[125][0] ), .B2(n38965), .ZN(n38958) );
  INV_X1 U39314 ( .A(n38958), .ZN(n1843) );
  OAI22_X1 U39315 ( .A1(n38966), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[125][1] ), .B2(n38965), .ZN(n38959) );
  INV_X1 U39316 ( .A(n38959), .ZN(n1842) );
  OAI22_X1 U39317 ( .A1(n38966), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[125][2] ), .B2(n38965), .ZN(n38960) );
  INV_X1 U39318 ( .A(n38960), .ZN(n1841) );
  OAI22_X1 U39319 ( .A1(n38966), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[125][3] ), .B2(n38965), .ZN(n38961) );
  INV_X1 U39320 ( .A(n38961), .ZN(n1840) );
  OAI22_X1 U39321 ( .A1(n38966), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[125][4] ), .B2(n38965), .ZN(n38962) );
  INV_X1 U39322 ( .A(n38962), .ZN(n1839) );
  OAI22_X1 U39323 ( .A1(n38966), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[125][5] ), .B2(n38965), .ZN(n38963) );
  INV_X1 U39324 ( .A(n38963), .ZN(n1838) );
  OAI22_X1 U39325 ( .A1(n38966), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[125][6] ), .B2(n38965), .ZN(n38964) );
  INV_X1 U39326 ( .A(n38964), .ZN(n1837) );
  OAI22_X1 U39327 ( .A1(n38966), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[125][7] ), .B2(n38965), .ZN(n38967) );
  INV_X1 U39328 ( .A(n38967), .ZN(n1836) );
  NOR2_X1 U39329 ( .A1(n38969), .A2(n38968), .ZN(n38977) );
  INV_X1 U39330 ( .A(n38977), .ZN(n38978) );
  OAI22_X1 U39331 ( .A1(n38978), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[126][0] ), .B2(n38977), .ZN(n38970) );
  INV_X1 U39332 ( .A(n38970), .ZN(n1835) );
  OAI22_X1 U39333 ( .A1(n38978), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[126][1] ), .B2(n38977), .ZN(n38971) );
  INV_X1 U39334 ( .A(n38971), .ZN(n1834) );
  OAI22_X1 U39335 ( .A1(n38978), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[126][2] ), .B2(n38977), .ZN(n38972) );
  INV_X1 U39336 ( .A(n38972), .ZN(n1833) );
  OAI22_X1 U39337 ( .A1(n38978), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[126][3] ), .B2(n38977), .ZN(n38973) );
  INV_X1 U39338 ( .A(n38973), .ZN(n1832) );
  OAI22_X1 U39339 ( .A1(n38978), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[126][4] ), .B2(n38977), .ZN(n38974) );
  INV_X1 U39340 ( .A(n38974), .ZN(n1831) );
  OAI22_X1 U39341 ( .A1(n38978), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[126][5] ), .B2(n38977), .ZN(n38975) );
  INV_X1 U39342 ( .A(n38975), .ZN(n1830) );
  OAI22_X1 U39343 ( .A1(n38978), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[126][6] ), .B2(n38977), .ZN(n38976) );
  INV_X1 U39344 ( .A(n38976), .ZN(n1829) );
  OAI22_X1 U39345 ( .A1(n38978), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[126][7] ), .B2(n38977), .ZN(n38979) );
  INV_X1 U39346 ( .A(n38979), .ZN(n1828) );
  INV_X1 U39347 ( .A(n38987), .ZN(n38988) );
  OAI22_X1 U39348 ( .A1(n38988), .A2(s_data_in_x[0]), .B1(
        \xmem_inst/mem[127][0] ), .B2(n38987), .ZN(n38980) );
  INV_X1 U39349 ( .A(n38980), .ZN(n1827) );
  OAI22_X1 U39350 ( .A1(n38988), .A2(s_data_in_x[1]), .B1(
        \xmem_inst/mem[127][1] ), .B2(n38987), .ZN(n38981) );
  INV_X1 U39351 ( .A(n38981), .ZN(n1826) );
  OAI22_X1 U39352 ( .A1(n38988), .A2(s_data_in_x[2]), .B1(
        \xmem_inst/mem[127][2] ), .B2(n38987), .ZN(n38982) );
  INV_X1 U39353 ( .A(n38982), .ZN(n1825) );
  OAI22_X1 U39354 ( .A1(n38988), .A2(s_data_in_x[3]), .B1(
        \xmem_inst/mem[127][3] ), .B2(n38987), .ZN(n38983) );
  INV_X1 U39355 ( .A(n38983), .ZN(n1824) );
  OAI22_X1 U39356 ( .A1(n38988), .A2(s_data_in_x[4]), .B1(
        \xmem_inst/mem[127][4] ), .B2(n38987), .ZN(n38984) );
  INV_X1 U39357 ( .A(n38984), .ZN(n1823) );
  OAI22_X1 U39358 ( .A1(n38988), .A2(s_data_in_x[5]), .B1(
        \xmem_inst/mem[127][5] ), .B2(n38987), .ZN(n38985) );
  INV_X1 U39359 ( .A(n38985), .ZN(n1822) );
  OAI22_X1 U39360 ( .A1(n38988), .A2(s_data_in_x[6]), .B1(
        \xmem_inst/mem[127][6] ), .B2(n38987), .ZN(n38986) );
  INV_X1 U39361 ( .A(n38986), .ZN(n1821) );
  OAI22_X1 U39362 ( .A1(n38988), .A2(s_data_in_x[7]), .B1(
        \xmem_inst/mem[127][7] ), .B2(n38987), .ZN(n38989) );
  INV_X1 U39363 ( .A(n38989), .ZN(n1820) );
  AOI22_X1 U39364 ( .A1(n6173), .A2(n38995), .B1(n38994), .B2(n3248), .ZN(
        n1819) );
  OAI22_X1 U39365 ( .A1(n8416), .A2(n38995), .B1(n38994), .B2(n38990), .ZN(
        n1817) );
  OAI22_X1 U39366 ( .A1(n8418), .A2(n38995), .B1(n38994), .B2(n3230), .ZN(
        n1816) );
  OAI22_X1 U39367 ( .A1(n8414), .A2(n38995), .B1(n38994), .B2(n38991), .ZN(
        n1815) );
  INV_X1 U39368 ( .A(n38992), .ZN(n38993) );
  OAI22_X1 U39369 ( .A1(n39041), .A2(n38995), .B1(n38994), .B2(n38993), .ZN(
        n1814) );
endmodule

