
module conv_128_32_opt_DW_mult_pipe_J1_0 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n361, n363, n365, n367, n369, n371, n373, n375, n377, n379,
         n381, n383, n385, n387, n389, n391, n393, n395, n397, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n412,
         n414, n416, n418, n420, n422, n424, n426, n428, n430, n432, n434,
         n436, n438, n440, n442, n444, n446, n448, n450, n452, n454, n456,
         n458, n460, n462, n464, n466, n468, n470, n472, n474, n476, n478,
         n480, n482, n484, n486, n488, n490, n492, n494, n496, n498, n500,
         n502, n504, n506, n508, n510, n512, n514, n516, n518, n520, n522,
         n523, n525, n526, n528, n529, n531, n532, n534, n535, n537, n538,
         n540, n542, n544, n546, n548, n550, n552, n554, n556, n558, n559,
         n560, n561;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n410), .SE(n520), .CK(clk), .Q(n560), 
        .QN(n22) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n410), .SE(n516), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n35) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n410), .SE(n514), .CK(clk), .Q(n559), 
        .QN(n27) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n410), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n338) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n410), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n34) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n410), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n23) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n410), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n410), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n31) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n410), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n32) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n410), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n33) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n28) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n410), .SE(n486), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n410), .SE(n484), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n410), .SE(n482), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(rst_n), .SE(n480), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n410), .SE(n478), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n410), .SE(n476), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n410), .SE(n474), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n410), .SE(n472), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(rst_n), .SE(n470), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n468), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n410), .SE(n466), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n410), .SE(n464), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(rst_n), .SE(n462), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n410), .SE(n460), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n410), .SE(n458), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n410), .SE(n456), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n410), .SE(n454), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n410), .SE(n450), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n410), .SE(n448), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n410), .SE(n446), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n410), .SE(n442), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n440), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n410), .SE(n438), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n410), .SE(n434), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n430), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n428), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n426), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n420), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n418), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n416), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n414), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n412), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n410), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n36) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n561), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n561), .SE(n395), .CK(
        clk), .Q(n403), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n561), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n561), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n355), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n561), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n354), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n561), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n561), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n352), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n561), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n351), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n561), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n350), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n561), .SE(n379), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n561), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n348), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n561), .SE(n375), .CK(
        clk), .Q(n408), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n561), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n346), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n561), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n345), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n561), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n344), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n561), .SE(n367), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n561), .SE(n365), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n561), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n561), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n561), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n339) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n410), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n337) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n410), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n26) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n410), .SE(n518), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n25) );
  MUX2_X1 U2 ( .A(n342), .B(n172), .S(n264), .Z(n365) );
  MUX2_X2 U3 ( .A(n340), .B(n128), .S(n264), .Z(n361) );
  BUF_X1 U4 ( .A(n168), .Z(n18) );
  BUF_X2 U5 ( .A(n91), .Z(n8) );
  BUF_X1 U6 ( .A(en), .Z(n296) );
  BUF_X1 U7 ( .A(n296), .Z(n264) );
  CLKBUF_X2 U8 ( .A(rst_n), .Z(n410) );
  CLKBUF_X1 U9 ( .A(n168), .Z(n16) );
  BUF_X1 U10 ( .A(\mult_x_1/n313 ), .Z(n91) );
  INV_X1 U11 ( .A(n25), .ZN(n19) );
  INV_X1 U12 ( .A(n9), .ZN(n178) );
  NAND2_X1 U13 ( .A1(n41), .A2(n42), .ZN(n157) );
  INV_X1 U14 ( .A(n166), .ZN(n6) );
  XOR2_X1 U15 ( .A(n337), .B(n338), .Z(n7) );
  OAI21_X1 U16 ( .B1(n114), .B2(n113), .A(n112), .ZN(n104) );
  XNOR2_X1 U17 ( .A(n77), .B(n206), .ZN(n223) );
  XNOR2_X1 U18 ( .A(n223), .B(n86), .ZN(n267) );
  XNOR2_X1 U19 ( .A(n225), .B(n224), .ZN(n86) );
  BUF_X1 U20 ( .A(n177), .Z(n11) );
  OR2_X1 U21 ( .A1(n133), .A2(n132), .ZN(n125) );
  NAND2_X1 U22 ( .A1(n133), .A2(n132), .ZN(n126) );
  XNOR2_X1 U23 ( .A(n133), .B(n132), .ZN(n134) );
  INV_X1 U24 ( .A(n250), .ZN(n246) );
  INV_X1 U25 ( .A(n249), .ZN(n245) );
  INV_X1 U26 ( .A(n224), .ZN(n220) );
  INV_X1 U27 ( .A(n225), .ZN(n221) );
  XNOR2_X1 U28 ( .A(n248), .B(n43), .ZN(n47) );
  XNOR2_X1 U29 ( .A(n250), .B(n249), .ZN(n43) );
  BUF_X2 U30 ( .A(\mult_x_1/n312 ), .Z(n20) );
  NAND2_X1 U31 ( .A1(n104), .A2(n103), .ZN(n111) );
  NAND2_X1 U32 ( .A1(n114), .A2(n113), .ZN(n103) );
  NAND2_X1 U33 ( .A1(n212), .A2(n211), .ZN(n214) );
  NAND2_X1 U34 ( .A1(n24), .A2(n217), .ZN(n211) );
  NAND2_X1 U35 ( .A1(n218), .A2(n210), .ZN(n212) );
  OR2_X1 U36 ( .A1(n24), .A2(n217), .ZN(n210) );
  NAND2_X1 U37 ( .A1(n252), .A2(n251), .ZN(n254) );
  NAND2_X1 U38 ( .A1(n250), .A2(n249), .ZN(n251) );
  NAND2_X1 U39 ( .A1(n248), .A2(n247), .ZN(n252) );
  NAND2_X1 U40 ( .A1(n246), .A2(n245), .ZN(n247) );
  NAND2_X1 U41 ( .A1(n227), .A2(n226), .ZN(n257) );
  NAND2_X1 U42 ( .A1(n225), .A2(n224), .ZN(n226) );
  NAND2_X1 U43 ( .A1(n223), .A2(n222), .ZN(n227) );
  NAND2_X1 U44 ( .A1(n221), .A2(n220), .ZN(n222) );
  INV_X1 U45 ( .A(n266), .ZN(n97) );
  MUX2_X1 U46 ( .A(n216), .B(n348), .S(n71), .Z(n377) );
  OAI22_X1 U47 ( .A1(n267), .A2(n98), .B1(n336), .B2(n407), .ZN(n381) );
  NAND2_X1 U48 ( .A1(n336), .A2(n97), .ZN(n98) );
  XOR2_X1 U49 ( .A(n559), .B(\mult_x_1/a[6] ), .Z(n9) );
  CLKBUF_X1 U50 ( .A(n177), .Z(n10) );
  CLKBUF_X1 U51 ( .A(n177), .Z(n12) );
  CLKBUF_X1 U52 ( .A(\mult_x_1/n281 ), .Z(n14) );
  NAND2_X1 U53 ( .A1(n74), .A2(n75), .ZN(n177) );
  XNOR2_X1 U54 ( .A(n117), .B(n91), .ZN(n13) );
  BUF_X4 U55 ( .A(n296), .Z(n15) );
  BUF_X2 U56 ( .A(n168), .Z(n17) );
  OR2_X1 U57 ( .A1(n36), .A2(\mult_x_1/n180 ), .ZN(n152) );
  OAI22_X1 U58 ( .A1(n157), .A2(n118), .B1(n119), .B2(n155), .ZN(n21) );
  AND2_X1 U59 ( .A1(n206), .A2(n205), .ZN(n24) );
  INV_X1 U60 ( .A(rst_n), .ZN(n561) );
  XOR2_X1 U61 ( .A(\mult_x_1/a[4] ), .B(n559), .Z(n37) );
  XNOR2_X1 U62 ( .A(n337), .B(n338), .ZN(n38) );
  NAND2_X1 U63 ( .A1(n37), .A2(n38), .ZN(n168) );
  BUF_X2 U64 ( .A(n559), .Z(n335) );
  OR2_X1 U65 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n39) );
  OAI22_X1 U66 ( .A1(n17), .A2(n27), .B1(n39), .B2(n166), .ZN(n164) );
  XNOR2_X1 U67 ( .A(n335), .B(\mult_x_1/n288 ), .ZN(n40) );
  INV_X2 U68 ( .A(n7), .ZN(n166) );
  XNOR2_X1 U69 ( .A(n335), .B(\mult_x_1/n287 ), .ZN(n167) );
  OAI22_X1 U70 ( .A1(n18), .A2(n40), .B1(n166), .B2(n167), .ZN(n163) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n312 ), .B(n34), .ZN(n41) );
  XNOR2_X1 U72 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n42) );
  XNOR2_X1 U73 ( .A(n20), .B(\mult_x_1/n286 ), .ZN(n45) );
  INV_X1 U74 ( .A(n42), .ZN(n58) );
  INV_X2 U75 ( .A(n58), .ZN(n155) );
  XNOR2_X1 U76 ( .A(n20), .B(\mult_x_1/n285 ), .ZN(n156) );
  OAI22_X1 U77 ( .A1(n157), .A2(n45), .B1(n155), .B2(n156), .ZN(n250) );
  XNOR2_X1 U78 ( .A(n91), .B(\mult_x_1/n284 ), .ZN(n44) );
  XNOR2_X1 U79 ( .A(n91), .B(\mult_x_1/n283 ), .ZN(n151) );
  OAI22_X1 U80 ( .A1(n152), .A2(n44), .B1(n151), .B2(n23), .ZN(n249) );
  XNOR2_X1 U81 ( .A(n8), .B(\mult_x_1/n285 ), .ZN(n53) );
  OAI22_X1 U82 ( .A1(n152), .A2(n53), .B1(n44), .B2(n23), .ZN(n50) );
  AND2_X1 U83 ( .A1(\mult_x_1/n288 ), .A2(n6), .ZN(n49) );
  XNOR2_X1 U84 ( .A(n20), .B(\mult_x_1/n287 ), .ZN(n51) );
  OAI22_X1 U85 ( .A1(n157), .A2(n51), .B1(n155), .B2(n45), .ZN(n48) );
  OR2_X1 U86 ( .A1(n47), .A2(n46), .ZN(n263) );
  NAND2_X1 U87 ( .A1(n47), .A2(n46), .ZN(n260) );
  NAND2_X1 U88 ( .A1(n263), .A2(n260), .ZN(n69) );
  FA_X1 U89 ( .A(n50), .B(n49), .CI(n48), .CO(n46), .S(n67) );
  XNOR2_X1 U90 ( .A(n20), .B(\mult_x_1/n288 ), .ZN(n52) );
  OAI22_X1 U91 ( .A1(n157), .A2(n52), .B1(n155), .B2(n51), .ZN(n55) );
  XNOR2_X1 U92 ( .A(n8), .B(\mult_x_1/n286 ), .ZN(n57) );
  OAI22_X1 U93 ( .A1(n152), .A2(n57), .B1(n53), .B2(n23), .ZN(n54) );
  NOR2_X1 U94 ( .A1(n67), .A2(n66), .ZN(n287) );
  HA_X1 U95 ( .A(n55), .B(n54), .CO(n66), .S(n64) );
  OR2_X1 U96 ( .A1(\mult_x_1/n288 ), .A2(n337), .ZN(n56) );
  OAI22_X1 U97 ( .A1(n157), .A2(n337), .B1(n56), .B2(n155), .ZN(n63) );
  OR2_X1 U98 ( .A1(n64), .A2(n63), .ZN(n283) );
  XNOR2_X1 U99 ( .A(n8), .B(\mult_x_1/n287 ), .ZN(n59) );
  OAI22_X1 U100 ( .A1(n152), .A2(n59), .B1(n57), .B2(n23), .ZN(n62) );
  AND2_X1 U101 ( .A1(\mult_x_1/n288 ), .A2(n58), .ZN(n61) );
  NOR2_X1 U102 ( .A1(n62), .A2(n61), .ZN(n276) );
  OAI22_X1 U103 ( .A1(n152), .A2(\mult_x_1/n288 ), .B1(n59), .B2(n23), .ZN(
        n273) );
  OR2_X1 U104 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n60) );
  NAND2_X1 U105 ( .A1(n60), .A2(n152), .ZN(n272) );
  NAND2_X1 U106 ( .A1(n273), .A2(n272), .ZN(n279) );
  NAND2_X1 U107 ( .A1(n62), .A2(n61), .ZN(n277) );
  OAI21_X1 U108 ( .B1(n276), .B2(n279), .A(n277), .ZN(n284) );
  NAND2_X1 U109 ( .A1(n64), .A2(n63), .ZN(n282) );
  INV_X1 U110 ( .A(n282), .ZN(n65) );
  AOI21_X1 U111 ( .B1(n283), .B2(n284), .A(n65), .ZN(n290) );
  NAND2_X1 U112 ( .A1(n67), .A2(n66), .ZN(n288) );
  OAI21_X1 U113 ( .B1(n287), .B2(n290), .A(n288), .ZN(n262) );
  INV_X1 U114 ( .A(n262), .ZN(n68) );
  XNOR2_X1 U115 ( .A(n69), .B(n68), .ZN(n72) );
  INV_X1 U116 ( .A(n15), .ZN(n71) );
  NAND2_X1 U117 ( .A1(n71), .A2(n538), .ZN(n70) );
  OAI21_X1 U118 ( .B1(n72), .B2(n71), .A(n70), .ZN(n446) );
  XNOR2_X1 U119 ( .A(n335), .B(\mult_x_1/n284 ), .ZN(n137) );
  XNOR2_X1 U120 ( .A(n335), .B(\mult_x_1/n283 ), .ZN(n136) );
  OAI22_X1 U121 ( .A1(n18), .A2(n137), .B1(n166), .B2(n136), .ZN(n73) );
  XNOR2_X1 U122 ( .A(n20), .B(\mult_x_1/n282 ), .ZN(n78) );
  XNOR2_X1 U123 ( .A(n20), .B(\mult_x_1/n281 ), .ZN(n118) );
  OAI22_X1 U124 ( .A1(n157), .A2(n78), .B1(n155), .B2(n118), .ZN(n138) );
  XNOR2_X1 U125 ( .A(n73), .B(n138), .ZN(n205) );
  INV_X1 U126 ( .A(n205), .ZN(n77) );
  XNOR2_X1 U127 ( .A(\mult_x_1/n310 ), .B(n35), .ZN(n74) );
  XNOR2_X1 U128 ( .A(n559), .B(\mult_x_1/a[6] ), .ZN(n75) );
  XNOR2_X1 U129 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n80) );
  XNOR2_X1 U130 ( .A(n19), .B(\mult_x_1/n286 ), .ZN(n85) );
  OAI22_X1 U131 ( .A1(n12), .A2(n80), .B1(n178), .B2(n85), .ZN(n89) );
  XNOR2_X1 U132 ( .A(n8), .B(n14), .ZN(n92) );
  AND2_X2 U133 ( .A1(n560), .A2(\mult_x_1/n281 ), .ZN(n117) );
  XNOR2_X1 U134 ( .A(n117), .B(n91), .ZN(n82) );
  OAI22_X1 U135 ( .A1(n152), .A2(n92), .B1(n82), .B2(n23), .ZN(n88) );
  NAND2_X1 U136 ( .A1(n22), .A2(\mult_x_1/n310 ), .ZN(n84) );
  INV_X1 U137 ( .A(n84), .ZN(n76) );
  AND2_X1 U138 ( .A1(\mult_x_1/n288 ), .A2(n76), .ZN(n87) );
  XNOR2_X1 U139 ( .A(n335), .B(\mult_x_1/n285 ), .ZN(n90) );
  OAI22_X1 U140 ( .A1(n17), .A2(n90), .B1(n166), .B2(n137), .ZN(n96) );
  XNOR2_X1 U141 ( .A(n20), .B(\mult_x_1/n283 ), .ZN(n93) );
  OAI22_X1 U142 ( .A1(n157), .A2(n93), .B1(n155), .B2(n78), .ZN(n95) );
  OR2_X1 U143 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n79) );
  OAI22_X1 U144 ( .A1(n11), .A2(n25), .B1(n79), .B2(n178), .ZN(n159) );
  XNOR2_X1 U145 ( .A(n19), .B(\mult_x_1/n288 ), .ZN(n81) );
  OAI22_X1 U146 ( .A1(n10), .A2(n81), .B1(n178), .B2(n80), .ZN(n158) );
  AOI21_X1 U147 ( .B1(n152), .B2(n23), .A(n13), .ZN(n83) );
  INV_X1 U148 ( .A(n83), .ZN(n142) );
  NOR2_X1 U149 ( .A1(n28), .A2(n84), .ZN(n141) );
  XNOR2_X1 U150 ( .A(n19), .B(\mult_x_1/n285 ), .ZN(n122) );
  OAI22_X1 U151 ( .A1(n12), .A2(n85), .B1(n178), .B2(n122), .ZN(n140) );
  FA_X1 U152 ( .A(n89), .B(n88), .CI(n87), .CO(n206), .S(n231) );
  XNOR2_X1 U153 ( .A(n335), .B(\mult_x_1/n286 ), .ZN(n165) );
  OAI22_X1 U154 ( .A1(n18), .A2(n165), .B1(n166), .B2(n90), .ZN(n162) );
  XNOR2_X1 U155 ( .A(n8), .B(\mult_x_1/n282 ), .ZN(n150) );
  OAI22_X1 U156 ( .A1(n152), .A2(n150), .B1(n92), .B2(n23), .ZN(n161) );
  XNOR2_X1 U157 ( .A(n20), .B(\mult_x_1/n284 ), .ZN(n154) );
  OAI22_X1 U158 ( .A1(n157), .A2(n154), .B1(n155), .B2(n93), .ZN(n160) );
  FA_X1 U159 ( .A(n96), .B(n95), .CI(n94), .CO(n225), .S(n229) );
  NOR2_X1 U180 ( .A1(n29), .A2(n84), .ZN(n175) );
  XNOR2_X1 U181 ( .A(n19), .B(n14), .ZN(n99) );
  XNOR2_X1 U182 ( .A(n117), .B(n19), .ZN(n176) );
  OAI22_X1 U183 ( .A1(n12), .A2(n99), .B1(n176), .B2(n178), .ZN(n183) );
  INV_X1 U184 ( .A(n183), .ZN(n174) );
  XNOR2_X1 U185 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n102) );
  OAI22_X1 U186 ( .A1(n12), .A2(n102), .B1(n178), .B2(n99), .ZN(n107) );
  XNOR2_X1 U187 ( .A(n117), .B(n335), .ZN(n101) );
  AOI21_X1 U188 ( .B1(n166), .B2(n16), .A(n101), .ZN(n100) );
  INV_X1 U189 ( .A(n100), .ZN(n106) );
  XNOR2_X1 U190 ( .A(n335), .B(n14), .ZN(n123) );
  OAI22_X1 U191 ( .A1(n18), .A2(n123), .B1(n101), .B2(n166), .ZN(n105) );
  INV_X1 U192 ( .A(n105), .ZN(n114) );
  XNOR2_X1 U193 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n116) );
  OAI22_X1 U194 ( .A1(n10), .A2(n116), .B1(n178), .B2(n102), .ZN(n113) );
  NOR2_X1 U195 ( .A1(n30), .A2(n84), .ZN(n112) );
  NOR2_X1 U196 ( .A1(n31), .A2(n84), .ZN(n110) );
  FA_X1 U197 ( .A(n107), .B(n106), .CI(n105), .CO(n173), .S(n109) );
  OR2_X1 U198 ( .A1(n190), .A2(n189), .ZN(n108) );
  MUX2_X1 U199 ( .A(n339), .B(n108), .S(n336), .Z(n359) );
  FA_X1 U200 ( .A(n111), .B(n110), .CI(n109), .CO(n189), .S(n193) );
  XNOR2_X1 U201 ( .A(n113), .B(n112), .ZN(n115) );
  XNOR2_X1 U202 ( .A(n115), .B(n114), .ZN(n131) );
  XNOR2_X1 U203 ( .A(n19), .B(\mult_x_1/n284 ), .ZN(n121) );
  OAI22_X1 U204 ( .A1(n11), .A2(n121), .B1(n178), .B2(n116), .ZN(n145) );
  XNOR2_X1 U205 ( .A(n117), .B(n20), .ZN(n119) );
  OAI22_X1 U206 ( .A1(n157), .A2(n118), .B1(n119), .B2(n155), .ZN(n144) );
  AOI21_X1 U207 ( .B1(n155), .B2(n157), .A(n119), .ZN(n120) );
  INV_X1 U208 ( .A(n120), .ZN(n143) );
  OAI22_X1 U209 ( .A1(n11), .A2(n122), .B1(n178), .B2(n121), .ZN(n209) );
  XNOR2_X1 U210 ( .A(n335), .B(\mult_x_1/n282 ), .ZN(n124) );
  OAI22_X1 U211 ( .A1(n17), .A2(n136), .B1(n166), .B2(n124), .ZN(n208) );
  INV_X1 U212 ( .A(n144), .ZN(n207) );
  OAI22_X1 U213 ( .A1(n17), .A2(n124), .B1(n166), .B2(n123), .ZN(n133) );
  NOR2_X1 U214 ( .A1(n32), .A2(n84), .ZN(n132) );
  NAND2_X1 U215 ( .A1(n135), .A2(n125), .ZN(n127) );
  NAND2_X1 U216 ( .A1(n127), .A2(n126), .ZN(n129) );
  OR2_X1 U217 ( .A1(n193), .A2(n192), .ZN(n128) );
  FA_X1 U218 ( .A(n131), .B(n130), .CI(n129), .CO(n192), .S(n196) );
  XNOR2_X1 U219 ( .A(n135), .B(n134), .ZN(n201) );
  OAI22_X1 U220 ( .A1(n18), .A2(n137), .B1(n166), .B2(n136), .ZN(n139) );
  OR2_X1 U221 ( .A1(n139), .A2(n138), .ZN(n204) );
  NOR2_X1 U222 ( .A1(n33), .A2(n84), .ZN(n203) );
  FA_X1 U223 ( .A(n142), .B(n141), .CI(n140), .CO(n202), .S(n224) );
  NAND2_X1 U224 ( .A1(n201), .A2(n199), .ZN(n148) );
  FA_X1 U225 ( .A(n145), .B(n21), .CI(n143), .CO(n130), .S(n198) );
  NAND2_X1 U226 ( .A1(n201), .A2(n198), .ZN(n147) );
  NAND2_X1 U227 ( .A1(n199), .A2(n198), .ZN(n146) );
  NAND3_X1 U228 ( .A1(n148), .A2(n147), .A3(n146), .ZN(n195) );
  OR2_X1 U229 ( .A1(n196), .A2(n195), .ZN(n149) );
  MUX2_X1 U230 ( .A(n341), .B(n149), .S(n336), .Z(n363) );
  OAI22_X1 U231 ( .A1(n152), .A2(n151), .B1(n150), .B2(n23), .ZN(n171) );
  INV_X1 U232 ( .A(n178), .ZN(n153) );
  AND2_X1 U233 ( .A1(\mult_x_1/n288 ), .A2(n153), .ZN(n170) );
  OAI22_X1 U234 ( .A1(n157), .A2(n156), .B1(n155), .B2(n154), .ZN(n169) );
  HA_X1 U235 ( .A(n159), .B(n158), .CO(n94), .S(n233) );
  FA_X1 U236 ( .A(n162), .B(n160), .CI(n161), .CO(n230), .S(n232) );
  HA_X1 U237 ( .A(n164), .B(n163), .CO(n244), .S(n248) );
  OAI22_X1 U238 ( .A1(n17), .A2(n167), .B1(n166), .B2(n165), .ZN(n243) );
  FA_X1 U239 ( .A(n171), .B(n170), .CI(n169), .CO(n234), .S(n242) );
  OR2_X1 U240 ( .A1(n240), .A2(n239), .ZN(n172) );
  FA_X1 U241 ( .A(n175), .B(n174), .CI(n173), .CO(n185), .S(n190) );
  AOI21_X1 U242 ( .B1(n178), .B2(n11), .A(n176), .ZN(n179) );
  INV_X1 U243 ( .A(n179), .ZN(n181) );
  NOR2_X1 U244 ( .A1(n26), .A2(n84), .ZN(n180) );
  XOR2_X1 U245 ( .A(n181), .B(n180), .Z(n182) );
  XOR2_X1 U246 ( .A(n183), .B(n182), .Z(n184) );
  OR2_X1 U247 ( .A1(n185), .A2(n184), .ZN(n187) );
  NAND2_X1 U248 ( .A1(n185), .A2(n184), .ZN(n186) );
  NAND2_X1 U249 ( .A1(n187), .A2(n186), .ZN(n188) );
  MUX2_X1 U250 ( .A(n343), .B(n188), .S(n336), .Z(n367) );
  NAND2_X1 U251 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U252 ( .A(n344), .B(n191), .S(n264), .Z(n369) );
  NAND2_X1 U253 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U254 ( .A(n345), .B(n194), .S(n264), .Z(n371) );
  NAND2_X1 U255 ( .A1(n196), .A2(n195), .ZN(n197) );
  MUX2_X1 U256 ( .A(n346), .B(n197), .S(n336), .Z(n373) );
  XNOR2_X1 U257 ( .A(n199), .B(n198), .ZN(n200) );
  XNOR2_X1 U258 ( .A(n200), .B(n201), .ZN(n215) );
  FA_X1 U259 ( .A(n204), .B(n203), .CI(n202), .CO(n199), .S(n218) );
  FA_X1 U260 ( .A(n208), .B(n209), .CI(n207), .CO(n135), .S(n217) );
  NOR2_X1 U261 ( .A1(n214), .A2(n215), .ZN(n213) );
  MUX2_X1 U262 ( .A(n347), .B(n213), .S(n264), .Z(n375) );
  NAND2_X1 U263 ( .A1(n215), .A2(n214), .ZN(n216) );
  XNOR2_X1 U264 ( .A(n24), .B(n217), .ZN(n219) );
  XNOR2_X1 U265 ( .A(n219), .B(n218), .ZN(n258) );
  NAND2_X1 U266 ( .A1(n258), .A2(n257), .ZN(n228) );
  MUX2_X1 U267 ( .A(n349), .B(n228), .S(n264), .Z(n379) );
  FA_X1 U268 ( .A(n231), .B(n230), .CI(n229), .CO(n266), .S(n237) );
  FA_X1 U269 ( .A(n234), .B(n233), .CI(n232), .CO(n236), .S(n240) );
  NOR2_X1 U270 ( .A1(n237), .A2(n236), .ZN(n235) );
  MUX2_X1 U271 ( .A(n352), .B(n235), .S(n264), .Z(n385) );
  NAND2_X1 U272 ( .A1(n237), .A2(n236), .ZN(n238) );
  MUX2_X1 U273 ( .A(n353), .B(n238), .S(n336), .Z(n387) );
  NAND2_X1 U274 ( .A1(n240), .A2(n239), .ZN(n241) );
  MUX2_X1 U275 ( .A(n354), .B(n241), .S(n264), .Z(n389) );
  FA_X1 U276 ( .A(n244), .B(n243), .CI(n242), .CO(n239), .S(n255) );
  NOR2_X1 U277 ( .A1(n255), .A2(n254), .ZN(n253) );
  MUX2_X1 U278 ( .A(n355), .B(n253), .S(n336), .Z(n391) );
  NAND2_X1 U279 ( .A1(n255), .A2(n254), .ZN(n256) );
  MUX2_X1 U280 ( .A(n356), .B(n256), .S(n264), .Z(n393) );
  NOR2_X1 U281 ( .A1(n258), .A2(n257), .ZN(n259) );
  MUX2_X1 U282 ( .A(n357), .B(n259), .S(n336), .Z(n395) );
  INV_X1 U283 ( .A(n260), .ZN(n261) );
  AOI21_X1 U284 ( .B1(n263), .B2(n262), .A(n261), .ZN(n265) );
  MUX2_X1 U285 ( .A(n358), .B(n265), .S(n264), .Z(n397) );
  NAND2_X1 U286 ( .A1(n267), .A2(n266), .ZN(n268) );
  NAND2_X1 U287 ( .A1(n268), .A2(n336), .ZN(n270) );
  OR2_X1 U288 ( .A1(n336), .A2(n402), .ZN(n269) );
  NAND2_X1 U289 ( .A1(n270), .A2(n269), .ZN(n383) );
  MUX2_X1 U290 ( .A(product[0]), .B(n522), .S(n15), .Z(n412) );
  MUX2_X1 U291 ( .A(n522), .B(n523), .S(n15), .Z(n414) );
  AND2_X1 U292 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n271) );
  MUX2_X1 U293 ( .A(n523), .B(n271), .S(n15), .Z(n416) );
  MUX2_X1 U294 ( .A(product[1]), .B(n525), .S(n15), .Z(n418) );
  MUX2_X1 U295 ( .A(n525), .B(n526), .S(n15), .Z(n420) );
  OR2_X1 U296 ( .A1(n273), .A2(n272), .ZN(n274) );
  AND2_X1 U297 ( .A1(n274), .A2(n279), .ZN(n275) );
  MUX2_X1 U298 ( .A(n526), .B(n275), .S(n15), .Z(n422) );
  MUX2_X1 U299 ( .A(product[2]), .B(n528), .S(n15), .Z(n424) );
  MUX2_X1 U300 ( .A(n528), .B(n529), .S(n15), .Z(n426) );
  INV_X1 U301 ( .A(n276), .ZN(n278) );
  NAND2_X1 U302 ( .A1(n278), .A2(n277), .ZN(n280) );
  XOR2_X1 U303 ( .A(n280), .B(n279), .Z(n281) );
  MUX2_X1 U304 ( .A(n529), .B(n281), .S(n15), .Z(n428) );
  MUX2_X1 U305 ( .A(product[3]), .B(n531), .S(n15), .Z(n430) );
  MUX2_X1 U306 ( .A(n531), .B(n532), .S(n15), .Z(n432) );
  NAND2_X1 U307 ( .A1(n283), .A2(n282), .ZN(n285) );
  XNOR2_X1 U308 ( .A(n285), .B(n284), .ZN(n286) );
  MUX2_X1 U309 ( .A(n532), .B(n286), .S(n15), .Z(n434) );
  MUX2_X1 U310 ( .A(product[4]), .B(n534), .S(n15), .Z(n436) );
  MUX2_X1 U311 ( .A(n534), .B(n535), .S(n15), .Z(n438) );
  INV_X1 U312 ( .A(n287), .ZN(n289) );
  NAND2_X1 U313 ( .A1(n289), .A2(n288), .ZN(n291) );
  XOR2_X1 U314 ( .A(n291), .B(n290), .Z(n292) );
  MUX2_X1 U315 ( .A(n535), .B(n292), .S(n15), .Z(n440) );
  MUX2_X1 U316 ( .A(product[5]), .B(n537), .S(n15), .Z(n442) );
  MUX2_X1 U317 ( .A(n537), .B(n538), .S(n15), .Z(n444) );
  MUX2_X1 U318 ( .A(product[6]), .B(n540), .S(n15), .Z(n448) );
  NAND2_X1 U319 ( .A1(n404), .A2(n356), .ZN(n293) );
  XOR2_X1 U320 ( .A(n293), .B(n358), .Z(n294) );
  MUX2_X1 U321 ( .A(n540), .B(n294), .S(n15), .Z(n450) );
  MUX2_X1 U322 ( .A(product[7]), .B(n542), .S(n15), .Z(n452) );
  OAI21_X1 U323 ( .B1(n355), .B2(n358), .A(n356), .ZN(n298) );
  NAND2_X1 U324 ( .A1(n342), .A2(n354), .ZN(n295) );
  XNOR2_X1 U325 ( .A(n298), .B(n295), .ZN(n297) );
  MUX2_X1 U326 ( .A(n542), .B(n297), .S(n15), .Z(n454) );
  BUF_X4 U327 ( .A(en), .Z(n336) );
  MUX2_X1 U328 ( .A(product[8]), .B(n544), .S(n336), .Z(n456) );
  AOI21_X1 U329 ( .B1(n298), .B2(n342), .A(n405), .ZN(n301) );
  NAND2_X1 U330 ( .A1(n406), .A2(n353), .ZN(n299) );
  XOR2_X1 U331 ( .A(n301), .B(n299), .Z(n300) );
  MUX2_X1 U332 ( .A(n544), .B(n300), .S(n336), .Z(n458) );
  MUX2_X1 U333 ( .A(product[9]), .B(n546), .S(n336), .Z(n460) );
  OAI21_X1 U334 ( .B1(n301), .B2(n352), .A(n353), .ZN(n309) );
  INV_X1 U335 ( .A(n309), .ZN(n304) );
  NAND2_X1 U336 ( .A1(n407), .A2(n351), .ZN(n302) );
  XOR2_X1 U337 ( .A(n304), .B(n302), .Z(n303) );
  MUX2_X1 U338 ( .A(n546), .B(n303), .S(n336), .Z(n462) );
  MUX2_X1 U339 ( .A(product[10]), .B(n548), .S(n336), .Z(n464) );
  OAI21_X1 U340 ( .B1(n304), .B2(n350), .A(n351), .ZN(n306) );
  NAND2_X1 U341 ( .A1(n403), .A2(n349), .ZN(n305) );
  XNOR2_X1 U342 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U343 ( .A(n548), .B(n307), .S(n336), .Z(n466) );
  MUX2_X1 U344 ( .A(product[11]), .B(n550), .S(n336), .Z(n468) );
  NOR2_X1 U345 ( .A1(n357), .A2(n350), .ZN(n310) );
  OAI21_X1 U346 ( .B1(n357), .B2(n351), .A(n349), .ZN(n308) );
  AOI21_X1 U347 ( .B1(n310), .B2(n309), .A(n308), .ZN(n332) );
  NAND2_X1 U348 ( .A1(n408), .A2(n348), .ZN(n311) );
  XOR2_X1 U349 ( .A(n332), .B(n311), .Z(n312) );
  MUX2_X1 U350 ( .A(n550), .B(n312), .S(n336), .Z(n470) );
  MUX2_X1 U351 ( .A(product[12]), .B(n552), .S(n336), .Z(n472) );
  OAI21_X1 U352 ( .B1(n332), .B2(n347), .A(n348), .ZN(n314) );
  NAND2_X1 U353 ( .A1(n341), .A2(n346), .ZN(n313) );
  XNOR2_X1 U354 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U355 ( .A(n552), .B(n315), .S(n336), .Z(n474) );
  MUX2_X1 U356 ( .A(product[13]), .B(n554), .S(n336), .Z(n476) );
  NAND2_X1 U357 ( .A1(n408), .A2(n341), .ZN(n317) );
  AOI21_X1 U358 ( .B1(n401), .B2(n341), .A(n409), .ZN(n316) );
  OAI21_X1 U359 ( .B1(n332), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U360 ( .A1(n340), .A2(n345), .ZN(n318) );
  XNOR2_X1 U361 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U362 ( .A(n554), .B(n320), .S(n336), .Z(n478) );
  MUX2_X1 U363 ( .A(product[14]), .B(n556), .S(n336), .Z(n480) );
  NAND2_X1 U364 ( .A1(n341), .A2(n340), .ZN(n322) );
  NOR2_X1 U365 ( .A1(n347), .A2(n322), .ZN(n328) );
  INV_X1 U366 ( .A(n328), .ZN(n324) );
  AOI21_X1 U367 ( .B1(n409), .B2(n340), .A(n400), .ZN(n321) );
  OAI21_X1 U368 ( .B1(n322), .B2(n348), .A(n321), .ZN(n329) );
  INV_X1 U369 ( .A(n329), .ZN(n323) );
  OAI21_X1 U370 ( .B1(n332), .B2(n324), .A(n323), .ZN(n326) );
  NAND2_X1 U371 ( .A1(n339), .A2(n344), .ZN(n325) );
  XNOR2_X1 U372 ( .A(n326), .B(n325), .ZN(n327) );
  MUX2_X1 U373 ( .A(n556), .B(n327), .S(n336), .Z(n482) );
  MUX2_X1 U374 ( .A(product[15]), .B(n558), .S(n336), .Z(n484) );
  NAND2_X1 U375 ( .A1(n328), .A2(n339), .ZN(n331) );
  AOI21_X1 U376 ( .B1(n329), .B2(n339), .A(n399), .ZN(n330) );
  OAI21_X1 U377 ( .B1(n332), .B2(n331), .A(n330), .ZN(n333) );
  XNOR2_X1 U378 ( .A(n333), .B(n343), .ZN(n334) );
  MUX2_X1 U379 ( .A(n558), .B(n334), .S(n336), .Z(n486) );
  MUX2_X1 U380 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n336), .Z(n488) );
  MUX2_X1 U381 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n336), .Z(n490) );
  MUX2_X1 U382 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n336), .Z(n492) );
  MUX2_X1 U383 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n336), .Z(n494) );
  MUX2_X1 U384 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n336), .Z(n496) );
  MUX2_X1 U385 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n336), .Z(n498) );
  MUX2_X1 U386 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n336), .Z(n500) );
  MUX2_X1 U387 ( .A(n14), .B(B_extended[7]), .S(n336), .Z(n502) );
  MUX2_X1 U388 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n336), .Z(n504) );
  MUX2_X1 U389 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n336), .Z(n506) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n336), .Z(n508) );
  MUX2_X1 U391 ( .A(n20), .B(A_extended[3]), .S(n336), .Z(n510) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n336), .Z(n512) );
  MUX2_X1 U393 ( .A(n335), .B(A_extended[5]), .S(n336), .Z(n514) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n336), .Z(n516) );
  MUX2_X1 U395 ( .A(n19), .B(A_extended[7]), .S(n336), .Z(n518) );
  OR2_X1 U396 ( .A1(n336), .A2(n560), .ZN(n520) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_1 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n365, n367, n369,
         n371, n373, n375, n377, n379, n381, n383, n385, n387, n389, n391,
         n393, n395, n397, n399, n401, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n416, n418, n420, n422, n424,
         n426, n428, n430, n432, n434, n436, n438, n440, n442, n444, n446,
         n448, n450, n452, n454, n456, n458, n460, n462, n464, n466, n468,
         n470, n472, n474, n476, n478, n480, n482, n484, n486, n488, n490,
         n492, n494, n496, n498, n500, n502, n504, n506, n508, n510, n512,
         n514, n516, n518, n520, n522, n524, n526, n527, n529, n530, n532,
         n533, n535, n536, n538, n539, n541, n542, n544, n546, n548, n550,
         n552, n554, n556, n558, n560, n562, n563, n564;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n414), .SE(n524), .CK(clk), .Q(n563), 
        .QN(n12) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n414), .SE(n520), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n24) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n414), .SE(n516), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n23) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n414), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n340) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n414), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n339) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n414), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n13) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n414), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n16) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n414), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n19) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n414), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n21) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n20) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n414), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n22) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n414), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n17) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n414), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n18) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n414), .SE(n490), .CK(clk), .Q(n562)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n414), .SE(n488), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n414), .SE(n486), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n414), .SE(n482), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n414), .SE(n480), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n414), .SE(n478), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n414), .SE(n476), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n414), .SE(n474), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n414), .SE(n470), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n414), .SE(n468), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n414), .SE(n466), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(rst_n), .SE(n464), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n414), .SE(n462), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n414), .SE(n460), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n414), .SE(n458), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n414), .SE(n456), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n454), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n414), .SE(n452), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n414), .SE(n450), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n414), .SE(n448), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n414), .SE(n442), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n414), .SE(n440), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n438), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n434), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n430), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n428), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n426), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n420), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n418), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n416), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n564), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n564), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n564), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n360), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n564), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n359), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n564), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n358), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n564), .SE(n391), .CK(
        clk), .Q(n26), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n564), .SE(n389), .CK(
        clk), .Q(n412), .QN(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n564), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n564), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n354), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n564), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n353), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n564), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n564), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n351), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n564), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n350), .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n564), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n349), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n564), .SE(n373), .CK(
        clk), .Q(n404), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n564), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n347), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n564), .SE(n369), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n564), .SE(n367), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n564), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n564), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n343), .QN(n411) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n414), .SE(n518), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n341) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n414), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n342) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n414), .SE(n522), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n15) );
  INV_X1 U2 ( .A(n105), .ZN(n7) );
  INV_X1 U3 ( .A(rst_n), .ZN(n564) );
  XOR2_X1 U4 ( .A(n339), .B(n340), .Z(n5) );
  OR2_X1 U5 ( .A1(n29), .A2(\mult_x_1/n180 ), .ZN(n227) );
  INV_X1 U6 ( .A(n68), .ZN(n60) );
  INV_X1 U7 ( .A(n67), .ZN(n59) );
  NAND2_X1 U8 ( .A1(n55), .A2(n54), .ZN(n68) );
  NAND2_X1 U9 ( .A1(n78), .A2(n79), .ZN(n54) );
  OAI21_X1 U10 ( .B1(n79), .B2(n78), .A(n80), .ZN(n55) );
  INV_X1 U11 ( .A(n130), .ZN(n127) );
  CLKBUF_X1 U12 ( .A(n342), .Z(n6) );
  INV_X1 U13 ( .A(n201), .ZN(n202) );
  OAI21_X1 U14 ( .B1(n204), .B2(n163), .A(n162), .ZN(n165) );
  NAND2_X1 U15 ( .A1(n63), .A2(n62), .ZN(n168) );
  NAND2_X1 U16 ( .A1(n68), .A2(n67), .ZN(n62) );
  NAND2_X1 U17 ( .A1(n60), .A2(n59), .ZN(n61) );
  NAND2_X1 U18 ( .A1(n188), .A2(n187), .ZN(n249) );
  NAND2_X1 U19 ( .A1(n192), .A2(n190), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n190), .B2(n192), .A(n191), .ZN(n188) );
  NAND2_X1 U21 ( .A1(n137), .A2(n136), .ZN(n240) );
  NAND2_X1 U22 ( .A1(n14), .A2(n135), .ZN(n136) );
  OAI21_X1 U23 ( .B1(n14), .B2(n135), .A(n134), .ZN(n137) );
  NAND2_X1 U24 ( .A1(n131), .A2(n130), .ZN(n132) );
  NAND2_X1 U25 ( .A1(n140), .A2(n139), .ZN(n82) );
  INV_X1 U26 ( .A(n105), .ZN(n207) );
  OR2_X1 U27 ( .A1(n27), .A2(n28), .ZN(n8) );
  INV_X1 U28 ( .A(n15), .ZN(n9) );
  NAND2_X1 U29 ( .A1(n203), .A2(n201), .ZN(n162) );
  NOR2_X1 U30 ( .A1(n203), .A2(n201), .ZN(n163) );
  XNOR2_X1 U31 ( .A(n203), .B(n202), .ZN(n205) );
  NOR2_X2 U32 ( .A1(n12), .A2(n16), .ZN(n102) );
  INV_X1 U33 ( .A(n5), .ZN(n10) );
  XNOR2_X1 U34 ( .A(n339), .B(n340), .ZN(n11) );
  INV_X1 U35 ( .A(n5), .ZN(n224) );
  XNOR2_X1 U36 ( .A(n70), .B(n69), .ZN(n140) );
  XNOR2_X1 U37 ( .A(n68), .B(n67), .ZN(n69) );
  XNOR2_X1 U38 ( .A(n342), .B(n23), .ZN(n33) );
  OR2_X1 U39 ( .A1(n38), .A2(n37), .ZN(n131) );
  AND2_X1 U40 ( .A1(n47), .A2(n46), .ZN(n14) );
  INV_X1 U41 ( .A(n341), .ZN(n337) );
  XNOR2_X1 U42 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n27) );
  XNOR2_X1 U43 ( .A(\mult_x_1/n311 ), .B(n24), .ZN(n28) );
  OR2_X1 U44 ( .A1(n27), .A2(n28), .ZN(n256) );
  XNOR2_X1 U45 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n51) );
  INV_X2 U46 ( .A(n28), .ZN(n257) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n43) );
  OAI22_X1 U48 ( .A1(n8), .A2(n51), .B1(n257), .B2(n43), .ZN(n73) );
  INV_X1 U49 ( .A(\mult_x_1/n313 ), .ZN(n29) );
  XNOR2_X1 U50 ( .A(n222), .B(\mult_x_1/n281 ), .ZN(n75) );
  XNOR2_X1 U51 ( .A(n102), .B(\mult_x_1/n313 ), .ZN(n40) );
  OAI22_X1 U52 ( .A1(n227), .A2(n75), .B1(n40), .B2(n13), .ZN(n72) );
  NAND2_X1 U53 ( .A1(n12), .A2(\mult_x_1/n310 ), .ZN(n39) );
  INV_X1 U54 ( .A(n39), .ZN(n30) );
  AND2_X1 U55 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n71) );
  XNOR2_X1 U56 ( .A(\mult_x_1/a[2] ), .B(n342), .ZN(n31) );
  NAND2_X1 U57 ( .A1(n31), .A2(n11), .ZN(n76) );
  XNOR2_X1 U58 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n49) );
  XNOR2_X1 U59 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n34) );
  OAI22_X1 U60 ( .A1(n76), .A2(n49), .B1(n224), .B2(n34), .ZN(n37) );
  INV_X1 U61 ( .A(n33), .ZN(n105) );
  XNOR2_X1 U62 ( .A(n337), .B(\mult_x_1/n283 ), .ZN(n36) );
  XNOR2_X1 U63 ( .A(\mult_x_1/n311 ), .B(n23), .ZN(n32) );
  NAND2_X1 U64 ( .A1(n33), .A2(n32), .ZN(n119) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n50) );
  OAI22_X1 U66 ( .A1(n207), .A2(n36), .B1(n119), .B2(n50), .ZN(n38) );
  XNOR2_X1 U67 ( .A(n37), .B(n38), .ZN(n46) );
  XNOR2_X1 U68 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n42) );
  XNOR2_X1 U69 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n122) );
  OAI22_X1 U70 ( .A1(n256), .A2(n42), .B1(n257), .B2(n122), .ZN(n116) );
  XNOR2_X1 U71 ( .A(n102), .B(\mult_x_1/n312 ), .ZN(n124) );
  OAI22_X1 U72 ( .A1(n76), .A2(n34), .B1(n124), .B2(n224), .ZN(n35) );
  INV_X1 U73 ( .A(n35), .ZN(n123) );
  XNOR2_X1 U74 ( .A(n337), .B(\mult_x_1/n282 ), .ZN(n118) );
  OAI22_X1 U75 ( .A1(n119), .A2(n36), .B1(n207), .B2(n118), .ZN(n115) );
  XNOR2_X1 U76 ( .A(n14), .B(n135), .ZN(n45) );
  NOR2_X1 U77 ( .A1(n17), .A2(n39), .ZN(n130) );
  XNOR2_X1 U78 ( .A(n131), .B(n130), .ZN(n44) );
  AOI21_X1 U79 ( .B1(n227), .B2(n13), .A(n40), .ZN(n41) );
  INV_X1 U80 ( .A(n41), .ZN(n58) );
  OAI22_X1 U81 ( .A1(n256), .A2(n43), .B1(n257), .B2(n42), .ZN(n57) );
  NOR2_X1 U82 ( .A1(n18), .A2(n39), .ZN(n56) );
  XNOR2_X1 U83 ( .A(n44), .B(n128), .ZN(n134) );
  XNOR2_X1 U84 ( .A(n45), .B(n134), .ZN(n169) );
  INV_X1 U85 ( .A(n46), .ZN(n48) );
  XNOR2_X1 U86 ( .A(n48), .B(n47), .ZN(n70) );
  BUF_X2 U87 ( .A(n76), .Z(n217) );
  XNOR2_X1 U88 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n77) );
  OAI22_X1 U89 ( .A1(n217), .A2(n77), .B1(n10), .B2(n49), .ZN(n79) );
  XNOR2_X1 U90 ( .A(n337), .B(\mult_x_1/n285 ), .ZN(n74) );
  OAI22_X1 U91 ( .A1(n119), .A2(n74), .B1(n207), .B2(n50), .ZN(n78) );
  XNOR2_X1 U92 ( .A(n9), .B(\mult_x_1/n288 ), .ZN(n52) );
  OAI22_X1 U93 ( .A1(n256), .A2(n52), .B1(n257), .B2(n51), .ZN(n89) );
  OR2_X1 U94 ( .A1(\mult_x_1/n288 ), .A2(n15), .ZN(n53) );
  OAI22_X1 U95 ( .A1(n256), .A2(n15), .B1(n53), .B2(n257), .ZN(n88) );
  AND2_X1 U96 ( .A1(n89), .A2(n88), .ZN(n80) );
  FA_X1 U97 ( .A(n58), .B(n57), .CI(n56), .CO(n128), .S(n67) );
  NAND2_X1 U98 ( .A1(n70), .A2(n61), .ZN(n63) );
  NAND2_X1 U99 ( .A1(n169), .A2(n168), .ZN(n64) );
  BUF_X2 U100 ( .A(en), .Z(n268) );
  NAND2_X1 U101 ( .A1(n64), .A2(n268), .ZN(n66) );
  OR2_X1 U102 ( .A1(n338), .A2(n26), .ZN(n65) );
  NAND2_X1 U103 ( .A1(n66), .A2(n65), .ZN(n391) );
  FA_X1 U104 ( .A(n73), .B(n72), .CI(n71), .CO(n47), .S(n144) );
  XNOR2_X1 U105 ( .A(n337), .B(\mult_x_1/n286 ), .ZN(n95) );
  OAI22_X1 U106 ( .A1(n119), .A2(n95), .B1(n7), .B2(n74), .ZN(n92) );
  CLKBUF_X1 U107 ( .A(\mult_x_1/n313 ), .Z(n222) );
  XNOR2_X1 U108 ( .A(n222), .B(\mult_x_1/n282 ), .ZN(n85) );
  OAI22_X1 U109 ( .A1(n227), .A2(n85), .B1(n75), .B2(n13), .ZN(n91) );
  XNOR2_X1 U110 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n87) );
  OAI22_X1 U111 ( .A1(n217), .A2(n87), .B1(n10), .B2(n77), .ZN(n90) );
  XNOR2_X1 U112 ( .A(n79), .B(n78), .ZN(n81) );
  XNOR2_X1 U113 ( .A(n81), .B(n80), .ZN(n142) );
  NAND2_X1 U114 ( .A1(n82), .A2(n338), .ZN(n84) );
  OR2_X1 U115 ( .A1(n338), .A2(n25), .ZN(n83) );
  NAND2_X1 U116 ( .A1(n84), .A2(n83), .ZN(n377) );
  XNOR2_X1 U137 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n161) );
  OAI22_X1 U138 ( .A1(n227), .A2(n161), .B1(n85), .B2(n13), .ZN(n99) );
  INV_X1 U139 ( .A(n257), .ZN(n86) );
  AND2_X1 U140 ( .A1(\mult_x_1/n288 ), .A2(n86), .ZN(n98) );
  XNOR2_X1 U141 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n160) );
  OAI22_X1 U142 ( .A1(n217), .A2(n160), .B1(n10), .B2(n87), .ZN(n97) );
  XOR2_X1 U143 ( .A(n89), .B(n88), .Z(n146) );
  FA_X1 U144 ( .A(n92), .B(n91), .CI(n90), .CO(n143), .S(n145) );
  OR2_X1 U145 ( .A1(\mult_x_1/n288 ), .A2(n341), .ZN(n93) );
  OAI22_X1 U146 ( .A1(n119), .A2(n341), .B1(n93), .B2(n7), .ZN(n159) );
  XNOR2_X1 U147 ( .A(n337), .B(\mult_x_1/n288 ), .ZN(n94) );
  XNOR2_X1 U148 ( .A(n337), .B(\mult_x_1/n287 ), .ZN(n96) );
  OAI22_X1 U149 ( .A1(n119), .A2(n94), .B1(n7), .B2(n96), .ZN(n158) );
  AND2_X1 U150 ( .A1(n159), .A2(n158), .ZN(n157) );
  OAI22_X1 U151 ( .A1(n119), .A2(n96), .B1(n7), .B2(n95), .ZN(n156) );
  FA_X1 U152 ( .A(n99), .B(n98), .CI(n97), .CO(n147), .S(n155) );
  OR2_X1 U153 ( .A1(n153), .A2(n152), .ZN(n100) );
  MUX2_X1 U154 ( .A(n345), .B(n100), .S(n338), .Z(n367) );
  NOR2_X1 U155 ( .A1(n19), .A2(n39), .ZN(n254) );
  XNOR2_X1 U156 ( .A(n9), .B(\mult_x_1/n281 ), .ZN(n101) );
  XNOR2_X1 U157 ( .A(n102), .B(n9), .ZN(n255) );
  OAI22_X1 U158 ( .A1(n8), .A2(n101), .B1(n255), .B2(n257), .ZN(n262) );
  INV_X1 U159 ( .A(n262), .ZN(n253) );
  XNOR2_X1 U160 ( .A(n9), .B(\mult_x_1/n282 ), .ZN(n108) );
  OAI22_X1 U161 ( .A1(n8), .A2(n108), .B1(n257), .B2(n101), .ZN(n113) );
  XNOR2_X1 U162 ( .A(n102), .B(\mult_x_1/n311 ), .ZN(n104) );
  AOI21_X1 U163 ( .B1(n7), .B2(n119), .A(n104), .ZN(n103) );
  INV_X1 U164 ( .A(n103), .ZN(n112) );
  XNOR2_X1 U165 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n117) );
  INV_X1 U166 ( .A(n104), .ZN(n106) );
  NAND2_X1 U167 ( .A1(n106), .A2(n105), .ZN(n107) );
  OAI21_X1 U168 ( .B1(n119), .B2(n117), .A(n107), .ZN(n111) );
  INV_X1 U169 ( .A(n111), .ZN(n177) );
  XNOR2_X1 U170 ( .A(n9), .B(\mult_x_1/n283 ), .ZN(n121) );
  OAI22_X1 U171 ( .A1(n8), .A2(n121), .B1(n257), .B2(n108), .ZN(n178) );
  NOR2_X1 U172 ( .A1(n20), .A2(n39), .ZN(n179) );
  OAI21_X1 U173 ( .B1(n177), .B2(n178), .A(n179), .ZN(n110) );
  NAND2_X1 U174 ( .A1(n178), .A2(n177), .ZN(n109) );
  NAND2_X1 U175 ( .A1(n110), .A2(n109), .ZN(n173) );
  NOR2_X1 U176 ( .A1(n21), .A2(n39), .ZN(n172) );
  FA_X1 U177 ( .A(n113), .B(n112), .CI(n111), .CO(n252), .S(n171) );
  NAND2_X1 U178 ( .A1(n246), .A2(n245), .ZN(n114) );
  MUX2_X1 U179 ( .A(n347), .B(n114), .S(n268), .Z(n371) );
  FA_X1 U180 ( .A(n115), .B(n116), .CI(n123), .CO(n182), .S(n135) );
  NOR2_X1 U181 ( .A1(n22), .A2(n39), .ZN(n184) );
  OAI22_X1 U182 ( .A1(n119), .A2(n118), .B1(n7), .B2(n117), .ZN(n183) );
  XNOR2_X1 U183 ( .A(n184), .B(n183), .ZN(n120) );
  XNOR2_X1 U184 ( .A(n182), .B(n120), .ZN(n196) );
  OAI22_X1 U185 ( .A1(n8), .A2(n122), .B1(n257), .B2(n121), .ZN(n176) );
  INV_X1 U186 ( .A(n123), .ZN(n175) );
  AOI21_X1 U187 ( .B1(n10), .B2(n217), .A(n124), .ZN(n125) );
  INV_X1 U188 ( .A(n125), .ZN(n174) );
  INV_X1 U189 ( .A(n131), .ZN(n126) );
  NAND2_X1 U190 ( .A1(n127), .A2(n126), .ZN(n129) );
  NAND2_X1 U191 ( .A1(n129), .A2(n128), .ZN(n133) );
  NAND2_X1 U192 ( .A1(n133), .A2(n132), .ZN(n194) );
  NOR2_X1 U193 ( .A1(n241), .A2(n240), .ZN(n138) );
  MUX2_X1 U194 ( .A(n348), .B(n138), .S(n268), .Z(n373) );
  NOR2_X1 U195 ( .A1(n140), .A2(n139), .ZN(n141) );
  MUX2_X1 U196 ( .A(n349), .B(n141), .S(n268), .Z(n375) );
  FA_X1 U197 ( .A(n144), .B(n143), .CI(n142), .CO(n139), .S(n150) );
  FA_X1 U198 ( .A(n147), .B(n146), .CI(n145), .CO(n149), .S(n153) );
  NOR2_X1 U199 ( .A1(n150), .A2(n149), .ZN(n148) );
  MUX2_X1 U200 ( .A(n351), .B(n148), .S(n338), .Z(n379) );
  NAND2_X1 U201 ( .A1(n150), .A2(n149), .ZN(n151) );
  MUX2_X1 U202 ( .A(n352), .B(n151), .S(n338), .Z(n381) );
  NAND2_X1 U203 ( .A1(n153), .A2(n152), .ZN(n154) );
  MUX2_X1 U204 ( .A(n353), .B(n154), .S(n338), .Z(n383) );
  FA_X1 U205 ( .A(n157), .B(n156), .CI(n155), .CO(n152), .S(n166) );
  XNOR2_X1 U206 ( .A(n159), .B(n158), .ZN(n204) );
  XNOR2_X1 U207 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n209) );
  OAI22_X1 U208 ( .A1(n217), .A2(n209), .B1(n10), .B2(n160), .ZN(n203) );
  XNOR2_X1 U209 ( .A(n222), .B(\mult_x_1/n284 ), .ZN(n206) );
  OAI22_X1 U210 ( .A1(n227), .A2(n206), .B1(n161), .B2(n13), .ZN(n201) );
  NOR2_X1 U211 ( .A1(n166), .A2(n165), .ZN(n164) );
  MUX2_X1 U212 ( .A(n354), .B(n164), .S(n268), .Z(n385) );
  NAND2_X1 U213 ( .A1(n166), .A2(n165), .ZN(n167) );
  MUX2_X1 U214 ( .A(n355), .B(n167), .S(n268), .Z(n387) );
  NOR2_X1 U215 ( .A1(n169), .A2(n168), .ZN(n170) );
  MUX2_X1 U216 ( .A(n356), .B(n170), .S(n338), .Z(n389) );
  FA_X1 U217 ( .A(n173), .B(n172), .CI(n171), .CO(n245), .S(n248) );
  FA_X1 U218 ( .A(n176), .B(n175), .CI(n174), .CO(n190), .S(n195) );
  XNOR2_X1 U219 ( .A(n178), .B(n177), .ZN(n180) );
  XNOR2_X1 U220 ( .A(n180), .B(n179), .ZN(n192) );
  OR2_X1 U221 ( .A1(n184), .A2(n183), .ZN(n181) );
  NAND2_X1 U222 ( .A1(n182), .A2(n181), .ZN(n186) );
  NAND2_X1 U223 ( .A1(n184), .A2(n183), .ZN(n185) );
  NAND2_X1 U224 ( .A1(n186), .A2(n185), .ZN(n191) );
  NAND2_X1 U225 ( .A1(n248), .A2(n249), .ZN(n189) );
  MUX2_X1 U226 ( .A(n358), .B(n189), .S(n338), .Z(n393) );
  XNOR2_X1 U227 ( .A(n191), .B(n190), .ZN(n193) );
  XNOR2_X1 U228 ( .A(n193), .B(n192), .ZN(n199) );
  FA_X1 U229 ( .A(n196), .B(n195), .CI(n194), .CO(n198), .S(n241) );
  NAND2_X1 U230 ( .A1(n199), .A2(n198), .ZN(n197) );
  MUX2_X1 U231 ( .A(n359), .B(n197), .S(n338), .Z(n395) );
  OR2_X1 U232 ( .A1(n199), .A2(n198), .ZN(n200) );
  MUX2_X1 U233 ( .A(n361), .B(n200), .S(n338), .Z(n399) );
  XNOR2_X1 U234 ( .A(n205), .B(n204), .ZN(n237) );
  INV_X1 U235 ( .A(n237), .ZN(n211) );
  XNOR2_X1 U236 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n218) );
  OAI22_X1 U237 ( .A1(n227), .A2(n218), .B1(n206), .B2(n13), .ZN(n214) );
  INV_X1 U238 ( .A(n7), .ZN(n208) );
  AND2_X1 U239 ( .A1(\mult_x_1/n288 ), .A2(n208), .ZN(n213) );
  XNOR2_X1 U240 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n215) );
  OAI22_X1 U241 ( .A1(n76), .A2(n215), .B1(n10), .B2(n209), .ZN(n212) );
  INV_X1 U242 ( .A(n236), .ZN(n210) );
  NAND2_X1 U243 ( .A1(n211), .A2(n210), .ZN(n292) );
  FA_X1 U244 ( .A(n214), .B(n213), .CI(n212), .CO(n236), .S(n235) );
  XNOR2_X1 U245 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n216) );
  OAI22_X1 U246 ( .A1(n217), .A2(n216), .B1(n10), .B2(n215), .ZN(n220) );
  XNOR2_X1 U247 ( .A(n222), .B(\mult_x_1/n286 ), .ZN(n223) );
  OAI22_X1 U248 ( .A1(n227), .A2(n223), .B1(n218), .B2(n13), .ZN(n219) );
  NOR2_X1 U249 ( .A1(n235), .A2(n234), .ZN(n285) );
  HA_X1 U250 ( .A(n220), .B(n219), .CO(n234), .S(n232) );
  OR2_X1 U251 ( .A1(\mult_x_1/n288 ), .A2(n6), .ZN(n221) );
  OAI22_X1 U252 ( .A1(n76), .A2(n6), .B1(n221), .B2(n10), .ZN(n231) );
  OR2_X1 U253 ( .A1(n232), .A2(n231), .ZN(n281) );
  XNOR2_X1 U254 ( .A(n222), .B(\mult_x_1/n287 ), .ZN(n226) );
  OAI22_X1 U255 ( .A1(n227), .A2(n226), .B1(n223), .B2(n13), .ZN(n230) );
  INV_X1 U256 ( .A(n10), .ZN(n225) );
  AND2_X1 U257 ( .A1(\mult_x_1/n288 ), .A2(n225), .ZN(n229) );
  NOR2_X1 U258 ( .A1(n230), .A2(n229), .ZN(n274) );
  OAI22_X1 U259 ( .A1(n227), .A2(\mult_x_1/n288 ), .B1(n226), .B2(n13), .ZN(
        n271) );
  OR2_X1 U260 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n228) );
  NAND2_X1 U261 ( .A1(n228), .A2(n227), .ZN(n270) );
  NAND2_X1 U262 ( .A1(n271), .A2(n270), .ZN(n277) );
  NAND2_X1 U263 ( .A1(n230), .A2(n229), .ZN(n275) );
  OAI21_X1 U264 ( .B1(n274), .B2(n277), .A(n275), .ZN(n282) );
  NAND2_X1 U265 ( .A1(n232), .A2(n231), .ZN(n280) );
  INV_X1 U266 ( .A(n280), .ZN(n233) );
  AOI21_X1 U267 ( .B1(n281), .B2(n282), .A(n233), .ZN(n288) );
  NAND2_X1 U268 ( .A1(n235), .A2(n234), .ZN(n286) );
  OAI21_X1 U269 ( .B1(n285), .B2(n288), .A(n286), .ZN(n293) );
  NAND2_X1 U270 ( .A1(n237), .A2(n236), .ZN(n291) );
  INV_X1 U271 ( .A(n291), .ZN(n238) );
  AOI21_X1 U272 ( .B1(n292), .B2(n293), .A(n238), .ZN(n239) );
  MUX2_X1 U273 ( .A(n362), .B(n239), .S(n268), .Z(n401) );
  INV_X1 U274 ( .A(n268), .ZN(n266) );
  NAND2_X1 U275 ( .A1(n360), .A2(n266), .ZN(n244) );
  NAND2_X1 U276 ( .A1(n241), .A2(n240), .ZN(n242) );
  NAND2_X1 U277 ( .A1(n242), .A2(n338), .ZN(n243) );
  NAND2_X1 U278 ( .A1(n244), .A2(n243), .ZN(n397) );
  OAI21_X1 U279 ( .B1(n246), .B2(n245), .A(n338), .ZN(n247) );
  OAI21_X1 U280 ( .B1(n338), .B2(n411), .A(n247), .ZN(n363) );
  NOR2_X1 U281 ( .A1(n249), .A2(n248), .ZN(n251) );
  NAND2_X1 U282 ( .A1(n266), .A2(n344), .ZN(n250) );
  OAI21_X1 U283 ( .B1(n251), .B2(n266), .A(n250), .ZN(n365) );
  FA_X1 U284 ( .A(n254), .B(n253), .CI(n252), .CO(n264), .S(n246) );
  AOI21_X1 U285 ( .B1(n257), .B2(n8), .A(n255), .ZN(n258) );
  INV_X1 U286 ( .A(n258), .ZN(n260) );
  NOR2_X1 U287 ( .A1(n16), .A2(n39), .ZN(n259) );
  XOR2_X1 U288 ( .A(n260), .B(n259), .Z(n261) );
  XNOR2_X1 U289 ( .A(n262), .B(n261), .ZN(n263) );
  XNOR2_X1 U290 ( .A(n264), .B(n263), .ZN(n267) );
  NAND2_X1 U291 ( .A1(n266), .A2(n346), .ZN(n265) );
  OAI21_X1 U292 ( .B1(n267), .B2(n266), .A(n265), .ZN(n369) );
  BUF_X2 U293 ( .A(rst_n), .Z(n414) );
  MUX2_X1 U294 ( .A(product[0]), .B(n526), .S(n338), .Z(n416) );
  MUX2_X1 U295 ( .A(n526), .B(n527), .S(n338), .Z(n418) );
  AND2_X1 U296 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n269) );
  MUX2_X1 U297 ( .A(n527), .B(n269), .S(n338), .Z(n420) );
  MUX2_X1 U298 ( .A(product[1]), .B(n529), .S(n338), .Z(n422) );
  MUX2_X1 U299 ( .A(n529), .B(n530), .S(n338), .Z(n424) );
  OR2_X1 U300 ( .A1(n271), .A2(n270), .ZN(n272) );
  AND2_X1 U301 ( .A1(n272), .A2(n277), .ZN(n273) );
  MUX2_X1 U302 ( .A(n530), .B(n273), .S(n268), .Z(n426) );
  MUX2_X1 U303 ( .A(product[2]), .B(n532), .S(n338), .Z(n428) );
  MUX2_X1 U304 ( .A(n532), .B(n533), .S(n338), .Z(n430) );
  INV_X1 U305 ( .A(n274), .ZN(n276) );
  NAND2_X1 U306 ( .A1(n276), .A2(n275), .ZN(n278) );
  XOR2_X1 U307 ( .A(n278), .B(n277), .Z(n279) );
  MUX2_X1 U308 ( .A(n533), .B(n279), .S(n338), .Z(n432) );
  MUX2_X1 U309 ( .A(product[3]), .B(n535), .S(n268), .Z(n434) );
  MUX2_X1 U310 ( .A(n535), .B(n536), .S(n338), .Z(n436) );
  NAND2_X1 U311 ( .A1(n281), .A2(n280), .ZN(n283) );
  XNOR2_X1 U312 ( .A(n283), .B(n282), .ZN(n284) );
  MUX2_X1 U313 ( .A(n536), .B(n284), .S(n268), .Z(n438) );
  MUX2_X1 U314 ( .A(product[4]), .B(n538), .S(n338), .Z(n440) );
  MUX2_X1 U315 ( .A(n538), .B(n539), .S(n268), .Z(n442) );
  INV_X1 U316 ( .A(n285), .ZN(n287) );
  NAND2_X1 U317 ( .A1(n287), .A2(n286), .ZN(n289) );
  XOR2_X1 U318 ( .A(n289), .B(n288), .Z(n290) );
  MUX2_X1 U319 ( .A(n539), .B(n290), .S(n338), .Z(n444) );
  MUX2_X1 U320 ( .A(product[5]), .B(n541), .S(n268), .Z(n446) );
  MUX2_X1 U321 ( .A(n541), .B(n542), .S(n338), .Z(n448) );
  NAND2_X1 U322 ( .A1(n292), .A2(n291), .ZN(n294) );
  XNOR2_X1 U323 ( .A(n294), .B(n293), .ZN(n295) );
  MUX2_X1 U324 ( .A(n542), .B(n295), .S(n268), .Z(n450) );
  MUX2_X1 U325 ( .A(product[6]), .B(n544), .S(n338), .Z(n452) );
  NAND2_X1 U326 ( .A1(n406), .A2(n355), .ZN(n296) );
  XOR2_X1 U327 ( .A(n296), .B(n362), .Z(n297) );
  MUX2_X1 U328 ( .A(n544), .B(n297), .S(n338), .Z(n454) );
  MUX2_X1 U329 ( .A(product[7]), .B(n546), .S(n268), .Z(n456) );
  OAI21_X1 U330 ( .B1(n354), .B2(n362), .A(n355), .ZN(n300) );
  NAND2_X1 U331 ( .A1(n345), .A2(n353), .ZN(n298) );
  XNOR2_X1 U332 ( .A(n300), .B(n298), .ZN(n299) );
  MUX2_X1 U333 ( .A(n546), .B(n299), .S(n338), .Z(n458) );
  BUF_X4 U334 ( .A(en), .Z(n338) );
  MUX2_X1 U335 ( .A(product[8]), .B(n548), .S(n268), .Z(n460) );
  AOI21_X1 U336 ( .B1(n300), .B2(n345), .A(n408), .ZN(n303) );
  NAND2_X1 U337 ( .A1(n409), .A2(n352), .ZN(n301) );
  XOR2_X1 U338 ( .A(n303), .B(n301), .Z(n302) );
  MUX2_X1 U339 ( .A(n548), .B(n302), .S(n338), .Z(n462) );
  MUX2_X1 U340 ( .A(product[9]), .B(n550), .S(n338), .Z(n464) );
  OAI21_X1 U341 ( .B1(n303), .B2(n351), .A(n352), .ZN(n311) );
  INV_X1 U342 ( .A(n311), .ZN(n306) );
  NAND2_X1 U343 ( .A1(n410), .A2(n350), .ZN(n304) );
  XOR2_X1 U344 ( .A(n306), .B(n304), .Z(n305) );
  MUX2_X1 U345 ( .A(n550), .B(n305), .S(n268), .Z(n466) );
  MUX2_X1 U346 ( .A(product[10]), .B(n552), .S(n338), .Z(n468) );
  OAI21_X1 U347 ( .B1(n306), .B2(n349), .A(n350), .ZN(n308) );
  NAND2_X1 U348 ( .A1(n412), .A2(n357), .ZN(n307) );
  XNOR2_X1 U349 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U350 ( .A(n552), .B(n309), .S(n338), .Z(n470) );
  MUX2_X1 U351 ( .A(product[11]), .B(n554), .S(n268), .Z(n472) );
  NOR2_X1 U352 ( .A1(n356), .A2(n349), .ZN(n312) );
  OAI21_X1 U353 ( .B1(n356), .B2(n350), .A(n357), .ZN(n310) );
  AOI21_X1 U354 ( .B1(n312), .B2(n311), .A(n310), .ZN(n334) );
  NAND2_X1 U355 ( .A1(n404), .A2(n360), .ZN(n313) );
  XOR2_X1 U356 ( .A(n334), .B(n313), .Z(n314) );
  MUX2_X1 U357 ( .A(n554), .B(n314), .S(n338), .Z(n474) );
  MUX2_X1 U358 ( .A(product[12]), .B(n556), .S(n338), .Z(n476) );
  OAI21_X1 U359 ( .B1(n334), .B2(n348), .A(n360), .ZN(n316) );
  NAND2_X1 U360 ( .A1(n361), .A2(n359), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n316), .B(n315), .ZN(n317) );
  MUX2_X1 U362 ( .A(n556), .B(n317), .S(n338), .Z(n478) );
  MUX2_X1 U363 ( .A(product[13]), .B(n558), .S(n268), .Z(n480) );
  NAND2_X1 U364 ( .A1(n404), .A2(n361), .ZN(n319) );
  AOI21_X1 U365 ( .B1(n405), .B2(n361), .A(n413), .ZN(n318) );
  OAI21_X1 U366 ( .B1(n334), .B2(n319), .A(n318), .ZN(n321) );
  NAND2_X1 U367 ( .A1(n344), .A2(n358), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U369 ( .A(n558), .B(n322), .S(n338), .Z(n482) );
  MUX2_X1 U370 ( .A(product[14]), .B(n560), .S(n338), .Z(n484) );
  NAND2_X1 U371 ( .A1(n361), .A2(n344), .ZN(n324) );
  NOR2_X1 U372 ( .A1(n348), .A2(n324), .ZN(n330) );
  INV_X1 U373 ( .A(n330), .ZN(n326) );
  AOI21_X1 U374 ( .B1(n413), .B2(n344), .A(n403), .ZN(n323) );
  OAI21_X1 U375 ( .B1(n324), .B2(n360), .A(n323), .ZN(n331) );
  INV_X1 U376 ( .A(n331), .ZN(n325) );
  OAI21_X1 U377 ( .B1(n334), .B2(n326), .A(n325), .ZN(n328) );
  NAND2_X1 U378 ( .A1(n343), .A2(n347), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  MUX2_X1 U380 ( .A(n560), .B(n329), .S(n268), .Z(n486) );
  MUX2_X1 U381 ( .A(product[15]), .B(n562), .S(n338), .Z(n488) );
  NAND2_X1 U382 ( .A1(n330), .A2(n343), .ZN(n333) );
  AOI21_X1 U383 ( .B1(n331), .B2(n343), .A(n407), .ZN(n332) );
  OAI21_X1 U384 ( .B1(n334), .B2(n333), .A(n332), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n335), .B(n346), .ZN(n336) );
  MUX2_X1 U386 ( .A(n562), .B(n336), .S(n338), .Z(n490) );
  MUX2_X1 U387 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n268), .Z(n492) );
  MUX2_X1 U388 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n338), .Z(n494) );
  MUX2_X1 U389 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n338), .Z(n496) );
  MUX2_X1 U390 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n268), .Z(n498) );
  MUX2_X1 U391 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n338), .Z(n500) );
  MUX2_X1 U392 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n338), .Z(n502) );
  MUX2_X1 U393 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n338), .Z(n504) );
  MUX2_X1 U394 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n268), .Z(n506) );
  MUX2_X1 U395 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n338), .Z(n508) );
  MUX2_X1 U396 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n338), .Z(n510) );
  MUX2_X1 U397 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n268), .Z(n512) );
  MUX2_X1 U398 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n338), .Z(n514) );
  MUX2_X1 U399 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n338), .Z(n516) );
  MUX2_X1 U400 ( .A(n337), .B(A_extended[5]), .S(n268), .Z(n518) );
  MUX2_X1 U401 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n338), .Z(n520) );
  MUX2_X1 U402 ( .A(n9), .B(A_extended[7]), .S(n338), .Z(n522) );
  OR2_X1 U403 ( .A1(n338), .A2(n563), .ZN(n524) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_2 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n367, n369, n371, n373,
         n375, n377, n379, n381, n383, n385, n387, n389, n391, n393, n395,
         n397, n399, n401, n403, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n419, n421, n423, n425, n427,
         n429, n431, n433, n435, n437, n439, n441, n443, n445, n447, n449,
         n451, n453, n455, n457, n459, n461, n463, n465, n467, n469, n471,
         n473, n475, n477, n479, n481, n483, n485, n487, n489, n491, n493,
         n495, n497, n499, n501, n503, n505, n507, n509, n511, n513, n515,
         n517, n519, n521, n523, n525, n527, n529, n530, n532, n533, n535,
         n536, n538, n539, n541, n542, n544, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n566, n567, n568;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n417), .SE(n527), .CK(clk), .Q(n567)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n523), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n344) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n417), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n342) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n417), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n31) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n417), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n20) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n417), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n28) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n417), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n27) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n24) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n417), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n25) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n26) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n417), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n21) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n493), .CK(clk), .Q(n565)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n491), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n417), .SE(n489), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n417), .SE(n487), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(rst_n), .SE(n485), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n417), .SE(n483), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(rst_n), .SE(n481), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n417), .SE(n479), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(rst_n), .SE(n477), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n417), .SE(n475), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG23_S3 ( .D(1'b0), .SI(rst_n), .SE(n473), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG24_S4 ( .D(1'b0), .SI(rst_n), .SE(n471), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG21_S3 ( .D(1'b0), .SI(rst_n), .SE(n469), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG22_S4 ( .D(1'b0), .SI(rst_n), .SE(n467), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n465), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(rst_n), .SE(n463), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n461), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n459), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n457), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n455), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n453), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n451), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n449), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n447), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n445), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n443), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n441), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n417), .SE(n439), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n417), .SE(n437), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n417), .SE(n435), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n417), .SE(n433), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n417), .SE(n431), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n417), .SE(n429), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n417), .SE(n427), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n417), .SE(n425), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n417), .SE(n423), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n417), .SE(n421), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n417), .SE(n419), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n417), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n33) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n417), .SE(n525), .CK(clk), .Q(n566), 
        .QN(n22) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n568), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n364) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n568), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n363), .QN(n416) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n568), .SE(n399), .CK(
        clk), .Q(n415), .QN(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n568), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n361), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n568), .SE(n395), .CK(
        clk), .Q(n405), .QN(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n568), .SE(n393), .CK(
        clk), .Q(n406), .QN(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n568), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n568), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n357), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n568), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n356), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n568), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n568), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n354), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n568), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n568), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n352), .QN(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n568), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n351), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n568), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n350), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n568), .SE(n373), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n568), .SE(n371), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n568), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n568), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n568), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n345), .QN(n409) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n343) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n417), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n341) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n23) );
  INV_X1 U2 ( .A(n7), .ZN(n215) );
  XNOR2_X2 U3 ( .A(n341), .B(n342), .ZN(n36) );
  XNOR2_X1 U4 ( .A(n66), .B(n65), .ZN(n67) );
  NAND2_X1 U5 ( .A1(n6), .A2(n5), .ZN(n66) );
  INV_X1 U6 ( .A(n56), .ZN(n5) );
  INV_X1 U7 ( .A(n55), .ZN(n6) );
  XOR2_X1 U8 ( .A(n343), .B(n344), .Z(n7) );
  CLKBUF_X2 U9 ( .A(n119), .Z(n229) );
  CLKBUF_X2 U10 ( .A(n46), .Z(n8) );
  BUF_X1 U11 ( .A(n39), .Z(n10) );
  AND2_X1 U12 ( .A1(n567), .A2(\mult_x_1/n281 ), .ZN(n176) );
  INV_X1 U13 ( .A(n33), .ZN(n9) );
  XNOR2_X1 U14 ( .A(n127), .B(n126), .ZN(n147) );
  INV_X1 U15 ( .A(n147), .ZN(n139) );
  AND2_X1 U16 ( .A1(n566), .A2(n567), .ZN(n41) );
  NAND2_X1 U17 ( .A1(n109), .A2(n108), .ZN(n110) );
  INV_X1 U18 ( .A(n113), .ZN(n109) );
  INV_X1 U19 ( .A(n112), .ZN(n108) );
  XNOR2_X1 U20 ( .A(n30), .B(n149), .ZN(n263) );
  XNOR2_X1 U21 ( .A(n161), .B(n160), .ZN(n231) );
  NAND2_X1 U22 ( .A1(n142), .A2(n141), .ZN(n271) );
  NAND2_X1 U23 ( .A1(n113), .A2(n112), .ZN(n114) );
  OR2_X1 U24 ( .A1(n77), .A2(n76), .ZN(n260) );
  NAND2_X1 U25 ( .A1(n77), .A2(n76), .ZN(n257) );
  BUF_X1 U26 ( .A(\mult_x_1/n312 ), .Z(n15) );
  BUF_X1 U27 ( .A(\mult_x_1/n311 ), .Z(n16) );
  NAND2_X1 U28 ( .A1(n229), .A2(n162), .ZN(n164) );
  INV_X1 U29 ( .A(n262), .ZN(n162) );
  INV_X1 U30 ( .A(n15), .ZN(n11) );
  OAI22_X1 U31 ( .A1(n57), .A2(n214), .B1(n215), .B2(n49), .ZN(n126) );
  NAND2_X1 U32 ( .A1(n35), .A2(n17), .ZN(n12) );
  NAND2_X1 U33 ( .A1(n35), .A2(n17), .ZN(n13) );
  NAND2_X1 U34 ( .A1(n35), .A2(n17), .ZN(n205) );
  XNOR2_X1 U35 ( .A(n125), .B(n124), .ZN(n127) );
  BUF_X1 U36 ( .A(n111), .Z(n14) );
  BUF_X4 U37 ( .A(n566), .Z(n339) );
  XNOR2_X1 U38 ( .A(n341), .B(n342), .ZN(n17) );
  BUF_X1 U39 ( .A(n255), .Z(n18) );
  XNOR2_X1 U40 ( .A(n343), .B(n344), .ZN(n19) );
  OAI21_X1 U41 ( .B1(n18), .B2(n254), .A(en), .ZN(n121) );
  BUF_X1 U42 ( .A(en), .Z(n119) );
  BUF_X1 U43 ( .A(rst_n), .Z(n417) );
  INV_X1 U44 ( .A(rst_n), .ZN(n568) );
  XOR2_X1 U45 ( .A(n123), .B(n122), .Z(n30) );
  AND2_X1 U46 ( .A1(n123), .A2(n122), .ZN(n32) );
  XNOR2_X1 U47 ( .A(n339), .B(n344), .ZN(n34) );
  NAND2_X2 U48 ( .A1(n34), .A2(n19), .ZN(n214) );
  XNOR2_X1 U49 ( .A(n339), .B(\mult_x_1/n285 ), .ZN(n49) );
  XNOR2_X1 U50 ( .A(n339), .B(\mult_x_1/n284 ), .ZN(n43) );
  OAI22_X1 U51 ( .A1(n214), .A2(n49), .B1(n215), .B2(n43), .ZN(n64) );
  XOR2_X1 U52 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n35) );
  XNOR2_X1 U53 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n48) );
  INV_X1 U54 ( .A(n36), .ZN(n37) );
  XNOR2_X1 U55 ( .A(n16), .B(\mult_x_1/n282 ), .ZN(n40) );
  OAI22_X1 U56 ( .A1(n12), .A2(n48), .B1(n36), .B2(n40), .ZN(n63) );
  XNOR2_X1 U57 ( .A(n176), .B(\mult_x_1/n312 ), .ZN(n44) );
  XNOR2_X1 U58 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n39) );
  XNOR2_X1 U59 ( .A(n31), .B(\mult_x_1/n312 ), .ZN(n38) );
  NAND2_X1 U60 ( .A1(n39), .A2(n38), .ZN(n46) );
  XNOR2_X1 U61 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n47) );
  OAI22_X1 U62 ( .A1(n44), .A2(n10), .B1(n46), .B2(n47), .ZN(n106) );
  INV_X1 U63 ( .A(n106), .ZN(n62) );
  XNOR2_X1 U64 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n174) );
  OAI22_X1 U65 ( .A1(n12), .A2(n40), .B1(n17), .B2(n174), .ZN(n113) );
  XNOR2_X1 U66 ( .A(n41), .B(n339), .ZN(n217) );
  NOR2_X1 U67 ( .A1(n24), .A2(n217), .ZN(n112) );
  XNOR2_X1 U68 ( .A(n113), .B(n112), .ZN(n42) );
  XNOR2_X1 U69 ( .A(n14), .B(n42), .ZN(n118) );
  XNOR2_X1 U70 ( .A(n339), .B(\mult_x_1/n283 ), .ZN(n103) );
  OAI22_X1 U71 ( .A1(n214), .A2(n43), .B1(n215), .B2(n103), .ZN(n107) );
  AOI21_X1 U72 ( .B1(n10), .B2(n8), .A(n44), .ZN(n45) );
  INV_X1 U73 ( .A(n45), .ZN(n105) );
  XNOR2_X1 U74 ( .A(n15), .B(\mult_x_1/n282 ), .ZN(n132) );
  OAI22_X1 U75 ( .A1(n8), .A2(n132), .B1(n10), .B2(n47), .ZN(n55) );
  XNOR2_X1 U76 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n131) );
  OAI22_X1 U77 ( .A1(n36), .A2(n48), .B1(n13), .B2(n131), .ZN(n56) );
  NOR2_X1 U78 ( .A1(n25), .A2(n217), .ZN(n65) );
  XNOR2_X1 U79 ( .A(n339), .B(\mult_x_1/n286 ), .ZN(n57) );
  NAND2_X1 U80 ( .A1(n20), .A2(n9), .ZN(n193) );
  CLKBUF_X1 U81 ( .A(\mult_x_1/n313 ), .Z(n73) );
  XNOR2_X1 U82 ( .A(n176), .B(n73), .ZN(n58) );
  AOI21_X1 U83 ( .B1(n193), .B2(n20), .A(n58), .ZN(n50) );
  INV_X1 U84 ( .A(n50), .ZN(n124) );
  NOR2_X1 U85 ( .A1(n26), .A2(n217), .ZN(n125) );
  OAI21_X1 U86 ( .B1(n126), .B2(n124), .A(n125), .ZN(n52) );
  NAND2_X1 U87 ( .A1(n124), .A2(n126), .ZN(n51) );
  NAND2_X1 U88 ( .A1(n52), .A2(n51), .ZN(n68) );
  OAI21_X1 U89 ( .B1(n66), .B2(n65), .A(n68), .ZN(n54) );
  NAND2_X1 U90 ( .A1(n66), .A2(n65), .ZN(n53) );
  NAND2_X1 U91 ( .A1(n54), .A2(n53), .ZN(n116) );
  NAND2_X1 U92 ( .A1(n274), .A2(n351), .ZN(n70) );
  XNOR2_X1 U93 ( .A(n56), .B(n55), .ZN(n123) );
  XNOR2_X1 U94 ( .A(n339), .B(\mult_x_1/n287 ), .ZN(n129) );
  OAI22_X1 U95 ( .A1(n214), .A2(n129), .B1(n215), .B2(n57), .ZN(n154) );
  XNOR2_X1 U96 ( .A(n73), .B(\mult_x_1/n281 ), .ZN(n156) );
  OAI22_X1 U97 ( .A1(n193), .A2(n156), .B1(n58), .B2(n20), .ZN(n150) );
  NAND2_X1 U98 ( .A1(n154), .A2(n150), .ZN(n61) );
  OR2_X1 U99 ( .A1(n217), .A2(n21), .ZN(n152) );
  INV_X1 U100 ( .A(n152), .ZN(n59) );
  OAI21_X1 U101 ( .B1(n154), .B2(n150), .A(n59), .ZN(n60) );
  NAND2_X1 U102 ( .A1(n61), .A2(n60), .ZN(n122) );
  FA_X1 U103 ( .A(n64), .B(n63), .CI(n62), .CO(n111), .S(n145) );
  XNOR2_X1 U104 ( .A(n68), .B(n67), .ZN(n144) );
  NAND2_X1 U105 ( .A1(n166), .A2(n229), .ZN(n69) );
  OAI211_X1 U106 ( .C1(n168), .C2(n274), .A(n70), .B(n69), .ZN(n377) );
  XNOR2_X1 U107 ( .A(n15), .B(\mult_x_1/n286 ), .ZN(n75) );
  XNOR2_X1 U108 ( .A(n15), .B(\mult_x_1/n285 ), .ZN(n195) );
  OAI22_X1 U109 ( .A1(n8), .A2(n75), .B1(n10), .B2(n195), .ZN(n246) );
  XNOR2_X1 U110 ( .A(n9), .B(\mult_x_1/n284 ), .ZN(n74) );
  XNOR2_X1 U111 ( .A(n73), .B(\mult_x_1/n283 ), .ZN(n192) );
  OAI22_X1 U112 ( .A1(n193), .A2(n74), .B1(n192), .B2(n20), .ZN(n245) );
  OR2_X1 U113 ( .A1(\mult_x_1/n288 ), .A2(n343), .ZN(n71) );
  OAI22_X1 U114 ( .A1(n13), .A2(n343), .B1(n71), .B2(n36), .ZN(n202) );
  XNOR2_X1 U115 ( .A(n16), .B(\mult_x_1/n288 ), .ZN(n72) );
  XNOR2_X1 U116 ( .A(n16), .B(\mult_x_1/n287 ), .ZN(n204) );
  OAI22_X1 U117 ( .A1(n12), .A2(n72), .B1(n36), .B2(n204), .ZN(n201) );
  XNOR2_X1 U118 ( .A(n73), .B(\mult_x_1/n285 ), .ZN(n80) );
  OAI22_X1 U119 ( .A1(n193), .A2(n80), .B1(n74), .B2(n20), .ZN(n94) );
  AND2_X1 U120 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n93) );
  XNOR2_X1 U121 ( .A(n15), .B(\mult_x_1/n287 ), .ZN(n78) );
  OAI22_X1 U122 ( .A1(n8), .A2(n78), .B1(n10), .B2(n75), .ZN(n92) );
  NAND2_X1 U123 ( .A1(n260), .A2(n257), .ZN(n100) );
  XNOR2_X1 U124 ( .A(n15), .B(\mult_x_1/n288 ), .ZN(n79) );
  OAI22_X1 U125 ( .A1(n8), .A2(n79), .B1(n10), .B2(n78), .ZN(n96) );
  XNOR2_X1 U126 ( .A(n9), .B(\mult_x_1/n286 ), .ZN(n83) );
  OAI22_X1 U127 ( .A1(n193), .A2(n83), .B1(n80), .B2(n20), .ZN(n95) );
  INV_X1 U128 ( .A(n95), .ZN(n81) );
  XNOR2_X1 U129 ( .A(n96), .B(n81), .ZN(n90) );
  OR2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n11), .ZN(n82) );
  OAI22_X1 U131 ( .A1(n8), .A2(n11), .B1(n82), .B2(n10), .ZN(n89) );
  OR2_X1 U132 ( .A1(n90), .A2(n89), .ZN(n288) );
  XNOR2_X1 U133 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n85) );
  OAI22_X1 U134 ( .A1(n193), .A2(n85), .B1(n83), .B2(n20), .ZN(n88) );
  INV_X1 U135 ( .A(n10), .ZN(n84) );
  AND2_X1 U136 ( .A1(\mult_x_1/n288 ), .A2(n84), .ZN(n87) );
  NOR2_X1 U137 ( .A1(n88), .A2(n87), .ZN(n281) );
  OAI22_X1 U138 ( .A1(n193), .A2(\mult_x_1/n288 ), .B1(n85), .B2(n20), .ZN(
        n278) );
  OR2_X1 U139 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n86) );
  NAND2_X1 U140 ( .A1(n86), .A2(n193), .ZN(n277) );
  NAND2_X1 U141 ( .A1(n278), .A2(n277), .ZN(n284) );
  NAND2_X1 U142 ( .A1(n88), .A2(n87), .ZN(n282) );
  OAI21_X1 U143 ( .B1(n281), .B2(n284), .A(n282), .ZN(n289) );
  NAND2_X1 U144 ( .A1(n90), .A2(n89), .ZN(n287) );
  INV_X1 U145 ( .A(n287), .ZN(n91) );
  AOI21_X1 U146 ( .B1(n288), .B2(n289), .A(n91), .ZN(n295) );
  FA_X1 U147 ( .A(n94), .B(n93), .CI(n92), .CO(n76), .S(n98) );
  AND2_X1 U148 ( .A1(n96), .A2(n95), .ZN(n97) );
  NOR2_X1 U149 ( .A1(n98), .A2(n97), .ZN(n292) );
  NAND2_X1 U150 ( .A1(n98), .A2(n97), .ZN(n293) );
  OAI21_X1 U151 ( .B1(n295), .B2(n292), .A(n293), .ZN(n259) );
  INV_X1 U152 ( .A(n259), .ZN(n99) );
  XNOR2_X1 U153 ( .A(n100), .B(n99), .ZN(n102) );
  NAND2_X1 U154 ( .A1(n274), .A2(n545), .ZN(n101) );
  OAI21_X1 U155 ( .B1(n102), .B2(n274), .A(n101), .ZN(n453) );
  XNOR2_X1 U156 ( .A(n339), .B(\mult_x_1/n282 ), .ZN(n172) );
  OAI22_X1 U157 ( .A1(n214), .A2(n103), .B1(n215), .B2(n172), .ZN(n171) );
  XNOR2_X1 U158 ( .A(n176), .B(\mult_x_1/n311 ), .ZN(n175) );
  OAI22_X1 U159 ( .A1(n36), .A2(n175), .B1(n205), .B2(n174), .ZN(n104) );
  INV_X1 U160 ( .A(n104), .ZN(n170) );
  NOR2_X1 U161 ( .A1(n27), .A2(n217), .ZN(n169) );
  FA_X1 U162 ( .A(n107), .B(n106), .CI(n105), .CO(n188), .S(n117) );
  NAND2_X1 U163 ( .A1(n111), .A2(n110), .ZN(n115) );
  NAND2_X1 U164 ( .A1(n115), .A2(n114), .ZN(n187) );
  FA_X1 U165 ( .A(n118), .B(n117), .CI(n116), .CO(n254), .S(n168) );
  NAND2_X1 U166 ( .A1(n274), .A2(n347), .ZN(n120) );
  NAND2_X1 U167 ( .A1(n121), .A2(n120), .ZN(n369) );
  OR2_X1 U168 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n128) );
  OAI22_X1 U169 ( .A1(n214), .A2(n22), .B1(n128), .B2(n215), .ZN(n197) );
  XNOR2_X1 U170 ( .A(n339), .B(\mult_x_1/n288 ), .ZN(n130) );
  OAI22_X1 U171 ( .A1(n214), .A2(n130), .B1(n215), .B2(n129), .ZN(n196) );
  XNOR2_X1 U172 ( .A(n16), .B(\mult_x_1/n285 ), .ZN(n155) );
  OAI22_X1 U173 ( .A1(n12), .A2(n155), .B1(n36), .B2(n131), .ZN(n159) );
  INV_X1 U174 ( .A(n159), .ZN(n134) );
  XNOR2_X1 U175 ( .A(n15), .B(\mult_x_1/n283 ), .ZN(n157) );
  OAI22_X1 U176 ( .A1(n8), .A2(n157), .B1(n10), .B2(n132), .ZN(n158) );
  INV_X1 U177 ( .A(n158), .ZN(n133) );
  NAND2_X1 U178 ( .A1(n134), .A2(n133), .ZN(n135) );
  NAND2_X1 U179 ( .A1(n161), .A2(n135), .ZN(n137) );
  NAND2_X1 U180 ( .A1(n159), .A2(n158), .ZN(n136) );
  NAND2_X1 U181 ( .A1(n137), .A2(n136), .ZN(n148) );
  INV_X1 U182 ( .A(n148), .ZN(n138) );
  NAND2_X1 U183 ( .A1(n139), .A2(n138), .ZN(n140) );
  NAND2_X1 U184 ( .A1(n30), .A2(n140), .ZN(n142) );
  NAND2_X1 U185 ( .A1(n147), .A2(n148), .ZN(n141) );
  INV_X1 U186 ( .A(n271), .ZN(n143) );
  NAND2_X1 U187 ( .A1(n143), .A2(n229), .ZN(n146) );
  FA_X1 U188 ( .A(n32), .B(n145), .CI(n144), .CO(n165), .S(n275) );
  OAI22_X1 U189 ( .A1(n146), .A2(n275), .B1(n340), .B2(n406), .ZN(n393) );
  XNOR2_X1 U190 ( .A(n148), .B(n147), .ZN(n149) );
  INV_X1 U191 ( .A(n150), .ZN(n151) );
  XNOR2_X1 U192 ( .A(n152), .B(n151), .ZN(n153) );
  XNOR2_X1 U193 ( .A(n154), .B(n153), .ZN(n233) );
  XNOR2_X1 U194 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n203) );
  OAI22_X1 U195 ( .A1(n13), .A2(n203), .B1(n36), .B2(n155), .ZN(n200) );
  XNOR2_X1 U196 ( .A(n9), .B(\mult_x_1/n282 ), .ZN(n191) );
  OAI22_X1 U197 ( .A1(n193), .A2(n191), .B1(n156), .B2(n20), .ZN(n199) );
  XNOR2_X1 U198 ( .A(n15), .B(\mult_x_1/n284 ), .ZN(n194) );
  OAI22_X1 U199 ( .A1(n8), .A2(n194), .B1(n10), .B2(n157), .ZN(n198) );
  XNOR2_X1 U200 ( .A(n159), .B(n158), .ZN(n160) );
  NAND2_X1 U201 ( .A1(n274), .A2(n352), .ZN(n163) );
  OAI21_X1 U202 ( .B1(n263), .B2(n164), .A(n163), .ZN(n379) );
  INV_X1 U203 ( .A(n165), .ZN(n166) );
  NAND2_X1 U204 ( .A1(n166), .A2(n229), .ZN(n167) );
  OAI22_X1 U205 ( .A1(n168), .A2(n167), .B1(n340), .B2(n415), .ZN(n399) );
  FA_X1 U226 ( .A(n171), .B(n170), .CI(n169), .CO(n186), .S(n189) );
  NOR2_X1 U227 ( .A1(n28), .A2(n217), .ZN(n185) );
  XNOR2_X1 U228 ( .A(n339), .B(\mult_x_1/n281 ), .ZN(n177) );
  OAI22_X1 U229 ( .A1(n214), .A2(n172), .B1(n215), .B2(n177), .ZN(n180) );
  AOI21_X1 U230 ( .B1(n36), .B2(n205), .A(n175), .ZN(n173) );
  INV_X1 U231 ( .A(n173), .ZN(n179) );
  OAI22_X1 U232 ( .A1(n36), .A2(n175), .B1(n12), .B2(n174), .ZN(n178) );
  INV_X1 U233 ( .A(n227), .ZN(n182) );
  NOR2_X1 U234 ( .A1(n29), .A2(n217), .ZN(n212) );
  XNOR2_X1 U235 ( .A(n176), .B(n339), .ZN(n213) );
  OAI22_X1 U236 ( .A1(n214), .A2(n177), .B1(n213), .B2(n215), .ZN(n221) );
  INV_X1 U237 ( .A(n221), .ZN(n211) );
  FA_X1 U238 ( .A(n180), .B(n179), .CI(n178), .CO(n210), .S(n184) );
  INV_X1 U239 ( .A(n228), .ZN(n181) );
  NAND2_X1 U240 ( .A1(n182), .A2(n181), .ZN(n183) );
  MUX2_X1 U241 ( .A(n345), .B(n183), .S(n229), .Z(n365) );
  FA_X1 U242 ( .A(n186), .B(n185), .CI(n184), .CO(n227), .S(n252) );
  FA_X1 U243 ( .A(n189), .B(n188), .CI(n187), .CO(n251), .S(n255) );
  OR2_X1 U244 ( .A1(n252), .A2(n251), .ZN(n190) );
  MUX2_X1 U245 ( .A(n346), .B(n190), .S(n340), .Z(n367) );
  OAI22_X1 U246 ( .A1(n193), .A2(n192), .B1(n191), .B2(n20), .ZN(n208) );
  AND2_X1 U247 ( .A1(\mult_x_1/n288 ), .A2(n7), .ZN(n207) );
  OAI22_X1 U248 ( .A1(n8), .A2(n195), .B1(n10), .B2(n194), .ZN(n206) );
  HA_X1 U249 ( .A(n197), .B(n196), .CO(n161), .S(n235) );
  FA_X1 U250 ( .A(n200), .B(n199), .CI(n198), .CO(n232), .S(n234) );
  HA_X1 U251 ( .A(n202), .B(n201), .CO(n243), .S(n244) );
  OAI22_X1 U252 ( .A1(n13), .A2(n204), .B1(n17), .B2(n203), .ZN(n242) );
  FA_X1 U253 ( .A(n208), .B(n207), .CI(n206), .CO(n236), .S(n241) );
  OR2_X1 U254 ( .A1(n239), .A2(n238), .ZN(n209) );
  MUX2_X1 U255 ( .A(n348), .B(n209), .S(n229), .Z(n371) );
  FA_X1 U256 ( .A(n212), .B(n211), .CI(n210), .CO(n223), .S(n228) );
  AOI21_X1 U257 ( .B1(n215), .B2(n214), .A(n213), .ZN(n216) );
  INV_X1 U258 ( .A(n216), .ZN(n219) );
  NOR2_X1 U259 ( .A1(n23), .A2(n217), .ZN(n218) );
  XOR2_X1 U260 ( .A(n219), .B(n218), .Z(n220) );
  XOR2_X1 U261 ( .A(n221), .B(n220), .Z(n222) );
  OR2_X1 U262 ( .A1(n223), .A2(n222), .ZN(n225) );
  NAND2_X1 U263 ( .A1(n223), .A2(n222), .ZN(n224) );
  NAND2_X1 U264 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U265 ( .A(n349), .B(n226), .S(n119), .Z(n373) );
  NAND2_X1 U266 ( .A1(n228), .A2(n227), .ZN(n230) );
  MUX2_X1 U267 ( .A(n350), .B(n230), .S(n229), .Z(n375) );
  FA_X1 U268 ( .A(n233), .B(n232), .CI(n231), .CO(n262), .S(n268) );
  FA_X1 U269 ( .A(n236), .B(n235), .CI(n234), .CO(n267), .S(n239) );
  NOR2_X1 U270 ( .A1(n268), .A2(n267), .ZN(n237) );
  MUX2_X1 U271 ( .A(n354), .B(n237), .S(n119), .Z(n383) );
  NAND2_X1 U272 ( .A1(n239), .A2(n238), .ZN(n240) );
  MUX2_X1 U273 ( .A(n356), .B(n240), .S(n119), .Z(n387) );
  FA_X1 U274 ( .A(n243), .B(n242), .CI(n241), .CO(n238), .S(n249) );
  FA_X1 U275 ( .A(n246), .B(n245), .CI(n244), .CO(n248), .S(n77) );
  NOR2_X1 U276 ( .A1(n249), .A2(n248), .ZN(n247) );
  MUX2_X1 U277 ( .A(n357), .B(n247), .S(n340), .Z(n389) );
  NAND2_X1 U278 ( .A1(n249), .A2(n248), .ZN(n250) );
  MUX2_X1 U279 ( .A(n358), .B(n250), .S(n340), .Z(n391) );
  NAND2_X1 U280 ( .A1(n252), .A2(n251), .ZN(n253) );
  MUX2_X1 U281 ( .A(n361), .B(n253), .S(n229), .Z(n397) );
  NAND2_X1 U282 ( .A1(n255), .A2(n254), .ZN(n256) );
  MUX2_X1 U283 ( .A(n363), .B(n256), .S(n340), .Z(n401) );
  INV_X1 U284 ( .A(n257), .ZN(n258) );
  AOI21_X1 U285 ( .B1(n260), .B2(n259), .A(n258), .ZN(n261) );
  MUX2_X1 U286 ( .A(n364), .B(n261), .S(n340), .Z(n403) );
  NAND2_X1 U287 ( .A1(n263), .A2(n262), .ZN(n264) );
  NAND2_X1 U288 ( .A1(n264), .A2(n340), .ZN(n266) );
  NAND2_X1 U289 ( .A1(n274), .A2(n353), .ZN(n265) );
  NAND2_X1 U290 ( .A1(n266), .A2(n265), .ZN(n381) );
  NAND2_X1 U291 ( .A1(n268), .A2(n267), .ZN(n269) );
  MUX2_X1 U292 ( .A(n269), .B(n355), .S(n274), .Z(n385) );
  INV_X1 U293 ( .A(n119), .ZN(n274) );
  OR2_X1 U294 ( .A1(n119), .A2(n405), .ZN(n270) );
  OAI21_X1 U295 ( .B1(n271), .B2(n274), .A(n270), .ZN(n272) );
  INV_X1 U296 ( .A(n272), .ZN(n273) );
  OAI21_X1 U297 ( .B1(n275), .B2(n274), .A(n273), .ZN(n395) );
  MUX2_X1 U298 ( .A(product[0]), .B(n529), .S(n340), .Z(n419) );
  MUX2_X1 U299 ( .A(n529), .B(n530), .S(n119), .Z(n421) );
  AND2_X1 U300 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n276) );
  MUX2_X1 U301 ( .A(n530), .B(n276), .S(n340), .Z(n423) );
  MUX2_X1 U302 ( .A(product[1]), .B(n532), .S(n340), .Z(n425) );
  MUX2_X1 U303 ( .A(n532), .B(n533), .S(n229), .Z(n427) );
  OR2_X1 U304 ( .A1(n278), .A2(n277), .ZN(n279) );
  AND2_X1 U305 ( .A1(n279), .A2(n284), .ZN(n280) );
  MUX2_X1 U306 ( .A(n533), .B(n280), .S(n340), .Z(n429) );
  MUX2_X1 U307 ( .A(product[2]), .B(n535), .S(n340), .Z(n431) );
  MUX2_X1 U308 ( .A(n535), .B(n536), .S(n340), .Z(n433) );
  INV_X1 U309 ( .A(n281), .ZN(n283) );
  NAND2_X1 U310 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U311 ( .A(n285), .B(n284), .Z(n286) );
  MUX2_X1 U312 ( .A(n536), .B(n286), .S(n340), .Z(n435) );
  MUX2_X1 U313 ( .A(product[3]), .B(n538), .S(n340), .Z(n437) );
  MUX2_X1 U314 ( .A(n538), .B(n539), .S(n340), .Z(n439) );
  NAND2_X1 U315 ( .A1(n288), .A2(n287), .ZN(n290) );
  XNOR2_X1 U316 ( .A(n290), .B(n289), .ZN(n291) );
  MUX2_X1 U317 ( .A(n539), .B(n291), .S(n340), .Z(n441) );
  MUX2_X1 U318 ( .A(product[4]), .B(n541), .S(n340), .Z(n443) );
  MUX2_X1 U319 ( .A(n541), .B(n542), .S(n229), .Z(n445) );
  INV_X1 U320 ( .A(n292), .ZN(n294) );
  NAND2_X1 U321 ( .A1(n294), .A2(n293), .ZN(n296) );
  XOR2_X1 U322 ( .A(n296), .B(n295), .Z(n297) );
  MUX2_X1 U323 ( .A(n542), .B(n297), .S(n229), .Z(n447) );
  MUX2_X1 U324 ( .A(product[5]), .B(n544), .S(n229), .Z(n449) );
  MUX2_X1 U325 ( .A(n544), .B(n545), .S(n340), .Z(n451) );
  MUX2_X1 U326 ( .A(product[6]), .B(n547), .S(n229), .Z(n455) );
  NAND2_X1 U327 ( .A1(n410), .A2(n358), .ZN(n298) );
  XOR2_X1 U328 ( .A(n298), .B(n364), .Z(n299) );
  MUX2_X1 U329 ( .A(n547), .B(n299), .S(n340), .Z(n457) );
  MUX2_X1 U330 ( .A(product[7]), .B(n549), .S(n119), .Z(n459) );
  OAI21_X1 U331 ( .B1(n357), .B2(n364), .A(n358), .ZN(n302) );
  NAND2_X1 U332 ( .A1(n348), .A2(n356), .ZN(n300) );
  XNOR2_X1 U333 ( .A(n302), .B(n300), .ZN(n301) );
  MUX2_X1 U334 ( .A(n549), .B(n301), .S(n340), .Z(n461) );
  BUF_X4 U335 ( .A(en), .Z(n340) );
  MUX2_X1 U336 ( .A(product[8]), .B(n551), .S(n340), .Z(n463) );
  AOI21_X1 U337 ( .B1(n302), .B2(n348), .A(n412), .ZN(n305) );
  NAND2_X1 U338 ( .A1(n413), .A2(n355), .ZN(n303) );
  XOR2_X1 U339 ( .A(n305), .B(n303), .Z(n304) );
  MUX2_X1 U340 ( .A(n551), .B(n304), .S(n340), .Z(n465) );
  MUX2_X1 U341 ( .A(product[9]), .B(n553), .S(n340), .Z(n467) );
  OAI21_X1 U342 ( .B1(n305), .B2(n354), .A(n355), .ZN(n313) );
  INV_X1 U343 ( .A(n313), .ZN(n308) );
  NAND2_X1 U344 ( .A1(n414), .A2(n353), .ZN(n306) );
  XOR2_X1 U345 ( .A(n308), .B(n306), .Z(n307) );
  MUX2_X1 U346 ( .A(n553), .B(n307), .S(n340), .Z(n469) );
  MUX2_X1 U347 ( .A(product[10]), .B(n555), .S(n340), .Z(n471) );
  OAI21_X1 U348 ( .B1(n308), .B2(n352), .A(n353), .ZN(n310) );
  NAND2_X1 U349 ( .A1(n406), .A2(n360), .ZN(n309) );
  XNOR2_X1 U350 ( .A(n310), .B(n309), .ZN(n311) );
  MUX2_X1 U351 ( .A(n555), .B(n311), .S(n340), .Z(n473) );
  MUX2_X1 U352 ( .A(product[11]), .B(n557), .S(n340), .Z(n475) );
  NOR2_X1 U353 ( .A1(n359), .A2(n352), .ZN(n314) );
  OAI21_X1 U354 ( .B1(n359), .B2(n353), .A(n360), .ZN(n312) );
  AOI21_X1 U355 ( .B1(n314), .B2(n313), .A(n312), .ZN(n336) );
  NAND2_X1 U356 ( .A1(n415), .A2(n351), .ZN(n315) );
  XOR2_X1 U357 ( .A(n336), .B(n315), .Z(n316) );
  MUX2_X1 U358 ( .A(n557), .B(n316), .S(n340), .Z(n477) );
  MUX2_X1 U359 ( .A(product[12]), .B(n559), .S(n340), .Z(n479) );
  OAI21_X1 U360 ( .B1(n336), .B2(n362), .A(n351), .ZN(n318) );
  NAND2_X1 U361 ( .A1(n347), .A2(n363), .ZN(n317) );
  XNOR2_X1 U362 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U363 ( .A(n559), .B(n319), .S(n340), .Z(n481) );
  MUX2_X1 U364 ( .A(product[13]), .B(n561), .S(n340), .Z(n483) );
  NAND2_X1 U365 ( .A1(n415), .A2(n347), .ZN(n321) );
  AOI21_X1 U366 ( .B1(n408), .B2(n347), .A(n416), .ZN(n320) );
  OAI21_X1 U367 ( .B1(n336), .B2(n321), .A(n320), .ZN(n323) );
  NAND2_X1 U368 ( .A1(n346), .A2(n361), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n324) );
  MUX2_X1 U370 ( .A(n561), .B(n324), .S(n340), .Z(n485) );
  MUX2_X1 U371 ( .A(product[14]), .B(n563), .S(n340), .Z(n487) );
  NAND2_X1 U372 ( .A1(n347), .A2(n346), .ZN(n331) );
  OR2_X1 U373 ( .A1(n362), .A2(n331), .ZN(n327) );
  AOI21_X1 U374 ( .B1(n416), .B2(n346), .A(n411), .ZN(n325) );
  OAI21_X1 U375 ( .B1(n331), .B2(n351), .A(n325), .ZN(n333) );
  INV_X1 U376 ( .A(n333), .ZN(n326) );
  OAI21_X1 U377 ( .B1(n336), .B2(n327), .A(n326), .ZN(n329) );
  NAND2_X1 U378 ( .A1(n345), .A2(n350), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  MUX2_X1 U380 ( .A(n563), .B(n330), .S(n340), .Z(n489) );
  MUX2_X1 U381 ( .A(product[15]), .B(n565), .S(n340), .Z(n491) );
  NOR2_X1 U382 ( .A1(n331), .A2(n409), .ZN(n332) );
  NAND2_X1 U383 ( .A1(n415), .A2(n332), .ZN(n335) );
  AOI21_X1 U384 ( .B1(n333), .B2(n345), .A(n407), .ZN(n334) );
  OAI21_X1 U385 ( .B1(n336), .B2(n335), .A(n334), .ZN(n337) );
  XNOR2_X1 U386 ( .A(n337), .B(n349), .ZN(n338) );
  MUX2_X1 U387 ( .A(n565), .B(n338), .S(n340), .Z(n493) );
  MUX2_X1 U388 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n340), .Z(n495) );
  MUX2_X1 U389 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n340), .Z(n497) );
  MUX2_X1 U390 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n340), .Z(n499) );
  MUX2_X1 U391 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n340), .Z(n501) );
  MUX2_X1 U392 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n340), .Z(n503) );
  MUX2_X1 U393 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n340), .Z(n505) );
  MUX2_X1 U394 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n340), .Z(n507) );
  MUX2_X1 U395 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n340), .Z(n509) );
  MUX2_X1 U396 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n340), .Z(n511) );
  MUX2_X1 U397 ( .A(n9), .B(A_extended[1]), .S(n340), .Z(n513) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n340), .Z(n515) );
  MUX2_X1 U399 ( .A(n15), .B(A_extended[3]), .S(n340), .Z(n517) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n340), .Z(n519) );
  MUX2_X1 U401 ( .A(n16), .B(A_extended[5]), .S(n340), .Z(n521) );
  MUX2_X1 U402 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n340), .Z(n523) );
  MUX2_X1 U403 ( .A(n339), .B(A_extended[7]), .S(n340), .Z(n525) );
  OR2_X1 U404 ( .A1(n340), .A2(n567), .ZN(n527) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_3 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n311 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n357, n359, n361, n363, n365, n367, n369, n371, n373, n375,
         n377, n379, n381, n383, n385, n387, n389, n391, n393, n395, n397,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n410,
         n412, n414, n416, n418, n420, n422, n424, n426, n428, n430, n432,
         n434, n436, n438, n440, n442, n444, n446, n448, n450, n452, n454,
         n456, n458, n460, n462, n464, n466, n468, n470, n472, n474, n476,
         n478, n480, n482, n484, n486, n488, n490, n492, n494, n496, n498,
         n500, n502, n504, n506, n508, n510, n512, n514, n516, n518, n519,
         n521, n522, n524, n525, n527, n528, n530, n531, n533, n535, n537,
         n539, n541, n543, n545, n547, n549, n551, n553, n554, n555, n556,
         n557, n558;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n407), .SE(n516), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n408), .SE(n514), .CK(clk), .Q(n556), 
        .QN(n28) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n408), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n30) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n407), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n331) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n408), .SE(n506), .CK(clk), .Q(n555), 
        .QN(n330) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n407), .SE(n504), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n29) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n408), .SE(n502), .CK(clk), .Q(n554), 
        .QN(n31) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n407), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n19) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n407), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n21) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n407), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n24) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n407), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n407), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n25) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n407), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n27) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n407), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n22) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n408), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n23) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n407), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n407), .SE(n482), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n408), .SE(n480), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n407), .SE(n478), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n407), .SE(n476), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n408), .SE(n474), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n407), .SE(n472), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n407), .SE(n470), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n408), .SE(n468), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n407), .SE(n466), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n407), .SE(n464), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n408), .SE(n462), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n407), .SE(n460), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n407), .SE(n458), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n408), .SE(n456), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n407), .SE(n454), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n408), .SE(n452), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n408), .SE(n450), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n408), .SE(n448), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n408), .SE(n446), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n408), .SE(n444), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n408), .SE(n442), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n408), .SE(n440), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n408), .SE(n438), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n408), .SE(n436), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n408), .SE(n434), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n408), .SE(n432), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n407), .SE(n430), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n407), .SE(n428), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n407), .SE(n426), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n407), .SE(n424), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n407), .SE(n422), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n407), .SE(n420), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n407), .SE(n418), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n407), .SE(n416), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n407), .SE(n414), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n407), .SE(n412), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n407), .SE(n410), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n558), .SE(n397), .CK(
        clk), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2_IP  ( .D(1'b1), .SI(n558), .SE(n395), .CK(
        clk), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n558), .SE(n393), .CK(
        clk), .QN(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n558), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n558), .SE(n389), .CK(
        clk), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n558), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n558), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n558), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n347), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n558), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n346), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n558), .SE(n379), .CK(
        clk), .Q(n33), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n558), .SE(n377), .CK(
        clk), .Q(n405), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n558), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n558), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n558), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n341), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n558), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n340), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n558), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n558), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n338), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n558), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n337), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n558), .SE(n361), .CK(
        clk), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n558), .SE(n359), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n558), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n334), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n558), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n333) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n407), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n332) );
  BUF_X2 U2 ( .A(en), .Z(n279) );
  BUF_X2 U3 ( .A(en), .Z(n329) );
  NAND2_X1 U4 ( .A1(n34), .A2(n35), .ZN(n210) );
  INV_X1 U5 ( .A(n36), .ZN(n212) );
  NAND2_X1 U6 ( .A1(n7), .A2(n5), .ZN(n383) );
  NAND2_X1 U7 ( .A1(n6), .A2(n347), .ZN(n5) );
  INV_X1 U8 ( .A(n16), .ZN(n6) );
  NAND2_X1 U9 ( .A1(n8), .A2(n16), .ZN(n7) );
  NAND2_X1 U10 ( .A1(n251), .A2(n250), .ZN(n8) );
  XNOR2_X2 U11 ( .A(n332), .B(n30), .ZN(n164) );
  CLKBUF_X2 U12 ( .A(rst_n), .Z(n407) );
  CLKBUF_X2 U13 ( .A(n554), .Z(n326) );
  BUF_X1 U14 ( .A(n555), .Z(n14) );
  BUF_X1 U15 ( .A(\mult_x_1/n311 ), .Z(n15) );
  INV_X1 U16 ( .A(n14), .ZN(n9) );
  INV_X1 U17 ( .A(n184), .ZN(n189) );
  NOR2_X1 U18 ( .A1(n186), .A2(n185), .ZN(n188) );
  NAND2_X1 U19 ( .A1(n186), .A2(n185), .ZN(n187) );
  OR2_X1 U20 ( .A1(n59), .A2(n58), .ZN(n186) );
  INV_X1 U21 ( .A(n329), .ZN(n47) );
  XNOR2_X1 U22 ( .A(n64), .B(n184), .ZN(n233) );
  XNOR2_X1 U23 ( .A(n185), .B(n186), .ZN(n64) );
  NAND2_X1 U24 ( .A1(n242), .A2(n241), .ZN(n243) );
  INV_X1 U25 ( .A(n245), .ZN(n241) );
  INV_X1 U26 ( .A(n246), .ZN(n242) );
  OAI22_X1 U27 ( .A1(n174), .A2(n55), .B1(n176), .B2(n69), .ZN(n58) );
  CLKBUF_X1 U28 ( .A(n555), .Z(n327) );
  OAI21_X1 U29 ( .B1(n189), .B2(n188), .A(n187), .ZN(n231) );
  NAND2_X1 U30 ( .A1(n46), .A2(n329), .ZN(n49) );
  NAND2_X1 U31 ( .A1(n47), .A2(n343), .ZN(n48) );
  NAND2_X1 U32 ( .A1(n236), .A2(n235), .ZN(n237) );
  NAND2_X1 U33 ( .A1(n20), .A2(n234), .ZN(n235) );
  OAI21_X1 U34 ( .B1(n20), .B2(n234), .A(n233), .ZN(n236) );
  NAND2_X1 U35 ( .A1(n248), .A2(n247), .ZN(n249) );
  NAND2_X1 U36 ( .A1(n246), .A2(n245), .ZN(n247) );
  NAND2_X1 U37 ( .A1(n244), .A2(n243), .ZN(n248) );
  NAND2_X1 U38 ( .A1(n13), .A2(n50), .ZN(n10) );
  NAND2_X1 U39 ( .A1(n13), .A2(n50), .ZN(n11) );
  NAND2_X1 U40 ( .A1(n13), .A2(n50), .ZN(n166) );
  XNOR2_X1 U41 ( .A(n330), .B(n331), .ZN(n12) );
  XNOR2_X1 U42 ( .A(n244), .B(n136), .ZN(n142) );
  XNOR2_X1 U43 ( .A(n332), .B(n30), .ZN(n13) );
  XNOR2_X1 U44 ( .A(n246), .B(n245), .ZN(n136) );
  BUF_X4 U45 ( .A(en), .Z(n16) );
  INV_X1 U46 ( .A(n169), .ZN(n17) );
  OAI22_X1 U47 ( .A1(n174), .A2(n85), .B1(n176), .B2(n173), .ZN(n18) );
  BUF_X1 U48 ( .A(rst_n), .Z(n408) );
  INV_X1 U49 ( .A(rst_n), .ZN(n558) );
  AND2_X1 U50 ( .A1(n75), .A2(n74), .ZN(n20) );
  XOR2_X1 U51 ( .A(n75), .B(n74), .Z(n32) );
  XNOR2_X1 U52 ( .A(n327), .B(n29), .ZN(n34) );
  XNOR2_X1 U53 ( .A(n554), .B(\mult_x_1/a[2] ), .ZN(n35) );
  XNOR2_X1 U54 ( .A(n14), .B(\mult_x_1/n286 ), .ZN(n43) );
  INV_X1 U55 ( .A(n35), .ZN(n36) );
  XNOR2_X1 U56 ( .A(n14), .B(\mult_x_1/n285 ), .ZN(n93) );
  OAI22_X1 U57 ( .A1(n210), .A2(n43), .B1(n212), .B2(n93), .ZN(n152) );
  NAND2_X1 U58 ( .A1(n326), .A2(n19), .ZN(n215) );
  XNOR2_X1 U59 ( .A(n326), .B(\mult_x_1/n284 ), .ZN(n42) );
  XNOR2_X1 U60 ( .A(n326), .B(\mult_x_1/n283 ), .ZN(n91) );
  OAI22_X1 U61 ( .A1(n215), .A2(n42), .B1(n91), .B2(n19), .ZN(n151) );
  XOR2_X1 U62 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n37) );
  XNOR2_X1 U63 ( .A(n330), .B(n331), .ZN(n38) );
  NAND2_X2 U64 ( .A1(n37), .A2(n12), .ZN(n176) );
  OR2_X1 U65 ( .A1(\mult_x_1/n288 ), .A2(n332), .ZN(n40) );
  INV_X1 U66 ( .A(n38), .ZN(n39) );
  INV_X2 U67 ( .A(n39), .ZN(n174) );
  OAI22_X1 U68 ( .A1(n176), .A2(n332), .B1(n40), .B2(n174), .ZN(n103) );
  XNOR2_X1 U69 ( .A(n15), .B(\mult_x_1/n288 ), .ZN(n41) );
  XNOR2_X1 U70 ( .A(n15), .B(\mult_x_1/n287 ), .ZN(n105) );
  OAI22_X1 U71 ( .A1(n176), .A2(n41), .B1(n174), .B2(n105), .ZN(n102) );
  XNOR2_X1 U72 ( .A(n326), .B(\mult_x_1/n285 ), .ZN(n206) );
  OAI22_X1 U73 ( .A1(n215), .A2(n206), .B1(n42), .B2(n19), .ZN(n203) );
  AND2_X1 U74 ( .A1(\mult_x_1/n288 ), .A2(n39), .ZN(n202) );
  XNOR2_X1 U75 ( .A(n14), .B(\mult_x_1/n287 ), .ZN(n204) );
  OAI22_X1 U76 ( .A1(n210), .A2(n204), .B1(n212), .B2(n43), .ZN(n201) );
  OR2_X1 U77 ( .A1(n45), .A2(n44), .ZN(n226) );
  NAND2_X1 U78 ( .A1(n45), .A2(n44), .ZN(n224) );
  NAND2_X1 U79 ( .A1(n226), .A2(n224), .ZN(n46) );
  NAND2_X1 U80 ( .A1(n49), .A2(n48), .ZN(n375) );
  XNOR2_X1 U81 ( .A(n15), .B(\mult_x_1/n283 ), .ZN(n55) );
  XNOR2_X1 U82 ( .A(n15), .B(\mult_x_1/n284 ), .ZN(n69) );
  XNOR2_X1 U83 ( .A(n14), .B(\mult_x_1/n282 ), .ZN(n70) );
  XNOR2_X1 U84 ( .A(n14), .B(\mult_x_1/n281 ), .ZN(n56) );
  OAI22_X1 U85 ( .A1(n210), .A2(n70), .B1(n212), .B2(n56), .ZN(n59) );
  XNOR2_X1 U86 ( .A(n58), .B(n59), .ZN(n75) );
  BUF_X4 U87 ( .A(n556), .Z(n328) );
  XNOR2_X1 U88 ( .A(n328), .B(n30), .ZN(n50) );
  XNOR2_X1 U89 ( .A(n328), .B(\mult_x_1/n287 ), .ZN(n71) );
  XNOR2_X1 U90 ( .A(n328), .B(\mult_x_1/n286 ), .ZN(n63) );
  OAI22_X1 U91 ( .A1(n166), .A2(n71), .B1(n13), .B2(n63), .ZN(n132) );
  XNOR2_X1 U92 ( .A(n326), .B(\mult_x_1/n281 ), .ZN(n98) );
  AND2_X1 U93 ( .A1(n557), .A2(\mult_x_1/n281 ), .ZN(n83) );
  XNOR2_X1 U94 ( .A(n83), .B(n326), .ZN(n60) );
  OAI22_X1 U95 ( .A1(n215), .A2(n98), .B1(n60), .B2(n19), .ZN(n131) );
  AND2_X1 U96 ( .A1(n557), .A2(n328), .ZN(n51) );
  XNOR2_X1 U97 ( .A(n51), .B(n328), .ZN(n57) );
  INV_X1 U98 ( .A(n57), .ZN(n52) );
  AND2_X1 U99 ( .A1(\mult_x_1/n288 ), .A2(n52), .ZN(n130) );
  XNOR2_X1 U100 ( .A(n328), .B(\mult_x_1/n285 ), .ZN(n62) );
  XNOR2_X1 U101 ( .A(n328), .B(\mult_x_1/n284 ), .ZN(n165) );
  OAI22_X1 U102 ( .A1(n166), .A2(n62), .B1(n164), .B2(n165), .ZN(n171) );
  XNOR2_X1 U103 ( .A(n15), .B(\mult_x_1/n282 ), .ZN(n175) );
  OAI22_X1 U104 ( .A1(n176), .A2(n55), .B1(n174), .B2(n175), .ZN(n170) );
  XNOR2_X1 U105 ( .A(n83), .B(n14), .ZN(n167) );
  OAI22_X1 U106 ( .A1(n210), .A2(n56), .B1(n167), .B2(n212), .ZN(n190) );
  INV_X1 U107 ( .A(n190), .ZN(n169) );
  XNOR2_X1 U108 ( .A(n20), .B(n234), .ZN(n65) );
  BUF_X2 U109 ( .A(n57), .Z(n172) );
  NOR2_X1 U110 ( .A1(n22), .A2(n172), .ZN(n185) );
  AOI21_X1 U111 ( .B1(n215), .B2(n19), .A(n60), .ZN(n61) );
  INV_X1 U112 ( .A(n61), .ZN(n68) );
  OAI22_X1 U113 ( .A1(n10), .A2(n63), .B1(n164), .B2(n62), .ZN(n67) );
  NOR2_X1 U114 ( .A1(n23), .A2(n172), .ZN(n66) );
  XNOR2_X1 U115 ( .A(n65), .B(n233), .ZN(n78) );
  FA_X1 U116 ( .A(n68), .B(n67), .CI(n66), .CO(n184), .S(n239) );
  XNOR2_X1 U117 ( .A(n15), .B(\mult_x_1/n285 ), .ZN(n97) );
  OAI22_X1 U118 ( .A1(n176), .A2(n97), .B1(n174), .B2(n69), .ZN(n129) );
  XNOR2_X1 U119 ( .A(n14), .B(\mult_x_1/n283 ), .ZN(n100) );
  OAI22_X1 U120 ( .A1(n210), .A2(n100), .B1(n212), .B2(n70), .ZN(n128) );
  XNOR2_X1 U121 ( .A(n328), .B(\mult_x_1/n288 ), .ZN(n72) );
  OAI22_X1 U122 ( .A1(n11), .A2(n72), .B1(n164), .B2(n71), .ZN(n96) );
  OR2_X1 U123 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n73) );
  OAI22_X1 U124 ( .A1(n164), .A2(n73), .B1(n11), .B2(n28), .ZN(n94) );
  AND2_X1 U125 ( .A1(n96), .A2(n94), .ZN(n127) );
  NOR2_X1 U126 ( .A1(n78), .A2(n77), .ZN(n76) );
  MUX2_X1 U127 ( .A(n344), .B(n76), .S(n279), .Z(n377) );
  NAND2_X1 U128 ( .A1(n78), .A2(n77), .ZN(n79) );
  NAND2_X1 U129 ( .A1(n79), .A2(n279), .ZN(n81) );
  OR2_X1 U130 ( .A1(n279), .A2(n33), .ZN(n80) );
  NAND2_X1 U131 ( .A1(n81), .A2(n80), .ZN(n379) );
  NOR2_X1 U154 ( .A1(n24), .A2(n172), .ZN(n112) );
  XNOR2_X1 U155 ( .A(n328), .B(\mult_x_1/n281 ), .ZN(n82) );
  XNOR2_X1 U156 ( .A(n83), .B(n328), .ZN(n113) );
  OAI22_X1 U157 ( .A1(n11), .A2(n82), .B1(n113), .B2(n164), .ZN(n118) );
  INV_X1 U158 ( .A(n118), .ZN(n111) );
  XNOR2_X1 U159 ( .A(n328), .B(\mult_x_1/n282 ), .ZN(n86) );
  OAI22_X1 U160 ( .A1(n10), .A2(n86), .B1(n164), .B2(n82), .ZN(n89) );
  XNOR2_X1 U161 ( .A(n83), .B(\mult_x_1/n311 ), .ZN(n85) );
  AOI21_X1 U162 ( .B1(n174), .B2(n176), .A(n85), .ZN(n84) );
  INV_X1 U163 ( .A(n84), .ZN(n88) );
  XNOR2_X1 U164 ( .A(n15), .B(\mult_x_1/n281 ), .ZN(n173) );
  OAI22_X1 U165 ( .A1(n174), .A2(n85), .B1(n176), .B2(n173), .ZN(n87) );
  XNOR2_X1 U166 ( .A(n328), .B(\mult_x_1/n283 ), .ZN(n163) );
  OAI22_X1 U167 ( .A1(n11), .A2(n163), .B1(n164), .B2(n86), .ZN(n162) );
  INV_X1 U168 ( .A(n87), .ZN(n161) );
  NOR2_X1 U169 ( .A1(n25), .A2(n172), .ZN(n160) );
  NOR2_X1 U170 ( .A1(n26), .A2(n172), .ZN(n158) );
  FA_X1 U171 ( .A(n89), .B(n88), .CI(n18), .CO(n110), .S(n157) );
  OR2_X1 U172 ( .A1(n125), .A2(n124), .ZN(n90) );
  MUX2_X1 U173 ( .A(n333), .B(n90), .S(n16), .Z(n355) );
  XNOR2_X1 U174 ( .A(n326), .B(\mult_x_1/n282 ), .ZN(n99) );
  OAI22_X1 U175 ( .A1(n215), .A2(n91), .B1(n99), .B2(n19), .ZN(n108) );
  INV_X1 U176 ( .A(n164), .ZN(n92) );
  AND2_X1 U177 ( .A1(\mult_x_1/n288 ), .A2(n92), .ZN(n107) );
  XNOR2_X1 U178 ( .A(n14), .B(\mult_x_1/n284 ), .ZN(n101) );
  OAI22_X1 U179 ( .A1(n210), .A2(n93), .B1(n212), .B2(n101), .ZN(n106) );
  INV_X1 U180 ( .A(n94), .ZN(n95) );
  XNOR2_X1 U181 ( .A(n96), .B(n95), .ZN(n138) );
  XNOR2_X1 U182 ( .A(n15), .B(\mult_x_1/n286 ), .ZN(n104) );
  OAI22_X1 U183 ( .A1(n176), .A2(n104), .B1(n174), .B2(n97), .ZN(n135) );
  OAI22_X1 U184 ( .A1(n215), .A2(n99), .B1(n98), .B2(n19), .ZN(n134) );
  OAI22_X1 U185 ( .A1(n210), .A2(n101), .B1(n212), .B2(n100), .ZN(n133) );
  HA_X1 U186 ( .A(n103), .B(n102), .CO(n149), .S(n150) );
  OAI22_X1 U187 ( .A1(n176), .A2(n105), .B1(n174), .B2(n104), .ZN(n148) );
  FA_X1 U188 ( .A(n108), .B(n107), .CI(n106), .CO(n139), .S(n147) );
  OR2_X1 U189 ( .A1(n145), .A2(n144), .ZN(n109) );
  MUX2_X1 U190 ( .A(n335), .B(n109), .S(n16), .Z(n359) );
  FA_X1 U191 ( .A(n112), .B(n111), .CI(n110), .CO(n120), .S(n125) );
  AOI21_X1 U192 ( .B1(n164), .B2(n10), .A(n113), .ZN(n114) );
  INV_X1 U193 ( .A(n114), .ZN(n116) );
  NOR2_X1 U194 ( .A1(n21), .A2(n172), .ZN(n115) );
  XOR2_X1 U195 ( .A(n116), .B(n115), .Z(n117) );
  XOR2_X1 U196 ( .A(n118), .B(n117), .Z(n119) );
  OR2_X1 U197 ( .A1(n120), .A2(n119), .ZN(n122) );
  NAND2_X1 U198 ( .A1(n120), .A2(n119), .ZN(n121) );
  NAND2_X1 U199 ( .A1(n122), .A2(n121), .ZN(n123) );
  MUX2_X1 U200 ( .A(n336), .B(n123), .S(n16), .Z(n361) );
  NAND2_X1 U201 ( .A1(n125), .A2(n124), .ZN(n126) );
  MUX2_X1 U202 ( .A(n337), .B(n126), .S(n16), .Z(n363) );
  FA_X1 U203 ( .A(n129), .B(n128), .CI(n127), .CO(n238), .S(n244) );
  FA_X1 U204 ( .A(n132), .B(n131), .CI(n130), .CO(n74), .S(n246) );
  FA_X1 U205 ( .A(n135), .B(n134), .CI(n133), .CO(n245), .S(n137) );
  FA_X1 U206 ( .A(n139), .B(n138), .CI(n137), .CO(n141), .S(n145) );
  NOR2_X1 U207 ( .A1(n142), .A2(n141), .ZN(n140) );
  MUX2_X1 U208 ( .A(n338), .B(n140), .S(n16), .Z(n365) );
  NAND2_X1 U209 ( .A1(n142), .A2(n141), .ZN(n143) );
  MUX2_X1 U210 ( .A(n339), .B(n143), .S(n16), .Z(n367) );
  NAND2_X1 U211 ( .A1(n145), .A2(n144), .ZN(n146) );
  MUX2_X1 U212 ( .A(n340), .B(n146), .S(n16), .Z(n369) );
  FA_X1 U213 ( .A(n149), .B(n148), .CI(n147), .CO(n144), .S(n155) );
  FA_X1 U214 ( .A(n152), .B(n151), .CI(n150), .CO(n154), .S(n45) );
  NOR2_X1 U215 ( .A1(n155), .A2(n154), .ZN(n153) );
  MUX2_X1 U216 ( .A(n341), .B(n153), .S(n16), .Z(n371) );
  NAND2_X1 U217 ( .A1(n155), .A2(n154), .ZN(n156) );
  MUX2_X1 U218 ( .A(n342), .B(n156), .S(n16), .Z(n373) );
  FA_X1 U219 ( .A(n159), .B(n158), .CI(n157), .CO(n124), .S(n199) );
  FA_X1 U220 ( .A(n162), .B(n161), .CI(n160), .CO(n159), .S(n183) );
  OAI22_X1 U221 ( .A1(n10), .A2(n165), .B1(n164), .B2(n163), .ZN(n192) );
  AOI21_X1 U222 ( .B1(n212), .B2(n210), .A(n167), .ZN(n168) );
  INV_X1 U223 ( .A(n168), .ZN(n191) );
  FA_X1 U224 ( .A(n170), .B(n171), .CI(n169), .CO(n196), .S(n234) );
  INV_X1 U225 ( .A(n196), .ZN(n179) );
  NOR2_X1 U226 ( .A1(n27), .A2(n172), .ZN(n194) );
  OAI22_X1 U227 ( .A1(n176), .A2(n175), .B1(n174), .B2(n173), .ZN(n193) );
  NOR2_X1 U228 ( .A1(n194), .A2(n193), .ZN(n178) );
  NAND2_X1 U229 ( .A1(n194), .A2(n193), .ZN(n177) );
  OAI21_X1 U230 ( .B1(n179), .B2(n178), .A(n177), .ZN(n181) );
  NAND2_X1 U231 ( .A1(n199), .A2(n198), .ZN(n180) );
  MUX2_X1 U232 ( .A(n346), .B(n180), .S(n329), .Z(n381) );
  FA_X1 U233 ( .A(n183), .B(n182), .CI(n181), .CO(n198), .S(n251) );
  FA_X1 U234 ( .A(n192), .B(n191), .CI(n17), .CO(n182), .S(n230) );
  XOR2_X1 U235 ( .A(n194), .B(n193), .Z(n195) );
  XOR2_X1 U236 ( .A(n196), .B(n195), .Z(n229) );
  OR2_X1 U237 ( .A1(n199), .A2(n198), .ZN(n200) );
  MUX2_X1 U238 ( .A(n348), .B(n200), .S(n16), .Z(n385) );
  FA_X1 U239 ( .A(n203), .B(n202), .CI(n201), .CO(n44), .S(n223) );
  XNOR2_X1 U240 ( .A(n14), .B(\mult_x_1/n288 ), .ZN(n205) );
  OAI22_X1 U241 ( .A1(n210), .A2(n205), .B1(n212), .B2(n204), .ZN(n208) );
  XNOR2_X1 U242 ( .A(n326), .B(\mult_x_1/n286 ), .ZN(n211) );
  OAI22_X1 U243 ( .A1(n215), .A2(n211), .B1(n206), .B2(n19), .ZN(n207) );
  NOR2_X1 U244 ( .A1(n223), .A2(n222), .ZN(n270) );
  HA_X1 U245 ( .A(n208), .B(n207), .CO(n222), .S(n220) );
  OR2_X1 U246 ( .A1(\mult_x_1/n288 ), .A2(n330), .ZN(n209) );
  OAI22_X1 U247 ( .A1(n210), .A2(n9), .B1(n209), .B2(n212), .ZN(n219) );
  OR2_X1 U248 ( .A1(n220), .A2(n219), .ZN(n266) );
  XNOR2_X1 U249 ( .A(n326), .B(\mult_x_1/n287 ), .ZN(n214) );
  OAI22_X1 U250 ( .A1(n215), .A2(n214), .B1(n211), .B2(n19), .ZN(n218) );
  INV_X1 U251 ( .A(n212), .ZN(n213) );
  AND2_X1 U252 ( .A1(\mult_x_1/n288 ), .A2(n213), .ZN(n217) );
  NOR2_X1 U253 ( .A1(n218), .A2(n217), .ZN(n259) );
  OAI22_X1 U254 ( .A1(n215), .A2(\mult_x_1/n288 ), .B1(n214), .B2(n19), .ZN(
        n256) );
  OR2_X1 U255 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n216) );
  NAND2_X1 U256 ( .A1(n216), .A2(n215), .ZN(n255) );
  NAND2_X1 U257 ( .A1(n256), .A2(n255), .ZN(n262) );
  NAND2_X1 U258 ( .A1(n218), .A2(n217), .ZN(n260) );
  OAI21_X1 U259 ( .B1(n259), .B2(n262), .A(n260), .ZN(n267) );
  NAND2_X1 U260 ( .A1(n220), .A2(n219), .ZN(n265) );
  INV_X1 U261 ( .A(n265), .ZN(n221) );
  AOI21_X1 U262 ( .B1(n266), .B2(n267), .A(n221), .ZN(n273) );
  NAND2_X1 U263 ( .A1(n223), .A2(n222), .ZN(n271) );
  OAI21_X1 U264 ( .B1(n270), .B2(n273), .A(n271), .ZN(n228) );
  INV_X1 U265 ( .A(n224), .ZN(n225) );
  AOI21_X1 U266 ( .B1(n226), .B2(n228), .A(n225), .ZN(n227) );
  MUX2_X1 U267 ( .A(n349), .B(n227), .S(n329), .Z(n387) );
  MUX2_X1 U268 ( .A(n350), .B(n228), .S(n279), .Z(n389) );
  FA_X1 U269 ( .A(n231), .B(n230), .CI(n229), .CO(n250), .S(n232) );
  MUX2_X1 U270 ( .A(n351), .B(n232), .S(n16), .Z(n391) );
  MUX2_X1 U271 ( .A(n352), .B(n237), .S(n329), .Z(n393) );
  FA_X1 U272 ( .A(n239), .B(n238), .CI(n32), .CO(n77), .S(n240) );
  MUX2_X1 U273 ( .A(n353), .B(n240), .S(n279), .Z(n395) );
  MUX2_X1 U274 ( .A(n354), .B(n249), .S(n16), .Z(n397) );
  OAI21_X1 U275 ( .B1(n251), .B2(n250), .A(n329), .ZN(n253) );
  OR2_X1 U276 ( .A1(n16), .A2(n401), .ZN(n252) );
  NAND2_X1 U277 ( .A1(n253), .A2(n252), .ZN(n357) );
  MUX2_X1 U278 ( .A(product[0]), .B(n518), .S(n329), .Z(n410) );
  MUX2_X1 U279 ( .A(n518), .B(n519), .S(n279), .Z(n412) );
  AND2_X1 U280 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n254) );
  MUX2_X1 U281 ( .A(n519), .B(n254), .S(n16), .Z(n414) );
  MUX2_X1 U282 ( .A(product[1]), .B(n521), .S(n329), .Z(n416) );
  MUX2_X1 U283 ( .A(n521), .B(n522), .S(n279), .Z(n418) );
  OR2_X1 U284 ( .A1(n256), .A2(n255), .ZN(n257) );
  AND2_X1 U285 ( .A1(n257), .A2(n262), .ZN(n258) );
  MUX2_X1 U286 ( .A(n522), .B(n258), .S(n16), .Z(n420) );
  MUX2_X1 U287 ( .A(product[2]), .B(n524), .S(n329), .Z(n422) );
  MUX2_X1 U288 ( .A(n524), .B(n525), .S(n279), .Z(n424) );
  INV_X1 U289 ( .A(n259), .ZN(n261) );
  NAND2_X1 U290 ( .A1(n261), .A2(n260), .ZN(n263) );
  XOR2_X1 U291 ( .A(n263), .B(n262), .Z(n264) );
  MUX2_X1 U292 ( .A(n525), .B(n264), .S(n16), .Z(n426) );
  MUX2_X1 U293 ( .A(product[3]), .B(n527), .S(n329), .Z(n428) );
  MUX2_X1 U294 ( .A(n527), .B(n528), .S(n16), .Z(n430) );
  NAND2_X1 U295 ( .A1(n266), .A2(n265), .ZN(n268) );
  XNOR2_X1 U296 ( .A(n268), .B(n267), .ZN(n269) );
  MUX2_X1 U297 ( .A(n528), .B(n269), .S(n329), .Z(n432) );
  MUX2_X1 U298 ( .A(product[4]), .B(n530), .S(n329), .Z(n434) );
  MUX2_X1 U299 ( .A(n530), .B(n531), .S(n329), .Z(n436) );
  INV_X1 U300 ( .A(n270), .ZN(n272) );
  NAND2_X1 U301 ( .A1(n272), .A2(n271), .ZN(n274) );
  XOR2_X1 U302 ( .A(n274), .B(n273), .Z(n275) );
  MUX2_X1 U303 ( .A(n531), .B(n275), .S(n279), .Z(n438) );
  MUX2_X1 U304 ( .A(product[5]), .B(n533), .S(n329), .Z(n440) );
  XNOR2_X1 U305 ( .A(n343), .B(n350), .ZN(n276) );
  MUX2_X1 U306 ( .A(n533), .B(n276), .S(n279), .Z(n442) );
  MUX2_X1 U307 ( .A(product[6]), .B(n535), .S(n279), .Z(n444) );
  NAND2_X1 U308 ( .A1(n402), .A2(n342), .ZN(n277) );
  XOR2_X1 U309 ( .A(n277), .B(n349), .Z(n278) );
  MUX2_X1 U310 ( .A(n535), .B(n278), .S(n279), .Z(n446) );
  MUX2_X1 U311 ( .A(product[7]), .B(n537), .S(n16), .Z(n448) );
  OAI21_X1 U312 ( .B1(n341), .B2(n349), .A(n342), .ZN(n282) );
  NAND2_X1 U313 ( .A1(n335), .A2(n340), .ZN(n280) );
  XNOR2_X1 U314 ( .A(n282), .B(n280), .ZN(n281) );
  MUX2_X1 U315 ( .A(n537), .B(n281), .S(n16), .Z(n450) );
  MUX2_X1 U316 ( .A(product[8]), .B(n539), .S(n279), .Z(n452) );
  AOI21_X1 U317 ( .B1(n282), .B2(n335), .A(n403), .ZN(n285) );
  NAND2_X1 U318 ( .A1(n404), .A2(n339), .ZN(n283) );
  XOR2_X1 U319 ( .A(n285), .B(n283), .Z(n284) );
  MUX2_X1 U320 ( .A(n539), .B(n284), .S(n16), .Z(n454) );
  MUX2_X1 U321 ( .A(product[9]), .B(n541), .S(n329), .Z(n456) );
  OAI21_X1 U322 ( .B1(n285), .B2(n338), .A(n339), .ZN(n296) );
  INV_X1 U323 ( .A(n296), .ZN(n289) );
  NOR2_X1 U324 ( .A1(n353), .A2(n354), .ZN(n293) );
  INV_X1 U325 ( .A(n293), .ZN(n286) );
  NAND2_X1 U326 ( .A1(n353), .A2(n354), .ZN(n294) );
  NAND2_X1 U327 ( .A1(n286), .A2(n294), .ZN(n287) );
  XOR2_X1 U328 ( .A(n289), .B(n287), .Z(n288) );
  MUX2_X1 U329 ( .A(n541), .B(n288), .S(n279), .Z(n458) );
  MUX2_X1 U330 ( .A(product[10]), .B(n543), .S(n16), .Z(n460) );
  OAI21_X1 U331 ( .B1(n289), .B2(n293), .A(n294), .ZN(n291) );
  NAND2_X1 U332 ( .A1(n405), .A2(n345), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n292) );
  MUX2_X1 U334 ( .A(n543), .B(n292), .S(n329), .Z(n462) );
  MUX2_X1 U335 ( .A(product[11]), .B(n545), .S(n16), .Z(n464) );
  NOR2_X1 U336 ( .A1(n344), .A2(n293), .ZN(n297) );
  OAI21_X1 U337 ( .B1(n344), .B2(n294), .A(n345), .ZN(n295) );
  AOI21_X1 U338 ( .B1(n297), .B2(n296), .A(n295), .ZN(n323) );
  NOR2_X1 U339 ( .A1(n351), .A2(n352), .ZN(n310) );
  INV_X1 U340 ( .A(n310), .ZN(n303) );
  NAND2_X1 U341 ( .A1(n351), .A2(n352), .ZN(n312) );
  NAND2_X1 U342 ( .A1(n303), .A2(n312), .ZN(n298) );
  XOR2_X1 U343 ( .A(n323), .B(n298), .Z(n299) );
  MUX2_X1 U344 ( .A(n545), .B(n299), .S(n279), .Z(n466) );
  MUX2_X1 U345 ( .A(product[12]), .B(n547), .S(n16), .Z(n468) );
  OAI21_X1 U346 ( .B1(n323), .B2(n310), .A(n312), .ZN(n301) );
  NAND2_X1 U347 ( .A1(n334), .A2(n347), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  MUX2_X1 U349 ( .A(n547), .B(n302), .S(n329), .Z(n470) );
  MUX2_X1 U350 ( .A(product[13]), .B(n549), .S(n279), .Z(n472) );
  NAND2_X1 U351 ( .A1(n303), .A2(n334), .ZN(n306) );
  INV_X1 U352 ( .A(n312), .ZN(n304) );
  AOI21_X1 U353 ( .B1(n304), .B2(n334), .A(n406), .ZN(n305) );
  OAI21_X1 U354 ( .B1(n323), .B2(n306), .A(n305), .ZN(n308) );
  NAND2_X1 U355 ( .A1(n348), .A2(n346), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U357 ( .A(n549), .B(n309), .S(n16), .Z(n474) );
  MUX2_X1 U358 ( .A(product[14]), .B(n551), .S(n329), .Z(n476) );
  NAND2_X1 U359 ( .A1(n334), .A2(n348), .ZN(n313) );
  NOR2_X1 U360 ( .A1(n310), .A2(n313), .ZN(n319) );
  INV_X1 U361 ( .A(n319), .ZN(n315) );
  AOI21_X1 U362 ( .B1(n406), .B2(n348), .A(n400), .ZN(n311) );
  OAI21_X1 U363 ( .B1(n313), .B2(n312), .A(n311), .ZN(n320) );
  INV_X1 U364 ( .A(n320), .ZN(n314) );
  OAI21_X1 U365 ( .B1(n323), .B2(n315), .A(n314), .ZN(n317) );
  NAND2_X1 U366 ( .A1(n333), .A2(n337), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U368 ( .A(n551), .B(n318), .S(n16), .Z(n478) );
  MUX2_X1 U369 ( .A(product[15]), .B(n553), .S(n279), .Z(n480) );
  NAND2_X1 U370 ( .A1(n319), .A2(n333), .ZN(n322) );
  AOI21_X1 U371 ( .B1(n320), .B2(n333), .A(n399), .ZN(n321) );
  OAI21_X1 U372 ( .B1(n323), .B2(n322), .A(n321), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(n336), .ZN(n325) );
  MUX2_X1 U374 ( .A(n553), .B(n325), .S(n16), .Z(n482) );
  MUX2_X1 U375 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n16), .Z(n484) );
  MUX2_X1 U376 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n16), .Z(n486) );
  MUX2_X1 U377 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n279), .Z(n488) );
  MUX2_X1 U378 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n16), .Z(n490) );
  MUX2_X1 U379 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n329), .Z(n492) );
  MUX2_X1 U380 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n279), .Z(n494) );
  MUX2_X1 U381 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n16), .Z(n496) );
  MUX2_X1 U382 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n329), .Z(n498) );
  MUX2_X1 U383 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n329), .Z(n500) );
  MUX2_X1 U384 ( .A(n326), .B(A_extended[1]), .S(n279), .Z(n502) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n16), .Z(n504) );
  MUX2_X1 U386 ( .A(n14), .B(A_extended[3]), .S(n329), .Z(n506) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n279), .Z(n508) );
  MUX2_X1 U388 ( .A(n15), .B(A_extended[5]), .S(n279), .Z(n510) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n329), .Z(n512) );
  MUX2_X1 U390 ( .A(n328), .B(A_extended[7]), .S(n16), .Z(n514) );
  OR2_X1 U391 ( .A1(n16), .A2(n557), .ZN(n516) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_4 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n311 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n365, n367, n369, n371, n373, n375, n377, n379, n381,
         n383, n385, n387, n389, n391, n393, n395, n397, n399, n401, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n417, n419, n421, n423, n425, n427, n429, n431, n433, n435,
         n437, n439, n441, n443, n445, n447, n449, n451, n453, n455, n457,
         n459, n461, n463, n465, n467, n469, n471, n473, n475, n477, n479,
         n481, n483, n485, n487, n489, n491, n493, n495, n497, n499, n501,
         n503, n505, n507, n509, n511, n513, n515, n517, n519, n521, n523,
         n525, n527, n528, n530, n531, n533, n534, n536, n537, n539, n540,
         n542, n543, n545, n547, n549, n551, n553, n555, n557, n559, n561,
         n563, n564, n565, n566, n567;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n414), .SE(n525), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n415), .SE(n521), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n31) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n414), .SE(n517), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n14) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n414), .SE(n513), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n27) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n415), .SE(n511), .CK(clk), .Q(n564), 
        .QN(n32) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n16) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n415), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n414), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n24) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n414), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n23) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n415), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n20) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n415), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n21) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n414), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n22) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n415), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n18) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n414), .SE(n491), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n414), .SE(n489), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n415), .SE(n487), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n415), .SE(n485), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n414), .SE(n483), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n414), .SE(n481), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n415), .SE(n479), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n414), .SE(n477), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n415), .SE(n475), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n414), .SE(n473), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n415), .SE(n471), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n414), .SE(n469), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n415), .SE(n467), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n465), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n463), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n461), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n415), .SE(n459), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n415), .SE(n457), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n415), .SE(n455), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n415), .SE(n453), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n415), .SE(n451), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n415), .SE(n449), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n415), .SE(n447), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n415), .SE(n445), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n415), .SE(n443), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n415), .SE(n441), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n415), .SE(n439), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n414), .SE(n437), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n414), .SE(n435), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n414), .SE(n433), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n414), .SE(n431), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n414), .SE(n429), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n414), .SE(n427), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n414), .SE(n425), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n414), .SE(n423), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n414), .SE(n421), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n414), .SE(n419), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n414), .SE(n417), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n515), .CK(clk), .Q(n565), 
        .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n567), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n567), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n567), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n567), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n359), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n567), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n358), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n567), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n567), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n356), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n567), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n355), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n567), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n567), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n353), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n567), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n352), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n567), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n351), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n567), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n350), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n567), .SE(n375), .CK(
        clk), .Q(n412), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n567), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n348), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n567), .SE(n371), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n567), .SE(n369), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n567), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n345), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n567), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n344), .QN(n29) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n567), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n343) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n415), .SE(n519), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n342) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n415), .SE(n523), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n17) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n414), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n19) );
  NAND2_X1 U2 ( .A1(n37), .A2(n38), .ZN(n230) );
  BUF_X1 U3 ( .A(n565), .Z(n339) );
  BUF_X1 U4 ( .A(n296), .Z(n255) );
  BUF_X2 U5 ( .A(en), .Z(n341) );
  BUF_X2 U6 ( .A(en), .Z(n12) );
  BUF_X2 U7 ( .A(n296), .Z(n5) );
  CLKBUF_X1 U8 ( .A(n55), .Z(n174) );
  XNOR2_X1 U9 ( .A(n7), .B(n42), .ZN(n136) );
  CLKBUF_X1 U10 ( .A(n137), .Z(n6) );
  BUF_X1 U11 ( .A(n117), .Z(n7) );
  XNOR2_X1 U12 ( .A(n200), .B(n199), .ZN(n216) );
  NOR2_X1 U13 ( .A1(n55), .A2(n18), .ZN(n79) );
  BUF_X1 U14 ( .A(en), .Z(n296) );
  OR2_X1 U15 ( .A1(n251), .A2(n252), .ZN(n250) );
  AND2_X1 U16 ( .A1(\mult_x_1/n310 ), .A2(n566), .ZN(n40) );
  XNOR2_X1 U17 ( .A(n216), .B(n215), .ZN(n244) );
  INV_X1 U18 ( .A(n212), .ZN(n213) );
  XNOR2_X1 U19 ( .A(n252), .B(n251), .ZN(n78) );
  XNOR2_X1 U20 ( .A(n88), .B(n87), .ZN(n92) );
  OAI21_X1 U21 ( .B1(n216), .B2(n204), .A(n203), .ZN(n206) );
  NAND2_X1 U22 ( .A1(n254), .A2(n253), .ZN(n256) );
  NAND2_X1 U23 ( .A1(n252), .A2(n251), .ZN(n253) );
  NAND2_X1 U24 ( .A1(n26), .A2(n250), .ZN(n254) );
  NAND2_X1 U25 ( .A1(n214), .A2(n212), .ZN(n203) );
  NOR2_X1 U26 ( .A1(n214), .A2(n212), .ZN(n204) );
  XNOR2_X1 U27 ( .A(n214), .B(n213), .ZN(n215) );
  XNOR2_X1 U28 ( .A(n146), .B(n338), .ZN(n8) );
  AND2_X1 U29 ( .A1(n566), .A2(\mult_x_1/n281 ), .ZN(n146) );
  CLKBUF_X1 U30 ( .A(n234), .Z(n9) );
  INV_X1 U31 ( .A(n19), .ZN(n10) );
  OAI22_X1 U32 ( .A1(n230), .A2(n44), .B1(n48), .B2(n232), .ZN(n11) );
  INV_X1 U33 ( .A(n17), .ZN(n13) );
  XNOR2_X1 U34 ( .A(n28), .B(n14), .ZN(n36) );
  OAI22_X1 U35 ( .A1(n162), .A2(n70), .B1(n218), .B2(n43), .ZN(n15) );
  BUF_X1 U36 ( .A(rst_n), .Z(n415) );
  BUF_X1 U37 ( .A(rst_n), .Z(n414) );
  INV_X1 U38 ( .A(rst_n), .ZN(n567) );
  INV_X1 U39 ( .A(n342), .ZN(n340) );
  XOR2_X1 U40 ( .A(n66), .B(n65), .Z(n26) );
  AND2_X1 U41 ( .A1(n66), .A2(n65), .ZN(n30) );
  INV_X1 U42 ( .A(n39), .ZN(n232) );
  NAND2_X1 U43 ( .A1(n143), .A2(n350), .ZN(n64) );
  XNOR2_X1 U44 ( .A(\mult_x_1/n311 ), .B(n31), .ZN(n34) );
  XNOR2_X1 U45 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n33) );
  OR2_X2 U46 ( .A1(n34), .A2(n33), .ZN(n171) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n46) );
  INV_X2 U48 ( .A(n34), .ZN(n172) );
  XNOR2_X1 U49 ( .A(n13), .B(\mult_x_1/n284 ), .ZN(n47) );
  OAI22_X1 U50 ( .A1(n171), .A2(n46), .B1(n172), .B2(n47), .ZN(n58) );
  XOR2_X1 U51 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n35) );
  NAND2_X2 U52 ( .A1(n36), .A2(n35), .ZN(n162) );
  XNOR2_X1 U53 ( .A(n340), .B(\mult_x_1/n283 ), .ZN(n43) );
  INV_X1 U54 ( .A(n36), .ZN(n107) );
  INV_X2 U55 ( .A(n107), .ZN(n218) );
  XNOR2_X1 U56 ( .A(n340), .B(\mult_x_1/n282 ), .ZN(n41) );
  OAI22_X1 U57 ( .A1(n162), .A2(n43), .B1(n218), .B2(n41), .ZN(n57) );
  XNOR2_X1 U58 ( .A(n565), .B(n27), .ZN(n37) );
  XNOR2_X1 U59 ( .A(n564), .B(\mult_x_1/a[2] ), .ZN(n38) );
  XNOR2_X1 U60 ( .A(n339), .B(n10), .ZN(n44) );
  XNOR2_X1 U61 ( .A(n146), .B(n339), .ZN(n48) );
  INV_X1 U62 ( .A(n38), .ZN(n39) );
  OAI22_X1 U63 ( .A1(n230), .A2(n44), .B1(n48), .B2(n232), .ZN(n113) );
  INV_X1 U64 ( .A(n113), .ZN(n56) );
  XNOR2_X1 U65 ( .A(n40), .B(\mult_x_1/n310 ), .ZN(n55) );
  NOR2_X1 U66 ( .A1(n20), .A2(n174), .ZN(n120) );
  XNOR2_X1 U67 ( .A(n340), .B(n10), .ZN(n110) );
  OAI22_X1 U68 ( .A1(n162), .A2(n41), .B1(n218), .B2(n110), .ZN(n119) );
  XNOR2_X1 U69 ( .A(n120), .B(n119), .ZN(n42) );
  XNOR2_X1 U70 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n70) );
  OAI22_X1 U71 ( .A1(n162), .A2(n70), .B1(n218), .B2(n43), .ZN(n52) );
  XNOR2_X1 U72 ( .A(n339), .B(\mult_x_1/n282 ), .ZN(n71) );
  OAI22_X1 U73 ( .A1(n230), .A2(n71), .B1(n232), .B2(n44), .ZN(n51) );
  OR2_X1 U74 ( .A1(n15), .A2(n51), .ZN(n61) );
  NOR2_X1 U75 ( .A1(n21), .A2(n174), .ZN(n60) );
  BUF_X2 U76 ( .A(n564), .Z(n338) );
  NAND2_X1 U77 ( .A1(n338), .A2(n16), .ZN(n234) );
  XNOR2_X1 U78 ( .A(n146), .B(n338), .ZN(n54) );
  AOI21_X1 U79 ( .B1(n234), .B2(n16), .A(n8), .ZN(n45) );
  INV_X1 U80 ( .A(n45), .ZN(n77) );
  XNOR2_X1 U81 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n53) );
  OAI22_X1 U82 ( .A1(n171), .A2(n53), .B1(n172), .B2(n46), .ZN(n76) );
  NOR2_X1 U83 ( .A1(n22), .A2(n55), .ZN(n75) );
  XNOR2_X1 U84 ( .A(n13), .B(\mult_x_1/n283 ), .ZN(n106) );
  OAI22_X1 U85 ( .A1(n171), .A2(n47), .B1(n172), .B2(n106), .ZN(n114) );
  AOI21_X1 U86 ( .B1(n232), .B2(n230), .A(n48), .ZN(n49) );
  INV_X1 U87 ( .A(n49), .ZN(n112) );
  XNOR2_X1 U88 ( .A(n138), .B(n137), .ZN(n50) );
  XNOR2_X1 U89 ( .A(n50), .B(n136), .ZN(n187) );
  XNOR2_X1 U90 ( .A(n52), .B(n51), .ZN(n66) );
  XNOR2_X1 U91 ( .A(n13), .B(\mult_x_1/n287 ), .ZN(n68) );
  OAI22_X1 U92 ( .A1(n171), .A2(n68), .B1(n172), .B2(n53), .ZN(n81) );
  XNOR2_X1 U93 ( .A(n338), .B(n10), .ZN(n83) );
  OAI22_X1 U94 ( .A1(n234), .A2(n83), .B1(n54), .B2(n16), .ZN(n80) );
  FA_X1 U95 ( .A(n58), .B(n57), .CI(n56), .CO(n117), .S(n248) );
  FA_X1 U96 ( .A(n61), .B(n60), .CI(n59), .CO(n138), .S(n247) );
  NAND2_X1 U97 ( .A1(n187), .A2(n188), .ZN(n62) );
  NAND2_X1 U98 ( .A1(n62), .A2(n5), .ZN(n63) );
  NAND2_X1 U99 ( .A1(n64), .A2(n63), .ZN(n377) );
  OR2_X1 U100 ( .A1(\mult_x_1/n288 ), .A2(n17), .ZN(n67) );
  OAI22_X1 U101 ( .A1(n171), .A2(n17), .B1(n67), .B2(n172), .ZN(n99) );
  XNOR2_X1 U102 ( .A(n13), .B(\mult_x_1/n288 ), .ZN(n69) );
  OAI22_X1 U103 ( .A1(n171), .A2(n69), .B1(n172), .B2(n68), .ZN(n98) );
  XNOR2_X1 U104 ( .A(n340), .B(\mult_x_1/n285 ), .ZN(n82) );
  OAI22_X1 U105 ( .A1(n162), .A2(n82), .B1(n218), .B2(n70), .ZN(n86) );
  XNOR2_X1 U106 ( .A(n339), .B(\mult_x_1/n283 ), .ZN(n84) );
  OAI22_X1 U107 ( .A1(n230), .A2(n84), .B1(n232), .B2(n71), .ZN(n85) );
  OR2_X1 U108 ( .A1(n86), .A2(n85), .ZN(n72) );
  NAND2_X1 U109 ( .A1(n88), .A2(n72), .ZN(n74) );
  NAND2_X1 U110 ( .A1(n86), .A2(n85), .ZN(n73) );
  NAND2_X1 U111 ( .A1(n74), .A2(n73), .ZN(n252) );
  FA_X1 U112 ( .A(n77), .B(n76), .CI(n75), .CO(n59), .S(n251) );
  XNOR2_X1 U113 ( .A(n26), .B(n78), .ZN(n258) );
  INV_X1 U114 ( .A(n258), .ZN(n90) );
  FA_X1 U115 ( .A(n81), .B(n80), .CI(n79), .CO(n65), .S(n94) );
  XNOR2_X1 U116 ( .A(n340), .B(\mult_x_1/n286 ), .ZN(n160) );
  OAI22_X1 U117 ( .A1(n162), .A2(n160), .B1(n218), .B2(n82), .ZN(n102) );
  XNOR2_X1 U118 ( .A(n338), .B(\mult_x_1/n282 ), .ZN(n95) );
  OAI22_X1 U119 ( .A1(n234), .A2(n95), .B1(n83), .B2(n16), .ZN(n101) );
  XNOR2_X1 U120 ( .A(n339), .B(\mult_x_1/n284 ), .ZN(n97) );
  OAI22_X1 U121 ( .A1(n230), .A2(n97), .B1(n232), .B2(n84), .ZN(n100) );
  XNOR2_X1 U122 ( .A(n86), .B(n85), .ZN(n87) );
  INV_X1 U123 ( .A(n257), .ZN(n89) );
  NAND3_X1 U124 ( .A1(n5), .A2(n90), .A3(n89), .ZN(n91) );
  OAI21_X1 U125 ( .B1(n5), .B2(n411), .A(n91), .ZN(n379) );
  NAND2_X1 U126 ( .A1(n143), .A2(n354), .ZN(n105) );
  FA_X1 U127 ( .A(n94), .B(n93), .CI(n92), .CO(n257), .S(n191) );
  XNOR2_X1 U128 ( .A(n338), .B(\mult_x_1/n283 ), .ZN(n202) );
  OAI22_X1 U129 ( .A1(n234), .A2(n202), .B1(n95), .B2(n16), .ZN(n165) );
  INV_X1 U130 ( .A(n172), .ZN(n96) );
  AND2_X1 U131 ( .A1(\mult_x_1/n288 ), .A2(n96), .ZN(n164) );
  XNOR2_X1 U132 ( .A(n339), .B(\mult_x_1/n285 ), .ZN(n201) );
  OAI22_X1 U133 ( .A1(n230), .A2(n201), .B1(n232), .B2(n97), .ZN(n163) );
  HA_X1 U134 ( .A(n99), .B(n98), .CO(n88), .S(n156) );
  FA_X1 U135 ( .A(n102), .B(n101), .CI(n100), .CO(n93), .S(n155) );
  NAND2_X1 U136 ( .A1(n191), .A2(n190), .ZN(n103) );
  NAND2_X1 U137 ( .A1(n103), .A2(n5), .ZN(n104) );
  NAND2_X1 U138 ( .A1(n105), .A2(n104), .ZN(n385) );
  XNOR2_X1 U139 ( .A(n13), .B(\mult_x_1/n282 ), .ZN(n129) );
  OAI22_X1 U140 ( .A1(n171), .A2(n106), .B1(n172), .B2(n129), .ZN(n125) );
  XNOR2_X1 U141 ( .A(n146), .B(\mult_x_1/n311 ), .ZN(n130) );
  INV_X1 U142 ( .A(n130), .ZN(n108) );
  NAND2_X1 U143 ( .A1(n108), .A2(n107), .ZN(n109) );
  OAI21_X1 U144 ( .B1(n162), .B2(n110), .A(n109), .ZN(n149) );
  INV_X1 U145 ( .A(n149), .ZN(n124) );
  XNOR2_X1 U146 ( .A(n125), .B(n124), .ZN(n111) );
  NOR2_X1 U147 ( .A1(n23), .A2(n174), .ZN(n123) );
  XNOR2_X1 U148 ( .A(n111), .B(n123), .ZN(n135) );
  FA_X1 U149 ( .A(n114), .B(n11), .CI(n112), .CO(n134), .S(n137) );
  INV_X1 U150 ( .A(n120), .ZN(n116) );
  INV_X1 U151 ( .A(n119), .ZN(n115) );
  NAND2_X1 U152 ( .A1(n116), .A2(n115), .ZN(n118) );
  NAND2_X1 U153 ( .A1(n117), .A2(n118), .ZN(n122) );
  NAND2_X1 U154 ( .A1(n120), .A2(n119), .ZN(n121) );
  NAND2_X1 U155 ( .A1(n122), .A2(n121), .ZN(n133) );
  INV_X1 U156 ( .A(n123), .ZN(n128) );
  NOR2_X1 U157 ( .A1(n125), .A2(n124), .ZN(n127) );
  NAND2_X1 U158 ( .A1(n125), .A2(n124), .ZN(n126) );
  OAI21_X1 U159 ( .B1(n128), .B2(n127), .A(n126), .ZN(n153) );
  NOR2_X1 U160 ( .A1(n24), .A2(n174), .ZN(n152) );
  XNOR2_X1 U161 ( .A(n13), .B(n10), .ZN(n147) );
  OAI22_X1 U162 ( .A1(n171), .A2(n129), .B1(n172), .B2(n147), .ZN(n150) );
  AOI21_X1 U163 ( .B1(n218), .B2(n162), .A(n130), .ZN(n131) );
  INV_X1 U164 ( .A(n131), .ZN(n148) );
  OAI21_X1 U165 ( .B1(n209), .B2(n210), .A(n5), .ZN(n132) );
  OAI21_X1 U166 ( .B1(n5), .B2(n29), .A(n132), .ZN(n365) );
  FA_X1 U167 ( .A(n135), .B(n134), .CI(n133), .CO(n209), .S(n263) );
  NAND2_X1 U168 ( .A1(n136), .A2(n6), .ZN(n141) );
  NAND2_X1 U169 ( .A1(n136), .A2(n138), .ZN(n140) );
  NAND2_X1 U170 ( .A1(n138), .A2(n6), .ZN(n139) );
  NAND3_X1 U171 ( .A1(n141), .A2(n140), .A3(n139), .ZN(n262) );
  NAND2_X1 U172 ( .A1(n263), .A2(n262), .ZN(n142) );
  NAND2_X1 U173 ( .A1(n142), .A2(n255), .ZN(n145) );
  INV_X1 U174 ( .A(n255), .ZN(n143) );
  NAND2_X1 U175 ( .A1(n143), .A2(n359), .ZN(n144) );
  NAND2_X1 U176 ( .A1(n145), .A2(n144), .ZN(n395) );
  NOR2_X1 U197 ( .A1(n25), .A2(n174), .ZN(n169) );
  XNOR2_X1 U198 ( .A(n146), .B(n13), .ZN(n170) );
  OAI22_X1 U199 ( .A1(n171), .A2(n147), .B1(n170), .B2(n172), .ZN(n178) );
  INV_X1 U200 ( .A(n178), .ZN(n168) );
  FA_X1 U201 ( .A(n150), .B(n149), .CI(n148), .CO(n167), .S(n151) );
  FA_X1 U202 ( .A(n153), .B(n152), .CI(n151), .CO(n184), .S(n210) );
  OR2_X1 U203 ( .A1(n185), .A2(n184), .ZN(n154) );
  MUX2_X1 U204 ( .A(n343), .B(n154), .S(n5), .Z(n363) );
  FA_X1 U205 ( .A(n157), .B(n156), .CI(n155), .CO(n190), .S(n194) );
  OR2_X1 U206 ( .A1(\mult_x_1/n288 ), .A2(n342), .ZN(n158) );
  OAI22_X1 U207 ( .A1(n162), .A2(n342), .B1(n158), .B2(n218), .ZN(n200) );
  XNOR2_X1 U208 ( .A(n340), .B(\mult_x_1/n288 ), .ZN(n159) );
  XNOR2_X1 U209 ( .A(n340), .B(\mult_x_1/n287 ), .ZN(n161) );
  OAI22_X1 U210 ( .A1(n162), .A2(n159), .B1(n218), .B2(n161), .ZN(n199) );
  AND2_X1 U211 ( .A1(n200), .A2(n199), .ZN(n198) );
  OAI22_X1 U212 ( .A1(n162), .A2(n161), .B1(n218), .B2(n160), .ZN(n197) );
  FA_X1 U213 ( .A(n165), .B(n164), .CI(n163), .CO(n157), .S(n196) );
  OR2_X1 U214 ( .A1(n194), .A2(n193), .ZN(n166) );
  MUX2_X1 U215 ( .A(n346), .B(n166), .S(n5), .Z(n369) );
  FA_X1 U216 ( .A(n169), .B(n168), .CI(n167), .CO(n180), .S(n185) );
  AOI21_X1 U217 ( .B1(n172), .B2(n171), .A(n170), .ZN(n173) );
  INV_X1 U218 ( .A(n173), .ZN(n176) );
  NOR2_X1 U219 ( .A1(n19), .A2(n174), .ZN(n175) );
  XOR2_X1 U220 ( .A(n176), .B(n175), .Z(n177) );
  XOR2_X1 U221 ( .A(n178), .B(n177), .Z(n179) );
  OR2_X1 U222 ( .A1(n180), .A2(n179), .ZN(n182) );
  NAND2_X1 U223 ( .A1(n180), .A2(n179), .ZN(n181) );
  NAND2_X1 U224 ( .A1(n182), .A2(n181), .ZN(n183) );
  MUX2_X1 U225 ( .A(n347), .B(n183), .S(n5), .Z(n371) );
  NAND2_X1 U226 ( .A1(n185), .A2(n184), .ZN(n186) );
  MUX2_X1 U227 ( .A(n348), .B(n186), .S(n5), .Z(n373) );
  NOR2_X1 U228 ( .A1(n187), .A2(n188), .ZN(n189) );
  MUX2_X1 U229 ( .A(n349), .B(n189), .S(n5), .Z(n375) );
  NOR2_X1 U230 ( .A1(n191), .A2(n190), .ZN(n192) );
  MUX2_X1 U231 ( .A(n353), .B(n192), .S(n5), .Z(n383) );
  NAND2_X1 U232 ( .A1(n194), .A2(n193), .ZN(n195) );
  MUX2_X1 U233 ( .A(n355), .B(n195), .S(n255), .Z(n387) );
  FA_X1 U234 ( .A(n198), .B(n197), .CI(n196), .CO(n193), .S(n207) );
  XNOR2_X1 U235 ( .A(n339), .B(\mult_x_1/n286 ), .ZN(n220) );
  OAI22_X1 U236 ( .A1(n230), .A2(n220), .B1(n232), .B2(n201), .ZN(n214) );
  XNOR2_X1 U237 ( .A(n338), .B(\mult_x_1/n284 ), .ZN(n217) );
  OAI22_X1 U238 ( .A1(n9), .A2(n217), .B1(n202), .B2(n16), .ZN(n212) );
  NOR2_X1 U239 ( .A1(n207), .A2(n206), .ZN(n205) );
  MUX2_X1 U240 ( .A(n356), .B(n205), .S(n255), .Z(n389) );
  NAND2_X1 U241 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U242 ( .A(n357), .B(n208), .S(n255), .Z(n391) );
  NAND2_X1 U243 ( .A1(n210), .A2(n209), .ZN(n211) );
  MUX2_X1 U244 ( .A(n358), .B(n211), .S(n255), .Z(n393) );
  XNOR2_X1 U245 ( .A(n338), .B(\mult_x_1/n285 ), .ZN(n226) );
  OAI22_X1 U246 ( .A1(n9), .A2(n226), .B1(n217), .B2(n16), .ZN(n223) );
  INV_X1 U247 ( .A(n218), .ZN(n219) );
  AND2_X1 U248 ( .A1(\mult_x_1/n288 ), .A2(n219), .ZN(n222) );
  XNOR2_X1 U249 ( .A(n339), .B(\mult_x_1/n287 ), .ZN(n224) );
  OAI22_X1 U250 ( .A1(n230), .A2(n224), .B1(n232), .B2(n220), .ZN(n221) );
  OR2_X1 U251 ( .A1(n244), .A2(n243), .ZN(n289) );
  FA_X1 U252 ( .A(n223), .B(n222), .CI(n221), .CO(n243), .S(n242) );
  XNOR2_X1 U253 ( .A(n339), .B(\mult_x_1/n288 ), .ZN(n225) );
  OAI22_X1 U254 ( .A1(n230), .A2(n225), .B1(n232), .B2(n224), .ZN(n228) );
  XNOR2_X1 U255 ( .A(n338), .B(\mult_x_1/n286 ), .ZN(n231) );
  OAI22_X1 U256 ( .A1(n234), .A2(n231), .B1(n226), .B2(n16), .ZN(n227) );
  NOR2_X1 U257 ( .A1(n242), .A2(n241), .ZN(n282) );
  HA_X1 U258 ( .A(n228), .B(n227), .CO(n241), .S(n239) );
  OR2_X1 U259 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n229) );
  OAI22_X1 U260 ( .A1(n230), .A2(n28), .B1(n229), .B2(n232), .ZN(n238) );
  OR2_X1 U261 ( .A1(n239), .A2(n238), .ZN(n278) );
  XNOR2_X1 U262 ( .A(n338), .B(\mult_x_1/n287 ), .ZN(n233) );
  OAI22_X1 U263 ( .A1(n9), .A2(n233), .B1(n231), .B2(n16), .ZN(n237) );
  AND2_X1 U264 ( .A1(\mult_x_1/n288 ), .A2(n39), .ZN(n236) );
  NOR2_X1 U265 ( .A1(n237), .A2(n236), .ZN(n271) );
  OAI22_X1 U266 ( .A1(n9), .A2(\mult_x_1/n288 ), .B1(n233), .B2(n16), .ZN(n268) );
  OR2_X1 U267 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n235) );
  NAND2_X1 U268 ( .A1(n235), .A2(n9), .ZN(n267) );
  NAND2_X1 U269 ( .A1(n268), .A2(n267), .ZN(n274) );
  NAND2_X1 U270 ( .A1(n237), .A2(n236), .ZN(n272) );
  OAI21_X1 U271 ( .B1(n271), .B2(n274), .A(n272), .ZN(n279) );
  NAND2_X1 U272 ( .A1(n239), .A2(n238), .ZN(n277) );
  INV_X1 U273 ( .A(n277), .ZN(n240) );
  AOI21_X1 U274 ( .B1(n278), .B2(n279), .A(n240), .ZN(n285) );
  NAND2_X1 U275 ( .A1(n242), .A2(n241), .ZN(n283) );
  OAI21_X1 U276 ( .B1(n282), .B2(n285), .A(n283), .ZN(n290) );
  NAND2_X1 U277 ( .A1(n244), .A2(n243), .ZN(n288) );
  INV_X1 U278 ( .A(n288), .ZN(n245) );
  AOI21_X1 U279 ( .B1(n289), .B2(n290), .A(n245), .ZN(n246) );
  MUX2_X1 U280 ( .A(n360), .B(n246), .S(n255), .Z(n397) );
  FA_X1 U281 ( .A(n30), .B(n248), .CI(n247), .CO(n188), .S(n249) );
  MUX2_X1 U282 ( .A(n361), .B(n249), .S(n255), .Z(n399) );
  MUX2_X1 U283 ( .A(n362), .B(n256), .S(n255), .Z(n401) );
  NAND2_X1 U284 ( .A1(n258), .A2(n257), .ZN(n259) );
  NAND2_X1 U285 ( .A1(n259), .A2(n5), .ZN(n261) );
  OR2_X1 U286 ( .A1(n5), .A2(n406), .ZN(n260) );
  NAND2_X1 U287 ( .A1(n261), .A2(n260), .ZN(n381) );
  OAI21_X1 U288 ( .B1(n262), .B2(n263), .A(n5), .ZN(n265) );
  OR2_X1 U289 ( .A1(n5), .A2(n404), .ZN(n264) );
  NAND2_X1 U290 ( .A1(n265), .A2(n264), .ZN(n367) );
  MUX2_X1 U291 ( .A(product[0]), .B(n527), .S(n341), .Z(n417) );
  MUX2_X1 U292 ( .A(n527), .B(n528), .S(n12), .Z(n419) );
  AND2_X1 U293 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n266) );
  MUX2_X1 U294 ( .A(n528), .B(n266), .S(n341), .Z(n421) );
  MUX2_X1 U295 ( .A(product[1]), .B(n530), .S(n12), .Z(n423) );
  MUX2_X1 U296 ( .A(n530), .B(n531), .S(n341), .Z(n425) );
  OR2_X1 U297 ( .A1(n268), .A2(n267), .ZN(n269) );
  AND2_X1 U298 ( .A1(n269), .A2(n274), .ZN(n270) );
  MUX2_X1 U299 ( .A(n531), .B(n270), .S(n12), .Z(n427) );
  MUX2_X1 U300 ( .A(product[2]), .B(n533), .S(n341), .Z(n429) );
  MUX2_X1 U301 ( .A(n533), .B(n534), .S(n12), .Z(n431) );
  INV_X1 U302 ( .A(n271), .ZN(n273) );
  NAND2_X1 U303 ( .A1(n273), .A2(n272), .ZN(n275) );
  XOR2_X1 U304 ( .A(n275), .B(n274), .Z(n276) );
  MUX2_X1 U305 ( .A(n534), .B(n276), .S(n341), .Z(n433) );
  MUX2_X1 U306 ( .A(product[3]), .B(n536), .S(n12), .Z(n435) );
  MUX2_X1 U307 ( .A(n536), .B(n537), .S(n341), .Z(n437) );
  NAND2_X1 U308 ( .A1(n278), .A2(n277), .ZN(n280) );
  XNOR2_X1 U309 ( .A(n280), .B(n279), .ZN(n281) );
  MUX2_X1 U310 ( .A(n537), .B(n281), .S(n12), .Z(n439) );
  MUX2_X1 U311 ( .A(product[4]), .B(n539), .S(n341), .Z(n441) );
  MUX2_X1 U312 ( .A(n539), .B(n540), .S(n12), .Z(n443) );
  INV_X1 U313 ( .A(n282), .ZN(n284) );
  NAND2_X1 U314 ( .A1(n284), .A2(n283), .ZN(n286) );
  XOR2_X1 U315 ( .A(n286), .B(n285), .Z(n287) );
  MUX2_X1 U316 ( .A(n540), .B(n287), .S(n341), .Z(n445) );
  MUX2_X1 U317 ( .A(product[5]), .B(n542), .S(n12), .Z(n447) );
  MUX2_X1 U318 ( .A(n542), .B(n543), .S(n341), .Z(n449) );
  NAND2_X1 U319 ( .A1(n289), .A2(n288), .ZN(n291) );
  XNOR2_X1 U320 ( .A(n291), .B(n290), .ZN(n292) );
  MUX2_X1 U321 ( .A(n543), .B(n292), .S(n12), .Z(n451) );
  MUX2_X1 U322 ( .A(product[6]), .B(n545), .S(n341), .Z(n453) );
  NAND2_X1 U323 ( .A1(n407), .A2(n357), .ZN(n293) );
  XOR2_X1 U324 ( .A(n293), .B(n360), .Z(n294) );
  MUX2_X1 U325 ( .A(n545), .B(n294), .S(n12), .Z(n455) );
  MUX2_X1 U326 ( .A(product[7]), .B(n547), .S(n341), .Z(n457) );
  OAI21_X1 U327 ( .B1(n356), .B2(n360), .A(n357), .ZN(n298) );
  NAND2_X1 U328 ( .A1(n346), .A2(n355), .ZN(n295) );
  XNOR2_X1 U329 ( .A(n298), .B(n295), .ZN(n297) );
  MUX2_X1 U330 ( .A(n547), .B(n297), .S(n12), .Z(n459) );
  MUX2_X1 U331 ( .A(product[8]), .B(n549), .S(n12), .Z(n461) );
  AOI21_X1 U332 ( .B1(n298), .B2(n346), .A(n409), .ZN(n301) );
  NAND2_X1 U333 ( .A1(n410), .A2(n354), .ZN(n299) );
  XOR2_X1 U334 ( .A(n301), .B(n299), .Z(n300) );
  MUX2_X1 U335 ( .A(n549), .B(n300), .S(n12), .Z(n463) );
  MUX2_X1 U336 ( .A(product[9]), .B(n551), .S(n12), .Z(n465) );
  OAI21_X1 U337 ( .B1(n301), .B2(n353), .A(n354), .ZN(n312) );
  INV_X1 U338 ( .A(n312), .ZN(n304) );
  NAND2_X1 U339 ( .A1(n411), .A2(n352), .ZN(n302) );
  XOR2_X1 U340 ( .A(n304), .B(n302), .Z(n303) );
  MUX2_X1 U341 ( .A(n551), .B(n303), .S(n341), .Z(n467) );
  MUX2_X1 U342 ( .A(product[10]), .B(n553), .S(n341), .Z(n469) );
  OAI21_X1 U343 ( .B1(n304), .B2(n351), .A(n352), .ZN(n307) );
  NOR2_X1 U344 ( .A1(n361), .A2(n362), .ZN(n310) );
  INV_X1 U345 ( .A(n310), .ZN(n305) );
  NAND2_X1 U346 ( .A1(n361), .A2(n362), .ZN(n309) );
  NAND2_X1 U347 ( .A1(n305), .A2(n309), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n307), .B(n306), .ZN(n308) );
  MUX2_X1 U349 ( .A(n553), .B(n308), .S(n341), .Z(n471) );
  MUX2_X1 U350 ( .A(product[11]), .B(n555), .S(n12), .Z(n473) );
  NOR2_X1 U351 ( .A1(n310), .A2(n351), .ZN(n313) );
  OAI21_X1 U352 ( .B1(n310), .B2(n352), .A(n309), .ZN(n311) );
  AOI21_X1 U353 ( .B1(n313), .B2(n312), .A(n311), .ZN(n335) );
  NAND2_X1 U354 ( .A1(n412), .A2(n350), .ZN(n314) );
  XOR2_X1 U355 ( .A(n335), .B(n314), .Z(n315) );
  MUX2_X1 U356 ( .A(n555), .B(n315), .S(n341), .Z(n475) );
  MUX2_X1 U357 ( .A(product[12]), .B(n557), .S(n12), .Z(n477) );
  OAI21_X1 U358 ( .B1(n335), .B2(n349), .A(n350), .ZN(n317) );
  NAND2_X1 U359 ( .A1(n345), .A2(n359), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U361 ( .A(n557), .B(n318), .S(n341), .Z(n479) );
  MUX2_X1 U362 ( .A(product[13]), .B(n559), .S(n12), .Z(n481) );
  NAND2_X1 U363 ( .A1(n412), .A2(n345), .ZN(n320) );
  AOI21_X1 U364 ( .B1(n405), .B2(n345), .A(n413), .ZN(n319) );
  OAI21_X1 U365 ( .B1(n335), .B2(n320), .A(n319), .ZN(n322) );
  NAND2_X1 U366 ( .A1(n344), .A2(n358), .ZN(n321) );
  XNOR2_X1 U367 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U368 ( .A(n559), .B(n323), .S(n341), .Z(n483) );
  MUX2_X1 U369 ( .A(product[14]), .B(n561), .S(n12), .Z(n485) );
  NAND2_X1 U370 ( .A1(n345), .A2(n344), .ZN(n325) );
  NOR2_X1 U371 ( .A1(n349), .A2(n325), .ZN(n331) );
  INV_X1 U372 ( .A(n331), .ZN(n327) );
  AOI21_X1 U373 ( .B1(n413), .B2(n344), .A(n408), .ZN(n324) );
  OAI21_X1 U374 ( .B1(n325), .B2(n350), .A(n324), .ZN(n332) );
  INV_X1 U375 ( .A(n332), .ZN(n326) );
  OAI21_X1 U376 ( .B1(n335), .B2(n327), .A(n326), .ZN(n329) );
  NAND2_X1 U377 ( .A1(n343), .A2(n348), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n330) );
  MUX2_X1 U379 ( .A(n561), .B(n330), .S(n341), .Z(n487) );
  MUX2_X1 U380 ( .A(product[15]), .B(n563), .S(n12), .Z(n489) );
  NAND2_X1 U381 ( .A1(n331), .A2(n343), .ZN(n334) );
  AOI21_X1 U382 ( .B1(n332), .B2(n343), .A(n403), .ZN(n333) );
  OAI21_X1 U383 ( .B1(n335), .B2(n334), .A(n333), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n336), .B(n347), .ZN(n337) );
  MUX2_X1 U385 ( .A(n563), .B(n337), .S(n341), .Z(n491) );
  MUX2_X1 U386 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n12), .Z(n493) );
  MUX2_X1 U387 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n12), .Z(n495) );
  MUX2_X1 U388 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n341), .Z(n497) );
  MUX2_X1 U389 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n12), .Z(n499) );
  MUX2_X1 U390 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n341), .Z(n501) );
  MUX2_X1 U391 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n12), .Z(n503) );
  MUX2_X1 U392 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n341), .Z(n505) );
  MUX2_X1 U393 ( .A(n10), .B(B_extended[7]), .S(n341), .Z(n507) );
  MUX2_X1 U394 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n12), .Z(n509) );
  MUX2_X1 U395 ( .A(n338), .B(A_extended[1]), .S(n341), .Z(n511) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n12), .Z(n513) );
  MUX2_X1 U397 ( .A(n339), .B(A_extended[3]), .S(n341), .Z(n515) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n341), .Z(n517) );
  MUX2_X1 U399 ( .A(n340), .B(A_extended[5]), .S(n12), .Z(n519) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n12), .Z(n521) );
  MUX2_X1 U401 ( .A(n13), .B(A_extended[7]), .S(n341), .Z(n523) );
  OR2_X1 U402 ( .A1(n341), .A2(n566), .ZN(n525) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_5 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n345, n347, n349, n351, n353, n355, n357,
         n359, n361, n363, n365, n367, n369, n371, n373, n375, n377, n379,
         n381, n383, n385, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n398, n400, n402, n404, n406, n408, n410, n412, n414,
         n416, n418, n420, n422, n424, n426, n428, n430, n432, n434, n436,
         n438, n440, n442, n444, n446, n448, n450, n452, n454, n456, n458,
         n460, n462, n464, n466, n468, n470, n472, n474, n476, n478, n480,
         n482, n484, n486, n488, n490, n492, n494, n496, n498, n500, n502,
         n504, n506, n507, n509, n510, n512, n513, n515, n516, n518, n519,
         n521, n523, n525, n527, n529, n531, n533, n535, n537, n539, n541,
         n542, n543, n544, n545;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n396), .SE(n504), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n396), .SE(n500), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n396), .SE(n498), .CK(clk), .Q(n543), 
        .QN(n319) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n395), .SE(n496), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n318) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(n542), 
        .QN(n18) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n396), .SE(n492), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n13) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n396), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n16) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n395), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n10) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n395), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n395), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n396), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n396), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n395), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n396), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n395), .SE(n472), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n17) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n395), .SE(n470), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n396), .SE(n468), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n396), .SE(n466), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n395), .SE(n464), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n395), .SE(n462), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n396), .SE(n460), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n395), .SE(n458), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n396), .SE(n456), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n395), .SE(n454), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n396), .SE(n452), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n395), .SE(n450), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n396), .SE(n448), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n395), .SE(n446), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n396), .SE(n444), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n395), .SE(n442), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n396), .SE(n440), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n396), .SE(n438), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n396), .SE(n436), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n396), .SE(n434), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n396), .SE(n432), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n396), .SE(n430), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n396), .SE(n428), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n396), .SE(n426), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n396), .SE(n424), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n396), .SE(n422), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n396), .SE(n420), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n395), .SE(n418), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n395), .SE(n416), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n395), .SE(n414), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n395), .SE(n412), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n395), .SE(n410), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n395), .SE(n408), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n395), .SE(n406), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n395), .SE(n404), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n395), .SE(n402), .CK(clk), .Q(n507)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n395), .SE(n400), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n395), .SE(n398), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(rst_n), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n19) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n545), .SE(n385), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2_IP  ( .D(1'b1), .SI(n545), .SE(n383), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n545), .SE(n381), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n545), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n545), .SE(n377), .CK(
        clk), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n545), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n545), .SE(n373), .CK(
        clk), .Q(n393), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n545), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n335), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n545), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n334), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n545), .SE(n367), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n545), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n545), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n545), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n330), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n545), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n329), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2  ( .D(n545), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n545), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n327), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n545), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n326), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n545), .SI(1'b1), .SE(n351), .CK(clk), 
        .Q(n325), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n545), .SE(n349), .CK(
        clk), .QN(n324) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n545), .SE(n347), .CK(
        clk), .QN(n323) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n545), .SI(1'b1), .SE(n345), .CK(clk), 
        .Q(n322) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n545), .SI(1'b1), .SE(n343), .CK(clk), 
        .Q(n321) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n395), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n320) );
  BUF_X2 U2 ( .A(n60), .Z(n5) );
  XOR2_X1 U3 ( .A(n235), .B(n234), .Z(n6) );
  XOR2_X1 U4 ( .A(n233), .B(n6), .Z(n157) );
  NAND2_X1 U5 ( .A1(n233), .A2(n235), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n233), .A2(n234), .ZN(n8) );
  NAND2_X1 U7 ( .A1(n235), .A2(n234), .ZN(n9) );
  NAND3_X1 U8 ( .A1(n7), .A2(n8), .A3(n9), .ZN(n236) );
  INV_X1 U9 ( .A(n320), .ZN(n316) );
  XNOR2_X1 U10 ( .A(n542), .B(\mult_x_1/a[4] ), .ZN(n27) );
  OAI22_X1 U11 ( .A1(n177), .A2(n44), .B1(n104), .B2(n32), .ZN(n48) );
  XNOR2_X1 U12 ( .A(n25), .B(n52), .ZN(n231) );
  XNOR2_X1 U13 ( .A(n50), .B(n51), .ZN(n25) );
  BUF_X2 U14 ( .A(n543), .Z(n315) );
  INV_X1 U15 ( .A(n10), .ZN(n11) );
  NAND2_X1 U16 ( .A1(n22), .A2(n23), .ZN(n113) );
  INV_X2 U17 ( .A(n320), .ZN(n12) );
  XNOR2_X1 U18 ( .A(n13), .B(\mult_x_1/n313 ), .ZN(n29) );
  NAND2_X2 U19 ( .A1(n203), .A2(n16), .ZN(n204) );
  OAI21_X1 U20 ( .B1(n104), .B2(n44), .A(n43), .ZN(n14) );
  AND2_X2 U21 ( .A1(n544), .A2(\mult_x_1/n281 ), .ZN(n63) );
  OAI22_X1 U22 ( .A1(n198), .A2(n45), .B1(n81), .B2(n200), .ZN(n15) );
  BUF_X1 U23 ( .A(rst_n), .Z(n396) );
  BUF_X1 U24 ( .A(rst_n), .Z(n395) );
  INV_X1 U25 ( .A(rst_n), .ZN(n545) );
  BUF_X2 U26 ( .A(n542), .Z(n314) );
  AND2_X2 U27 ( .A1(n544), .A2(\mult_x_1/n310 ), .ZN(n116) );
  XNOR2_X1 U28 ( .A(n116), .B(n316), .ZN(n60) );
  XNOR2_X1 U29 ( .A(n116), .B(\mult_x_1/n287 ), .ZN(n20) );
  NOR2_X1 U30 ( .A1(n5), .A2(n20), .ZN(n50) );
  BUF_X2 U31 ( .A(\mult_x_1/n313 ), .Z(n203) );
  XNOR2_X1 U32 ( .A(n63), .B(n203), .ZN(n38) );
  AOI21_X1 U33 ( .B1(n204), .B2(n16), .A(n38), .ZN(n21) );
  INV_X1 U34 ( .A(n21), .ZN(n51) );
  XOR2_X1 U35 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n22) );
  XNOR2_X1 U36 ( .A(n543), .B(\mult_x_1/a[6] ), .ZN(n23) );
  XNOR2_X1 U37 ( .A(n12), .B(\mult_x_1/n286 ), .ZN(n36) );
  INV_X1 U38 ( .A(n23), .ZN(n24) );
  INV_X2 U39 ( .A(n24), .ZN(n114) );
  XNOR2_X1 U40 ( .A(n12), .B(\mult_x_1/n285 ), .ZN(n42) );
  OAI22_X1 U41 ( .A1(n113), .A2(n36), .B1(n114), .B2(n42), .ZN(n52) );
  XOR2_X1 U42 ( .A(n318), .B(n319), .Z(n26) );
  NAND2_X2 U43 ( .A1(n26), .A2(n27), .ZN(n104) );
  XNOR2_X1 U44 ( .A(n315), .B(\mult_x_1/n285 ), .ZN(n95) );
  BUF_X2 U45 ( .A(n27), .Z(n177) );
  XNOR2_X1 U46 ( .A(n315), .B(\mult_x_1/n284 ), .ZN(n32) );
  OAI22_X1 U47 ( .A1(n104), .A2(n95), .B1(n177), .B2(n32), .ZN(n151) );
  XNOR2_X1 U48 ( .A(\mult_x_1/a[2] ), .B(n542), .ZN(n28) );
  OR2_X2 U49 ( .A1(n28), .A2(n29), .ZN(n198) );
  XNOR2_X1 U50 ( .A(n314), .B(\mult_x_1/n283 ), .ZN(n98) );
  INV_X2 U51 ( .A(n29), .ZN(n200) );
  XNOR2_X1 U52 ( .A(n314), .B(\mult_x_1/n282 ), .ZN(n33) );
  OAI22_X1 U53 ( .A1(n198), .A2(n98), .B1(n200), .B2(n33), .ZN(n150) );
  OR2_X1 U54 ( .A1(\mult_x_1/n288 ), .A2(n320), .ZN(n30) );
  OAI22_X1 U55 ( .A1(n113), .A2(n320), .B1(n30), .B2(n114), .ZN(n94) );
  XNOR2_X1 U56 ( .A(n316), .B(\mult_x_1/n288 ), .ZN(n31) );
  XNOR2_X1 U57 ( .A(n316), .B(\mult_x_1/n287 ), .ZN(n37) );
  OAI22_X1 U58 ( .A1(n113), .A2(n31), .B1(n114), .B2(n37), .ZN(n93) );
  XNOR2_X1 U59 ( .A(n315), .B(\mult_x_1/n283 ), .ZN(n44) );
  XNOR2_X1 U60 ( .A(n314), .B(\mult_x_1/n281 ), .ZN(n45) );
  OAI22_X1 U61 ( .A1(n198), .A2(n33), .B1(n200), .B2(n45), .ZN(n47) );
  XNOR2_X1 U62 ( .A(n48), .B(n47), .ZN(n41) );
  INV_X1 U63 ( .A(n116), .ZN(n34) );
  OR2_X1 U64 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n35) );
  NOR2_X1 U65 ( .A1(n35), .A2(n5), .ZN(n40) );
  OAI22_X1 U66 ( .A1(n113), .A2(n37), .B1(n114), .B2(n36), .ZN(n145) );
  XNOR2_X1 U67 ( .A(n203), .B(\mult_x_1/n281 ), .ZN(n96) );
  OAI22_X1 U68 ( .A1(n204), .A2(n96), .B1(n38), .B2(n16), .ZN(n144) );
  NOR2_X1 U69 ( .A1(n60), .A2(n17), .ZN(n143) );
  FA_X1 U70 ( .A(n41), .B(n40), .CI(n39), .CO(n224), .S(n229) );
  XNOR2_X1 U71 ( .A(n12), .B(\mult_x_1/n284 ), .ZN(n80) );
  OAI22_X1 U72 ( .A1(n113), .A2(n42), .B1(n114), .B2(n80), .ZN(n87) );
  XNOR2_X1 U73 ( .A(n315), .B(\mult_x_1/n282 ), .ZN(n85) );
  OR2_X1 U74 ( .A1(n177), .A2(n85), .ZN(n43) );
  OAI21_X1 U75 ( .B1(n104), .B2(n44), .A(n43), .ZN(n88) );
  XNOR2_X1 U76 ( .A(n87), .B(n14), .ZN(n46) );
  XNOR2_X1 U77 ( .A(n63), .B(n314), .ZN(n81) );
  OAI22_X1 U78 ( .A1(n198), .A2(n45), .B1(n81), .B2(n200), .ZN(n137) );
  INV_X1 U79 ( .A(n137), .ZN(n86) );
  XNOR2_X1 U80 ( .A(n46), .B(n86), .ZN(n223) );
  XNOR2_X1 U81 ( .A(n224), .B(n223), .ZN(n55) );
  OR2_X1 U82 ( .A1(n48), .A2(n47), .ZN(n135) );
  XNOR2_X1 U83 ( .A(n116), .B(\mult_x_1/n286 ), .ZN(n49) );
  NOR2_X1 U84 ( .A1(n49), .A2(n5), .ZN(n134) );
  OAI21_X1 U85 ( .B1(n52), .B2(n51), .A(n50), .ZN(n54) );
  NAND2_X1 U86 ( .A1(n52), .A2(n51), .ZN(n53) );
  NAND2_X1 U87 ( .A1(n54), .A2(n53), .ZN(n133) );
  XNOR2_X1 U88 ( .A(n55), .B(n222), .ZN(n187) );
  NAND2_X1 U89 ( .A1(n187), .A2(n186), .ZN(n56) );
  BUF_X4 U90 ( .A(en), .Z(n266) );
  NAND2_X1 U91 ( .A1(n56), .A2(n266), .ZN(n59) );
  INV_X1 U92 ( .A(n266), .ZN(n57) );
  NAND2_X1 U93 ( .A1(n57), .A2(n333), .ZN(n58) );
  NAND2_X1 U94 ( .A1(n59), .A2(n58), .ZN(n367) );
  XNOR2_X1 U117 ( .A(n116), .B(\mult_x_1/n282 ), .ZN(n61) );
  NOR2_X1 U118 ( .A1(n61), .A2(n5), .ZN(n111) );
  XNOR2_X1 U119 ( .A(n12), .B(\mult_x_1/n281 ), .ZN(n62) );
  XNOR2_X1 U120 ( .A(n63), .B(n12), .ZN(n112) );
  OAI22_X1 U121 ( .A1(n113), .A2(n62), .B1(n112), .B2(n114), .ZN(n121) );
  INV_X1 U122 ( .A(n121), .ZN(n110) );
  XNOR2_X1 U123 ( .A(n12), .B(\mult_x_1/n282 ), .ZN(n67) );
  OAI22_X1 U124 ( .A1(n113), .A2(n67), .B1(n114), .B2(n62), .ZN(n71) );
  XNOR2_X1 U125 ( .A(n63), .B(n315), .ZN(n65) );
  AOI21_X1 U126 ( .B1(n104), .B2(n177), .A(n65), .ZN(n64) );
  INV_X1 U127 ( .A(n64), .ZN(n70) );
  XNOR2_X1 U128 ( .A(n315), .B(\mult_x_1/n281 ), .ZN(n84) );
  OAI22_X1 U129 ( .A1(n104), .A2(n84), .B1(n65), .B2(n177), .ZN(n69) );
  XNOR2_X1 U130 ( .A(n116), .B(\mult_x_1/n284 ), .ZN(n66) );
  NOR2_X1 U131 ( .A1(n66), .A2(n5), .ZN(n78) );
  XNOR2_X1 U132 ( .A(n12), .B(\mult_x_1/n283 ), .ZN(n79) );
  OAI22_X1 U133 ( .A1(n113), .A2(n79), .B1(n114), .B2(n67), .ZN(n77) );
  INV_X1 U134 ( .A(n69), .ZN(n76) );
  XNOR2_X1 U135 ( .A(n116), .B(\mult_x_1/n283 ), .ZN(n68) );
  NOR2_X1 U136 ( .A1(n68), .A2(n5), .ZN(n74) );
  FA_X1 U137 ( .A(n71), .B(n70), .CI(n69), .CO(n109), .S(n73) );
  OR2_X1 U138 ( .A1(n128), .A2(n127), .ZN(n72) );
  MUX2_X1 U139 ( .A(n321), .B(n72), .S(n266), .Z(n343) );
  FA_X1 U140 ( .A(n75), .B(n74), .CI(n73), .CO(n127), .S(n184) );
  FA_X1 U141 ( .A(n78), .B(n77), .CI(n76), .CO(n75), .S(n132) );
  OAI22_X1 U142 ( .A1(n113), .A2(n80), .B1(n114), .B2(n79), .ZN(n138) );
  AOI21_X1 U143 ( .B1(n200), .B2(n198), .A(n81), .ZN(n82) );
  INV_X1 U144 ( .A(n82), .ZN(n136) );
  XNOR2_X1 U145 ( .A(n116), .B(\mult_x_1/n285 ), .ZN(n83) );
  NOR2_X1 U146 ( .A1(n83), .A2(n5), .ZN(n141) );
  OAI22_X1 U147 ( .A1(n104), .A2(n85), .B1(n177), .B2(n84), .ZN(n140) );
  OAI21_X1 U148 ( .B1(n88), .B2(n87), .A(n86), .ZN(n90) );
  NAND2_X1 U149 ( .A1(n14), .A2(n87), .ZN(n89) );
  NAND2_X1 U150 ( .A1(n90), .A2(n89), .ZN(n139) );
  OR2_X1 U151 ( .A1(n184), .A2(n183), .ZN(n91) );
  MUX2_X1 U152 ( .A(n322), .B(n91), .S(n266), .Z(n345) );
  XNOR2_X1 U153 ( .A(n203), .B(\mult_x_1/n283 ), .ZN(n166) );
  XNOR2_X1 U154 ( .A(n203), .B(\mult_x_1/n282 ), .ZN(n97) );
  OAI22_X1 U155 ( .A1(n204), .A2(n166), .B1(n97), .B2(n16), .ZN(n107) );
  INV_X1 U156 ( .A(n114), .ZN(n92) );
  AND2_X1 U157 ( .A1(\mult_x_1/n288 ), .A2(n92), .ZN(n106) );
  XNOR2_X1 U158 ( .A(n314), .B(\mult_x_1/n285 ), .ZN(n165) );
  XNOR2_X1 U159 ( .A(n314), .B(\mult_x_1/n284 ), .ZN(n99) );
  OAI22_X1 U160 ( .A1(n198), .A2(n165), .B1(n200), .B2(n99), .ZN(n105) );
  HA_X1 U161 ( .A(n94), .B(n93), .CO(n149), .S(n153) );
  XNOR2_X1 U162 ( .A(n315), .B(\mult_x_1/n286 ), .ZN(n102) );
  OAI22_X1 U163 ( .A1(n104), .A2(n102), .B1(n177), .B2(n95), .ZN(n148) );
  OAI22_X1 U164 ( .A1(n204), .A2(n97), .B1(n96), .B2(n16), .ZN(n147) );
  OAI22_X1 U165 ( .A1(n198), .A2(n99), .B1(n200), .B2(n98), .ZN(n146) );
  OR2_X1 U166 ( .A1(\mult_x_1/n288 ), .A2(n319), .ZN(n100) );
  OAI22_X1 U167 ( .A1(n104), .A2(n319), .B1(n100), .B2(n177), .ZN(n168) );
  XNOR2_X1 U168 ( .A(n315), .B(\mult_x_1/n288 ), .ZN(n101) );
  XNOR2_X1 U169 ( .A(n315), .B(\mult_x_1/n287 ), .ZN(n103) );
  OAI22_X1 U170 ( .A1(n104), .A2(n101), .B1(n177), .B2(n103), .ZN(n167) );
  OAI22_X1 U171 ( .A1(n104), .A2(n103), .B1(n177), .B2(n102), .ZN(n163) );
  FA_X1 U172 ( .A(n107), .B(n106), .CI(n105), .CO(n154), .S(n162) );
  OR2_X1 U173 ( .A1(n160), .A2(n159), .ZN(n108) );
  MUX2_X1 U174 ( .A(n323), .B(n108), .S(n266), .Z(n347) );
  FA_X1 U175 ( .A(n111), .B(n110), .CI(n109), .CO(n123), .S(n128) );
  AOI21_X1 U176 ( .B1(n114), .B2(n113), .A(n112), .ZN(n115) );
  INV_X1 U177 ( .A(n115), .ZN(n119) );
  XNOR2_X1 U178 ( .A(n116), .B(n11), .ZN(n117) );
  NOR2_X1 U179 ( .A1(n117), .A2(n5), .ZN(n118) );
  XOR2_X1 U180 ( .A(n119), .B(n118), .Z(n120) );
  XOR2_X1 U181 ( .A(n121), .B(n120), .Z(n122) );
  OR2_X1 U182 ( .A1(n123), .A2(n122), .ZN(n125) );
  NAND2_X1 U183 ( .A1(n123), .A2(n122), .ZN(n124) );
  NAND2_X1 U184 ( .A1(n125), .A2(n124), .ZN(n126) );
  MUX2_X1 U185 ( .A(n324), .B(n126), .S(n266), .Z(n349) );
  NAND2_X1 U186 ( .A1(n128), .A2(n127), .ZN(n129) );
  MUX2_X1 U187 ( .A(n325), .B(n129), .S(n266), .Z(n351) );
  FA_X1 U188 ( .A(n132), .B(n131), .CI(n130), .CO(n183), .S(n238) );
  FA_X1 U189 ( .A(n135), .B(n134), .CI(n133), .CO(n220), .S(n222) );
  FA_X1 U190 ( .A(n138), .B(n15), .CI(n136), .CO(n131), .S(n219) );
  FA_X1 U191 ( .A(n141), .B(n140), .CI(n139), .CO(n130), .S(n218) );
  NAND2_X1 U192 ( .A1(n238), .A2(n237), .ZN(n142) );
  MUX2_X1 U193 ( .A(n326), .B(n142), .S(n266), .Z(n353) );
  FA_X1 U194 ( .A(n143), .B(n144), .CI(n145), .CO(n39), .S(n235) );
  FA_X1 U195 ( .A(n148), .B(n147), .CI(n146), .CO(n234), .S(n152) );
  FA_X1 U196 ( .A(n151), .B(n150), .CI(n149), .CO(n230), .S(n233) );
  FA_X1 U197 ( .A(n154), .B(n153), .CI(n152), .CO(n156), .S(n160) );
  NOR2_X1 U198 ( .A1(n157), .A2(n156), .ZN(n155) );
  MUX2_X1 U199 ( .A(n327), .B(n155), .S(n266), .Z(n355) );
  NAND2_X1 U200 ( .A1(n157), .A2(n156), .ZN(n158) );
  MUX2_X1 U201 ( .A(n328), .B(n158), .S(n266), .Z(n357) );
  NAND2_X1 U202 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2_X1 U203 ( .A(n329), .B(n161), .S(n266), .Z(n359) );
  FA_X1 U204 ( .A(n164), .B(n163), .CI(n162), .CO(n159), .S(n171) );
  XNOR2_X1 U205 ( .A(n314), .B(\mult_x_1/n286 ), .ZN(n179) );
  OAI22_X1 U206 ( .A1(n198), .A2(n179), .B1(n200), .B2(n165), .ZN(n175) );
  XNOR2_X1 U207 ( .A(n203), .B(\mult_x_1/n284 ), .ZN(n176) );
  OAI22_X1 U208 ( .A1(n204), .A2(n176), .B1(n166), .B2(n16), .ZN(n174) );
  HA_X1 U209 ( .A(n168), .B(n167), .CO(n164), .S(n173) );
  NOR2_X1 U210 ( .A1(n171), .A2(n170), .ZN(n169) );
  MUX2_X1 U211 ( .A(n330), .B(n169), .S(n266), .Z(n361) );
  NAND2_X1 U212 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U213 ( .A(n331), .B(n172), .S(n266), .Z(n363) );
  FA_X1 U214 ( .A(n175), .B(n174), .CI(n173), .CO(n170), .S(n181) );
  XNOR2_X1 U215 ( .A(n203), .B(\mult_x_1/n285 ), .ZN(n194) );
  OAI22_X1 U216 ( .A1(n204), .A2(n194), .B1(n176), .B2(n16), .ZN(n191) );
  INV_X1 U217 ( .A(n177), .ZN(n178) );
  AND2_X1 U218 ( .A1(\mult_x_1/n288 ), .A2(n178), .ZN(n190) );
  XNOR2_X1 U219 ( .A(n314), .B(\mult_x_1/n287 ), .ZN(n192) );
  OAI22_X1 U220 ( .A1(n198), .A2(n192), .B1(n200), .B2(n179), .ZN(n189) );
  OR2_X1 U221 ( .A1(n181), .A2(n180), .ZN(n215) );
  NAND2_X1 U222 ( .A1(n181), .A2(n180), .ZN(n213) );
  NAND2_X1 U223 ( .A1(n215), .A2(n213), .ZN(n182) );
  MUX2_X1 U224 ( .A(n332), .B(n182), .S(n266), .Z(n365) );
  NAND2_X1 U225 ( .A1(n184), .A2(n183), .ZN(n185) );
  MUX2_X1 U226 ( .A(n334), .B(n185), .S(n266), .Z(n369) );
  NOR2_X1 U227 ( .A1(n187), .A2(n186), .ZN(n188) );
  MUX2_X1 U228 ( .A(n336), .B(n188), .S(n266), .Z(n373) );
  FA_X1 U229 ( .A(n191), .B(n190), .CI(n189), .CO(n180), .S(n212) );
  XNOR2_X1 U230 ( .A(n314), .B(\mult_x_1/n288 ), .ZN(n193) );
  OAI22_X1 U231 ( .A1(n198), .A2(n193), .B1(n200), .B2(n192), .ZN(n196) );
  XNOR2_X1 U232 ( .A(n203), .B(\mult_x_1/n286 ), .ZN(n199) );
  OAI22_X1 U233 ( .A1(n204), .A2(n199), .B1(n194), .B2(n16), .ZN(n195) );
  NOR2_X1 U234 ( .A1(n212), .A2(n211), .ZN(n257) );
  HA_X1 U235 ( .A(n196), .B(n195), .CO(n211), .S(n209) );
  OR2_X1 U236 ( .A1(\mult_x_1/n288 ), .A2(n18), .ZN(n197) );
  OAI22_X1 U237 ( .A1(n198), .A2(n18), .B1(n197), .B2(n200), .ZN(n208) );
  OR2_X1 U238 ( .A1(n209), .A2(n208), .ZN(n253) );
  XNOR2_X1 U239 ( .A(n203), .B(\mult_x_1/n287 ), .ZN(n202) );
  OAI22_X1 U240 ( .A1(n204), .A2(n202), .B1(n199), .B2(n16), .ZN(n207) );
  INV_X1 U241 ( .A(n200), .ZN(n201) );
  AND2_X1 U242 ( .A1(\mult_x_1/n288 ), .A2(n201), .ZN(n206) );
  NOR2_X1 U243 ( .A1(n207), .A2(n206), .ZN(n246) );
  OAI22_X1 U244 ( .A1(n204), .A2(\mult_x_1/n288 ), .B1(n202), .B2(n16), .ZN(
        n243) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n205) );
  NAND2_X1 U246 ( .A1(n205), .A2(n204), .ZN(n242) );
  NAND2_X1 U247 ( .A1(n243), .A2(n242), .ZN(n249) );
  NAND2_X1 U248 ( .A1(n207), .A2(n206), .ZN(n247) );
  OAI21_X1 U249 ( .B1(n246), .B2(n249), .A(n247), .ZN(n254) );
  NAND2_X1 U250 ( .A1(n209), .A2(n208), .ZN(n252) );
  INV_X1 U251 ( .A(n252), .ZN(n210) );
  AOI21_X1 U252 ( .B1(n253), .B2(n254), .A(n210), .ZN(n260) );
  NAND2_X1 U253 ( .A1(n212), .A2(n211), .ZN(n258) );
  OAI21_X1 U254 ( .B1(n257), .B2(n260), .A(n258), .ZN(n217) );
  INV_X1 U255 ( .A(n213), .ZN(n214) );
  AOI21_X1 U256 ( .B1(n215), .B2(n217), .A(n214), .ZN(n216) );
  MUX2_X1 U257 ( .A(n337), .B(n216), .S(n266), .Z(n375) );
  MUX2_X1 U258 ( .A(n338), .B(n217), .S(n266), .Z(n377) );
  FA_X1 U259 ( .A(n220), .B(n219), .CI(n218), .CO(n237), .S(n221) );
  MUX2_X1 U260 ( .A(n339), .B(n221), .S(n266), .Z(n379) );
  NAND2_X1 U261 ( .A1(n222), .A2(n224), .ZN(n227) );
  NAND2_X1 U262 ( .A1(n222), .A2(n223), .ZN(n226) );
  NAND2_X1 U263 ( .A1(n224), .A2(n223), .ZN(n225) );
  NAND3_X1 U264 ( .A1(n227), .A2(n226), .A3(n225), .ZN(n228) );
  MUX2_X1 U265 ( .A(n340), .B(n228), .S(n266), .Z(n381) );
  FA_X1 U266 ( .A(n231), .B(n230), .CI(n229), .CO(n186), .S(n232) );
  MUX2_X1 U267 ( .A(n341), .B(n232), .S(n266), .Z(n383) );
  MUX2_X1 U268 ( .A(n342), .B(n236), .S(n266), .Z(n385) );
  OAI21_X1 U269 ( .B1(n238), .B2(n237), .A(n266), .ZN(n240) );
  OR2_X1 U270 ( .A1(n266), .A2(n389), .ZN(n239) );
  NAND2_X1 U271 ( .A1(n240), .A2(n239), .ZN(n371) );
  MUX2_X1 U272 ( .A(product[0]), .B(n506), .S(n266), .Z(n398) );
  MUX2_X1 U273 ( .A(n506), .B(n507), .S(n266), .Z(n400) );
  AND2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n241) );
  MUX2_X1 U275 ( .A(n507), .B(n241), .S(n266), .Z(n402) );
  MUX2_X1 U276 ( .A(product[1]), .B(n509), .S(n266), .Z(n404) );
  MUX2_X1 U277 ( .A(n509), .B(n510), .S(n266), .Z(n406) );
  OR2_X1 U278 ( .A1(n243), .A2(n242), .ZN(n244) );
  AND2_X1 U279 ( .A1(n244), .A2(n249), .ZN(n245) );
  MUX2_X1 U280 ( .A(n510), .B(n245), .S(n266), .Z(n408) );
  MUX2_X1 U281 ( .A(product[2]), .B(n512), .S(n266), .Z(n410) );
  MUX2_X1 U282 ( .A(n512), .B(n513), .S(n266), .Z(n412) );
  INV_X1 U283 ( .A(n246), .ZN(n248) );
  NAND2_X1 U284 ( .A1(n248), .A2(n247), .ZN(n250) );
  XOR2_X1 U285 ( .A(n250), .B(n249), .Z(n251) );
  MUX2_X1 U286 ( .A(n513), .B(n251), .S(n266), .Z(n414) );
  MUX2_X1 U287 ( .A(product[3]), .B(n515), .S(n266), .Z(n416) );
  MUX2_X1 U288 ( .A(n515), .B(n516), .S(n266), .Z(n418) );
  NAND2_X1 U289 ( .A1(n253), .A2(n252), .ZN(n255) );
  XNOR2_X1 U290 ( .A(n255), .B(n254), .ZN(n256) );
  MUX2_X1 U291 ( .A(n516), .B(n256), .S(n266), .Z(n420) );
  MUX2_X1 U292 ( .A(product[4]), .B(n518), .S(n266), .Z(n422) );
  MUX2_X1 U293 ( .A(n518), .B(n519), .S(n266), .Z(n424) );
  INV_X1 U294 ( .A(n257), .ZN(n259) );
  NAND2_X1 U295 ( .A1(n259), .A2(n258), .ZN(n261) );
  XOR2_X1 U296 ( .A(n261), .B(n260), .Z(n262) );
  MUX2_X1 U297 ( .A(n519), .B(n262), .S(n266), .Z(n426) );
  MUX2_X1 U298 ( .A(product[5]), .B(n521), .S(n266), .Z(n428) );
  XNOR2_X1 U299 ( .A(n332), .B(n338), .ZN(n263) );
  MUX2_X1 U300 ( .A(n521), .B(n263), .S(n266), .Z(n430) );
  MUX2_X1 U301 ( .A(product[6]), .B(n523), .S(n266), .Z(n432) );
  NAND2_X1 U302 ( .A1(n390), .A2(n331), .ZN(n264) );
  XOR2_X1 U303 ( .A(n264), .B(n337), .Z(n265) );
  MUX2_X1 U304 ( .A(n523), .B(n265), .S(n266), .Z(n434) );
  MUX2_X1 U305 ( .A(product[7]), .B(n525), .S(n266), .Z(n436) );
  OAI21_X1 U306 ( .B1(n330), .B2(n337), .A(n331), .ZN(n269) );
  NAND2_X1 U307 ( .A1(n323), .A2(n329), .ZN(n267) );
  XNOR2_X1 U308 ( .A(n269), .B(n267), .ZN(n268) );
  BUF_X2 U309 ( .A(en), .Z(n317) );
  MUX2_X1 U310 ( .A(n525), .B(n268), .S(n317), .Z(n438) );
  MUX2_X1 U311 ( .A(product[8]), .B(n527), .S(n317), .Z(n440) );
  AOI21_X1 U312 ( .B1(n269), .B2(n323), .A(n391), .ZN(n272) );
  NAND2_X1 U313 ( .A1(n392), .A2(n328), .ZN(n270) );
  XOR2_X1 U314 ( .A(n272), .B(n270), .Z(n271) );
  MUX2_X1 U315 ( .A(n527), .B(n271), .S(n317), .Z(n442) );
  MUX2_X1 U316 ( .A(product[9]), .B(n529), .S(n317), .Z(n444) );
  OAI21_X1 U317 ( .B1(n272), .B2(n327), .A(n328), .ZN(n283) );
  INV_X1 U318 ( .A(n283), .ZN(n276) );
  NOR2_X1 U319 ( .A1(n341), .A2(n342), .ZN(n280) );
  INV_X1 U320 ( .A(n280), .ZN(n273) );
  NAND2_X1 U321 ( .A1(n341), .A2(n342), .ZN(n281) );
  NAND2_X1 U322 ( .A1(n273), .A2(n281), .ZN(n274) );
  XOR2_X1 U323 ( .A(n276), .B(n274), .Z(n275) );
  MUX2_X1 U324 ( .A(n529), .B(n275), .S(n317), .Z(n446) );
  MUX2_X1 U325 ( .A(product[10]), .B(n531), .S(n317), .Z(n448) );
  OAI21_X1 U326 ( .B1(n276), .B2(n280), .A(n281), .ZN(n278) );
  NAND2_X1 U327 ( .A1(n393), .A2(n333), .ZN(n277) );
  XNOR2_X1 U328 ( .A(n278), .B(n277), .ZN(n279) );
  MUX2_X1 U329 ( .A(n531), .B(n279), .S(n317), .Z(n450) );
  MUX2_X1 U330 ( .A(product[11]), .B(n533), .S(n317), .Z(n452) );
  NOR2_X1 U331 ( .A1(n336), .A2(n280), .ZN(n284) );
  OAI21_X1 U332 ( .B1(n336), .B2(n281), .A(n333), .ZN(n282) );
  AOI21_X1 U333 ( .B1(n284), .B2(n283), .A(n282), .ZN(n311) );
  NOR2_X1 U334 ( .A1(n339), .A2(n340), .ZN(n287) );
  INV_X1 U335 ( .A(n287), .ZN(n306) );
  NAND2_X1 U336 ( .A1(n339), .A2(n340), .ZN(n298) );
  NAND2_X1 U337 ( .A1(n306), .A2(n298), .ZN(n285) );
  XOR2_X1 U338 ( .A(n311), .B(n285), .Z(n286) );
  MUX2_X1 U339 ( .A(n533), .B(n286), .S(n317), .Z(n454) );
  MUX2_X1 U340 ( .A(product[12]), .B(n535), .S(n317), .Z(n456) );
  OAI21_X1 U341 ( .B1(n311), .B2(n287), .A(n298), .ZN(n289) );
  NAND2_X1 U342 ( .A1(n335), .A2(n326), .ZN(n288) );
  XNOR2_X1 U343 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U344 ( .A(n535), .B(n290), .S(n317), .Z(n458) );
  MUX2_X1 U345 ( .A(product[13]), .B(n537), .S(n317), .Z(n460) );
  NAND2_X1 U346 ( .A1(n306), .A2(n335), .ZN(n293) );
  INV_X1 U347 ( .A(n298), .ZN(n291) );
  AOI21_X1 U348 ( .B1(n291), .B2(n335), .A(n394), .ZN(n292) );
  OAI21_X1 U349 ( .B1(n311), .B2(n293), .A(n292), .ZN(n295) );
  NAND2_X1 U350 ( .A1(n322), .A2(n334), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n296) );
  MUX2_X1 U352 ( .A(n537), .B(n296), .S(n317), .Z(n462) );
  MUX2_X1 U353 ( .A(product[14]), .B(n539), .S(n317), .Z(n464) );
  NAND2_X1 U354 ( .A1(n335), .A2(n322), .ZN(n299) );
  INV_X1 U355 ( .A(n299), .ZN(n305) );
  NAND2_X1 U356 ( .A1(n306), .A2(n305), .ZN(n301) );
  AOI21_X1 U357 ( .B1(n394), .B2(n322), .A(n388), .ZN(n297) );
  OAI21_X1 U358 ( .B1(n299), .B2(n298), .A(n297), .ZN(n308) );
  INV_X1 U359 ( .A(n308), .ZN(n300) );
  OAI21_X1 U360 ( .B1(n311), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U361 ( .A1(n321), .A2(n325), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U363 ( .A(n539), .B(n304), .S(n317), .Z(n466) );
  MUX2_X1 U364 ( .A(product[15]), .B(n541), .S(n317), .Z(n468) );
  AND2_X1 U365 ( .A1(n321), .A2(n305), .ZN(n307) );
  NAND2_X1 U366 ( .A1(n307), .A2(n306), .ZN(n310) );
  AOI21_X1 U367 ( .B1(n308), .B2(n321), .A(n387), .ZN(n309) );
  OAI21_X1 U368 ( .B1(n311), .B2(n310), .A(n309), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n312), .B(n324), .ZN(n313) );
  MUX2_X1 U370 ( .A(n541), .B(n313), .S(n317), .Z(n470) );
  MUX2_X1 U371 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n317), .Z(n472) );
  MUX2_X1 U372 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n317), .Z(n474) );
  MUX2_X1 U373 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n317), .Z(n476) );
  MUX2_X1 U374 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n317), .Z(n478) );
  MUX2_X1 U375 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n317), .Z(n480) );
  MUX2_X1 U376 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n317), .Z(n482) );
  MUX2_X1 U377 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n317), .Z(n484) );
  MUX2_X1 U378 ( .A(n11), .B(B_extended[7]), .S(n317), .Z(n486) );
  MUX2_X1 U379 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n317), .Z(n488) );
  MUX2_X1 U380 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n317), .Z(n490) );
  MUX2_X1 U381 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n317), .Z(n492) );
  MUX2_X1 U382 ( .A(n314), .B(A_extended[3]), .S(n317), .Z(n494) );
  MUX2_X1 U383 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n317), .Z(n496) );
  MUX2_X1 U384 ( .A(n315), .B(A_extended[5]), .S(n317), .Z(n498) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n317), .Z(n500) );
  MUX2_X1 U386 ( .A(n12), .B(A_extended[7]), .S(n317), .Z(n502) );
  OR2_X1 U387 ( .A1(n317), .A2(n544), .ZN(n504) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_6 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n342, n344, n346, n348, n350, n352, n354,
         n356, n358, n360, n362, n364, n366, n368, n370, n372, n374, n376,
         n378, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n393, n395, n397, n399, n401, n403, n405, n407, n409,
         n411, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n504, n506, n507, n509, n510, n512, n513, n515,
         n516, n518, n519, n521, n523, n525, n527, n529, n531, n533, n535,
         n537, n539, n540, n541, n542;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n391), .SE(n501), .CK(clk), .Q(n541), 
        .QN(n35) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n391), .SE(n497), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n32) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n391), .SE(n495), .CK(clk), .Q(n540), 
        .QN(n24) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n391), .SE(n493), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n391), .SE(n489), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n391), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n21) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n391), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n23) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n391), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n391), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n27) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n390), .SE(n477), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n391), .SE(n475), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n28) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n391), .SE(n473), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n30) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n390), .SE(n471), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n29) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n390), .SE(n469), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n22) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n391), .SE(n467), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n391), .SE(n465), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n391), .SE(n463), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n390), .SE(n461), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n391), .SE(n459), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n391), .SE(n457), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n391), .SE(n455), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n391), .SE(n453), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n391), .SE(n451), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n390), .SE(n449), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG23_S3 ( .D(1'b0), .SI(n390), .SE(n447), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG24_S4 ( .D(1'b0), .SI(n391), .SE(n445), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG21_S3 ( .D(1'b0), .SI(n391), .SE(n443), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG22_S4 ( .D(1'b0), .SI(n390), .SE(n441), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n391), .SE(n439), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n391), .SE(n437), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n391), .SE(n435), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n391), .SE(n433), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n391), .SE(n431), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n390), .SE(n429), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n391), .SE(n427), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n391), .SE(n425), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n390), .SE(n423), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n391), .SE(n421), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n391), .SE(n419), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n390), .SE(n417), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n391), .SE(n415), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n390), .SE(n413), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n390), .SE(n411), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n390), .SE(n409), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n390), .SE(n407), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n390), .SE(n405), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n390), .SE(n403), .CK(clk), .Q(n507)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n390), .SE(n401), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n390), .SE(n399), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n390), .SE(n397), .CK(clk), .Q(n504)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n390), .SE(n395), .CK(clk), .Q(n503)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n390), .SE(n393), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n391), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n34) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n391), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n319) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n542), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n542), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n338), .QN(n382) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n542), .SE(n374), .CK(
        clk), .Q(n386), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n542), .SE(n372), .CK(
        clk), .Q(n388), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n542), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n542), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n334), .QN(n381) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n542), .SE(n366), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n542), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n542), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n331), .QN(n383) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n542), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n330), .QN(n384) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n542), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n542), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n328), .QN(n385) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n542), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n542), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n326), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n542), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n325), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n542), .SI(1'b1), .SE(n348), .CK(clk), 
        .Q(n324), .QN(n380) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n542), .SE(n346), .CK(
        clk), .QN(n323) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n542), .SE(n344), .CK(
        clk), .QN(n322) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n542), .SI(1'b1), .SE(n342), .CK(clk), 
        .Q(n321) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n542), .SI(1'b1), .SE(n340), .CK(clk), 
        .Q(n320) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n391), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n318) );
  NAND2_X2 U2 ( .A1(n41), .A2(n40), .ZN(n124) );
  AND3_X1 U3 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n223) );
  BUF_X1 U4 ( .A(n100), .Z(n6) );
  NAND2_X1 U5 ( .A1(n36), .A2(n37), .ZN(n118) );
  NAND2_X2 U6 ( .A1(n21), .A2(\mult_x_1/n313 ), .ZN(n199) );
  AND2_X2 U7 ( .A1(n541), .A2(\mult_x_1/n281 ), .ZN(n95) );
  NOR2_X1 U8 ( .A1(n172), .A2(n171), .ZN(n102) );
  NAND2_X1 U9 ( .A1(n172), .A2(n171), .ZN(n101) );
  XNOR2_X1 U10 ( .A(n108), .B(n107), .ZN(n109) );
  BUF_X2 U11 ( .A(n51), .Z(n5) );
  XOR2_X1 U12 ( .A(n222), .B(n221), .Z(n7) );
  XOR2_X1 U13 ( .A(n220), .B(n7), .Z(n134) );
  NAND2_X1 U14 ( .A1(n220), .A2(n222), .ZN(n8) );
  NAND2_X1 U15 ( .A1(n220), .A2(n221), .ZN(n9) );
  NAND2_X1 U16 ( .A1(n222), .A2(n221), .ZN(n10) );
  BUF_X8 U17 ( .A(en), .Z(n317) );
  BUF_X2 U18 ( .A(n40), .Z(n11) );
  OAI22_X1 U19 ( .A1(n124), .A2(n85), .B1(n43), .B2(n11), .ZN(n12) );
  XNOR2_X1 U20 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n40) );
  OAI22_X1 U21 ( .A1(n20), .A2(n125), .B1(n5), .B2(n99), .ZN(n13) );
  XNOR2_X1 U22 ( .A(n319), .B(\mult_x_1/a[2] ), .ZN(n50) );
  OR2_X1 U23 ( .A1(n164), .A2(n13), .ZN(n172) );
  XOR2_X1 U24 ( .A(n169), .B(n170), .Z(n14) );
  XOR2_X1 U25 ( .A(n168), .B(n14), .Z(n231) );
  NAND2_X1 U26 ( .A1(n168), .A2(n169), .ZN(n15) );
  NAND2_X1 U27 ( .A1(n168), .A2(n170), .ZN(n16) );
  NAND2_X1 U28 ( .A1(n169), .A2(n170), .ZN(n17) );
  NAND3_X1 U29 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n110) );
  OAI22_X1 U30 ( .A1(n6), .A2(n99), .B1(n82), .B2(n5), .ZN(n18) );
  INV_X1 U31 ( .A(n100), .ZN(n19) );
  INV_X1 U32 ( .A(n19), .ZN(n20) );
  BUF_X1 U33 ( .A(rst_n), .Z(n390) );
  INV_X1 U34 ( .A(rst_n), .ZN(n542) );
  AND2_X1 U35 ( .A1(n219), .A2(n218), .ZN(n31) );
  XOR2_X1 U36 ( .A(n219), .B(n218), .Z(n33) );
  INV_X2 U57 ( .A(n318), .ZN(n316) );
  NAND2_X1 U58 ( .A1(n35), .A2(n316), .ZN(n112) );
  NOR2_X1 U59 ( .A1(n25), .A2(n112), .ZN(n66) );
  XNOR2_X1 U60 ( .A(n32), .B(\mult_x_1/n310 ), .ZN(n36) );
  XNOR2_X1 U61 ( .A(\mult_x_1/a[6] ), .B(n540), .ZN(n37) );
  XNOR2_X1 U62 ( .A(n316), .B(\mult_x_1/n281 ), .ZN(n39) );
  XNOR2_X1 U63 ( .A(n95), .B(n316), .ZN(n67) );
  INV_X1 U64 ( .A(n37), .ZN(n38) );
  INV_X2 U65 ( .A(n38), .ZN(n116) );
  OAI22_X1 U66 ( .A1(n118), .A2(n39), .B1(n67), .B2(n116), .ZN(n72) );
  INV_X1 U67 ( .A(n72), .ZN(n65) );
  XNOR2_X1 U68 ( .A(n316), .B(\mult_x_1/n282 ), .ZN(n44) );
  OAI22_X1 U69 ( .A1(n118), .A2(n44), .B1(n116), .B2(n39), .ZN(n47) );
  XOR2_X1 U70 ( .A(\mult_x_1/a[4] ), .B(n540), .Z(n41) );
  BUF_X2 U71 ( .A(n540), .Z(n315) );
  XNOR2_X1 U72 ( .A(n95), .B(n315), .ZN(n43) );
  AOI21_X1 U73 ( .B1(n11), .B2(n124), .A(n43), .ZN(n42) );
  INV_X1 U74 ( .A(n42), .ZN(n46) );
  XNOR2_X1 U75 ( .A(n315), .B(\mult_x_1/n281 ), .ZN(n85) );
  OAI22_X1 U76 ( .A1(n124), .A2(n85), .B1(n43), .B2(n11), .ZN(n45) );
  INV_X1 U77 ( .A(n45), .ZN(n94) );
  XNOR2_X1 U78 ( .A(n316), .B(\mult_x_1/n283 ), .ZN(n81) );
  OAI22_X1 U79 ( .A1(n118), .A2(n81), .B1(n116), .B2(n44), .ZN(n93) );
  NOR2_X1 U80 ( .A1(n26), .A2(n112), .ZN(n92) );
  NOR2_X1 U81 ( .A1(n27), .A2(n112), .ZN(n151) );
  FA_X1 U82 ( .A(n47), .B(n46), .CI(n12), .CO(n64), .S(n150) );
  OR2_X1 U83 ( .A1(n79), .A2(n78), .ZN(n48) );
  MUX2_X1 U84 ( .A(n320), .B(n48), .S(n317), .Z(n340) );
  BUF_X2 U85 ( .A(\mult_x_1/n313 ), .Z(n198) );
  XNOR2_X1 U86 ( .A(n198), .B(\mult_x_1/n283 ), .ZN(n143) );
  XNOR2_X1 U87 ( .A(n198), .B(\mult_x_1/n282 ), .ZN(n54) );
  OAI22_X1 U88 ( .A1(n199), .A2(n143), .B1(n54), .B2(n21), .ZN(n62) );
  INV_X1 U89 ( .A(n116), .ZN(n49) );
  AND2_X1 U90 ( .A1(\mult_x_1/n288 ), .A2(n49), .ZN(n61) );
  XNOR2_X1 U91 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n51) );
  NAND2_X1 U92 ( .A1(n51), .A2(n50), .ZN(n100) );
  BUF_X2 U93 ( .A(\mult_x_1/n312 ), .Z(n193) );
  XNOR2_X1 U94 ( .A(n193), .B(\mult_x_1/n285 ), .ZN(n142) );
  XNOR2_X1 U95 ( .A(n193), .B(\mult_x_1/n284 ), .ZN(n55) );
  OAI22_X1 U96 ( .A1(n6), .A2(n142), .B1(n5), .B2(n55), .ZN(n60) );
  OR2_X1 U97 ( .A1(\mult_x_1/n288 ), .A2(n318), .ZN(n52) );
  OAI22_X1 U98 ( .A1(n118), .A2(n318), .B1(n52), .B2(n116), .ZN(n128) );
  XNOR2_X1 U99 ( .A(n316), .B(\mult_x_1/n288 ), .ZN(n53) );
  XNOR2_X1 U100 ( .A(n316), .B(\mult_x_1/n287 ), .ZN(n117) );
  OAI22_X1 U101 ( .A1(n118), .A2(n53), .B1(n116), .B2(n117), .ZN(n127) );
  XNOR2_X1 U102 ( .A(n315), .B(\mult_x_1/n286 ), .ZN(n58) );
  XNOR2_X1 U103 ( .A(n315), .B(\mult_x_1/n285 ), .ZN(n123) );
  OAI22_X1 U104 ( .A1(n124), .A2(n58), .B1(n11), .B2(n123), .ZN(n121) );
  XNOR2_X1 U105 ( .A(n198), .B(\mult_x_1/n281 ), .ZN(n114) );
  OAI22_X1 U106 ( .A1(n199), .A2(n54), .B1(n114), .B2(n21), .ZN(n120) );
  XNOR2_X1 U107 ( .A(n193), .B(\mult_x_1/n283 ), .ZN(n126) );
  OAI22_X1 U108 ( .A1(n6), .A2(n55), .B1(n5), .B2(n126), .ZN(n119) );
  OR2_X1 U109 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n56) );
  OAI22_X1 U110 ( .A1(n124), .A2(n24), .B1(n56), .B2(n11), .ZN(n145) );
  XNOR2_X1 U111 ( .A(n315), .B(\mult_x_1/n288 ), .ZN(n57) );
  XNOR2_X1 U112 ( .A(n315), .B(\mult_x_1/n287 ), .ZN(n59) );
  OAI22_X1 U113 ( .A1(n124), .A2(n57), .B1(n11), .B2(n59), .ZN(n144) );
  AND2_X1 U114 ( .A1(n145), .A2(n144), .ZN(n141) );
  OAI22_X1 U115 ( .A1(n124), .A2(n59), .B1(n11), .B2(n58), .ZN(n140) );
  FA_X1 U116 ( .A(n62), .B(n61), .CI(n60), .CO(n131), .S(n139) );
  OR2_X1 U117 ( .A1(n137), .A2(n136), .ZN(n63) );
  MUX2_X1 U118 ( .A(n322), .B(n63), .S(n317), .Z(n344) );
  FA_X1 U119 ( .A(n66), .B(n65), .CI(n64), .CO(n74), .S(n79) );
  AOI21_X1 U120 ( .B1(n116), .B2(n118), .A(n67), .ZN(n68) );
  INV_X1 U121 ( .A(n68), .ZN(n70) );
  NOR2_X1 U122 ( .A1(n23), .A2(n112), .ZN(n69) );
  XOR2_X1 U123 ( .A(n70), .B(n69), .Z(n71) );
  XOR2_X1 U124 ( .A(n72), .B(n71), .Z(n73) );
  OR2_X1 U125 ( .A1(n74), .A2(n73), .ZN(n76) );
  NAND2_X1 U126 ( .A1(n74), .A2(n73), .ZN(n75) );
  NAND2_X1 U127 ( .A1(n76), .A2(n75), .ZN(n77) );
  MUX2_X1 U128 ( .A(n323), .B(n77), .S(n317), .Z(n346) );
  NAND2_X1 U129 ( .A1(n79), .A2(n78), .ZN(n80) );
  MUX2_X1 U130 ( .A(n324), .B(n80), .S(n317), .Z(n348) );
  XNOR2_X1 U131 ( .A(n316), .B(\mult_x_1/n284 ), .ZN(n84) );
  OAI22_X1 U132 ( .A1(n118), .A2(n84), .B1(n116), .B2(n81), .ZN(n106) );
  XNOR2_X1 U133 ( .A(n193), .B(\mult_x_1/n281 ), .ZN(n99) );
  XNOR2_X1 U134 ( .A(n95), .B(n193), .ZN(n82) );
  OAI22_X1 U135 ( .A1(n20), .A2(n99), .B1(n82), .B2(n5), .ZN(n105) );
  AOI21_X1 U136 ( .B1(n5), .B2(n6), .A(n82), .ZN(n83) );
  INV_X1 U137 ( .A(n83), .ZN(n104) );
  XNOR2_X1 U138 ( .A(n316), .B(\mult_x_1/n285 ), .ZN(n97) );
  OAI22_X1 U139 ( .A1(n118), .A2(n97), .B1(n116), .B2(n84), .ZN(n170) );
  XNOR2_X1 U140 ( .A(n315), .B(\mult_x_1/n283 ), .ZN(n98) );
  XNOR2_X1 U141 ( .A(n315), .B(\mult_x_1/n282 ), .ZN(n86) );
  OAI22_X1 U142 ( .A1(n124), .A2(n98), .B1(n11), .B2(n86), .ZN(n169) );
  INV_X1 U143 ( .A(n105), .ZN(n168) );
  NOR2_X1 U144 ( .A1(n28), .A2(n112), .ZN(n108) );
  INV_X1 U145 ( .A(n108), .ZN(n88) );
  OAI22_X1 U146 ( .A1(n124), .A2(n86), .B1(n11), .B2(n85), .ZN(n107) );
  INV_X1 U147 ( .A(n107), .ZN(n87) );
  NAND2_X1 U148 ( .A1(n88), .A2(n87), .ZN(n89) );
  NAND2_X1 U149 ( .A1(n110), .A2(n89), .ZN(n91) );
  NAND2_X1 U150 ( .A1(n108), .A2(n107), .ZN(n90) );
  NAND2_X1 U151 ( .A1(n91), .A2(n90), .ZN(n154) );
  FA_X1 U152 ( .A(n94), .B(n93), .CI(n92), .CO(n152), .S(n153) );
  XNOR2_X1 U153 ( .A(n95), .B(n198), .ZN(n113) );
  AOI21_X1 U154 ( .B1(n199), .B2(n21), .A(n113), .ZN(n96) );
  INV_X1 U155 ( .A(n96), .ZN(n214) );
  XNOR2_X1 U156 ( .A(n316), .B(\mult_x_1/n286 ), .ZN(n115) );
  OAI22_X1 U157 ( .A1(n118), .A2(n115), .B1(n116), .B2(n97), .ZN(n213) );
  NOR2_X1 U158 ( .A1(n29), .A2(n112), .ZN(n212) );
  INV_X1 U159 ( .A(n173), .ZN(n103) );
  XNOR2_X1 U160 ( .A(n315), .B(\mult_x_1/n284 ), .ZN(n122) );
  OAI22_X1 U161 ( .A1(n124), .A2(n122), .B1(n11), .B2(n98), .ZN(n164) );
  XNOR2_X1 U162 ( .A(n193), .B(\mult_x_1/n282 ), .ZN(n125) );
  OAI22_X1 U163 ( .A1(n6), .A2(n125), .B1(n5), .B2(n99), .ZN(n163) );
  NOR2_X1 U164 ( .A1(n30), .A2(n112), .ZN(n171) );
  OAI21_X1 U165 ( .B1(n103), .B2(n102), .A(n101), .ZN(n162) );
  FA_X1 U166 ( .A(n106), .B(n18), .CI(n104), .CO(n155), .S(n161) );
  XNOR2_X1 U167 ( .A(n110), .B(n109), .ZN(n160) );
  NAND2_X1 U168 ( .A1(n158), .A2(n157), .ZN(n111) );
  MUX2_X1 U169 ( .A(n325), .B(n111), .S(n317), .Z(n350) );
  NOR2_X1 U170 ( .A1(n112), .A2(n22), .ZN(n167) );
  OAI22_X1 U171 ( .A1(n199), .A2(n114), .B1(n113), .B2(n21), .ZN(n166) );
  OAI22_X1 U172 ( .A1(n118), .A2(n117), .B1(n116), .B2(n115), .ZN(n165) );
  FA_X1 U173 ( .A(n121), .B(n120), .CI(n119), .CO(n221), .S(n129) );
  OAI22_X1 U174 ( .A1(n124), .A2(n123), .B1(n11), .B2(n122), .ZN(n217) );
  OAI22_X1 U175 ( .A1(n6), .A2(n126), .B1(n5), .B2(n125), .ZN(n216) );
  HA_X1 U176 ( .A(n128), .B(n127), .CO(n215), .S(n130) );
  FA_X1 U177 ( .A(n131), .B(n130), .CI(n129), .CO(n133), .S(n137) );
  NOR2_X1 U178 ( .A1(n134), .A2(n133), .ZN(n132) );
  MUX2_X1 U179 ( .A(n328), .B(n132), .S(n317), .Z(n356) );
  NAND2_X1 U180 ( .A1(n134), .A2(n133), .ZN(n135) );
  MUX2_X1 U181 ( .A(n329), .B(n135), .S(n317), .Z(n358) );
  NAND2_X1 U182 ( .A1(n137), .A2(n136), .ZN(n138) );
  MUX2_X1 U183 ( .A(n330), .B(n138), .S(n317), .Z(n360) );
  FA_X1 U184 ( .A(n141), .B(n140), .CI(n139), .CO(n136), .S(n148) );
  XNOR2_X1 U185 ( .A(n193), .B(\mult_x_1/n286 ), .ZN(n184) );
  OAI22_X1 U186 ( .A1(n6), .A2(n184), .B1(n5), .B2(n142), .ZN(n181) );
  XNOR2_X1 U187 ( .A(n198), .B(\mult_x_1/n284 ), .ZN(n182) );
  OAI22_X1 U188 ( .A1(n199), .A2(n182), .B1(n143), .B2(n21), .ZN(n180) );
  XOR2_X1 U189 ( .A(n145), .B(n144), .Z(n179) );
  NOR2_X1 U190 ( .A1(n148), .A2(n147), .ZN(n146) );
  MUX2_X1 U191 ( .A(n331), .B(n146), .S(n317), .Z(n362) );
  NAND2_X1 U192 ( .A1(n148), .A2(n147), .ZN(n149) );
  BUF_X4 U193 ( .A(en), .Z(n276) );
  MUX2_X1 U194 ( .A(n332), .B(n149), .S(n276), .Z(n364) );
  FA_X1 U195 ( .A(n152), .B(n151), .CI(n150), .CO(n78), .S(n237) );
  FA_X1 U196 ( .A(n155), .B(n154), .CI(n153), .CO(n238), .S(n158) );
  NAND2_X1 U197 ( .A1(n237), .A2(n238), .ZN(n156) );
  MUX2_X1 U198 ( .A(n334), .B(n156), .S(n276), .Z(n368) );
  OR2_X1 U199 ( .A1(n158), .A2(n157), .ZN(n159) );
  MUX2_X1 U200 ( .A(n335), .B(n159), .S(n276), .Z(n370) );
  FA_X1 U201 ( .A(n160), .B(n161), .CI(n162), .CO(n157), .S(n177) );
  XNOR2_X1 U202 ( .A(n164), .B(n163), .ZN(n219) );
  FA_X1 U203 ( .A(n167), .B(n166), .CI(n165), .CO(n218), .S(n222) );
  XNOR2_X1 U204 ( .A(n172), .B(n171), .ZN(n174) );
  XNOR2_X1 U205 ( .A(n174), .B(n173), .ZN(n230) );
  NOR2_X1 U206 ( .A1(n177), .A2(n176), .ZN(n175) );
  MUX2_X1 U207 ( .A(n337), .B(n175), .S(n276), .Z(n374) );
  NAND2_X1 U208 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2_X1 U209 ( .A(n338), .B(n178), .S(n276), .Z(n376) );
  FA_X1 U210 ( .A(n181), .B(n180), .CI(n179), .CO(n147), .S(n209) );
  XNOR2_X1 U211 ( .A(n198), .B(\mult_x_1/n285 ), .ZN(n190) );
  OAI22_X1 U212 ( .A1(n199), .A2(n190), .B1(n182), .B2(n21), .ZN(n187) );
  INV_X1 U213 ( .A(n11), .ZN(n183) );
  AND2_X1 U214 ( .A1(\mult_x_1/n288 ), .A2(n183), .ZN(n186) );
  XNOR2_X1 U215 ( .A(n193), .B(\mult_x_1/n287 ), .ZN(n188) );
  OAI22_X1 U216 ( .A1(n6), .A2(n188), .B1(n5), .B2(n184), .ZN(n185) );
  OR2_X1 U217 ( .A1(n209), .A2(n208), .ZN(n269) );
  FA_X1 U218 ( .A(n187), .B(n186), .CI(n185), .CO(n208), .S(n207) );
  XNOR2_X1 U219 ( .A(n193), .B(\mult_x_1/n288 ), .ZN(n189) );
  OAI22_X1 U220 ( .A1(n6), .A2(n189), .B1(n5), .B2(n188), .ZN(n192) );
  XNOR2_X1 U221 ( .A(n198), .B(\mult_x_1/n286 ), .ZN(n195) );
  OAI22_X1 U222 ( .A1(n199), .A2(n195), .B1(n190), .B2(n21), .ZN(n191) );
  NOR2_X1 U223 ( .A1(n207), .A2(n206), .ZN(n262) );
  HA_X1 U224 ( .A(n192), .B(n191), .CO(n206), .S(n204) );
  OR2_X1 U225 ( .A1(\mult_x_1/n288 ), .A2(n319), .ZN(n194) );
  OAI22_X1 U226 ( .A1(n319), .A2(n6), .B1(n194), .B2(n5), .ZN(n203) );
  OR2_X1 U227 ( .A1(n204), .A2(n203), .ZN(n258) );
  XNOR2_X1 U228 ( .A(n198), .B(\mult_x_1/n287 ), .ZN(n197) );
  OAI22_X1 U229 ( .A1(n199), .A2(n197), .B1(n195), .B2(n21), .ZN(n202) );
  INV_X1 U230 ( .A(n5), .ZN(n196) );
  AND2_X1 U231 ( .A1(\mult_x_1/n288 ), .A2(n196), .ZN(n201) );
  NOR2_X1 U232 ( .A1(n202), .A2(n201), .ZN(n251) );
  OAI22_X1 U233 ( .A1(n199), .A2(\mult_x_1/n288 ), .B1(n197), .B2(n21), .ZN(
        n248) );
  OR2_X1 U234 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n200) );
  NAND2_X1 U235 ( .A1(n200), .A2(n199), .ZN(n247) );
  NAND2_X1 U236 ( .A1(n248), .A2(n247), .ZN(n254) );
  NAND2_X1 U237 ( .A1(n202), .A2(n201), .ZN(n252) );
  OAI21_X1 U238 ( .B1(n251), .B2(n254), .A(n252), .ZN(n259) );
  NAND2_X1 U239 ( .A1(n204), .A2(n203), .ZN(n257) );
  INV_X1 U240 ( .A(n257), .ZN(n205) );
  AOI21_X1 U241 ( .B1(n258), .B2(n259), .A(n205), .ZN(n265) );
  NAND2_X1 U242 ( .A1(n207), .A2(n206), .ZN(n263) );
  OAI21_X1 U243 ( .B1(n262), .B2(n265), .A(n263), .ZN(n270) );
  NAND2_X1 U244 ( .A1(n209), .A2(n208), .ZN(n268) );
  INV_X1 U245 ( .A(n268), .ZN(n210) );
  AOI21_X1 U246 ( .B1(n269), .B2(n270), .A(n210), .ZN(n211) );
  MUX2_X1 U247 ( .A(n339), .B(n211), .S(n276), .Z(n378) );
  FA_X1 U248 ( .A(n214), .B(n213), .CI(n212), .CO(n173), .S(n233) );
  FA_X1 U249 ( .A(n217), .B(n216), .CI(n215), .CO(n232), .S(n220) );
  NAND2_X1 U250 ( .A1(n223), .A2(n317), .ZN(n225) );
  INV_X1 U251 ( .A(en), .ZN(n226) );
  NAND2_X1 U252 ( .A1(n226), .A2(n326), .ZN(n224) );
  OAI21_X1 U253 ( .B1(n229), .B2(n225), .A(n224), .ZN(n352) );
  NAND2_X1 U254 ( .A1(n226), .A2(n327), .ZN(n228) );
  NAND2_X1 U255 ( .A1(n223), .A2(n317), .ZN(n227) );
  OAI211_X1 U256 ( .C1(n229), .C2(n226), .A(n228), .B(n227), .ZN(n354) );
  FA_X1 U257 ( .A(n31), .B(n231), .CI(n230), .CO(n176), .S(n245) );
  FA_X1 U258 ( .A(n233), .B(n232), .CI(n33), .CO(n241), .S(n229) );
  NAND2_X1 U259 ( .A1(n245), .A2(n241), .ZN(n234) );
  NAND2_X1 U260 ( .A1(n234), .A2(n276), .ZN(n236) );
  NAND2_X1 U261 ( .A1(n226), .A2(n333), .ZN(n235) );
  NAND2_X1 U262 ( .A1(n236), .A2(n235), .ZN(n366) );
  OAI21_X1 U263 ( .B1(n238), .B2(n237), .A(n317), .ZN(n240) );
  NAND2_X1 U264 ( .A1(n226), .A2(n321), .ZN(n239) );
  NAND2_X1 U265 ( .A1(n240), .A2(n239), .ZN(n342) );
  INV_X1 U266 ( .A(n241), .ZN(n242) );
  NAND2_X1 U267 ( .A1(n242), .A2(n276), .ZN(n244) );
  NAND2_X1 U268 ( .A1(n226), .A2(n336), .ZN(n243) );
  OAI21_X1 U269 ( .B1(n245), .B2(n244), .A(n243), .ZN(n372) );
  BUF_X2 U270 ( .A(rst_n), .Z(n391) );
  MUX2_X1 U271 ( .A(product[0]), .B(n503), .S(n276), .Z(n393) );
  MUX2_X1 U272 ( .A(n503), .B(n504), .S(n276), .Z(n395) );
  AND2_X1 U273 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n246) );
  MUX2_X1 U274 ( .A(n504), .B(n246), .S(n276), .Z(n397) );
  MUX2_X1 U275 ( .A(product[1]), .B(n506), .S(n276), .Z(n399) );
  MUX2_X1 U276 ( .A(n506), .B(n507), .S(n276), .Z(n401) );
  OR2_X1 U277 ( .A1(n248), .A2(n247), .ZN(n249) );
  AND2_X1 U278 ( .A1(n249), .A2(n254), .ZN(n250) );
  MUX2_X1 U279 ( .A(n507), .B(n250), .S(n276), .Z(n403) );
  MUX2_X1 U280 ( .A(product[2]), .B(n509), .S(n276), .Z(n405) );
  MUX2_X1 U281 ( .A(n509), .B(n510), .S(n276), .Z(n407) );
  INV_X1 U282 ( .A(n251), .ZN(n253) );
  NAND2_X1 U283 ( .A1(n253), .A2(n252), .ZN(n255) );
  XOR2_X1 U284 ( .A(n255), .B(n254), .Z(n256) );
  MUX2_X1 U285 ( .A(n510), .B(n256), .S(n276), .Z(n409) );
  MUX2_X1 U286 ( .A(product[3]), .B(n512), .S(n276), .Z(n411) );
  MUX2_X1 U287 ( .A(n512), .B(n513), .S(n276), .Z(n413) );
  NAND2_X1 U288 ( .A1(n258), .A2(n257), .ZN(n260) );
  XNOR2_X1 U289 ( .A(n260), .B(n259), .ZN(n261) );
  MUX2_X1 U290 ( .A(n513), .B(n261), .S(n276), .Z(n415) );
  MUX2_X1 U291 ( .A(product[4]), .B(n515), .S(n276), .Z(n417) );
  MUX2_X1 U292 ( .A(n515), .B(n516), .S(n276), .Z(n419) );
  INV_X1 U293 ( .A(n262), .ZN(n264) );
  NAND2_X1 U294 ( .A1(n264), .A2(n263), .ZN(n266) );
  XOR2_X1 U295 ( .A(n266), .B(n265), .Z(n267) );
  MUX2_X1 U296 ( .A(n516), .B(n267), .S(n276), .Z(n421) );
  MUX2_X1 U297 ( .A(product[5]), .B(n518), .S(n276), .Z(n423) );
  MUX2_X1 U298 ( .A(n518), .B(n519), .S(n276), .Z(n425) );
  NAND2_X1 U299 ( .A1(n269), .A2(n268), .ZN(n271) );
  XNOR2_X1 U300 ( .A(n271), .B(n270), .ZN(n272) );
  MUX2_X1 U301 ( .A(n519), .B(n272), .S(n276), .Z(n427) );
  MUX2_X1 U302 ( .A(product[6]), .B(n521), .S(n276), .Z(n429) );
  NAND2_X1 U303 ( .A1(n383), .A2(n332), .ZN(n273) );
  XOR2_X1 U304 ( .A(n273), .B(n339), .Z(n274) );
  MUX2_X1 U305 ( .A(n521), .B(n274), .S(n276), .Z(n431) );
  MUX2_X1 U306 ( .A(product[7]), .B(n523), .S(n276), .Z(n433) );
  OAI21_X1 U307 ( .B1(n331), .B2(n339), .A(n332), .ZN(n278) );
  NAND2_X1 U308 ( .A1(n322), .A2(n330), .ZN(n275) );
  XNOR2_X1 U309 ( .A(n278), .B(n275), .ZN(n277) );
  MUX2_X1 U310 ( .A(n523), .B(n277), .S(n276), .Z(n435) );
  MUX2_X1 U311 ( .A(product[8]), .B(n525), .S(n317), .Z(n437) );
  AOI21_X1 U312 ( .B1(n278), .B2(n322), .A(n384), .ZN(n281) );
  NAND2_X1 U313 ( .A1(n385), .A2(n329), .ZN(n279) );
  XOR2_X1 U314 ( .A(n281), .B(n279), .Z(n280) );
  MUX2_X1 U315 ( .A(n525), .B(n280), .S(n317), .Z(n439) );
  MUX2_X1 U316 ( .A(product[9]), .B(n527), .S(n317), .Z(n441) );
  OAI21_X1 U317 ( .B1(n281), .B2(n328), .A(n329), .ZN(n289) );
  INV_X1 U318 ( .A(n289), .ZN(n284) );
  NAND2_X1 U319 ( .A1(n387), .A2(n327), .ZN(n282) );
  XOR2_X1 U320 ( .A(n284), .B(n282), .Z(n283) );
  MUX2_X1 U321 ( .A(n527), .B(n283), .S(n317), .Z(n443) );
  MUX2_X1 U322 ( .A(product[10]), .B(n529), .S(n317), .Z(n445) );
  OAI21_X1 U323 ( .B1(n284), .B2(n326), .A(n327), .ZN(n286) );
  NAND2_X1 U324 ( .A1(n388), .A2(n333), .ZN(n285) );
  XNOR2_X1 U325 ( .A(n286), .B(n285), .ZN(n287) );
  MUX2_X1 U326 ( .A(n529), .B(n287), .S(n317), .Z(n447) );
  MUX2_X1 U327 ( .A(product[11]), .B(n531), .S(n317), .Z(n449) );
  NOR2_X1 U328 ( .A1(n336), .A2(n326), .ZN(n290) );
  OAI21_X1 U329 ( .B1(n336), .B2(n327), .A(n333), .ZN(n288) );
  AOI21_X1 U330 ( .B1(n290), .B2(n289), .A(n288), .ZN(n312) );
  NAND2_X1 U331 ( .A1(n386), .A2(n338), .ZN(n291) );
  XOR2_X1 U332 ( .A(n312), .B(n291), .Z(n292) );
  MUX2_X1 U333 ( .A(n531), .B(n292), .S(n317), .Z(n451) );
  MUX2_X1 U334 ( .A(product[12]), .B(n533), .S(n317), .Z(n453) );
  OAI21_X1 U335 ( .B1(n312), .B2(n337), .A(n338), .ZN(n294) );
  NAND2_X1 U336 ( .A1(n335), .A2(n325), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  MUX2_X1 U338 ( .A(n533), .B(n295), .S(n317), .Z(n455) );
  MUX2_X1 U339 ( .A(product[13]), .B(n535), .S(n317), .Z(n457) );
  NAND2_X1 U340 ( .A1(n386), .A2(n335), .ZN(n297) );
  AOI21_X1 U341 ( .B1(n382), .B2(n335), .A(n389), .ZN(n296) );
  OAI21_X1 U342 ( .B1(n312), .B2(n297), .A(n296), .ZN(n299) );
  NAND2_X1 U343 ( .A1(n321), .A2(n334), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U345 ( .A(n535), .B(n300), .S(n317), .Z(n459) );
  MUX2_X1 U346 ( .A(product[14]), .B(n537), .S(n317), .Z(n461) );
  NAND2_X1 U347 ( .A1(n335), .A2(n321), .ZN(n302) );
  NOR2_X1 U348 ( .A1(n337), .A2(n302), .ZN(n308) );
  INV_X1 U349 ( .A(n308), .ZN(n304) );
  AOI21_X1 U350 ( .B1(n389), .B2(n321), .A(n381), .ZN(n301) );
  OAI21_X1 U351 ( .B1(n302), .B2(n338), .A(n301), .ZN(n309) );
  INV_X1 U352 ( .A(n309), .ZN(n303) );
  OAI21_X1 U353 ( .B1(n312), .B2(n304), .A(n303), .ZN(n306) );
  NAND2_X1 U354 ( .A1(n320), .A2(n324), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U356 ( .A(n537), .B(n307), .S(n317), .Z(n463) );
  MUX2_X1 U357 ( .A(product[15]), .B(n539), .S(n317), .Z(n465) );
  NAND2_X1 U358 ( .A1(n308), .A2(n320), .ZN(n311) );
  AOI21_X1 U359 ( .B1(n309), .B2(n320), .A(n380), .ZN(n310) );
  OAI21_X1 U360 ( .B1(n312), .B2(n311), .A(n310), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n313), .B(n323), .ZN(n314) );
  MUX2_X1 U362 ( .A(n539), .B(n314), .S(n317), .Z(n467) );
  MUX2_X1 U363 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n317), .Z(n469) );
  MUX2_X1 U364 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n317), .Z(n471) );
  MUX2_X1 U365 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n317), .Z(n473) );
  MUX2_X1 U366 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n317), .Z(n475) );
  MUX2_X1 U367 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n317), .Z(n477) );
  MUX2_X1 U368 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n317), .Z(n479) );
  MUX2_X1 U369 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n317), .Z(n481) );
  MUX2_X1 U370 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n317), .Z(n483) );
  MUX2_X1 U371 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n317), .Z(n485) );
  MUX2_X1 U372 ( .A(n198), .B(A_extended[1]), .S(n317), .Z(n487) );
  MUX2_X1 U373 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n317), .Z(n489) );
  MUX2_X1 U374 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n317), .Z(n491) );
  MUX2_X1 U375 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n317), .Z(n493) );
  MUX2_X1 U376 ( .A(n315), .B(A_extended[5]), .S(n317), .Z(n495) );
  MUX2_X1 U377 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n317), .Z(n497) );
  MUX2_X1 U378 ( .A(n316), .B(A_extended[7]), .S(n317), .Z(n499) );
  OR2_X1 U379 ( .A1(n317), .A2(n541), .ZN(n501) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_7 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n363, n365, n367, n369, n371, n373, n375, n377,
         n379, n381, n383, n385, n387, n389, n391, n393, n395, n397, n399,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n412, n414,
         n416, n418, n420, n422, n424, n426, n428, n430, n432, n434, n436,
         n438, n440, n442, n444, n446, n448, n450, n452, n454, n456, n458,
         n460, n462, n464, n466, n468, n470, n472, n474, n476, n478, n480,
         n482, n484, n486, n488, n490, n492, n494, n496, n498, n500, n502,
         n504, n506, n508, n510, n512, n514, n516, n518, n520, n522, n523,
         n525, n526, n528, n529, n531, n532, n534, n535, n537, n538, n540,
         n542, n544, n546, n548, n550, n552, n554, n556, n558, n559, n560,
         n561;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n520), .CK(clk), .Q(n560), 
        .QN(n17) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n516), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n30) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n514), .CK(clk), .Q(n559), 
        .QN(n21) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(rst_n), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(rst_n), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n32) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n18) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n27) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n28) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n23) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n486), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(rst_n), .SE(n482), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(rst_n), .SE(n480), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(rst_n), .SE(n478), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(rst_n), .SE(n476), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(rst_n), .SE(n474), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(rst_n), .SE(n470), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(rst_n), .SE(n468), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(rst_n), .SE(n466), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(rst_n), .SE(n464), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(rst_n), .SE(n462), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(rst_n), .SE(n460), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n458), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(rst_n), .SE(n456), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n454), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n450), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n448), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n442), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n440), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n438), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n434), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n430), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n428), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n426), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n420), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n418), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n416), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n414), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n412), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n22) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n561), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n561), .SE(n397), .CK(
        clk), .QN(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n561), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n358), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n561), .SE(n393), .CK(
        clk), .Q(n408), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n561), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n356), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n561), .SE(n389), .CK(
        clk), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n561), .SE(n387), .CK(
        clk), .Q(n407), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n561), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n561), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n352), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n561), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n561), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n350), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n561), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n561), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n348), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n561), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n347), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n561), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n346), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n561), .SE(n369), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n561), .SE(n367), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n561), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n561), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n561), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n341) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n518), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n19) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n20) );
  BUF_X2 U2 ( .A(en), .Z(n8) );
  OR2_X1 U3 ( .A1(n103), .A2(n102), .ZN(n157) );
  BUF_X1 U4 ( .A(\mult_x_1/n281 ), .Z(n6) );
  CLKBUF_X1 U5 ( .A(n182), .Z(n7) );
  INV_X1 U6 ( .A(n209), .ZN(n117) );
  OAI21_X1 U7 ( .B1(n160), .B2(n159), .A(n158), .ZN(n254) );
  NAND2_X1 U8 ( .A1(n157), .A2(n156), .ZN(n158) );
  NOR2_X1 U9 ( .A1(n157), .A2(n156), .ZN(n159) );
  AND2_X1 U10 ( .A1(n560), .A2(\mult_x_1/n281 ), .ZN(n14) );
  AND2_X1 U11 ( .A1(n560), .A2(\mult_x_1/n281 ), .ZN(n125) );
  XNOR2_X1 U12 ( .A(n75), .B(n40), .ZN(n67) );
  XNOR2_X1 U13 ( .A(n77), .B(n76), .ZN(n40) );
  NAND2_X1 U14 ( .A1(n79), .A2(n78), .ZN(n80) );
  NAND2_X1 U15 ( .A1(n77), .A2(n76), .ZN(n78) );
  NAND2_X1 U16 ( .A1(n75), .A2(n74), .ZN(n79) );
  OR2_X1 U17 ( .A1(n76), .A2(n77), .ZN(n74) );
  NAND2_X1 U18 ( .A1(n223), .A2(n222), .ZN(n225) );
  NAND2_X1 U19 ( .A1(n229), .A2(n228), .ZN(n222) );
  NAND2_X1 U20 ( .A1(n231), .A2(n221), .ZN(n223) );
  OR2_X1 U21 ( .A1(n229), .A2(n228), .ZN(n221) );
  XNOR2_X1 U22 ( .A(n231), .B(n230), .ZN(n237) );
  XNOR2_X1 U23 ( .A(n229), .B(n228), .ZN(n230) );
  NAND2_X1 U24 ( .A1(n120), .A2(n119), .ZN(n246) );
  NAND2_X1 U25 ( .A1(n29), .A2(n118), .ZN(n120) );
  NAND2_X1 U26 ( .A1(n117), .A2(n116), .ZN(n118) );
  NAND2_X1 U27 ( .A1(n169), .A2(n168), .ZN(n259) );
  NAND2_X1 U28 ( .A1(n254), .A2(n252), .ZN(n168) );
  NAND2_X1 U29 ( .A1(n94), .A2(n93), .ZN(n9) );
  NAND2_X1 U30 ( .A1(n94), .A2(n93), .ZN(n194) );
  XNOR2_X1 U31 ( .A(n30), .B(n559), .ZN(n10) );
  BUF_X1 U32 ( .A(n162), .Z(n11) );
  CLKBUF_X1 U33 ( .A(n112), .Z(n12) );
  BUF_X2 U34 ( .A(n112), .Z(n13) );
  MUX2_X1 U35 ( .A(n170), .B(n343), .S(n83), .Z(n365) );
  OAI22_X1 U36 ( .A1(n179), .A2(n146), .B1(n127), .B2(n177), .ZN(n15) );
  INV_X1 U37 ( .A(n10), .ZN(n195) );
  OAI21_X1 U38 ( .B1(n254), .B2(n252), .A(n253), .ZN(n169) );
  INV_X1 U39 ( .A(n19), .ZN(n16) );
  BUF_X2 U40 ( .A(en), .Z(n299) );
  INV_X1 U41 ( .A(rst_n), .ZN(n561) );
  XOR2_X1 U42 ( .A(n106), .B(n105), .Z(n29) );
  AND2_X1 U43 ( .A1(n105), .A2(n106), .ZN(n31) );
  XNOR2_X1 U44 ( .A(\mult_x_1/a[4] ), .B(n559), .ZN(n33) );
  XOR2_X1 U45 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .Z(n34) );
  OR2_X2 U46 ( .A1(n34), .A2(n33), .ZN(n179) );
  BUF_X2 U47 ( .A(n559), .Z(n339) );
  OR2_X1 U48 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n35) );
  INV_X2 U49 ( .A(n34), .ZN(n177) );
  OAI22_X1 U50 ( .A1(n179), .A2(n21), .B1(n35), .B2(n177), .ZN(n70) );
  XNOR2_X1 U51 ( .A(n339), .B(\mult_x_1/n288 ), .ZN(n36) );
  XNOR2_X1 U52 ( .A(n339), .B(\mult_x_1/n287 ), .ZN(n71) );
  OAI22_X1 U53 ( .A1(n179), .A2(n36), .B1(n177), .B2(n71), .ZN(n69) );
  BUF_X2 U54 ( .A(\mult_x_1/n313 ), .Z(n91) );
  NAND2_X1 U55 ( .A1(n91), .A2(n18), .ZN(n182) );
  XNOR2_X1 U56 ( .A(n91), .B(\mult_x_1/n284 ), .ZN(n41) );
  XNOR2_X1 U57 ( .A(n91), .B(\mult_x_1/n283 ), .ZN(n72) );
  OAI22_X1 U58 ( .A1(n7), .A2(n41), .B1(n72), .B2(n18), .ZN(n77) );
  XOR2_X1 U59 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[2] ), .Z(n37) );
  XNOR2_X1 U60 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n38) );
  NAND2_X1 U61 ( .A1(n37), .A2(n38), .ZN(n112) );
  BUF_X2 U62 ( .A(\mult_x_1/n312 ), .Z(n338) );
  XNOR2_X1 U63 ( .A(n338), .B(\mult_x_1/n286 ), .ZN(n43) );
  INV_X1 U64 ( .A(n38), .ZN(n39) );
  INV_X2 U65 ( .A(n39), .ZN(n184) );
  XNOR2_X1 U66 ( .A(n338), .B(\mult_x_1/n285 ), .ZN(n73) );
  OAI22_X1 U67 ( .A1(n13), .A2(n43), .B1(n184), .B2(n73), .ZN(n76) );
  INV_X1 U68 ( .A(n67), .ZN(n45) );
  XNOR2_X1 U69 ( .A(n91), .B(\mult_x_1/n285 ), .ZN(n51) );
  OAI22_X1 U70 ( .A1(n182), .A2(n51), .B1(n41), .B2(n18), .ZN(n48) );
  INV_X1 U71 ( .A(n177), .ZN(n42) );
  AND2_X1 U72 ( .A1(\mult_x_1/n288 ), .A2(n42), .ZN(n47) );
  XNOR2_X1 U73 ( .A(n338), .B(\mult_x_1/n287 ), .ZN(n49) );
  OAI22_X1 U74 ( .A1(n13), .A2(n49), .B1(n184), .B2(n43), .ZN(n46) );
  INV_X1 U75 ( .A(n66), .ZN(n44) );
  NAND2_X1 U76 ( .A1(n45), .A2(n44), .ZN(n268) );
  FA_X1 U77 ( .A(n48), .B(n47), .CI(n46), .CO(n66), .S(n65) );
  XNOR2_X1 U78 ( .A(n338), .B(\mult_x_1/n288 ), .ZN(n50) );
  OAI22_X1 U79 ( .A1(n13), .A2(n50), .B1(n184), .B2(n49), .ZN(n53) );
  XNOR2_X1 U80 ( .A(n91), .B(\mult_x_1/n286 ), .ZN(n55) );
  OAI22_X1 U81 ( .A1(n182), .A2(n55), .B1(n51), .B2(n18), .ZN(n52) );
  NOR2_X1 U82 ( .A1(n65), .A2(n64), .ZN(n291) );
  HA_X1 U83 ( .A(n53), .B(n52), .CO(n64), .S(n62) );
  OR2_X1 U84 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n54) );
  OAI22_X1 U85 ( .A1(n13), .A2(n22), .B1(n54), .B2(n184), .ZN(n61) );
  OR2_X1 U86 ( .A1(n62), .A2(n61), .ZN(n287) );
  XNOR2_X1 U87 ( .A(n91), .B(\mult_x_1/n287 ), .ZN(n57) );
  OAI22_X1 U88 ( .A1(n7), .A2(n57), .B1(n55), .B2(n18), .ZN(n60) );
  INV_X1 U89 ( .A(n184), .ZN(n56) );
  AND2_X1 U90 ( .A1(\mult_x_1/n288 ), .A2(n56), .ZN(n59) );
  NOR2_X1 U91 ( .A1(n60), .A2(n59), .ZN(n280) );
  OAI22_X1 U92 ( .A1(n182), .A2(\mult_x_1/n288 ), .B1(n57), .B2(n18), .ZN(n277) );
  OR2_X1 U93 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n58) );
  NAND2_X1 U94 ( .A1(n58), .A2(n7), .ZN(n276) );
  NAND2_X1 U95 ( .A1(n277), .A2(n276), .ZN(n283) );
  NAND2_X1 U96 ( .A1(n60), .A2(n59), .ZN(n281) );
  OAI21_X1 U97 ( .B1(n280), .B2(n283), .A(n281), .ZN(n288) );
  NAND2_X1 U98 ( .A1(n62), .A2(n61), .ZN(n286) );
  INV_X1 U99 ( .A(n286), .ZN(n63) );
  AOI21_X1 U100 ( .B1(n287), .B2(n288), .A(n63), .ZN(n294) );
  NAND2_X1 U101 ( .A1(n65), .A2(n64), .ZN(n292) );
  OAI21_X1 U102 ( .B1(n291), .B2(n294), .A(n292), .ZN(n270) );
  NAND2_X1 U103 ( .A1(n67), .A2(n66), .ZN(n269) );
  INV_X1 U104 ( .A(n269), .ZN(n68) );
  AOI21_X1 U105 ( .B1(n268), .B2(n270), .A(n68), .ZN(n262) );
  HA_X1 U106 ( .A(n70), .B(n69), .CO(n188), .S(n75) );
  XNOR2_X1 U107 ( .A(n339), .B(\mult_x_1/n286 ), .ZN(n178) );
  OAI22_X1 U108 ( .A1(n179), .A2(n71), .B1(n177), .B2(n178), .ZN(n187) );
  XNOR2_X1 U109 ( .A(n91), .B(\mult_x_1/n282 ), .ZN(n181) );
  OAI22_X1 U110 ( .A1(n182), .A2(n72), .B1(n181), .B2(n18), .ZN(n173) );
  XNOR2_X1 U111 ( .A(n30), .B(n559), .ZN(n86) );
  AND2_X1 U112 ( .A1(\mult_x_1/n288 ), .A2(n10), .ZN(n172) );
  XNOR2_X1 U113 ( .A(n338), .B(\mult_x_1/n284 ), .ZN(n185) );
  OAI22_X1 U114 ( .A1(n13), .A2(n73), .B1(n184), .B2(n185), .ZN(n171) );
  NOR2_X1 U115 ( .A1(n81), .A2(n80), .ZN(n242) );
  NAND2_X1 U116 ( .A1(n81), .A2(n80), .ZN(n243) );
  OAI21_X1 U117 ( .B1(n262), .B2(n242), .A(n243), .ZN(n82) );
  NAND2_X1 U118 ( .A1(n82), .A2(n8), .ZN(n85) );
  INV_X1 U119 ( .A(n340), .ZN(n83) );
  NAND2_X1 U120 ( .A1(n83), .A2(n359), .ZN(n84) );
  NAND2_X1 U121 ( .A1(n85), .A2(n84), .ZN(n397) );
  XNOR2_X1 U122 ( .A(n339), .B(\mult_x_1/n284 ), .ZN(n110) );
  XNOR2_X1 U123 ( .A(n339), .B(\mult_x_1/n283 ), .ZN(n95) );
  OAI22_X1 U124 ( .A1(n179), .A2(n110), .B1(n177), .B2(n95), .ZN(n103) );
  XNOR2_X1 U125 ( .A(n338), .B(\mult_x_1/n282 ), .ZN(n111) );
  XNOR2_X1 U126 ( .A(n338), .B(n6), .ZN(n96) );
  OAI22_X1 U127 ( .A1(n12), .A2(n111), .B1(n184), .B2(n96), .ZN(n102) );
  XNOR2_X1 U128 ( .A(n103), .B(n102), .ZN(n106) );
  XNOR2_X1 U129 ( .A(\mult_x_1/n310 ), .B(n30), .ZN(n93) );
  INV_X1 U130 ( .A(n86), .ZN(n94) );
  XNOR2_X1 U131 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n114) );
  INV_X1 U132 ( .A(n114), .ZN(n87) );
  NAND3_X1 U133 ( .A1(n93), .A2(n94), .A3(n87), .ZN(n90) );
  XNOR2_X1 U134 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n100) );
  INV_X1 U135 ( .A(n100), .ZN(n88) );
  NAND2_X1 U136 ( .A1(n88), .A2(n10), .ZN(n89) );
  NAND2_X1 U137 ( .A1(n90), .A2(n89), .ZN(n217) );
  XNOR2_X1 U138 ( .A(n91), .B(n6), .ZN(n180) );
  XNOR2_X1 U139 ( .A(n14), .B(n91), .ZN(n97) );
  OAI22_X1 U140 ( .A1(n182), .A2(n180), .B1(n97), .B2(n18), .ZN(n216) );
  NAND2_X1 U141 ( .A1(n17), .A2(\mult_x_1/n310 ), .ZN(n101) );
  INV_X1 U142 ( .A(n101), .ZN(n92) );
  AND2_X1 U143 ( .A1(\mult_x_1/n288 ), .A2(n92), .ZN(n215) );
  XNOR2_X1 U144 ( .A(n16), .B(\mult_x_1/n285 ), .ZN(n99) );
  XNOR2_X1 U145 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n140) );
  OAI22_X1 U146 ( .A1(n194), .A2(n99), .B1(n195), .B2(n140), .ZN(n145) );
  XNOR2_X1 U147 ( .A(n339), .B(\mult_x_1/n282 ), .ZN(n147) );
  OAI22_X1 U148 ( .A1(n179), .A2(n95), .B1(n177), .B2(n147), .ZN(n144) );
  XNOR2_X1 U149 ( .A(n125), .B(n338), .ZN(n141) );
  OAI22_X1 U150 ( .A1(n12), .A2(n96), .B1(n184), .B2(n141), .ZN(n162) );
  INV_X1 U151 ( .A(n162), .ZN(n143) );
  AOI21_X1 U152 ( .B1(n182), .B2(n18), .A(n97), .ZN(n98) );
  INV_X1 U153 ( .A(n98), .ZN(n109) );
  OAI22_X1 U154 ( .A1(n9), .A2(n100), .B1(n195), .B2(n99), .ZN(n108) );
  NOR2_X1 U155 ( .A1(n23), .A2(n101), .ZN(n107) );
  NOR2_X1 U156 ( .A1(n24), .A2(n101), .ZN(n156) );
  XNOR2_X1 U157 ( .A(n157), .B(n156), .ZN(n104) );
  XNOR2_X1 U158 ( .A(n104), .B(n155), .ZN(n256) );
  FA_X1 U159 ( .A(n109), .B(n107), .CI(n108), .CO(n155), .S(n209) );
  XNOR2_X1 U160 ( .A(n339), .B(\mult_x_1/n285 ), .ZN(n176) );
  OAI22_X1 U161 ( .A1(n179), .A2(n176), .B1(n177), .B2(n110), .ZN(n214) );
  XNOR2_X1 U162 ( .A(n338), .B(\mult_x_1/n283 ), .ZN(n183) );
  OAI22_X1 U163 ( .A1(n13), .A2(n183), .B1(n184), .B2(n111), .ZN(n213) );
  OR2_X1 U164 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n113) );
  OAI22_X1 U165 ( .A1(n9), .A2(n19), .B1(n113), .B2(n195), .ZN(n175) );
  XNOR2_X1 U166 ( .A(n16), .B(\mult_x_1/n288 ), .ZN(n115) );
  OAI22_X1 U167 ( .A1(n194), .A2(n115), .B1(n195), .B2(n114), .ZN(n174) );
  INV_X1 U168 ( .A(n210), .ZN(n116) );
  NAND2_X1 U169 ( .A1(n209), .A2(n210), .ZN(n119) );
  NAND2_X1 U170 ( .A1(n247), .A2(n246), .ZN(n121) );
  NAND2_X1 U171 ( .A1(n121), .A2(n299), .ZN(n123) );
  NAND2_X1 U172 ( .A1(n83), .A2(n355), .ZN(n122) );
  NAND2_X1 U173 ( .A1(n123), .A2(n122), .ZN(n389) );
  NOR2_X1 U194 ( .A1(n25), .A2(n101), .ZN(n192) );
  XNOR2_X1 U195 ( .A(n16), .B(n6), .ZN(n124) );
  XNOR2_X1 U196 ( .A(n14), .B(n16), .ZN(n193) );
  OAI22_X1 U197 ( .A1(n9), .A2(n124), .B1(n193), .B2(n195), .ZN(n200) );
  INV_X1 U198 ( .A(n200), .ZN(n191) );
  XNOR2_X1 U199 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n128) );
  OAI22_X1 U200 ( .A1(n9), .A2(n128), .B1(n195), .B2(n124), .ZN(n131) );
  XNOR2_X1 U201 ( .A(n14), .B(n339), .ZN(n127) );
  AOI21_X1 U202 ( .B1(n177), .B2(n179), .A(n127), .ZN(n126) );
  INV_X1 U203 ( .A(n126), .ZN(n130) );
  XNOR2_X1 U204 ( .A(n339), .B(n6), .ZN(n146) );
  OAI22_X1 U205 ( .A1(n179), .A2(n146), .B1(n127), .B2(n177), .ZN(n129) );
  NOR2_X1 U206 ( .A1(n26), .A2(n101), .ZN(n138) );
  XNOR2_X1 U207 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n139) );
  OAI22_X1 U208 ( .A1(n194), .A2(n139), .B1(n195), .B2(n128), .ZN(n137) );
  INV_X1 U209 ( .A(n129), .ZN(n136) );
  NOR2_X1 U210 ( .A1(n27), .A2(n101), .ZN(n134) );
  FA_X1 U211 ( .A(n131), .B(n130), .CI(n15), .CO(n190), .S(n133) );
  OR2_X1 U212 ( .A1(n207), .A2(n206), .ZN(n132) );
  MUX2_X1 U213 ( .A(n341), .B(n132), .S(n8), .Z(n361) );
  FA_X1 U214 ( .A(n135), .B(n134), .CI(n133), .CO(n206), .S(n250) );
  FA_X1 U215 ( .A(n138), .B(n137), .CI(n136), .CO(n135), .S(n154) );
  OAI22_X1 U216 ( .A1(n9), .A2(n140), .B1(n195), .B2(n139), .ZN(n163) );
  AOI21_X1 U217 ( .B1(n184), .B2(n13), .A(n141), .ZN(n142) );
  INV_X1 U218 ( .A(n142), .ZN(n161) );
  FA_X1 U219 ( .A(n145), .B(n144), .CI(n143), .CO(n167), .S(n257) );
  NOR2_X1 U220 ( .A1(n28), .A2(n101), .ZN(n165) );
  OAI22_X1 U221 ( .A1(n179), .A2(n147), .B1(n177), .B2(n146), .ZN(n164) );
  OR2_X1 U222 ( .A1(n165), .A2(n164), .ZN(n148) );
  NAND2_X1 U223 ( .A1(n167), .A2(n148), .ZN(n150) );
  NAND2_X1 U224 ( .A1(n165), .A2(n164), .ZN(n149) );
  NAND2_X1 U225 ( .A1(n150), .A2(n149), .ZN(n152) );
  OR2_X1 U226 ( .A1(n250), .A2(n249), .ZN(n151) );
  MUX2_X1 U227 ( .A(n342), .B(n151), .S(n8), .Z(n363) );
  FA_X1 U228 ( .A(n154), .B(n153), .CI(n152), .CO(n249), .S(n260) );
  INV_X1 U229 ( .A(n155), .ZN(n160) );
  FA_X1 U230 ( .A(n163), .B(n11), .CI(n161), .CO(n153), .S(n252) );
  XNOR2_X1 U231 ( .A(n165), .B(n164), .ZN(n166) );
  XNOR2_X1 U232 ( .A(n167), .B(n166), .ZN(n253) );
  OR2_X1 U233 ( .A1(n260), .A2(n259), .ZN(n170) );
  FA_X1 U234 ( .A(n173), .B(n172), .CI(n171), .CO(n234), .S(n186) );
  HA_X1 U235 ( .A(n175), .B(n174), .CO(n212), .S(n233) );
  OAI22_X1 U236 ( .A1(n179), .A2(n178), .B1(n177), .B2(n176), .ZN(n220) );
  OAI22_X1 U237 ( .A1(n182), .A2(n181), .B1(n180), .B2(n18), .ZN(n219) );
  OAI22_X1 U238 ( .A1(n13), .A2(n185), .B1(n184), .B2(n183), .ZN(n218) );
  FA_X1 U239 ( .A(n188), .B(n187), .CI(n186), .CO(n239), .S(n81) );
  OR2_X1 U240 ( .A1(n240), .A2(n239), .ZN(n189) );
  MUX2_X1 U241 ( .A(n344), .B(n189), .S(n8), .Z(n367) );
  FA_X1 U242 ( .A(n192), .B(n191), .CI(n190), .CO(n202), .S(n207) );
  AOI21_X1 U243 ( .B1(n195), .B2(n9), .A(n193), .ZN(n196) );
  INV_X1 U244 ( .A(n196), .ZN(n198) );
  NOR2_X1 U245 ( .A1(n20), .A2(n101), .ZN(n197) );
  XOR2_X1 U246 ( .A(n198), .B(n197), .Z(n199) );
  XOR2_X1 U247 ( .A(n200), .B(n199), .Z(n201) );
  OR2_X1 U248 ( .A1(n202), .A2(n201), .ZN(n204) );
  NAND2_X1 U249 ( .A1(n202), .A2(n201), .ZN(n203) );
  NAND2_X1 U250 ( .A1(n204), .A2(n203), .ZN(n205) );
  MUX2_X1 U251 ( .A(n345), .B(n205), .S(n8), .Z(n369) );
  NAND2_X1 U252 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U253 ( .A(n346), .B(n208), .S(n8), .Z(n371) );
  XNOR2_X1 U254 ( .A(n210), .B(n209), .ZN(n211) );
  XNOR2_X1 U255 ( .A(n29), .B(n211), .ZN(n226) );
  FA_X1 U256 ( .A(n214), .B(n213), .CI(n212), .CO(n210), .S(n231) );
  FA_X1 U257 ( .A(n217), .B(n216), .CI(n215), .CO(n105), .S(n229) );
  FA_X1 U258 ( .A(n220), .B(n219), .CI(n218), .CO(n228), .S(n232) );
  NOR2_X1 U259 ( .A1(n226), .A2(n225), .ZN(n224) );
  MUX2_X1 U260 ( .A(n348), .B(n224), .S(n299), .Z(n375) );
  NAND2_X1 U261 ( .A1(n226), .A2(n225), .ZN(n227) );
  MUX2_X1 U262 ( .A(n349), .B(n227), .S(n299), .Z(n377) );
  FA_X1 U263 ( .A(n234), .B(n233), .CI(n232), .CO(n236), .S(n240) );
  NOR2_X1 U264 ( .A1(n237), .A2(n236), .ZN(n235) );
  MUX2_X1 U265 ( .A(n350), .B(n235), .S(n8), .Z(n379) );
  NAND2_X1 U266 ( .A1(n237), .A2(n236), .ZN(n238) );
  MUX2_X1 U267 ( .A(n351), .B(n238), .S(n299), .Z(n381) );
  NAND2_X1 U268 ( .A1(n240), .A2(n239), .ZN(n241) );
  MUX2_X1 U269 ( .A(n352), .B(n241), .S(n8), .Z(n383) );
  INV_X1 U270 ( .A(n242), .ZN(n244) );
  NAND2_X1 U271 ( .A1(n244), .A2(n243), .ZN(n245) );
  MUX2_X1 U272 ( .A(n353), .B(n245), .S(n299), .Z(n385) );
  NOR2_X1 U273 ( .A1(n247), .A2(n246), .ZN(n248) );
  MUX2_X1 U274 ( .A(n354), .B(n248), .S(n340), .Z(n387) );
  NAND2_X1 U275 ( .A1(n250), .A2(n249), .ZN(n251) );
  MUX2_X1 U276 ( .A(n356), .B(n251), .S(n299), .Z(n391) );
  XNOR2_X1 U277 ( .A(n253), .B(n252), .ZN(n255) );
  XNOR2_X1 U278 ( .A(n255), .B(n254), .ZN(n264) );
  FA_X1 U279 ( .A(n31), .B(n257), .CI(n256), .CO(n263), .S(n247) );
  NOR2_X1 U280 ( .A1(n264), .A2(n263), .ZN(n258) );
  MUX2_X1 U281 ( .A(n357), .B(n258), .S(n299), .Z(n393) );
  NAND2_X1 U282 ( .A1(n260), .A2(n259), .ZN(n261) );
  MUX2_X1 U283 ( .A(n358), .B(n261), .S(n340), .Z(n395) );
  MUX2_X1 U284 ( .A(n360), .B(n262), .S(n8), .Z(n399) );
  NAND2_X1 U285 ( .A1(n264), .A2(n263), .ZN(n265) );
  NAND2_X1 U286 ( .A1(n265), .A2(n299), .ZN(n267) );
  NAND2_X1 U287 ( .A1(n83), .A2(n347), .ZN(n266) );
  NAND2_X1 U288 ( .A1(n267), .A2(n266), .ZN(n373) );
  NAND2_X1 U289 ( .A1(n269), .A2(n268), .ZN(n271) );
  XNOR2_X1 U290 ( .A(n271), .B(n270), .ZN(n272) );
  NAND2_X1 U291 ( .A1(n272), .A2(n340), .ZN(n274) );
  NAND2_X1 U292 ( .A1(n83), .A2(n538), .ZN(n273) );
  NAND2_X1 U293 ( .A1(n274), .A2(n273), .ZN(n446) );
  MUX2_X1 U294 ( .A(product[0]), .B(n522), .S(n8), .Z(n412) );
  MUX2_X1 U295 ( .A(n522), .B(n523), .S(n340), .Z(n414) );
  AND2_X1 U296 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n275) );
  MUX2_X1 U297 ( .A(n523), .B(n275), .S(n299), .Z(n416) );
  MUX2_X1 U298 ( .A(product[1]), .B(n525), .S(n340), .Z(n418) );
  MUX2_X1 U299 ( .A(n525), .B(n526), .S(n8), .Z(n420) );
  OR2_X1 U300 ( .A1(n277), .A2(n276), .ZN(n278) );
  AND2_X1 U301 ( .A1(n278), .A2(n283), .ZN(n279) );
  MUX2_X1 U302 ( .A(n526), .B(n279), .S(n340), .Z(n422) );
  MUX2_X1 U303 ( .A(product[2]), .B(n528), .S(n299), .Z(n424) );
  MUX2_X1 U304 ( .A(n528), .B(n529), .S(n340), .Z(n426) );
  INV_X1 U305 ( .A(n280), .ZN(n282) );
  NAND2_X1 U306 ( .A1(n282), .A2(n281), .ZN(n284) );
  XOR2_X1 U307 ( .A(n284), .B(n283), .Z(n285) );
  MUX2_X1 U308 ( .A(n529), .B(n285), .S(n8), .Z(n428) );
  MUX2_X1 U309 ( .A(product[3]), .B(n531), .S(n340), .Z(n430) );
  MUX2_X1 U310 ( .A(n531), .B(n532), .S(n299), .Z(n432) );
  NAND2_X1 U311 ( .A1(n287), .A2(n286), .ZN(n289) );
  XNOR2_X1 U312 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U313 ( .A(n532), .B(n290), .S(n8), .Z(n434) );
  MUX2_X1 U314 ( .A(product[4]), .B(n534), .S(n340), .Z(n436) );
  MUX2_X1 U315 ( .A(n534), .B(n535), .S(n340), .Z(n438) );
  INV_X1 U316 ( .A(n291), .ZN(n293) );
  NAND2_X1 U317 ( .A1(n293), .A2(n292), .ZN(n295) );
  XOR2_X1 U318 ( .A(n295), .B(n294), .Z(n296) );
  MUX2_X1 U319 ( .A(n535), .B(n296), .S(n340), .Z(n440) );
  MUX2_X1 U320 ( .A(product[5]), .B(n537), .S(n340), .Z(n442) );
  MUX2_X1 U321 ( .A(n537), .B(n538), .S(n299), .Z(n444) );
  MUX2_X1 U322 ( .A(product[6]), .B(n540), .S(n340), .Z(n448) );
  XOR2_X1 U323 ( .A(n353), .B(n360), .Z(n297) );
  MUX2_X1 U324 ( .A(n540), .B(n297), .S(n8), .Z(n450) );
  MUX2_X1 U325 ( .A(product[7]), .B(n542), .S(n340), .Z(n452) );
  NAND2_X1 U326 ( .A1(n344), .A2(n352), .ZN(n298) );
  XNOR2_X1 U327 ( .A(n359), .B(n298), .ZN(n300) );
  MUX2_X1 U328 ( .A(n542), .B(n300), .S(n299), .Z(n454) );
  BUF_X4 U329 ( .A(en), .Z(n340) );
  MUX2_X1 U330 ( .A(product[8]), .B(n544), .S(n299), .Z(n456) );
  AOI21_X1 U331 ( .B1(n359), .B2(n344), .A(n404), .ZN(n303) );
  NAND2_X1 U332 ( .A1(n405), .A2(n351), .ZN(n301) );
  XOR2_X1 U333 ( .A(n303), .B(n301), .Z(n302) );
  MUX2_X1 U334 ( .A(n544), .B(n302), .S(n340), .Z(n458) );
  MUX2_X1 U335 ( .A(product[9]), .B(n546), .S(n340), .Z(n460) );
  OAI21_X1 U336 ( .B1(n303), .B2(n350), .A(n351), .ZN(n311) );
  INV_X1 U337 ( .A(n311), .ZN(n306) );
  NAND2_X1 U338 ( .A1(n406), .A2(n349), .ZN(n304) );
  XOR2_X1 U339 ( .A(n306), .B(n304), .Z(n305) );
  MUX2_X1 U340 ( .A(n546), .B(n305), .S(n299), .Z(n462) );
  MUX2_X1 U341 ( .A(product[10]), .B(n548), .S(n8), .Z(n464) );
  OAI21_X1 U342 ( .B1(n306), .B2(n348), .A(n349), .ZN(n308) );
  NAND2_X1 U343 ( .A1(n407), .A2(n355), .ZN(n307) );
  XNOR2_X1 U344 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U345 ( .A(n548), .B(n309), .S(n340), .Z(n466) );
  MUX2_X1 U346 ( .A(product[11]), .B(n550), .S(n340), .Z(n468) );
  NOR2_X1 U347 ( .A1(n354), .A2(n348), .ZN(n312) );
  OAI21_X1 U348 ( .B1(n354), .B2(n349), .A(n355), .ZN(n310) );
  AOI21_X1 U349 ( .B1(n312), .B2(n311), .A(n310), .ZN(n335) );
  NAND2_X1 U350 ( .A1(n408), .A2(n347), .ZN(n313) );
  XOR2_X1 U351 ( .A(n335), .B(n313), .Z(n314) );
  MUX2_X1 U352 ( .A(n550), .B(n314), .S(n299), .Z(n470) );
  MUX2_X1 U353 ( .A(product[12]), .B(n552), .S(n8), .Z(n472) );
  OAI21_X1 U354 ( .B1(n335), .B2(n357), .A(n347), .ZN(n316) );
  NAND2_X1 U355 ( .A1(n343), .A2(n358), .ZN(n315) );
  XNOR2_X1 U356 ( .A(n316), .B(n315), .ZN(n317) );
  MUX2_X1 U357 ( .A(n552), .B(n317), .S(n340), .Z(n474) );
  MUX2_X1 U358 ( .A(product[13]), .B(n554), .S(n340), .Z(n476) );
  NAND2_X1 U359 ( .A1(n408), .A2(n343), .ZN(n319) );
  AOI21_X1 U360 ( .B1(n403), .B2(n343), .A(n409), .ZN(n318) );
  OAI21_X1 U361 ( .B1(n335), .B2(n319), .A(n318), .ZN(n321) );
  NAND2_X1 U362 ( .A1(n342), .A2(n356), .ZN(n320) );
  XNOR2_X1 U363 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U364 ( .A(n554), .B(n322), .S(n299), .Z(n478) );
  MUX2_X1 U365 ( .A(product[14]), .B(n556), .S(n8), .Z(n480) );
  NAND2_X1 U366 ( .A1(n343), .A2(n342), .ZN(n324) );
  INV_X1 U367 ( .A(n324), .ZN(n330) );
  NAND2_X1 U368 ( .A1(n408), .A2(n330), .ZN(n326) );
  AOI21_X1 U369 ( .B1(n409), .B2(n342), .A(n402), .ZN(n323) );
  OAI21_X1 U370 ( .B1(n324), .B2(n347), .A(n323), .ZN(n332) );
  INV_X1 U371 ( .A(n332), .ZN(n325) );
  OAI21_X1 U372 ( .B1(n335), .B2(n326), .A(n325), .ZN(n328) );
  NAND2_X1 U373 ( .A1(n341), .A2(n346), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n329) );
  MUX2_X1 U375 ( .A(n556), .B(n329), .S(n340), .Z(n482) );
  MUX2_X1 U376 ( .A(product[15]), .B(n558), .S(n340), .Z(n484) );
  AND2_X1 U377 ( .A1(n408), .A2(n341), .ZN(n331) );
  NAND2_X1 U378 ( .A1(n331), .A2(n330), .ZN(n334) );
  AOI21_X1 U379 ( .B1(n332), .B2(n341), .A(n401), .ZN(n333) );
  OAI21_X1 U380 ( .B1(n335), .B2(n334), .A(n333), .ZN(n336) );
  XNOR2_X1 U381 ( .A(n336), .B(n345), .ZN(n337) );
  MUX2_X1 U382 ( .A(n558), .B(n337), .S(n299), .Z(n486) );
  MUX2_X1 U383 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n340), .Z(n488) );
  MUX2_X1 U384 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n299), .Z(n490) );
  MUX2_X1 U385 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n340), .Z(n492) );
  MUX2_X1 U386 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n8), .Z(n494) );
  MUX2_X1 U387 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n8), .Z(n496) );
  MUX2_X1 U388 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n340), .Z(n498) );
  MUX2_X1 U389 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n8), .Z(n500) );
  MUX2_X1 U390 ( .A(n6), .B(B_extended[7]), .S(n8), .Z(n502) );
  MUX2_X1 U391 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n8), .Z(n504) );
  MUX2_X1 U392 ( .A(n91), .B(A_extended[1]), .S(n340), .Z(n506) );
  MUX2_X1 U393 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n340), .Z(n508) );
  MUX2_X1 U394 ( .A(n338), .B(A_extended[3]), .S(n299), .Z(n510) );
  MUX2_X1 U395 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n340), .Z(n512) );
  MUX2_X1 U396 ( .A(n339), .B(A_extended[5]), .S(n8), .Z(n514) );
  MUX2_X1 U397 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n340), .Z(n516) );
  MUX2_X1 U398 ( .A(n16), .B(A_extended[7]), .S(n340), .Z(n518) );
  OR2_X1 U399 ( .A1(n299), .A2(n560), .ZN(n520) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_8 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n354, n356, n358, n360, n362, n364, n366, n368, n370,
         n372, n374, n376, n378, n380, n382, n384, n386, n388, n390, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n407, n409, n411, n413, n415, n417, n419, n421, n423,
         n425, n427, n429, n431, n433, n435, n437, n439, n441, n443, n445,
         n447, n449, n451, n453, n455, n457, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n515, n517, n518, n520, n521, n523, n524, n526, n527, n529,
         n530, n532, n533, n535, n537, n539, n541, n543, n545, n547, n549,
         n551, n553, n554, n555, n556, n557;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n404), .SE(n515), .CK(clk), .Q(n556), 
        .QN(n402) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n404), .SE(n511), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n22) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n405), .SE(n509), .CK(clk), .Q(n555), 
        .QN(n21) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n405), .SE(n507), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n23) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n404), .SE(n503), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n12) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n404), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n15) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n405), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n404), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n404), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n404), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n404), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n405), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n405), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n20) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n404), .SE(n481), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n404), .SE(n479), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n405), .SE(n477), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n404), .SE(n475), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n404), .SE(n473), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n404), .SE(n471), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n405), .SE(n469), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n404), .SE(n467), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n404), .SE(n465), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n405), .SE(n463), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n404), .SE(n461), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n404), .SE(n459), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n405), .SE(n457), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n404), .SE(n455), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n404), .SE(n453), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n404), .SE(n451), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n405), .SE(n449), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n405), .SE(n447), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n405), .SE(n445), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n405), .SE(n443), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n405), .SE(n441), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n405), .SE(n439), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n405), .SE(n437), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n405), .SE(n435), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n405), .SE(n433), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n405), .SE(n431), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n405), .SE(n429), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n404), .SE(n427), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n404), .SE(n425), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n404), .SE(n423), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n404), .SE(n421), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n404), .SE(n419), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n404), .SE(n417), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n404), .SE(n415), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n404), .SE(n413), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n404), .SE(n411), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n404), .SE(n409), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n404), .SE(n407), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n405), .SE(n505), .CK(clk), .Q(n554), 
        .QN(n24) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n404), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n26) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n557), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n557), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n350), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n557), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n349), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n557), .SE(n384), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n557), .SE(n382), .CK(
        clk), .Q(n400), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n557), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n557), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n345), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n557), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n344), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n557), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n557), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n342), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n557), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n341), .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n557), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n340), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n557), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n339), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n557), .SE(n364), .CK(
        clk), .Q(n399), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n557), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n337), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n557), .SE(n360), .CK(
        clk), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n557), .SE(n358), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n557), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n557), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n557), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n332) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n404), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n403) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n404), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n19) );
  INV_X1 U2 ( .A(n229), .ZN(n149) );
  BUF_X1 U3 ( .A(n289), .Z(n200) );
  BUF_X1 U4 ( .A(n289), .Z(n257) );
  BUF_X2 U5 ( .A(\mult_x_1/n310 ), .Z(n330) );
  OAI22_X1 U6 ( .A1(n151), .A2(n56), .B1(n149), .B2(n38), .ZN(n5) );
  INV_X1 U7 ( .A(n134), .ZN(n113) );
  OAI21_X1 U8 ( .B1(n128), .B2(n127), .A(n126), .ZN(n130) );
  NAND2_X1 U9 ( .A1(n128), .A2(n127), .ZN(n129) );
  AND2_X1 U10 ( .A1(n556), .A2(\mult_x_1/n281 ), .ZN(n13) );
  AND2_X1 U11 ( .A1(n556), .A2(\mult_x_1/n281 ), .ZN(n88) );
  NAND2_X1 U12 ( .A1(n135), .A2(n134), .ZN(n117) );
  OAI21_X1 U13 ( .B1(n37), .B2(n36), .A(n35), .ZN(n183) );
  NAND2_X1 U14 ( .A1(n120), .A2(n119), .ZN(n219) );
  NAND2_X1 U15 ( .A1(n124), .A2(n122), .ZN(n119) );
  OAI21_X1 U16 ( .B1(n124), .B2(n122), .A(n123), .ZN(n120) );
  NAND2_X1 U17 ( .A1(n130), .A2(n129), .ZN(n180) );
  XNOR2_X1 U18 ( .A(n135), .B(n134), .ZN(n136) );
  XNOR2_X1 U19 ( .A(n26), .B(n12), .ZN(n6) );
  XNOR2_X1 U20 ( .A(n53), .B(n52), .ZN(n55) );
  XOR2_X1 U21 ( .A(n192), .B(n193), .Z(n7) );
  XOR2_X1 U22 ( .A(n191), .B(n7), .Z(n199) );
  NAND2_X1 U23 ( .A1(n191), .A2(n192), .ZN(n8) );
  NAND2_X1 U24 ( .A1(n191), .A2(n193), .ZN(n9) );
  NAND2_X1 U25 ( .A1(n192), .A2(n193), .ZN(n10) );
  NAND3_X1 U26 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n188) );
  INV_X1 U27 ( .A(n32), .ZN(n11) );
  INV_X1 U28 ( .A(n32), .ZN(n242) );
  XNOR2_X1 U29 ( .A(n26), .B(n12), .ZN(n31) );
  XNOR2_X1 U30 ( .A(n24), .B(\mult_x_1/a[2] ), .ZN(n30) );
  BUF_X2 U31 ( .A(n554), .Z(n328) );
  XNOR2_X1 U32 ( .A(n88), .B(\mult_x_1/n313 ), .ZN(n14) );
  INV_X1 U33 ( .A(n15), .ZN(n16) );
  NAND2_X2 U34 ( .A1(n19), .A2(\mult_x_1/n313 ), .ZN(n245) );
  XNOR2_X1 U35 ( .A(n137), .B(n136), .ZN(n178) );
  NOR2_X1 U36 ( .A1(n63), .A2(n62), .ZN(n36) );
  NAND2_X1 U37 ( .A1(n63), .A2(n62), .ZN(n35) );
  NAND2_X1 U38 ( .A1(n118), .A2(n117), .ZN(n123) );
  XNOR2_X1 U39 ( .A(n163), .B(n330), .ZN(n17) );
  XNOR2_X1 U40 ( .A(n163), .B(n330), .ZN(n18) );
  XNOR2_X1 U41 ( .A(n163), .B(n330), .ZN(n164) );
  BUF_X2 U42 ( .A(en), .Z(n331) );
  BUF_X2 U43 ( .A(en), .Z(n289) );
  BUF_X1 U44 ( .A(rst_n), .Z(n405) );
  INV_X1 U45 ( .A(rst_n), .ZN(n557) );
  XNOR2_X1 U46 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n27) );
  XNOR2_X1 U47 ( .A(n555), .B(n22), .ZN(n28) );
  OR2_X2 U48 ( .A1(n27), .A2(n28), .ZN(n160) );
  XNOR2_X1 U49 ( .A(n330), .B(\mult_x_1/n287 ), .ZN(n60) );
  INV_X1 U50 ( .A(n28), .ZN(n161) );
  XNOR2_X1 U51 ( .A(n330), .B(\mult_x_1/n286 ), .ZN(n45) );
  OAI22_X1 U52 ( .A1(n160), .A2(n60), .B1(n161), .B2(n45), .ZN(n75) );
  XNOR2_X1 U53 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n77) );
  XNOR2_X1 U54 ( .A(n88), .B(\mult_x_1/n313 ), .ZN(n46) );
  OAI22_X1 U55 ( .A1(n245), .A2(n77), .B1(n46), .B2(n19), .ZN(n74) );
  NOR2_X4 U56 ( .A1(n403), .A2(n402), .ZN(n163) );
  NOR2_X1 U57 ( .A1(n18), .A2(n20), .ZN(n73) );
  INV_X1 U58 ( .A(n64), .ZN(n37) );
  XNOR2_X1 U59 ( .A(\mult_x_1/a[4] ), .B(n555), .ZN(n29) );
  XNOR2_X1 U60 ( .A(n23), .B(n554), .ZN(n229) );
  OR2_X2 U61 ( .A1(n29), .A2(n229), .ZN(n151) );
  BUF_X2 U62 ( .A(n555), .Z(n329) );
  XNOR2_X1 U63 ( .A(n329), .B(\mult_x_1/n284 ), .ZN(n56) );
  XNOR2_X1 U64 ( .A(n329), .B(\mult_x_1/n283 ), .ZN(n38) );
  OAI22_X1 U65 ( .A1(n151), .A2(n56), .B1(n149), .B2(n38), .ZN(n42) );
  NAND2_X1 U66 ( .A1(n6), .A2(n30), .ZN(n78) );
  XNOR2_X1 U67 ( .A(n328), .B(\mult_x_1/n282 ), .ZN(n57) );
  INV_X1 U68 ( .A(n31), .ZN(n32) );
  XNOR2_X1 U69 ( .A(n328), .B(\mult_x_1/n281 ), .ZN(n39) );
  OAI22_X1 U70 ( .A1(n78), .A2(n57), .B1(n242), .B2(n39), .ZN(n41) );
  XNOR2_X1 U71 ( .A(n42), .B(n41), .ZN(n63) );
  INV_X1 U72 ( .A(n163), .ZN(n33) );
  OR2_X1 U73 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n34) );
  NOR2_X1 U74 ( .A1(n34), .A2(n164), .ZN(n62) );
  XNOR2_X1 U75 ( .A(n330), .B(\mult_x_1/n285 ), .ZN(n44) );
  XNOR2_X1 U76 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n105) );
  OAI22_X1 U77 ( .A1(n160), .A2(n44), .B1(n161), .B2(n105), .ZN(n110) );
  XNOR2_X1 U78 ( .A(n329), .B(\mult_x_1/n282 ), .ZN(n112) );
  OAI22_X1 U79 ( .A1(n151), .A2(n38), .B1(n149), .B2(n112), .ZN(n109) );
  XNOR2_X1 U80 ( .A(n13), .B(n328), .ZN(n106) );
  OAI22_X1 U81 ( .A1(n78), .A2(n39), .B1(n106), .B2(n242), .ZN(n40) );
  INV_X1 U82 ( .A(n40), .ZN(n108) );
  OR2_X1 U83 ( .A1(n5), .A2(n41), .ZN(n128) );
  XNOR2_X1 U84 ( .A(n163), .B(\mult_x_1/n286 ), .ZN(n43) );
  NOR2_X1 U85 ( .A1(n43), .A2(n164), .ZN(n127) );
  XNOR2_X1 U86 ( .A(n128), .B(n127), .ZN(n51) );
  OAI22_X1 U87 ( .A1(n160), .A2(n45), .B1(n161), .B2(n44), .ZN(n53) );
  AOI21_X1 U88 ( .B1(n245), .B2(n19), .A(n14), .ZN(n47) );
  INV_X1 U89 ( .A(n47), .ZN(n52) );
  XNOR2_X1 U90 ( .A(n163), .B(\mult_x_1/n287 ), .ZN(n48) );
  NOR2_X1 U91 ( .A1(n48), .A2(n17), .ZN(n54) );
  OAI21_X1 U92 ( .B1(n53), .B2(n52), .A(n54), .ZN(n50) );
  NAND2_X1 U93 ( .A1(n53), .A2(n52), .ZN(n49) );
  NAND2_X1 U94 ( .A1(n50), .A2(n49), .ZN(n126) );
  XNOR2_X1 U95 ( .A(n51), .B(n126), .ZN(n181) );
  XNOR2_X1 U96 ( .A(n55), .B(n54), .ZN(n72) );
  XNOR2_X1 U97 ( .A(n329), .B(\mult_x_1/n285 ), .ZN(n76) );
  OAI22_X1 U98 ( .A1(n151), .A2(n76), .B1(n149), .B2(n56), .ZN(n82) );
  CLKBUF_X1 U99 ( .A(n78), .Z(n240) );
  XNOR2_X1 U100 ( .A(n328), .B(\mult_x_1/n283 ), .ZN(n79) );
  OAI22_X1 U101 ( .A1(n240), .A2(n79), .B1(n11), .B2(n57), .ZN(n81) );
  INV_X1 U102 ( .A(n330), .ZN(n59) );
  OR2_X1 U103 ( .A1(\mult_x_1/n288 ), .A2(n59), .ZN(n58) );
  OAI22_X1 U104 ( .A1(n160), .A2(n59), .B1(n58), .B2(n161), .ZN(n142) );
  XNOR2_X1 U105 ( .A(n330), .B(\mult_x_1/n288 ), .ZN(n61) );
  OAI22_X1 U106 ( .A1(n160), .A2(n61), .B1(n161), .B2(n60), .ZN(n141) );
  XNOR2_X1 U107 ( .A(n63), .B(n62), .ZN(n65) );
  XNOR2_X1 U108 ( .A(n65), .B(n64), .ZN(n70) );
  NAND2_X1 U109 ( .A1(n217), .A2(n216), .ZN(n66) );
  NAND2_X1 U110 ( .A1(n66), .A2(n257), .ZN(n69) );
  INV_X1 U111 ( .A(n257), .ZN(n67) );
  NAND2_X1 U112 ( .A1(n67), .A2(n348), .ZN(n68) );
  NAND2_X1 U113 ( .A1(n69), .A2(n68), .ZN(n384) );
  FA_X1 U114 ( .A(n72), .B(n71), .CI(n70), .CO(n216), .S(n189) );
  FA_X1 U115 ( .A(n75), .B(n74), .CI(n73), .CO(n64), .S(n193) );
  XNOR2_X1 U116 ( .A(n329), .B(\mult_x_1/n286 ), .ZN(n148) );
  OAI22_X1 U117 ( .A1(n151), .A2(n148), .B1(n149), .B2(n76), .ZN(n145) );
  XNOR2_X1 U118 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n139) );
  OAI22_X1 U119 ( .A1(n245), .A2(n139), .B1(n77), .B2(n19), .ZN(n144) );
  XNOR2_X1 U120 ( .A(n328), .B(\mult_x_1/n284 ), .ZN(n140) );
  OAI22_X1 U121 ( .A1(n240), .A2(n140), .B1(n11), .B2(n79), .ZN(n143) );
  FA_X1 U122 ( .A(n82), .B(n81), .CI(n80), .CO(n71), .S(n191) );
  NAND2_X1 U123 ( .A1(n189), .A2(n188), .ZN(n83) );
  NAND2_X1 U124 ( .A1(n83), .A2(n200), .ZN(n85) );
  OR2_X1 U125 ( .A1(n200), .A2(n25), .ZN(n84) );
  NAND2_X1 U126 ( .A1(n85), .A2(n84), .ZN(n370) );
  XNOR2_X1 U147 ( .A(n163), .B(\mult_x_1/n282 ), .ZN(n86) );
  NOR2_X1 U148 ( .A1(n86), .A2(n18), .ZN(n158) );
  XNOR2_X1 U149 ( .A(n330), .B(n16), .ZN(n87) );
  XNOR2_X1 U150 ( .A(n13), .B(n330), .ZN(n159) );
  OAI22_X1 U151 ( .A1(n160), .A2(n87), .B1(n159), .B2(n161), .ZN(n169) );
  INV_X1 U152 ( .A(n169), .ZN(n157) );
  XNOR2_X1 U153 ( .A(n330), .B(\mult_x_1/n282 ), .ZN(n91) );
  OAI22_X1 U154 ( .A1(n160), .A2(n91), .B1(n161), .B2(n87), .ZN(n96) );
  XNOR2_X1 U155 ( .A(n88), .B(n329), .ZN(n90) );
  AOI21_X1 U156 ( .B1(n149), .B2(n151), .A(n90), .ZN(n89) );
  INV_X1 U157 ( .A(n89), .ZN(n95) );
  XNOR2_X1 U158 ( .A(n329), .B(\mult_x_1/n281 ), .ZN(n111) );
  OAI22_X1 U159 ( .A1(n151), .A2(n111), .B1(n90), .B2(n149), .ZN(n94) );
  INV_X1 U160 ( .A(n94), .ZN(n103) );
  XNOR2_X1 U161 ( .A(n330), .B(\mult_x_1/n283 ), .ZN(n104) );
  OAI22_X1 U162 ( .A1(n160), .A2(n104), .B1(n161), .B2(n91), .ZN(n102) );
  XNOR2_X1 U163 ( .A(n163), .B(\mult_x_1/n284 ), .ZN(n92) );
  NOR2_X1 U164 ( .A1(n92), .A2(n17), .ZN(n101) );
  XNOR2_X1 U165 ( .A(n163), .B(\mult_x_1/n283 ), .ZN(n93) );
  NOR2_X1 U166 ( .A1(n93), .A2(n17), .ZN(n99) );
  FA_X1 U167 ( .A(n96), .B(n95), .CI(n94), .CO(n156), .S(n98) );
  OR2_X1 U168 ( .A1(n176), .A2(n175), .ZN(n97) );
  MUX2_X1 U169 ( .A(n332), .B(n97), .S(n257), .Z(n352) );
  FA_X1 U170 ( .A(n100), .B(n99), .CI(n98), .CO(n175), .S(n220) );
  FA_X1 U171 ( .A(n103), .B(n102), .CI(n101), .CO(n100), .S(n124) );
  OAI22_X1 U172 ( .A1(n160), .A2(n105), .B1(n161), .B2(n104), .ZN(n133) );
  INV_X1 U173 ( .A(n108), .ZN(n132) );
  AOI21_X1 U174 ( .B1(n11), .B2(n78), .A(n106), .ZN(n107) );
  INV_X1 U175 ( .A(n107), .ZN(n131) );
  FA_X1 U176 ( .A(n110), .B(n109), .CI(n108), .CO(n137), .S(n182) );
  XNOR2_X1 U177 ( .A(n163), .B(\mult_x_1/n285 ), .ZN(n116) );
  OR2_X1 U178 ( .A1(n116), .A2(n17), .ZN(n114) );
  OAI22_X1 U179 ( .A1(n151), .A2(n112), .B1(n149), .B2(n111), .ZN(n134) );
  NAND2_X1 U180 ( .A1(n114), .A2(n113), .ZN(n115) );
  NAND2_X1 U181 ( .A1(n137), .A2(n115), .ZN(n118) );
  NOR2_X1 U182 ( .A1(n116), .A2(n164), .ZN(n135) );
  OR2_X1 U183 ( .A1(n220), .A2(n219), .ZN(n121) );
  MUX2_X1 U184 ( .A(n333), .B(n121), .S(n257), .Z(n354) );
  XNOR2_X1 U185 ( .A(n123), .B(n122), .ZN(n125) );
  XNOR2_X1 U186 ( .A(n125), .B(n124), .ZN(n223) );
  FA_X1 U187 ( .A(n133), .B(n132), .CI(n131), .CO(n122), .S(n179) );
  OR2_X1 U188 ( .A1(n223), .A2(n222), .ZN(n138) );
  MUX2_X1 U189 ( .A(n334), .B(n138), .S(n200), .Z(n356) );
  XNOR2_X1 U190 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n209) );
  OAI22_X1 U191 ( .A1(n245), .A2(n209), .B1(n139), .B2(n19), .ZN(n154) );
  AND2_X1 U192 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n153) );
  XNOR2_X1 U193 ( .A(n328), .B(\mult_x_1/n285 ), .ZN(n208) );
  OAI22_X1 U194 ( .A1(n240), .A2(n208), .B1(n11), .B2(n140), .ZN(n152) );
  HA_X1 U195 ( .A(n142), .B(n141), .CO(n80), .S(n195) );
  FA_X1 U196 ( .A(n145), .B(n144), .CI(n143), .CO(n192), .S(n194) );
  OR2_X1 U197 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n146) );
  OAI22_X1 U198 ( .A1(n151), .A2(n21), .B1(n146), .B2(n149), .ZN(n211) );
  XNOR2_X1 U199 ( .A(n329), .B(\mult_x_1/n288 ), .ZN(n147) );
  XNOR2_X1 U200 ( .A(n329), .B(\mult_x_1/n287 ), .ZN(n150) );
  OAI22_X1 U201 ( .A1(n151), .A2(n147), .B1(n149), .B2(n150), .ZN(n210) );
  OAI22_X1 U202 ( .A1(n151), .A2(n150), .B1(n149), .B2(n148), .ZN(n206) );
  FA_X1 U203 ( .A(n154), .B(n153), .CI(n152), .CO(n196), .S(n205) );
  OR2_X1 U204 ( .A1(n203), .A2(n202), .ZN(n155) );
  MUX2_X1 U205 ( .A(n335), .B(n155), .S(n200), .Z(n358) );
  FA_X1 U206 ( .A(n158), .B(n157), .CI(n156), .CO(n171), .S(n176) );
  AOI21_X1 U207 ( .B1(n161), .B2(n160), .A(n159), .ZN(n162) );
  INV_X1 U208 ( .A(n162), .ZN(n167) );
  XNOR2_X1 U209 ( .A(n163), .B(n16), .ZN(n165) );
  NOR2_X1 U210 ( .A1(n165), .A2(n18), .ZN(n166) );
  XOR2_X1 U211 ( .A(n167), .B(n166), .Z(n168) );
  XOR2_X1 U212 ( .A(n169), .B(n168), .Z(n170) );
  OR2_X1 U213 ( .A1(n171), .A2(n170), .ZN(n173) );
  NAND2_X1 U214 ( .A1(n171), .A2(n170), .ZN(n172) );
  NAND2_X1 U215 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2_X1 U216 ( .A(n336), .B(n174), .S(n200), .Z(n360) );
  NAND2_X1 U217 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U218 ( .A(n337), .B(n177), .S(n200), .Z(n362) );
  FA_X1 U219 ( .A(n180), .B(n179), .CI(n178), .CO(n222), .S(n186) );
  FA_X1 U220 ( .A(n183), .B(n182), .CI(n181), .CO(n185), .S(n217) );
  NOR2_X1 U221 ( .A1(n186), .A2(n185), .ZN(n184) );
  MUX2_X1 U222 ( .A(n338), .B(n184), .S(n200), .Z(n364) );
  NAND2_X1 U223 ( .A1(n186), .A2(n185), .ZN(n187) );
  MUX2_X1 U224 ( .A(n339), .B(n187), .S(n200), .Z(n366) );
  NOR2_X1 U225 ( .A1(n189), .A2(n188), .ZN(n190) );
  MUX2_X1 U226 ( .A(n340), .B(n190), .S(n200), .Z(n368) );
  FA_X1 U227 ( .A(n196), .B(n195), .CI(n194), .CO(n198), .S(n203) );
  NOR2_X1 U228 ( .A1(n199), .A2(n198), .ZN(n197) );
  MUX2_X1 U229 ( .A(n342), .B(n197), .S(n200), .Z(n372) );
  NAND2_X1 U230 ( .A1(n199), .A2(n198), .ZN(n201) );
  MUX2_X1 U231 ( .A(n343), .B(n201), .S(n200), .Z(n374) );
  NAND2_X1 U232 ( .A1(n203), .A2(n202), .ZN(n204) );
  MUX2_X1 U233 ( .A(n344), .B(n204), .S(n257), .Z(n376) );
  FA_X1 U234 ( .A(n207), .B(n206), .CI(n205), .CO(n202), .S(n214) );
  XNOR2_X1 U235 ( .A(n328), .B(\mult_x_1/n286 ), .ZN(n230) );
  OAI22_X1 U236 ( .A1(n240), .A2(n230), .B1(n11), .B2(n208), .ZN(n227) );
  XNOR2_X1 U237 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n228) );
  OAI22_X1 U238 ( .A1(n245), .A2(n228), .B1(n209), .B2(n19), .ZN(n226) );
  HA_X1 U239 ( .A(n211), .B(n210), .CO(n207), .S(n225) );
  NOR2_X1 U240 ( .A1(n214), .A2(n213), .ZN(n212) );
  MUX2_X1 U241 ( .A(n345), .B(n212), .S(n257), .Z(n378) );
  NAND2_X1 U242 ( .A1(n214), .A2(n213), .ZN(n215) );
  MUX2_X1 U243 ( .A(n346), .B(n215), .S(n257), .Z(n380) );
  NOR2_X1 U244 ( .A1(n217), .A2(n216), .ZN(n218) );
  MUX2_X1 U245 ( .A(n347), .B(n218), .S(n257), .Z(n382) );
  NAND2_X1 U246 ( .A1(n220), .A2(n219), .ZN(n221) );
  MUX2_X1 U247 ( .A(n349), .B(n221), .S(n257), .Z(n386) );
  NAND2_X1 U248 ( .A1(n223), .A2(n222), .ZN(n224) );
  MUX2_X1 U249 ( .A(n350), .B(n224), .S(n257), .Z(n388) );
  FA_X1 U250 ( .A(n227), .B(n226), .CI(n225), .CO(n213), .S(n255) );
  XNOR2_X1 U251 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n236) );
  OAI22_X1 U252 ( .A1(n245), .A2(n236), .B1(n228), .B2(n19), .ZN(n233) );
  AND2_X1 U253 ( .A1(n229), .A2(\mult_x_1/n288 ), .ZN(n232) );
  XNOR2_X1 U254 ( .A(n328), .B(\mult_x_1/n287 ), .ZN(n234) );
  OAI22_X1 U255 ( .A1(n240), .A2(n234), .B1(n11), .B2(n230), .ZN(n231) );
  OR2_X1 U256 ( .A1(n255), .A2(n254), .ZN(n282) );
  FA_X1 U257 ( .A(n233), .B(n232), .CI(n231), .CO(n254), .S(n253) );
  XNOR2_X1 U258 ( .A(n328), .B(\mult_x_1/n288 ), .ZN(n235) );
  OAI22_X1 U259 ( .A1(n78), .A2(n235), .B1(n11), .B2(n234), .ZN(n238) );
  XNOR2_X1 U260 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n241) );
  OAI22_X1 U261 ( .A1(n245), .A2(n241), .B1(n236), .B2(n19), .ZN(n237) );
  NOR2_X1 U262 ( .A1(n253), .A2(n252), .ZN(n275) );
  HA_X1 U263 ( .A(n238), .B(n237), .CO(n252), .S(n250) );
  OR2_X1 U264 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n239) );
  OAI22_X1 U265 ( .A1(n240), .A2(n24), .B1(n239), .B2(n11), .ZN(n249) );
  OR2_X1 U266 ( .A1(n250), .A2(n249), .ZN(n271) );
  XNOR2_X1 U267 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n244) );
  OAI22_X1 U268 ( .A1(n245), .A2(n244), .B1(n241), .B2(n19), .ZN(n248) );
  INV_X1 U269 ( .A(n11), .ZN(n243) );
  AND2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(n243), .ZN(n247) );
  NOR2_X1 U271 ( .A1(n248), .A2(n247), .ZN(n264) );
  OAI22_X1 U272 ( .A1(n245), .A2(\mult_x_1/n288 ), .B1(n244), .B2(n19), .ZN(
        n261) );
  OR2_X1 U273 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n246) );
  NAND2_X1 U274 ( .A1(n246), .A2(n245), .ZN(n260) );
  NAND2_X1 U275 ( .A1(n261), .A2(n260), .ZN(n267) );
  NAND2_X1 U276 ( .A1(n248), .A2(n247), .ZN(n265) );
  OAI21_X1 U277 ( .B1(n264), .B2(n267), .A(n265), .ZN(n272) );
  NAND2_X1 U278 ( .A1(n250), .A2(n249), .ZN(n270) );
  INV_X1 U279 ( .A(n270), .ZN(n251) );
  AOI21_X1 U280 ( .B1(n271), .B2(n272), .A(n251), .ZN(n278) );
  NAND2_X1 U281 ( .A1(n253), .A2(n252), .ZN(n276) );
  OAI21_X1 U282 ( .B1(n275), .B2(n278), .A(n276), .ZN(n283) );
  NAND2_X1 U283 ( .A1(n255), .A2(n254), .ZN(n281) );
  INV_X1 U284 ( .A(n281), .ZN(n256) );
  AOI21_X1 U285 ( .B1(n282), .B2(n283), .A(n256), .ZN(n258) );
  MUX2_X1 U286 ( .A(n351), .B(n258), .S(n257), .Z(n390) );
  BUF_X2 U287 ( .A(rst_n), .Z(n404) );
  MUX2_X1 U288 ( .A(product[0]), .B(n517), .S(n331), .Z(n407) );
  MUX2_X1 U289 ( .A(n517), .B(n518), .S(n331), .Z(n409) );
  AND2_X1 U290 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n259) );
  MUX2_X1 U291 ( .A(n518), .B(n259), .S(n331), .Z(n411) );
  MUX2_X1 U292 ( .A(product[1]), .B(n520), .S(n331), .Z(n413) );
  MUX2_X1 U293 ( .A(n520), .B(n521), .S(n331), .Z(n415) );
  OR2_X1 U294 ( .A1(n261), .A2(n260), .ZN(n262) );
  AND2_X1 U295 ( .A1(n262), .A2(n267), .ZN(n263) );
  MUX2_X1 U296 ( .A(n521), .B(n263), .S(n331), .Z(n417) );
  MUX2_X1 U297 ( .A(product[2]), .B(n523), .S(n331), .Z(n419) );
  MUX2_X1 U298 ( .A(n523), .B(n524), .S(n331), .Z(n421) );
  INV_X1 U299 ( .A(n264), .ZN(n266) );
  NAND2_X1 U300 ( .A1(n266), .A2(n265), .ZN(n268) );
  XOR2_X1 U301 ( .A(n268), .B(n267), .Z(n269) );
  MUX2_X1 U302 ( .A(n524), .B(n269), .S(n331), .Z(n423) );
  MUX2_X1 U303 ( .A(product[3]), .B(n526), .S(n331), .Z(n425) );
  MUX2_X1 U304 ( .A(n526), .B(n527), .S(n331), .Z(n427) );
  NAND2_X1 U305 ( .A1(n271), .A2(n270), .ZN(n273) );
  XNOR2_X1 U306 ( .A(n273), .B(n272), .ZN(n274) );
  MUX2_X1 U307 ( .A(n527), .B(n274), .S(n331), .Z(n429) );
  MUX2_X1 U308 ( .A(product[4]), .B(n529), .S(n331), .Z(n431) );
  MUX2_X1 U309 ( .A(n529), .B(n530), .S(n331), .Z(n433) );
  INV_X1 U310 ( .A(n275), .ZN(n277) );
  NAND2_X1 U311 ( .A1(n277), .A2(n276), .ZN(n279) );
  XOR2_X1 U312 ( .A(n279), .B(n278), .Z(n280) );
  MUX2_X1 U313 ( .A(n530), .B(n280), .S(n331), .Z(n435) );
  MUX2_X1 U314 ( .A(product[5]), .B(n532), .S(n331), .Z(n437) );
  MUX2_X1 U315 ( .A(n532), .B(n533), .S(n331), .Z(n439) );
  NAND2_X1 U316 ( .A1(n282), .A2(n281), .ZN(n284) );
  XNOR2_X1 U317 ( .A(n284), .B(n283), .ZN(n285) );
  MUX2_X1 U318 ( .A(n533), .B(n285), .S(n331), .Z(n441) );
  MUX2_X1 U319 ( .A(product[6]), .B(n535), .S(n331), .Z(n443) );
  NAND2_X1 U320 ( .A1(n395), .A2(n346), .ZN(n286) );
  XOR2_X1 U321 ( .A(n286), .B(n351), .Z(n287) );
  MUX2_X1 U322 ( .A(n535), .B(n287), .S(n331), .Z(n445) );
  MUX2_X1 U323 ( .A(product[7]), .B(n537), .S(n331), .Z(n447) );
  OAI21_X1 U324 ( .B1(n345), .B2(n351), .A(n346), .ZN(n291) );
  NAND2_X1 U325 ( .A1(n335), .A2(n344), .ZN(n288) );
  XNOR2_X1 U326 ( .A(n291), .B(n288), .ZN(n290) );
  MUX2_X1 U327 ( .A(n537), .B(n290), .S(n331), .Z(n449) );
  MUX2_X1 U328 ( .A(product[8]), .B(n539), .S(n289), .Z(n451) );
  AOI21_X1 U329 ( .B1(n291), .B2(n335), .A(n396), .ZN(n294) );
  NAND2_X1 U330 ( .A1(n397), .A2(n343), .ZN(n292) );
  XOR2_X1 U331 ( .A(n294), .B(n292), .Z(n293) );
  MUX2_X1 U332 ( .A(n539), .B(n293), .S(n289), .Z(n453) );
  MUX2_X1 U333 ( .A(product[9]), .B(n541), .S(n289), .Z(n455) );
  OAI21_X1 U334 ( .B1(n294), .B2(n342), .A(n343), .ZN(n302) );
  INV_X1 U335 ( .A(n302), .ZN(n297) );
  NAND2_X1 U336 ( .A1(n398), .A2(n341), .ZN(n295) );
  XOR2_X1 U337 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U338 ( .A(n541), .B(n296), .S(n289), .Z(n457) );
  MUX2_X1 U339 ( .A(product[10]), .B(n543), .S(n289), .Z(n459) );
  OAI21_X1 U340 ( .B1(n297), .B2(n340), .A(n341), .ZN(n299) );
  NAND2_X1 U341 ( .A1(n400), .A2(n348), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U343 ( .A(n543), .B(n300), .S(n289), .Z(n461) );
  MUX2_X1 U344 ( .A(product[11]), .B(n545), .S(n289), .Z(n463) );
  NOR2_X1 U345 ( .A1(n347), .A2(n340), .ZN(n303) );
  OAI21_X1 U346 ( .B1(n347), .B2(n341), .A(n348), .ZN(n301) );
  AOI21_X1 U347 ( .B1(n303), .B2(n302), .A(n301), .ZN(n325) );
  NAND2_X1 U348 ( .A1(n399), .A2(n339), .ZN(n304) );
  XOR2_X1 U349 ( .A(n325), .B(n304), .Z(n305) );
  MUX2_X1 U350 ( .A(n545), .B(n305), .S(n289), .Z(n465) );
  MUX2_X1 U351 ( .A(product[12]), .B(n547), .S(n289), .Z(n467) );
  OAI21_X1 U352 ( .B1(n325), .B2(n338), .A(n339), .ZN(n307) );
  NAND2_X1 U353 ( .A1(n334), .A2(n350), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  MUX2_X1 U355 ( .A(n547), .B(n308), .S(n289), .Z(n469) );
  MUX2_X1 U356 ( .A(product[13]), .B(n549), .S(n289), .Z(n471) );
  NAND2_X1 U357 ( .A1(n399), .A2(n334), .ZN(n310) );
  AOI21_X1 U358 ( .B1(n394), .B2(n334), .A(n401), .ZN(n309) );
  OAI21_X1 U359 ( .B1(n325), .B2(n310), .A(n309), .ZN(n312) );
  NAND2_X1 U360 ( .A1(n333), .A2(n349), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U362 ( .A(n549), .B(n313), .S(n289), .Z(n473) );
  MUX2_X1 U363 ( .A(product[14]), .B(n551), .S(n289), .Z(n475) );
  NAND2_X1 U364 ( .A1(n334), .A2(n333), .ZN(n315) );
  NOR2_X1 U365 ( .A1(n338), .A2(n315), .ZN(n321) );
  INV_X1 U366 ( .A(n321), .ZN(n317) );
  AOI21_X1 U367 ( .B1(n401), .B2(n333), .A(n393), .ZN(n314) );
  OAI21_X1 U368 ( .B1(n315), .B2(n339), .A(n314), .ZN(n322) );
  INV_X1 U369 ( .A(n322), .ZN(n316) );
  OAI21_X1 U370 ( .B1(n325), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U371 ( .A1(n332), .A2(n337), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U373 ( .A(n551), .B(n320), .S(n289), .Z(n477) );
  MUX2_X1 U374 ( .A(product[15]), .B(n553), .S(n289), .Z(n479) );
  NAND2_X1 U375 ( .A1(n321), .A2(n332), .ZN(n324) );
  AOI21_X1 U376 ( .B1(n322), .B2(n332), .A(n392), .ZN(n323) );
  OAI21_X1 U377 ( .B1(n325), .B2(n324), .A(n323), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(n336), .ZN(n327) );
  MUX2_X1 U379 ( .A(n553), .B(n327), .S(n289), .Z(n481) );
  MUX2_X1 U380 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n331), .Z(n483) );
  MUX2_X1 U381 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n331), .Z(n485) );
  MUX2_X1 U382 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n331), .Z(n487) );
  MUX2_X1 U383 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n331), .Z(n489) );
  MUX2_X1 U384 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n331), .Z(n491) );
  MUX2_X1 U385 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n331), .Z(n493) );
  MUX2_X1 U386 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n331), .Z(n495) );
  MUX2_X1 U387 ( .A(n16), .B(B_extended[7]), .S(n331), .Z(n497) );
  MUX2_X1 U388 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n331), .Z(n499) );
  MUX2_X1 U389 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n331), .Z(n501) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n331), .Z(n503) );
  MUX2_X1 U391 ( .A(n328), .B(A_extended[3]), .S(n331), .Z(n505) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n331), .Z(n507) );
  MUX2_X1 U393 ( .A(n329), .B(A_extended[5]), .S(n331), .Z(n509) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n331), .Z(n511) );
  MUX2_X1 U395 ( .A(n330), .B(A_extended[7]), .S(n331), .Z(n513) );
  OR2_X1 U396 ( .A1(n331), .A2(n556), .ZN(n515) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_9 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n374, n376, n378, n380, n382, n384, n386, n388,
         n390, n392, n394, n396, n398, n400, n402, n404, n406, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n422, n424, n426, n428, n430, n432, n434, n436, n438, n440, n442,
         n444, n446, n448, n450, n452, n454, n456, n458, n460, n462, n464,
         n466, n468, n470, n472, n474, n476, n478, n480, n482, n484, n486,
         n488, n490, n492, n494, n496, n498, n500, n502, n504, n506, n508,
         n510, n512, n514, n516, n518, n520, n522, n524, n526, n528, n530,
         n532, n534, n535, n537, n538, n540, n541, n543, n544, n546, n547,
         n549, n550, n552, n553, n555, n557, n559, n561, n563, n565, n567,
         n569, n571, n572, n573, n574;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n420), .SE(n532), .CK(clk), .Q(n573)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n420), .SE(n528), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n34) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n420), .SE(n526), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n417) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n420), .SE(n524), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n29) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n420), .SE(n520), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n21) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n420), .SE(n516), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n420), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n18) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n420), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n420), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n419), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n419), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n419), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n419), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n419), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n419), .SE(n498), .CK(clk), .Q(n571)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n419), .SE(n496), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n419), .SE(n494), .CK(clk), .Q(n569)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n419), .SE(n492), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n419), .SE(n490), .CK(clk), .Q(n567)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n419), .SE(n488), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n418), .SE(n486), .CK(clk), .Q(n565)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n418), .SE(n484), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n418), .SE(n482), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n418), .SE(n480), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n418), .SE(n478), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n418), .SE(n476), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n418), .SE(n474), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n418), .SE(n472), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n418), .SE(n470), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n418), .SE(n468), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n418), .SE(n466), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n418), .SE(n464), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n418), .SE(n462), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n418), .SE(n460), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n418), .SE(n458), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n418), .SE(n456), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n420), .SE(n454), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n418), .SE(n452), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(rst_n), .SE(n450), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(rst_n), .SE(n448), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n419), .SE(n442), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n418), .SE(n440), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n418), .SE(n438), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n419), .SE(n436), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n418), .SE(n434), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n418), .SE(n432), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n420), .SE(n430), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n274), .SE(n428), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n274), .SE(n426), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n274), .SE(n424), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n420), .SE(n530), .CK(clk), .Q(n572), 
        .QN(n353) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n420), .SE(n518), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n33) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n420), .SE(n522), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n574), .SE(n406), .CK(
        clk), .QN(n371) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n574), .SI(1'b1), .SE(n404), .CK(clk), 
        .Q(n370), .QN(n32) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n574), .SI(1'b1), .SE(n402), .CK(clk), 
        .Q(n369), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n574), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n368) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n574), .SE(n398), .CK(
        clk), .QN(n367) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n574), .SE(n396), .CK(
        clk), .Q(n411), .QN(n366) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n574), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n365), .QN(n416) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n574), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n364), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n574), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n363), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n574), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n574), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n361), .QN(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n574), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n574), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n359), .QN(n415) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n574), .SE(n380), .CK(
        clk), .Q(n410), .QN(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n574), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n357), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n574), .SE(n376), .CK(
        clk), .QN(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n574), .SE(n374), .CK(
        clk), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n574), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n354) );
  BUF_X1 U2 ( .A(n40), .Z(n147) );
  NOR2_X1 U3 ( .A1(n57), .A2(n148), .ZN(n167) );
  BUF_X1 U4 ( .A(n54), .Z(n148) );
  BUF_X2 U5 ( .A(en), .Z(n352) );
  BUF_X4 U6 ( .A(en), .Z(n312) );
  CLKBUF_X2 U7 ( .A(n274), .Z(n418) );
  INV_X1 U8 ( .A(n249), .ZN(n27) );
  CLKBUF_X1 U9 ( .A(n302), .Z(n7) );
  XNOR2_X1 U10 ( .A(n108), .B(n349), .ZN(n8) );
  CLKBUF_X1 U11 ( .A(\mult_x_1/n281 ), .Z(n9) );
  BUF_X1 U12 ( .A(n206), .Z(n10) );
  NAND2_X1 U13 ( .A1(n70), .A2(n30), .ZN(n50) );
  CLKBUF_X1 U14 ( .A(n168), .Z(n16) );
  CLKBUF_X1 U15 ( .A(n353), .Z(n11) );
  AOI22_X1 U16 ( .A1(n177), .A2(n98), .B1(n175), .B2(n174), .ZN(n99) );
  OR2_X1 U17 ( .A1(n175), .A2(n174), .ZN(n98) );
  NAND2_X1 U18 ( .A1(n229), .A2(n228), .ZN(n265) );
  NAND2_X1 U19 ( .A1(n231), .A2(n230), .ZN(n228) );
  NAND2_X1 U20 ( .A1(n233), .A2(n31), .ZN(n229) );
  XNOR2_X1 U21 ( .A(n70), .B(n69), .ZN(n182) );
  NAND2_X1 U22 ( .A1(n50), .A2(n49), .ZN(n212) );
  NAND2_X1 U23 ( .A1(n170), .A2(n169), .ZN(n210) );
  XNOR2_X1 U24 ( .A(n68), .B(n67), .ZN(n69) );
  NAND2_X1 U25 ( .A1(n68), .A2(n67), .ZN(n49) );
  INV_X1 U26 ( .A(n56), .ZN(n12) );
  OAI22_X1 U27 ( .A1(n135), .A2(n59), .B1(n133), .B2(n78), .ZN(n13) );
  XNOR2_X1 U28 ( .A(n221), .B(n14), .ZN(n266) );
  XNOR2_X1 U29 ( .A(n223), .B(n222), .ZN(n14) );
  BUF_X1 U30 ( .A(n123), .Z(n15) );
  BUF_X1 U31 ( .A(n123), .Z(n247) );
  INV_X1 U32 ( .A(n55), .ZN(n17) );
  AND2_X1 U33 ( .A1(n573), .A2(n572), .ZN(n40) );
  INV_X1 U34 ( .A(n99), .ZN(n163) );
  XNOR2_X1 U35 ( .A(n28), .B(n18), .ZN(n85) );
  NAND2_X2 U36 ( .A1(n48), .A2(n47), .ZN(n135) );
  INV_X1 U37 ( .A(n235), .ZN(n19) );
  INV_X1 U38 ( .A(n235), .ZN(n20) );
  INV_X1 U39 ( .A(n235), .ZN(n133) );
  AND2_X2 U40 ( .A1(n573), .A2(\mult_x_1/n281 ), .ZN(n108) );
  XNOR2_X1 U41 ( .A(n21), .B(\mult_x_1/n312 ), .ZN(n45) );
  OAI22_X1 U42 ( .A1(n135), .A2(n80), .B1(n111), .B2(n19), .ZN(n22) );
  NAND2_X1 U43 ( .A1(n16), .A2(n167), .ZN(n169) );
  AOI21_X1 U44 ( .B1(n306), .B2(n307), .A(n264), .ZN(n23) );
  XNOR2_X1 U45 ( .A(n177), .B(n176), .ZN(n208) );
  XNOR2_X1 U46 ( .A(n175), .B(n174), .ZN(n176) );
  OR2_X1 U47 ( .A1(n13), .A2(n96), .ZN(n174) );
  NAND2_X1 U48 ( .A1(n221), .A2(n223), .ZN(n24) );
  NAND2_X1 U49 ( .A1(n221), .A2(n222), .ZN(n25) );
  NAND2_X1 U50 ( .A1(n223), .A2(n222), .ZN(n26) );
  NAND3_X1 U51 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n192) );
  INV_X1 U52 ( .A(n249), .ZN(n245) );
  BUF_X1 U53 ( .A(n274), .Z(n419) );
  BUF_X1 U54 ( .A(n274), .Z(n420) );
  BUF_X2 U55 ( .A(n572), .Z(n351) );
  INV_X1 U56 ( .A(rst_n), .ZN(n574) );
  OR2_X1 U57 ( .A1(n68), .A2(n67), .ZN(n30) );
  OR2_X1 U58 ( .A1(n231), .A2(n230), .ZN(n31) );
  AND2_X1 U59 ( .A1(n163), .A2(n162), .ZN(n35) );
  BUF_X2 U60 ( .A(\mult_x_1/n313 ), .Z(n349) );
  NAND2_X2 U61 ( .A1(n349), .A2(n5), .ZN(n251) );
  XNOR2_X1 U62 ( .A(n108), .B(n349), .ZN(n53) );
  AOI21_X1 U63 ( .B1(n251), .B2(n5), .A(n8), .ZN(n36) );
  INV_X1 U64 ( .A(n36), .ZN(n94) );
  XNOR2_X1 U65 ( .A(n572), .B(n34), .ZN(n37) );
  XNOR2_X1 U66 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n38) );
  NAND2_X1 U67 ( .A1(n37), .A2(n38), .ZN(n42) );
  BUF_X1 U68 ( .A(n42), .Z(n84) );
  XNOR2_X1 U69 ( .A(n351), .B(\mult_x_1/n286 ), .ZN(n51) );
  INV_X1 U70 ( .A(n38), .ZN(n39) );
  CLKBUF_X2 U71 ( .A(n38), .Z(n145) );
  XNOR2_X1 U72 ( .A(n351), .B(\mult_x_1/n285 ), .ZN(n76) );
  OAI22_X1 U73 ( .A1(n84), .A2(n51), .B1(n145), .B2(n76), .ZN(n93) );
  XNOR2_X1 U74 ( .A(n147), .B(\mult_x_1/n287 ), .ZN(n41) );
  XNOR2_X1 U75 ( .A(n40), .B(n351), .ZN(n54) );
  NOR2_X1 U76 ( .A1(n41), .A2(n148), .ZN(n92) );
  BUF_X2 U77 ( .A(n42), .Z(n144) );
  OR2_X1 U78 ( .A1(\mult_x_1/n288 ), .A2(n11), .ZN(n43) );
  OAI22_X1 U79 ( .A1(n144), .A2(n11), .B1(n43), .B2(n145), .ZN(n125) );
  XNOR2_X1 U80 ( .A(n351), .B(\mult_x_1/n288 ), .ZN(n44) );
  XNOR2_X1 U81 ( .A(n351), .B(\mult_x_1/n287 ), .ZN(n52) );
  OAI22_X1 U82 ( .A1(n144), .A2(n44), .B1(n145), .B2(n52), .ZN(n124) );
  XNOR2_X1 U83 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n46) );
  NAND2_X1 U84 ( .A1(n45), .A2(n46), .ZN(n123) );
  BUF_X2 U85 ( .A(\mult_x_1/n312 ), .Z(n350) );
  XNOR2_X1 U86 ( .A(n350), .B(\mult_x_1/n283 ), .ZN(n66) );
  INV_X1 U87 ( .A(n46), .ZN(n249) );
  XNOR2_X1 U88 ( .A(n350), .B(\mult_x_1/n282 ), .ZN(n58) );
  OAI22_X1 U89 ( .A1(n247), .A2(n66), .B1(n27), .B2(n58), .ZN(n68) );
  XNOR2_X1 U90 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n48) );
  XNOR2_X1 U91 ( .A(\mult_x_1/n311 ), .B(n29), .ZN(n47) );
  BUF_X2 U92 ( .A(\mult_x_1/n311 ), .Z(n130) );
  XNOR2_X1 U93 ( .A(n130), .B(\mult_x_1/n285 ), .ZN(n64) );
  INV_X1 U94 ( .A(n48), .ZN(n235) );
  XNOR2_X1 U95 ( .A(n130), .B(\mult_x_1/n284 ), .ZN(n59) );
  OAI22_X1 U96 ( .A1(n135), .A2(n64), .B1(n19), .B2(n59), .ZN(n67) );
  OAI22_X1 U97 ( .A1(n84), .A2(n52), .B1(n145), .B2(n51), .ZN(n63) );
  XNOR2_X1 U98 ( .A(n349), .B(\mult_x_1/n281 ), .ZN(n65) );
  OAI22_X1 U99 ( .A1(n251), .A2(n65), .B1(n53), .B2(n5), .ZN(n62) );
  INV_X1 U100 ( .A(n54), .ZN(n55) );
  AND2_X1 U101 ( .A1(\mult_x_1/n288 ), .A2(n55), .ZN(n61) );
  INV_X1 U102 ( .A(n147), .ZN(n56) );
  OR2_X1 U103 ( .A1(\mult_x_1/n288 ), .A2(n56), .ZN(n57) );
  OAI22_X1 U104 ( .A1(n123), .A2(n58), .B1(n245), .B2(n85), .ZN(n96) );
  XNOR2_X1 U105 ( .A(n130), .B(\mult_x_1/n283 ), .ZN(n78) );
  OAI22_X1 U106 ( .A1(n135), .A2(n59), .B1(n133), .B2(n78), .ZN(n97) );
  XNOR2_X1 U107 ( .A(n97), .B(n96), .ZN(n168) );
  XNOR2_X1 U108 ( .A(n168), .B(n167), .ZN(n60) );
  XNOR2_X1 U109 ( .A(n166), .B(n60), .ZN(n211) );
  FA_X1 U110 ( .A(n63), .B(n62), .CI(n61), .CO(n166), .S(n184) );
  XNOR2_X1 U111 ( .A(n130), .B(\mult_x_1/n286 ), .ZN(n132) );
  OAI22_X1 U112 ( .A1(n135), .A2(n132), .B1(n20), .B2(n64), .ZN(n128) );
  XNOR2_X1 U113 ( .A(n349), .B(\mult_x_1/n282 ), .ZN(n121) );
  OAI22_X1 U114 ( .A1(n251), .A2(n121), .B1(n65), .B2(n5), .ZN(n127) );
  XNOR2_X1 U115 ( .A(n350), .B(\mult_x_1/n284 ), .ZN(n122) );
  OAI22_X1 U116 ( .A1(n15), .A2(n122), .B1(n27), .B2(n66), .ZN(n126) );
  NAND2_X1 U117 ( .A1(n180), .A2(n179), .ZN(n71) );
  NAND2_X1 U118 ( .A1(n71), .A2(n312), .ZN(n74) );
  INV_X1 U119 ( .A(n312), .ZN(n72) );
  NAND2_X1 U120 ( .A1(n72), .A2(n360), .ZN(n73) );
  NAND2_X1 U121 ( .A1(n74), .A2(n73), .ZN(n384) );
  XNOR2_X1 U122 ( .A(n147), .B(\mult_x_1/n285 ), .ZN(n75) );
  NOR2_X1 U123 ( .A1(n75), .A2(n17), .ZN(n91) );
  XNOR2_X1 U124 ( .A(n130), .B(\mult_x_1/n282 ), .ZN(n77) );
  XNOR2_X1 U125 ( .A(n130), .B(\mult_x_1/n281 ), .ZN(n80) );
  OAI22_X1 U126 ( .A1(n135), .A2(n77), .B1(n19), .B2(n80), .ZN(n90) );
  XNOR2_X1 U127 ( .A(n351), .B(\mult_x_1/n284 ), .ZN(n83) );
  OAI22_X1 U128 ( .A1(n144), .A2(n76), .B1(n145), .B2(n83), .ZN(n173) );
  OAI22_X1 U129 ( .A1(n135), .A2(n78), .B1(n20), .B2(n77), .ZN(n172) );
  XNOR2_X1 U130 ( .A(n108), .B(n350), .ZN(n86) );
  OAI22_X1 U131 ( .A1(n123), .A2(n85), .B1(n86), .B2(n245), .ZN(n79) );
  INV_X1 U132 ( .A(n79), .ZN(n171) );
  XNOR2_X1 U133 ( .A(n108), .B(n130), .ZN(n111) );
  OAI22_X1 U134 ( .A1(n135), .A2(n80), .B1(n111), .B2(n19), .ZN(n118) );
  INV_X1 U135 ( .A(n118), .ZN(n115) );
  XNOR2_X1 U136 ( .A(n351), .B(\mult_x_1/n283 ), .ZN(n82) );
  XNOR2_X1 U137 ( .A(n351), .B(\mult_x_1/n282 ), .ZN(n110) );
  OAI22_X1 U138 ( .A1(n144), .A2(n82), .B1(n145), .B2(n110), .ZN(n114) );
  XNOR2_X1 U139 ( .A(n147), .B(\mult_x_1/n284 ), .ZN(n81) );
  NOR2_X1 U140 ( .A1(n81), .A2(n148), .ZN(n113) );
  OAI22_X1 U141 ( .A1(n84), .A2(n83), .B1(n145), .B2(n82), .ZN(n102) );
  OAI22_X1 U142 ( .A1(n123), .A2(n85), .B1(n86), .B2(n27), .ZN(n101) );
  AOI21_X1 U143 ( .B1(n27), .B2(n15), .A(n86), .ZN(n87) );
  INV_X1 U144 ( .A(n87), .ZN(n100) );
  XNOR2_X1 U145 ( .A(n200), .B(n199), .ZN(n88) );
  XNOR2_X1 U146 ( .A(n88), .B(n198), .ZN(n206) );
  FA_X1 U147 ( .A(n91), .B(n90), .CI(n89), .CO(n198), .S(n164) );
  FA_X1 U148 ( .A(n94), .B(n93), .CI(n92), .CO(n177), .S(n213) );
  XNOR2_X1 U149 ( .A(n147), .B(\mult_x_1/n286 ), .ZN(n95) );
  NOR2_X1 U150 ( .A1(n95), .A2(n148), .ZN(n175) );
  FA_X1 U151 ( .A(n102), .B(n101), .CI(n100), .CO(n199), .S(n162) );
  AOI21_X1 U152 ( .B1(n164), .B2(n163), .A(n35), .ZN(n104) );
  NAND2_X1 U153 ( .A1(n164), .A2(n162), .ZN(n103) );
  NAND2_X1 U154 ( .A1(n104), .A2(n103), .ZN(n205) );
  OAI21_X1 U155 ( .B1(n10), .B2(n205), .A(n312), .ZN(n106) );
  OR2_X1 U156 ( .A1(n312), .A2(n32), .ZN(n105) );
  NAND2_X1 U157 ( .A1(n106), .A2(n105), .ZN(n404) );
  XNOR2_X1 U176 ( .A(n12), .B(\mult_x_1/n282 ), .ZN(n107) );
  NOR2_X1 U177 ( .A1(n107), .A2(n17), .ZN(n142) );
  XNOR2_X1 U178 ( .A(n351), .B(\mult_x_1/n281 ), .ZN(n109) );
  XNOR2_X1 U179 ( .A(n108), .B(n351), .ZN(n143) );
  OAI22_X1 U180 ( .A1(n144), .A2(n109), .B1(n143), .B2(n145), .ZN(n153) );
  INV_X1 U181 ( .A(n153), .ZN(n141) );
  OAI22_X1 U182 ( .A1(n144), .A2(n110), .B1(n145), .B2(n109), .ZN(n119) );
  AOI21_X1 U183 ( .B1(n20), .B2(n135), .A(n111), .ZN(n112) );
  INV_X1 U184 ( .A(n112), .ZN(n117) );
  FA_X1 U185 ( .A(n115), .B(n114), .CI(n113), .CO(n197), .S(n200) );
  XNOR2_X1 U186 ( .A(n12), .B(\mult_x_1/n283 ), .ZN(n116) );
  NOR2_X1 U187 ( .A1(n116), .A2(n17), .ZN(n196) );
  FA_X1 U188 ( .A(n119), .B(n22), .CI(n117), .CO(n140), .S(n195) );
  OR2_X1 U189 ( .A1(n160), .A2(n159), .ZN(n120) );
  MUX2_X1 U190 ( .A(n354), .B(n120), .S(n312), .Z(n372) );
  XNOR2_X1 U191 ( .A(n349), .B(\mult_x_1/n283 ), .ZN(n227) );
  OAI22_X1 U192 ( .A1(n251), .A2(n227), .B1(n121), .B2(n5), .ZN(n138) );
  AND2_X1 U193 ( .A1(\mult_x_1/n288 ), .A2(n39), .ZN(n137) );
  XNOR2_X1 U194 ( .A(n350), .B(\mult_x_1/n285 ), .ZN(n226) );
  OAI22_X1 U195 ( .A1(n123), .A2(n226), .B1(n245), .B2(n122), .ZN(n136) );
  HA_X1 U196 ( .A(n125), .B(n124), .CO(n70), .S(n186) );
  FA_X1 U197 ( .A(n128), .B(n127), .CI(n126), .CO(n183), .S(n185) );
  OR2_X1 U198 ( .A1(\mult_x_1/n288 ), .A2(n417), .ZN(n129) );
  OAI22_X1 U199 ( .A1(n135), .A2(n417), .B1(n129), .B2(n133), .ZN(n225) );
  XNOR2_X1 U200 ( .A(n130), .B(\mult_x_1/n287 ), .ZN(n134) );
  XNOR2_X1 U201 ( .A(n130), .B(\mult_x_1/n288 ), .ZN(n131) );
  OAI22_X1 U202 ( .A1(n20), .A2(n134), .B1(n131), .B2(n135), .ZN(n224) );
  AND2_X1 U203 ( .A1(n225), .A2(n224), .ZN(n223) );
  OAI22_X1 U204 ( .A1(n135), .A2(n134), .B1(n19), .B2(n132), .ZN(n222) );
  FA_X1 U205 ( .A(n138), .B(n137), .CI(n136), .CO(n187), .S(n221) );
  OR2_X1 U206 ( .A1(n193), .A2(n192), .ZN(n139) );
  MUX2_X1 U207 ( .A(n355), .B(n139), .S(n312), .Z(n374) );
  FA_X1 U208 ( .A(n142), .B(n141), .CI(n140), .CO(n155), .S(n160) );
  AOI21_X1 U209 ( .B1(n145), .B2(n144), .A(n143), .ZN(n146) );
  INV_X1 U210 ( .A(n146), .ZN(n151) );
  XNOR2_X1 U211 ( .A(n147), .B(n9), .ZN(n149) );
  NOR2_X1 U212 ( .A1(n149), .A2(n17), .ZN(n150) );
  XOR2_X1 U213 ( .A(n151), .B(n150), .Z(n152) );
  XOR2_X1 U214 ( .A(n153), .B(n152), .Z(n154) );
  OR2_X1 U215 ( .A1(n155), .A2(n154), .ZN(n157) );
  NAND2_X1 U216 ( .A1(n155), .A2(n154), .ZN(n156) );
  NAND2_X1 U217 ( .A1(n157), .A2(n156), .ZN(n158) );
  MUX2_X1 U218 ( .A(n356), .B(n158), .S(n312), .Z(n376) );
  NAND2_X1 U219 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2_X1 U220 ( .A(n357), .B(n161), .S(n312), .Z(n378) );
  XNOR2_X1 U221 ( .A(n163), .B(n162), .ZN(n165) );
  XNOR2_X1 U222 ( .A(n164), .B(n165), .ZN(n269) );
  OAI21_X1 U223 ( .B1(n167), .B2(n168), .A(n166), .ZN(n170) );
  FA_X1 U224 ( .A(n173), .B(n172), .CI(n171), .CO(n89), .S(n209) );
  NOR2_X1 U225 ( .A1(n269), .A2(n270), .ZN(n178) );
  MUX2_X1 U226 ( .A(n358), .B(n178), .S(n312), .Z(n380) );
  NOR2_X1 U227 ( .A1(n180), .A2(n179), .ZN(n181) );
  MUX2_X1 U228 ( .A(n359), .B(n181), .S(n312), .Z(n382) );
  FA_X1 U229 ( .A(n184), .B(n183), .CI(n182), .CO(n179), .S(n190) );
  FA_X1 U230 ( .A(n187), .B(n186), .CI(n185), .CO(n189), .S(n193) );
  NOR2_X1 U231 ( .A1(n190), .A2(n189), .ZN(n188) );
  MUX2_X1 U232 ( .A(n361), .B(n188), .S(n312), .Z(n386) );
  NAND2_X1 U233 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U234 ( .A(n362), .B(n191), .S(n312), .Z(n388) );
  NAND2_X1 U235 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U236 ( .A(n363), .B(n194), .S(n312), .Z(n390) );
  FA_X1 U237 ( .A(n197), .B(n196), .CI(n195), .CO(n159), .S(n219) );
  NAND2_X1 U238 ( .A1(n198), .A2(n200), .ZN(n203) );
  NAND2_X1 U239 ( .A1(n198), .A2(n199), .ZN(n202) );
  NAND2_X1 U240 ( .A1(n200), .A2(n199), .ZN(n201) );
  NAND3_X1 U241 ( .A1(n203), .A2(n202), .A3(n201), .ZN(n218) );
  NAND2_X1 U242 ( .A1(n219), .A2(n218), .ZN(n204) );
  MUX2_X1 U243 ( .A(n364), .B(n204), .S(n312), .Z(n392) );
  NAND2_X1 U244 ( .A1(n206), .A2(n205), .ZN(n207) );
  MUX2_X1 U245 ( .A(n365), .B(n207), .S(n312), .Z(n394) );
  FA_X1 U246 ( .A(n210), .B(n209), .CI(n208), .CO(n270), .S(n216) );
  FA_X1 U247 ( .A(n213), .B(n212), .CI(n211), .CO(n215), .S(n180) );
  NOR2_X1 U248 ( .A1(n216), .A2(n215), .ZN(n214) );
  MUX2_X1 U249 ( .A(n366), .B(n214), .S(n312), .Z(n396) );
  NAND2_X1 U250 ( .A1(n216), .A2(n215), .ZN(n217) );
  MUX2_X1 U251 ( .A(n367), .B(n217), .S(n312), .Z(n398) );
  OR2_X1 U252 ( .A1(n219), .A2(n218), .ZN(n220) );
  MUX2_X1 U253 ( .A(n368), .B(n220), .S(n312), .Z(n400) );
  XOR2_X1 U254 ( .A(n225), .B(n224), .Z(n233) );
  XNOR2_X1 U255 ( .A(n350), .B(\mult_x_1/n286 ), .ZN(n236) );
  OAI22_X1 U256 ( .A1(n15), .A2(n236), .B1(n27), .B2(n226), .ZN(n231) );
  XNOR2_X1 U257 ( .A(n349), .B(\mult_x_1/n284 ), .ZN(n234) );
  OAI22_X1 U258 ( .A1(n251), .A2(n234), .B1(n227), .B2(n5), .ZN(n230) );
  OR2_X1 U259 ( .A1(n266), .A2(n265), .ZN(n277) );
  INV_X1 U260 ( .A(n277), .ZN(n267) );
  XNOR2_X1 U261 ( .A(n231), .B(n230), .ZN(n232) );
  XNOR2_X1 U262 ( .A(n233), .B(n232), .ZN(n263) );
  XNOR2_X1 U263 ( .A(n349), .B(\mult_x_1/n285 ), .ZN(n242) );
  OAI22_X1 U264 ( .A1(n251), .A2(n242), .B1(n234), .B2(n5), .ZN(n239) );
  AND2_X1 U265 ( .A1(\mult_x_1/n288 ), .A2(n235), .ZN(n238) );
  XNOR2_X1 U266 ( .A(n350), .B(\mult_x_1/n287 ), .ZN(n240) );
  OAI22_X1 U267 ( .A1(n15), .A2(n240), .B1(n27), .B2(n236), .ZN(n237) );
  OR2_X1 U268 ( .A1(n263), .A2(n262), .ZN(n306) );
  FA_X1 U269 ( .A(n239), .B(n238), .CI(n237), .CO(n262), .S(n261) );
  XNOR2_X1 U270 ( .A(n350), .B(\mult_x_1/n288 ), .ZN(n241) );
  OAI22_X1 U271 ( .A1(n247), .A2(n241), .B1(n27), .B2(n240), .ZN(n244) );
  XNOR2_X1 U272 ( .A(n349), .B(\mult_x_1/n286 ), .ZN(n248) );
  OAI22_X1 U273 ( .A1(n251), .A2(n248), .B1(n242), .B2(n5), .ZN(n243) );
  NOR2_X1 U274 ( .A1(n261), .A2(n260), .ZN(n299) );
  HA_X1 U275 ( .A(n244), .B(n243), .CO(n260), .S(n255) );
  OR2_X1 U276 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n246) );
  OAI22_X1 U277 ( .A1(n15), .A2(n28), .B1(n246), .B2(n27), .ZN(n256) );
  NAND2_X1 U278 ( .A1(n255), .A2(n256), .ZN(n294) );
  INV_X1 U279 ( .A(n294), .ZN(n259) );
  XNOR2_X1 U280 ( .A(n349), .B(\mult_x_1/n287 ), .ZN(n250) );
  OAI22_X1 U281 ( .A1(n251), .A2(n250), .B1(n248), .B2(n5), .ZN(n254) );
  AND2_X1 U282 ( .A1(\mult_x_1/n288 ), .A2(n249), .ZN(n253) );
  NOR2_X1 U283 ( .A1(n254), .A2(n253), .ZN(n288) );
  OAI22_X1 U284 ( .A1(n251), .A2(\mult_x_1/n288 ), .B1(n250), .B2(n5), .ZN(
        n285) );
  OR2_X1 U285 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n252) );
  NAND2_X1 U286 ( .A1(n252), .A2(n251), .ZN(n284) );
  NAND2_X1 U287 ( .A1(n285), .A2(n284), .ZN(n291) );
  NAND2_X1 U288 ( .A1(n254), .A2(n253), .ZN(n289) );
  OAI21_X1 U289 ( .B1(n288), .B2(n291), .A(n289), .ZN(n296) );
  INV_X1 U290 ( .A(n255), .ZN(n258) );
  INV_X1 U291 ( .A(n256), .ZN(n257) );
  NAND2_X1 U292 ( .A1(n258), .A2(n257), .ZN(n295) );
  OAI21_X1 U293 ( .B1(n259), .B2(n296), .A(n295), .ZN(n302) );
  NAND2_X1 U294 ( .A1(n261), .A2(n260), .ZN(n300) );
  OAI21_X1 U295 ( .B1(n302), .B2(n299), .A(n300), .ZN(n307) );
  NAND2_X1 U296 ( .A1(n263), .A2(n262), .ZN(n305) );
  INV_X1 U297 ( .A(n305), .ZN(n264) );
  AOI21_X1 U298 ( .B1(n306), .B2(n307), .A(n264), .ZN(n279) );
  NAND2_X1 U299 ( .A1(n266), .A2(n265), .ZN(n276) );
  OAI21_X1 U300 ( .B1(n267), .B2(n23), .A(n276), .ZN(n268) );
  MUX2_X1 U301 ( .A(n371), .B(n268), .S(n312), .Z(n406) );
  NAND2_X1 U302 ( .A1(n269), .A2(n270), .ZN(n271) );
  NAND2_X1 U303 ( .A1(n271), .A2(n312), .ZN(n273) );
  OR2_X1 U304 ( .A1(n312), .A2(n409), .ZN(n272) );
  NAND2_X1 U305 ( .A1(n273), .A2(n272), .ZN(n402) );
  BUF_X1 U306 ( .A(rst_n), .Z(n274) );
  NAND2_X1 U307 ( .A1(n352), .A2(A_extended[5]), .ZN(n275) );
  OAI21_X1 U308 ( .B1(n352), .B2(n417), .A(n275), .ZN(n526) );
  AND2_X1 U309 ( .A1(n277), .A2(n276), .ZN(n278) );
  XNOR2_X1 U310 ( .A(n279), .B(n278), .ZN(n280) );
  NAND2_X1 U311 ( .A1(n280), .A2(n312), .ZN(n282) );
  NAND2_X1 U312 ( .A1(n553), .A2(n72), .ZN(n281) );
  NAND2_X1 U313 ( .A1(n282), .A2(n281), .ZN(n462) );
  MUX2_X1 U314 ( .A(product[0]), .B(n534), .S(n312), .Z(n422) );
  MUX2_X1 U315 ( .A(n534), .B(n535), .S(n312), .Z(n424) );
  AND2_X1 U316 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n283) );
  MUX2_X1 U317 ( .A(n535), .B(n283), .S(n312), .Z(n426) );
  MUX2_X1 U318 ( .A(product[1]), .B(n537), .S(n312), .Z(n428) );
  MUX2_X1 U319 ( .A(n537), .B(n538), .S(n312), .Z(n430) );
  OR2_X1 U320 ( .A1(n285), .A2(n284), .ZN(n286) );
  AND2_X1 U321 ( .A1(n286), .A2(n291), .ZN(n287) );
  MUX2_X1 U322 ( .A(n538), .B(n287), .S(n312), .Z(n432) );
  MUX2_X1 U323 ( .A(product[2]), .B(n540), .S(n312), .Z(n434) );
  MUX2_X1 U324 ( .A(n540), .B(n541), .S(n312), .Z(n436) );
  INV_X1 U325 ( .A(n288), .ZN(n290) );
  NAND2_X1 U326 ( .A1(n290), .A2(n289), .ZN(n292) );
  XOR2_X1 U327 ( .A(n292), .B(n291), .Z(n293) );
  MUX2_X1 U328 ( .A(n541), .B(n293), .S(n312), .Z(n438) );
  MUX2_X1 U329 ( .A(product[3]), .B(n543), .S(n312), .Z(n440) );
  MUX2_X1 U330 ( .A(n543), .B(n544), .S(n312), .Z(n442) );
  NAND2_X1 U331 ( .A1(n295), .A2(n294), .ZN(n297) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n298) );
  MUX2_X1 U333 ( .A(n544), .B(n298), .S(n312), .Z(n444) );
  MUX2_X1 U334 ( .A(product[4]), .B(n546), .S(n312), .Z(n446) );
  MUX2_X1 U335 ( .A(n546), .B(n547), .S(n312), .Z(n448) );
  INV_X1 U336 ( .A(n299), .ZN(n301) );
  NAND2_X1 U337 ( .A1(n301), .A2(n300), .ZN(n303) );
  XOR2_X1 U338 ( .A(n303), .B(n7), .Z(n304) );
  MUX2_X1 U339 ( .A(n547), .B(n304), .S(n312), .Z(n450) );
  MUX2_X1 U340 ( .A(product[5]), .B(n549), .S(n312), .Z(n452) );
  MUX2_X1 U341 ( .A(n549), .B(n550), .S(n312), .Z(n454) );
  NAND2_X1 U342 ( .A1(n306), .A2(n305), .ZN(n308) );
  XNOR2_X1 U343 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U344 ( .A(n550), .B(n309), .S(n312), .Z(n456) );
  MUX2_X1 U345 ( .A(product[6]), .B(n552), .S(n312), .Z(n458) );
  MUX2_X1 U346 ( .A(n552), .B(n553), .S(n312), .Z(n460) );
  MUX2_X1 U347 ( .A(product[7]), .B(n555), .S(n312), .Z(n464) );
  NAND2_X1 U348 ( .A1(n355), .A2(n363), .ZN(n310) );
  XNOR2_X1 U349 ( .A(n371), .B(n310), .ZN(n311) );
  MUX2_X1 U350 ( .A(n555), .B(n311), .S(n312), .Z(n466) );
  MUX2_X1 U351 ( .A(product[8]), .B(n557), .S(n312), .Z(n468) );
  AOI21_X1 U352 ( .B1(n371), .B2(n355), .A(n413), .ZN(n315) );
  NAND2_X1 U353 ( .A1(n414), .A2(n362), .ZN(n313) );
  XOR2_X1 U354 ( .A(n315), .B(n313), .Z(n314) );
  MUX2_X1 U355 ( .A(n557), .B(n314), .S(n352), .Z(n470) );
  MUX2_X1 U356 ( .A(product[9]), .B(n559), .S(n352), .Z(n472) );
  OAI21_X1 U357 ( .B1(n315), .B2(n361), .A(n362), .ZN(n323) );
  INV_X1 U358 ( .A(n323), .ZN(n318) );
  NAND2_X1 U359 ( .A1(n415), .A2(n360), .ZN(n316) );
  XOR2_X1 U360 ( .A(n318), .B(n316), .Z(n317) );
  MUX2_X1 U361 ( .A(n559), .B(n317), .S(n352), .Z(n474) );
  MUX2_X1 U362 ( .A(product[10]), .B(n561), .S(n352), .Z(n476) );
  OAI21_X1 U363 ( .B1(n318), .B2(n359), .A(n360), .ZN(n320) );
  NAND2_X1 U364 ( .A1(n411), .A2(n367), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U366 ( .A(n561), .B(n321), .S(n352), .Z(n478) );
  MUX2_X1 U367 ( .A(product[11]), .B(n563), .S(n352), .Z(n480) );
  NOR2_X1 U368 ( .A1(n366), .A2(n359), .ZN(n324) );
  OAI21_X1 U369 ( .B1(n366), .B2(n360), .A(n367), .ZN(n322) );
  AOI21_X1 U370 ( .B1(n324), .B2(n323), .A(n322), .ZN(n346) );
  NAND2_X1 U371 ( .A1(n410), .A2(n369), .ZN(n325) );
  XOR2_X1 U372 ( .A(n346), .B(n325), .Z(n326) );
  MUX2_X1 U373 ( .A(n563), .B(n326), .S(n352), .Z(n482) );
  MUX2_X1 U374 ( .A(product[12]), .B(n565), .S(n352), .Z(n484) );
  OAI21_X1 U375 ( .B1(n346), .B2(n358), .A(n369), .ZN(n328) );
  NAND2_X1 U376 ( .A1(n370), .A2(n365), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  MUX2_X1 U378 ( .A(n565), .B(n329), .S(n352), .Z(n486) );
  MUX2_X1 U379 ( .A(product[13]), .B(n567), .S(n352), .Z(n488) );
  NAND2_X1 U380 ( .A1(n410), .A2(n370), .ZN(n331) );
  AOI21_X1 U381 ( .B1(n409), .B2(n370), .A(n416), .ZN(n330) );
  OAI21_X1 U382 ( .B1(n346), .B2(n331), .A(n330), .ZN(n333) );
  NAND2_X1 U383 ( .A1(n368), .A2(n364), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  MUX2_X1 U385 ( .A(n567), .B(n334), .S(n352), .Z(n490) );
  MUX2_X1 U386 ( .A(product[14]), .B(n569), .S(n352), .Z(n492) );
  NAND2_X1 U387 ( .A1(n370), .A2(n368), .ZN(n336) );
  NOR2_X1 U388 ( .A1(n358), .A2(n336), .ZN(n342) );
  INV_X1 U389 ( .A(n342), .ZN(n338) );
  AOI21_X1 U390 ( .B1(n416), .B2(n368), .A(n408), .ZN(n335) );
  OAI21_X1 U391 ( .B1(n336), .B2(n369), .A(n335), .ZN(n343) );
  INV_X1 U392 ( .A(n343), .ZN(n337) );
  OAI21_X1 U393 ( .B1(n346), .B2(n338), .A(n337), .ZN(n340) );
  NAND2_X1 U394 ( .A1(n354), .A2(n357), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  MUX2_X1 U396 ( .A(n569), .B(n341), .S(n352), .Z(n494) );
  MUX2_X1 U397 ( .A(product[15]), .B(n571), .S(n352), .Z(n496) );
  NAND2_X1 U398 ( .A1(n342), .A2(n354), .ZN(n345) );
  AOI21_X1 U399 ( .B1(n343), .B2(n354), .A(n412), .ZN(n344) );
  OAI21_X1 U400 ( .B1(n346), .B2(n345), .A(n344), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n347), .B(n356), .ZN(n348) );
  MUX2_X1 U402 ( .A(n571), .B(n348), .S(n352), .Z(n498) );
  MUX2_X1 U403 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n352), .Z(n500) );
  MUX2_X1 U404 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n352), .Z(n502) );
  MUX2_X1 U405 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n352), .Z(n504) );
  MUX2_X1 U406 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n352), .Z(n506) );
  MUX2_X1 U407 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n352), .Z(n508) );
  MUX2_X1 U408 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n352), .Z(n510) );
  MUX2_X1 U409 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n352), .Z(n512) );
  MUX2_X1 U410 ( .A(n9), .B(B_extended[7]), .S(n352), .Z(n514) );
  MUX2_X1 U411 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n352), .Z(n516) );
  MUX2_X1 U412 ( .A(n349), .B(A_extended[1]), .S(n352), .Z(n518) );
  MUX2_X1 U413 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n352), .Z(n520) );
  MUX2_X1 U414 ( .A(n350), .B(A_extended[3]), .S(n352), .Z(n522) );
  MUX2_X1 U415 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n352), .Z(n524) );
  MUX2_X1 U416 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n352), .Z(n528) );
  MUX2_X1 U417 ( .A(n351), .B(A_extended[7]), .S(n352), .Z(n530) );
  OR2_X1 U418 ( .A1(n352), .A2(n573), .ZN(n532) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_10 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n385, n387, n389, n391, n393, n395, n397, n399, n401,
         n403, n405, n407, n409, n411, n413, n415, n417, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n433,
         n435, n437, n439, n441, n443, n445, n447, n449, n451, n453, n455,
         n457, n459, n461, n463, n465, n467, n469, n471, n473, n475, n477,
         n479, n481, n483, n485, n487, n489, n491, n493, n495, n497, n499,
         n501, n503, n505, n507, n509, n511, n513, n515, n517, n519, n521,
         n523, n525, n527, n529, n531, n533, n535, n537, n539, n541, n543,
         n545, n546, n548, n549, n551, n552, n554, n555, n557, n558, n560,
         n561, n563, n564, n566, n568, n570, n572, n574, n576, n578, n580,
         n582, n583, n584, n585;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n430), .SE(n543), .CK(clk), .Q(n584), 
        .QN(n427) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n431), .SE(n539), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n431), .SE(n537), .CK(clk), .Q(n583), 
        .QN(n28) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n431), .SE(n535), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n26) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n431), .SE(n533), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n27) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n431), .SE(n531), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n431), .SE(n527), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n17) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n431), .SE(n525), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n19) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n431), .SE(n523), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n23) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n431), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n430), .SE(n519), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n24) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n430), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n22) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n430), .SE(n515), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n21) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n430), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n20) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n430), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n18) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n430), .SE(n509), .CK(clk), .Q(n582)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n430), .SE(n507), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n430), .SE(n505), .CK(clk), .Q(n580)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n430), .SE(n503), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n430), .SE(n501), .CK(clk), .Q(n578)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n430), .SE(n499), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n431), .SE(n497), .CK(clk), .Q(n576)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n429), .SE(n495), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n429), .SE(n493), .CK(clk), .Q(n574)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n431), .SE(n491), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n429), .SE(n489), .CK(clk), .Q(n572)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n430), .SE(n487), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n430), .SE(n485), .CK(clk), .Q(n570)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n483), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n481), .CK(clk), .Q(n568)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n479), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n477), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n475), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(rst_n), .SE(n473), .CK(clk), .Q(n564), 
        .QN(n31) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n471), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n469), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n429), .SE(n467), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n430), .SE(n465), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n463), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(rst_n), .SE(n461), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(rst_n), .SE(n459), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(rst_n), .SE(n457), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(rst_n), .SE(n455), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n429), .SE(n453), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n429), .SE(n451), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n429), .SE(n449), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n429), .SE(n447), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n429), .SE(n445), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n429), .SE(n443), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n429), .SE(n441), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n429), .SE(n439), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n429), .SE(n437), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n429), .SE(n435), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n429), .SE(n433), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n431), .SE(n529), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n33) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n431), .SE(n541), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n428) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n585), .SE(n417), .CK(
        clk), .QN(n382) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n585), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n381), .QN(n420) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n585), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n380), .QN(n426) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n585), .SE(n411), .CK(
        clk), .Q(n34), .QN(n379) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n585), .SE(n409), .CK(
        clk), .Q(n425), .QN(n378) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n585), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n377), .QN(n422) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n585), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n376) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n585), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n375), .QN(n423) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n585), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n374), .QN(n30) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n585), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n373), .QN(n424) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n585), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n372), .QN(n421) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n585), .SE(n395), .CK(
        clk), .Q(n364), .QN(n371) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n585), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n370), .QN(n419) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n585), .SE(n391), .CK(
        clk), .QN(n369) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n585), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n368) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n585), .SE(n387), .CK(
        clk), .QN(n367) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n585), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n366) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n585), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n365) );
  BUF_X1 U2 ( .A(n51), .Z(n5) );
  XNOR2_X1 U3 ( .A(n583), .B(\mult_x_1/a[6] ), .ZN(n51) );
  XNOR2_X1 U4 ( .A(\mult_x_1/a[2] ), .B(n33), .ZN(n6) );
  INV_X1 U5 ( .A(n19), .ZN(n7) );
  INV_X1 U6 ( .A(n428), .ZN(n8) );
  NAND2_X2 U7 ( .A1(n150), .A2(n17), .ZN(n151) );
  NAND2_X1 U8 ( .A1(n112), .A2(n111), .ZN(n97) );
  INV_X1 U9 ( .A(n112), .ZN(n99) );
  CLKBUF_X1 U10 ( .A(n260), .Z(n9) );
  XNOR2_X1 U11 ( .A(n16), .B(n24), .ZN(n206) );
  NAND2_X1 U12 ( .A1(n225), .A2(n224), .ZN(n246) );
  NAND2_X1 U13 ( .A1(n219), .A2(n218), .ZN(n220) );
  XNOR2_X1 U14 ( .A(n16), .B(n20), .ZN(n38) );
  INV_X1 U15 ( .A(n223), .ZN(n219) );
  XNOR2_X1 U16 ( .A(n16), .B(n19), .ZN(n261) );
  XNOR2_X1 U17 ( .A(n16), .B(n21), .ZN(n74) );
  XNOR2_X1 U18 ( .A(n16), .B(n22), .ZN(n185) );
  NAND2_X1 U19 ( .A1(n173), .A2(n172), .ZN(n174) );
  XNOR2_X1 U20 ( .A(n133), .B(n132), .ZN(n161) );
  XNOR2_X1 U21 ( .A(n131), .B(n130), .ZN(n132) );
  XNOR2_X1 U22 ( .A(n239), .B(n238), .ZN(n120) );
  NAND2_X1 U23 ( .A1(n127), .A2(n126), .ZN(n128) );
  NAND2_X1 U24 ( .A1(n131), .A2(n130), .ZN(n126) );
  NAND2_X1 U25 ( .A1(n133), .A2(n125), .ZN(n127) );
  OR2_X1 U26 ( .A1(n131), .A2(n130), .ZN(n125) );
  XNOR2_X1 U27 ( .A(n16), .B(n23), .ZN(n197) );
  NAND2_X1 U28 ( .A1(n101), .A2(n100), .ZN(n235) );
  NAND2_X1 U29 ( .A1(n113), .A2(n97), .ZN(n101) );
  NAND2_X1 U30 ( .A1(n241), .A2(n240), .ZN(n277) );
  NAND2_X1 U31 ( .A1(n239), .A2(n238), .ZN(n240) );
  NAND2_X1 U32 ( .A1(n237), .A2(n236), .ZN(n241) );
  OR2_X1 U33 ( .A1(n239), .A2(n238), .ZN(n236) );
  XNOR2_X1 U34 ( .A(n16), .B(n25), .ZN(n207) );
  NAND2_X1 U35 ( .A1(n250), .A2(n249), .ZN(n283) );
  NAND2_X1 U36 ( .A1(n15), .A2(n247), .ZN(n249) );
  OAI21_X1 U37 ( .B1(n15), .B2(n247), .A(n246), .ZN(n250) );
  OR2_X1 U38 ( .A1(n129), .A2(n128), .ZN(n286) );
  NAND2_X1 U39 ( .A1(n129), .A2(n128), .ZN(n287) );
  OAI211_X1 U40 ( .C1(n167), .C2(n108), .A(n166), .B(n165), .ZN(n401) );
  CLKBUF_X1 U41 ( .A(n208), .Z(n10) );
  CLKBUF_X1 U42 ( .A(n115), .Z(n11) );
  BUF_X1 U43 ( .A(n115), .Z(n12) );
  XNOR2_X1 U44 ( .A(\mult_x_1/a[2] ), .B(n33), .ZN(n42) );
  NAND2_X1 U45 ( .A1(n99), .A2(n98), .ZN(n100) );
  XNOR2_X1 U46 ( .A(n428), .B(n21), .ZN(n52) );
  OAI22_X1 U47 ( .A1(n178), .A2(n78), .B1(n177), .B2(n179), .ZN(n13) );
  INV_X1 U48 ( .A(n135), .ZN(n14) );
  INV_X1 U49 ( .A(n135), .ZN(n201) );
  INV_X1 U50 ( .A(n192), .ZN(n85) );
  BUF_X2 U51 ( .A(\mult_x_1/n312 ), .Z(n93) );
  FA_X1 U52 ( .A(n214), .B(n213), .CI(n212), .S(n15) );
  OR2_X2 U53 ( .A1(n72), .A2(n73), .ZN(n173) );
  OR2_X1 U54 ( .A1(n427), .A2(n428), .ZN(n16) );
  OR2_X1 U55 ( .A1(n427), .A2(n428), .ZN(n259) );
  XNOR2_X1 U56 ( .A(n237), .B(n120), .ZN(n129) );
  NAND2_X1 U57 ( .A1(n223), .A2(n222), .ZN(n224) );
  XNOR2_X1 U58 ( .A(n223), .B(n222), .ZN(n186) );
  INV_X1 U59 ( .A(n222), .ZN(n218) );
  BUF_X1 U60 ( .A(rst_n), .Z(n431) );
  BUF_X1 U61 ( .A(rst_n), .Z(n430) );
  BUF_X1 U62 ( .A(rst_n), .Z(n429) );
  INV_X1 U63 ( .A(rst_n), .ZN(n585) );
  BUF_X2 U64 ( .A(n583), .Z(n362) );
  AND3_X1 U65 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n29) );
  INV_X1 U66 ( .A(\mult_x_1/n310 ), .ZN(n44) );
  OR2_X1 U67 ( .A1(n325), .A2(n31), .ZN(n32) );
  BUF_X1 U68 ( .A(\mult_x_1/n313 ), .Z(n150) );
  AND2_X1 U69 ( .A1(n584), .A2(\mult_x_1/n281 ), .ZN(n199) );
  XNOR2_X1 U70 ( .A(n199), .B(n150), .ZN(n54) );
  AOI21_X1 U71 ( .B1(n151), .B2(n17), .A(n54), .ZN(n35) );
  INV_X1 U72 ( .A(n35), .ZN(n71) );
  XNOR2_X1 U73 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n76) );
  XNOR2_X1 U74 ( .A(n44), .B(\mult_x_1/a[6] ), .ZN(n36) );
  NAND2_X2 U75 ( .A1(n36), .A2(n51), .ZN(n257) );
  OAI22_X1 U76 ( .A1(n5), .A2(n76), .B1(n52), .B2(n257), .ZN(n70) );
  INV_X1 U77 ( .A(\mult_x_1/n310 ), .ZN(n37) );
  XNOR2_X2 U78 ( .A(n259), .B(n37), .ZN(n260) );
  NOR2_X1 U79 ( .A1(n38), .A2(n260), .ZN(n69) );
  XNOR2_X1 U80 ( .A(n583), .B(n26), .ZN(n39) );
  XNOR2_X1 U81 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n40) );
  NAND2_X1 U82 ( .A1(n39), .A2(n40), .ZN(n115) );
  XNOR2_X1 U83 ( .A(n362), .B(\mult_x_1/n285 ), .ZN(n61) );
  INV_X1 U84 ( .A(n40), .ZN(n135) );
  XNOR2_X1 U85 ( .A(n362), .B(\mult_x_1/n284 ), .ZN(n48) );
  OAI22_X1 U86 ( .A1(n12), .A2(n61), .B1(n14), .B2(n48), .ZN(n57) );
  XNOR2_X1 U87 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n41) );
  OR2_X2 U88 ( .A1(n41), .A2(n42), .ZN(n178) );
  XNOR2_X1 U89 ( .A(n93), .B(\mult_x_1/n283 ), .ZN(n63) );
  INV_X2 U90 ( .A(n6), .ZN(n179) );
  XNOR2_X1 U91 ( .A(n93), .B(\mult_x_1/n282 ), .ZN(n49) );
  OAI22_X1 U92 ( .A1(n178), .A2(n63), .B1(n179), .B2(n49), .ZN(n56) );
  OR2_X1 U93 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n43) );
  OAI22_X1 U94 ( .A1(n257), .A2(n37), .B1(n43), .B2(n5), .ZN(n103) );
  XNOR2_X1 U95 ( .A(n8), .B(\mult_x_1/n288 ), .ZN(n45) );
  OR2_X1 U96 ( .A1(n257), .A2(n45), .ZN(n47) );
  XNOR2_X1 U97 ( .A(n8), .B(\mult_x_1/n287 ), .ZN(n53) );
  OR2_X1 U98 ( .A1(n5), .A2(n53), .ZN(n46) );
  NAND2_X1 U99 ( .A1(n47), .A2(n46), .ZN(n102) );
  XNOR2_X1 U100 ( .A(n362), .B(\mult_x_1/n283 ), .ZN(n77) );
  OAI22_X1 U101 ( .A1(n11), .A2(n48), .B1(n201), .B2(n77), .ZN(n73) );
  XNOR2_X1 U102 ( .A(n93), .B(\mult_x_1/n281 ), .ZN(n78) );
  OAI22_X1 U103 ( .A1(n178), .A2(n49), .B1(n78), .B2(n179), .ZN(n72) );
  XNOR2_X1 U104 ( .A(n73), .B(n72), .ZN(n81) );
  OR2_X1 U105 ( .A1(\mult_x_1/n288 ), .A2(n16), .ZN(n50) );
  NOR2_X1 U106 ( .A1(n50), .A2(n260), .ZN(n80) );
  OAI22_X1 U107 ( .A1(n257), .A2(n53), .B1(n5), .B2(n52), .ZN(n60) );
  CLKBUF_X1 U108 ( .A(\mult_x_1/n313 ), .Z(n146) );
  XNOR2_X1 U109 ( .A(n146), .B(\mult_x_1/n281 ), .ZN(n62) );
  OAI22_X1 U110 ( .A1(n151), .A2(n62), .B1(n54), .B2(n17), .ZN(n59) );
  NOR2_X1 U111 ( .A1(n18), .A2(n260), .ZN(n58) );
  FA_X1 U112 ( .A(n57), .B(n56), .CI(n55), .CO(n83), .S(n92) );
  FA_X1 U113 ( .A(n58), .B(n59), .CI(n60), .CO(n79), .S(n90) );
  NAND2_X1 U114 ( .A1(n92), .A2(n90), .ZN(n66) );
  XNOR2_X1 U115 ( .A(n362), .B(\mult_x_1/n286 ), .ZN(n118) );
  OAI22_X1 U116 ( .A1(n12), .A2(n118), .B1(n14), .B2(n61), .ZN(n106) );
  XNOR2_X1 U117 ( .A(n150), .B(\mult_x_1/n282 ), .ZN(n96) );
  OAI22_X1 U118 ( .A1(n151), .A2(n96), .B1(n62), .B2(n17), .ZN(n105) );
  XNOR2_X1 U119 ( .A(n93), .B(\mult_x_1/n284 ), .ZN(n94) );
  OAI22_X1 U120 ( .A1(n178), .A2(n94), .B1(n179), .B2(n63), .ZN(n104) );
  NAND2_X1 U121 ( .A1(n92), .A2(n89), .ZN(n65) );
  NAND2_X1 U122 ( .A1(n90), .A2(n89), .ZN(n64) );
  BUF_X4 U123 ( .A(en), .Z(n325) );
  NAND2_X1 U124 ( .A1(n29), .A2(n363), .ZN(n68) );
  NAND2_X1 U125 ( .A1(n108), .A2(n373), .ZN(n67) );
  OAI21_X1 U126 ( .B1(n167), .B2(n68), .A(n67), .ZN(n399) );
  FA_X1 U127 ( .A(n71), .B(n70), .CI(n69), .CO(n171), .S(n84) );
  NOR2_X1 U128 ( .A1(n74), .A2(n260), .ZN(n172) );
  XNOR2_X1 U129 ( .A(n173), .B(n172), .ZN(n75) );
  XNOR2_X1 U130 ( .A(n75), .B(n171), .ZN(n189) );
  XNOR2_X1 U131 ( .A(n8), .B(\mult_x_1/n284 ), .ZN(n176) );
  OAI22_X1 U132 ( .A1(n5), .A2(n176), .B1(n76), .B2(n257), .ZN(n183) );
  XNOR2_X1 U133 ( .A(n362), .B(\mult_x_1/n282 ), .ZN(n184) );
  OAI22_X1 U134 ( .A1(n12), .A2(n77), .B1(n14), .B2(n184), .ZN(n182) );
  XNOR2_X1 U135 ( .A(n199), .B(n93), .ZN(n177) );
  OAI22_X1 U136 ( .A1(n178), .A2(n78), .B1(n177), .B2(n179), .ZN(n216) );
  INV_X1 U137 ( .A(n216), .ZN(n181) );
  FA_X1 U138 ( .A(n81), .B(n80), .CI(n79), .CO(n187), .S(n82) );
  INV_X1 U139 ( .A(n193), .ZN(n86) );
  FA_X1 U140 ( .A(n84), .B(n83), .CI(n82), .CO(n192), .S(n167) );
  NAND3_X1 U141 ( .A1(n86), .A2(n85), .A3(n363), .ZN(n88) );
  NAND2_X1 U142 ( .A1(n108), .A2(n378), .ZN(n87) );
  NAND2_X1 U143 ( .A1(n88), .A2(n87), .ZN(n409) );
  XOR2_X1 U144 ( .A(n90), .B(n89), .Z(n91) );
  XOR2_X1 U145 ( .A(n92), .B(n91), .Z(n275) );
  XNOR2_X1 U146 ( .A(n93), .B(\mult_x_1/n285 ), .ZN(n123) );
  OAI22_X1 U147 ( .A1(n178), .A2(n123), .B1(n179), .B2(n94), .ZN(n113) );
  INV_X1 U148 ( .A(n5), .ZN(n95) );
  NAND2_X1 U149 ( .A1(n95), .A2(\mult_x_1/n288 ), .ZN(n112) );
  XNOR2_X1 U150 ( .A(n146), .B(\mult_x_1/n283 ), .ZN(n124) );
  OAI22_X1 U151 ( .A1(n151), .A2(n124), .B1(n96), .B2(n17), .ZN(n98) );
  INV_X1 U152 ( .A(n98), .ZN(n111) );
  HA_X1 U153 ( .A(n103), .B(n102), .CO(n55), .S(n234) );
  FA_X1 U154 ( .A(n106), .B(n105), .CI(n104), .CO(n89), .S(n233) );
  NAND2_X1 U155 ( .A1(n275), .A2(n274), .ZN(n107) );
  NAND2_X1 U156 ( .A1(n107), .A2(n363), .ZN(n110) );
  INV_X1 U157 ( .A(n363), .ZN(n108) );
  NAND2_X1 U158 ( .A1(n108), .A2(n376), .ZN(n109) );
  NAND2_X1 U159 ( .A1(n110), .A2(n109), .ZN(n405) );
  XNOR2_X1 U160 ( .A(n112), .B(n111), .ZN(n114) );
  XNOR2_X1 U161 ( .A(n114), .B(n113), .ZN(n237) );
  OR2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n116) );
  OAI22_X1 U163 ( .A1(n12), .A2(n28), .B1(n116), .B2(n201), .ZN(n122) );
  XNOR2_X1 U164 ( .A(n362), .B(\mult_x_1/n288 ), .ZN(n117) );
  XNOR2_X1 U165 ( .A(n362), .B(\mult_x_1/n287 ), .ZN(n119) );
  OAI22_X1 U166 ( .A1(n12), .A2(n117), .B1(n201), .B2(n119), .ZN(n121) );
  OAI22_X1 U167 ( .A1(n12), .A2(n119), .B1(n14), .B2(n118), .ZN(n238) );
  HA_X1 U168 ( .A(n122), .B(n121), .CO(n239), .S(n133) );
  XNOR2_X1 U169 ( .A(n93), .B(\mult_x_1/n286 ), .ZN(n136) );
  OAI22_X1 U170 ( .A1(n178), .A2(n136), .B1(n179), .B2(n123), .ZN(n131) );
  XNOR2_X1 U171 ( .A(n150), .B(\mult_x_1/n284 ), .ZN(n134) );
  OAI22_X1 U172 ( .A1(n151), .A2(n134), .B1(n124), .B2(n17), .ZN(n130) );
  NAND2_X1 U173 ( .A1(n286), .A2(n287), .ZN(n163) );
  XNOR2_X1 U174 ( .A(n146), .B(\mult_x_1/n285 ), .ZN(n142) );
  OAI22_X1 U175 ( .A1(n151), .A2(n142), .B1(n134), .B2(n17), .ZN(n139) );
  AND2_X1 U176 ( .A1(\mult_x_1/n288 ), .A2(n135), .ZN(n138) );
  XNOR2_X1 U177 ( .A(n93), .B(\mult_x_1/n287 ), .ZN(n140) );
  OAI22_X1 U178 ( .A1(n178), .A2(n140), .B1(n179), .B2(n136), .ZN(n137) );
  OR2_X1 U179 ( .A1(n161), .A2(n160), .ZN(n319) );
  FA_X1 U180 ( .A(n139), .B(n138), .CI(n137), .CO(n160), .S(n159) );
  XNOR2_X1 U181 ( .A(n93), .B(\mult_x_1/n288 ), .ZN(n141) );
  OAI22_X1 U182 ( .A1(n178), .A2(n141), .B1(n179), .B2(n140), .ZN(n144) );
  XNOR2_X1 U183 ( .A(n150), .B(\mult_x_1/n286 ), .ZN(n147) );
  OAI22_X1 U184 ( .A1(n151), .A2(n147), .B1(n142), .B2(n17), .ZN(n143) );
  NOR2_X1 U185 ( .A1(n159), .A2(n158), .ZN(n312) );
  HA_X1 U186 ( .A(n144), .B(n143), .CO(n158), .S(n156) );
  OR2_X1 U187 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n145) );
  OAI22_X1 U188 ( .A1(n178), .A2(n27), .B1(n145), .B2(n179), .ZN(n155) );
  OR2_X1 U189 ( .A1(n156), .A2(n155), .ZN(n308) );
  XNOR2_X1 U190 ( .A(n146), .B(\mult_x_1/n287 ), .ZN(n149) );
  OAI22_X1 U191 ( .A1(n151), .A2(n149), .B1(n147), .B2(n17), .ZN(n154) );
  INV_X1 U192 ( .A(n179), .ZN(n148) );
  AND2_X1 U193 ( .A1(\mult_x_1/n288 ), .A2(n148), .ZN(n153) );
  NOR2_X1 U194 ( .A1(n154), .A2(n153), .ZN(n301) );
  OAI22_X1 U195 ( .A1(n151), .A2(\mult_x_1/n288 ), .B1(n149), .B2(n17), .ZN(
        n298) );
  OR2_X1 U196 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n152) );
  NAND2_X1 U197 ( .A1(n152), .A2(n151), .ZN(n297) );
  NAND2_X1 U198 ( .A1(n298), .A2(n297), .ZN(n304) );
  NAND2_X1 U199 ( .A1(n154), .A2(n153), .ZN(n302) );
  OAI21_X1 U200 ( .B1(n301), .B2(n304), .A(n302), .ZN(n309) );
  NAND2_X1 U201 ( .A1(n156), .A2(n155), .ZN(n307) );
  INV_X1 U202 ( .A(n307), .ZN(n157) );
  AOI21_X1 U203 ( .B1(n308), .B2(n309), .A(n157), .ZN(n315) );
  NAND2_X1 U204 ( .A1(n159), .A2(n158), .ZN(n313) );
  OAI21_X1 U205 ( .B1(n312), .B2(n315), .A(n313), .ZN(n320) );
  NAND2_X1 U206 ( .A1(n161), .A2(n160), .ZN(n318) );
  INV_X1 U207 ( .A(n318), .ZN(n162) );
  AOI21_X1 U208 ( .B1(n319), .B2(n320), .A(n162), .ZN(n288) );
  XNOR2_X1 U209 ( .A(n163), .B(n288), .ZN(n164) );
  OAI21_X1 U210 ( .B1(n164), .B2(n108), .A(n32), .ZN(n473) );
  OR2_X1 U211 ( .A1(n363), .A2(n30), .ZN(n166) );
  NAND2_X1 U212 ( .A1(n363), .A2(n29), .ZN(n165) );
  INV_X1 U213 ( .A(n173), .ZN(n169) );
  INV_X1 U214 ( .A(n172), .ZN(n168) );
  NAND2_X1 U215 ( .A1(n169), .A2(n168), .ZN(n170) );
  NAND2_X1 U216 ( .A1(n171), .A2(n170), .ZN(n175) );
  NAND2_X1 U217 ( .A1(n175), .A2(n174), .ZN(n229) );
  XNOR2_X1 U218 ( .A(n8), .B(\mult_x_1/n283 ), .ZN(n205) );
  OAI22_X1 U219 ( .A1(n257), .A2(n176), .B1(n5), .B2(n205), .ZN(n217) );
  AOI21_X1 U220 ( .B1(n179), .B2(n178), .A(n177), .ZN(n180) );
  INV_X1 U221 ( .A(n180), .ZN(n215) );
  FA_X1 U222 ( .A(n183), .B(n182), .CI(n181), .CO(n221), .S(n188) );
  XNOR2_X1 U223 ( .A(n362), .B(\mult_x_1/n281 ), .ZN(n203) );
  OAI22_X1 U224 ( .A1(n12), .A2(n184), .B1(n14), .B2(n203), .ZN(n223) );
  NOR2_X1 U225 ( .A1(n185), .A2(n260), .ZN(n222) );
  XNOR2_X1 U226 ( .A(n221), .B(n186), .ZN(n227) );
  FA_X1 U227 ( .A(n189), .B(n188), .CI(n187), .CO(n291), .S(n193) );
  INV_X1 U228 ( .A(n291), .ZN(n190) );
  NAND2_X1 U229 ( .A1(n190), .A2(n325), .ZN(n191) );
  OAI22_X1 U230 ( .A1(n292), .A2(n191), .B1(n325), .B2(n364), .ZN(n395) );
  NAND2_X1 U231 ( .A1(n193), .A2(n192), .ZN(n194) );
  NAND2_X1 U232 ( .A1(n194), .A2(n325), .ZN(n196) );
  OR2_X1 U233 ( .A1(n325), .A2(n34), .ZN(n195) );
  NAND2_X1 U234 ( .A1(n196), .A2(n195), .ZN(n411) );
  NOR2_X1 U253 ( .A1(n197), .A2(n9), .ZN(n255) );
  XNOR2_X1 U254 ( .A(\mult_x_1/n310 ), .B(n7), .ZN(n198) );
  XNOR2_X1 U255 ( .A(n199), .B(n8), .ZN(n256) );
  OAI22_X1 U256 ( .A1(n257), .A2(n198), .B1(n256), .B2(n5), .ZN(n265) );
  INV_X1 U257 ( .A(n265), .ZN(n254) );
  XNOR2_X1 U258 ( .A(n8), .B(\mult_x_1/n282 ), .ZN(n204) );
  OAI22_X1 U259 ( .A1(n257), .A2(n204), .B1(n5), .B2(n198), .ZN(n210) );
  XNOR2_X1 U260 ( .A(n199), .B(n362), .ZN(n202) );
  AOI21_X1 U261 ( .B1(n14), .B2(n11), .A(n202), .ZN(n200) );
  INV_X1 U262 ( .A(n200), .ZN(n209) );
  OAI22_X1 U263 ( .A1(n11), .A2(n203), .B1(n202), .B2(n201), .ZN(n208) );
  INV_X1 U264 ( .A(n208), .ZN(n214) );
  OAI22_X1 U265 ( .A1(n257), .A2(n205), .B1(n5), .B2(n204), .ZN(n213) );
  NOR2_X1 U266 ( .A1(n206), .A2(n260), .ZN(n212) );
  NOR2_X1 U267 ( .A1(n207), .A2(n9), .ZN(n244) );
  FA_X1 U268 ( .A(n210), .B(n209), .CI(n10), .CO(n253), .S(n243) );
  OR2_X1 U269 ( .A1(n272), .A2(n271), .ZN(n211) );
  MUX2_X1 U270 ( .A(n365), .B(n211), .S(n325), .Z(n383) );
  FA_X1 U271 ( .A(n214), .B(n213), .CI(n212), .CO(n245), .S(n248) );
  FA_X1 U272 ( .A(n217), .B(n13), .CI(n215), .CO(n247), .S(n228) );
  XNOR2_X1 U273 ( .A(n248), .B(n247), .ZN(n226) );
  NAND2_X1 U274 ( .A1(n221), .A2(n220), .ZN(n225) );
  XNOR2_X1 U275 ( .A(n226), .B(n246), .ZN(n281) );
  INV_X1 U276 ( .A(n281), .ZN(n231) );
  FA_X1 U277 ( .A(n229), .B(n228), .CI(n227), .CO(n280), .S(n292) );
  INV_X1 U278 ( .A(n280), .ZN(n230) );
  NAND2_X1 U279 ( .A1(n231), .A2(n230), .ZN(n232) );
  MUX2_X1 U280 ( .A(n366), .B(n232), .S(n325), .Z(n385) );
  FA_X1 U281 ( .A(n235), .B(n234), .CI(n233), .CO(n274), .S(n278) );
  OR2_X1 U282 ( .A1(n278), .A2(n277), .ZN(n242) );
  MUX2_X1 U283 ( .A(n367), .B(n242), .S(n325), .Z(n387) );
  FA_X1 U284 ( .A(n245), .B(n244), .CI(n243), .CO(n271), .S(n284) );
  OR2_X1 U285 ( .A1(n284), .A2(n283), .ZN(n252) );
  MUX2_X1 U286 ( .A(n368), .B(n252), .S(n325), .Z(n389) );
  FA_X1 U287 ( .A(n255), .B(n254), .CI(n253), .CO(n267), .S(n272) );
  AOI21_X1 U288 ( .B1(n5), .B2(n257), .A(n256), .ZN(n258) );
  INV_X1 U289 ( .A(n258), .ZN(n263) );
  NOR2_X1 U290 ( .A1(n261), .A2(n9), .ZN(n262) );
  XOR2_X1 U291 ( .A(n263), .B(n262), .Z(n264) );
  XOR2_X1 U292 ( .A(n265), .B(n264), .Z(n266) );
  OR2_X1 U293 ( .A1(n267), .A2(n266), .ZN(n269) );
  NAND2_X1 U294 ( .A1(n267), .A2(n266), .ZN(n268) );
  NAND2_X1 U295 ( .A1(n269), .A2(n268), .ZN(n270) );
  MUX2_X1 U296 ( .A(n369), .B(n270), .S(n363), .Z(n391) );
  NAND2_X1 U297 ( .A1(n272), .A2(n271), .ZN(n273) );
  MUX2_X1 U298 ( .A(n370), .B(n273), .S(n363), .Z(n393) );
  NOR2_X1 U299 ( .A1(n275), .A2(n274), .ZN(n276) );
  MUX2_X1 U300 ( .A(n375), .B(n276), .S(n363), .Z(n403) );
  NAND2_X1 U301 ( .A1(n278), .A2(n277), .ZN(n279) );
  MUX2_X1 U302 ( .A(n377), .B(n279), .S(n325), .Z(n407) );
  NAND2_X1 U303 ( .A1(n281), .A2(n280), .ZN(n282) );
  MUX2_X1 U304 ( .A(n380), .B(n282), .S(n325), .Z(n413) );
  NAND2_X1 U305 ( .A1(n284), .A2(n283), .ZN(n285) );
  MUX2_X1 U306 ( .A(n381), .B(n285), .S(n325), .Z(n415) );
  INV_X1 U307 ( .A(n286), .ZN(n289) );
  OAI21_X1 U308 ( .B1(n289), .B2(n288), .A(n287), .ZN(n290) );
  MUX2_X1 U309 ( .A(n382), .B(n290), .S(n363), .Z(n417) );
  NAND2_X1 U310 ( .A1(n292), .A2(n291), .ZN(n293) );
  NAND2_X1 U311 ( .A1(n293), .A2(n363), .ZN(n295) );
  OR2_X1 U312 ( .A1(n363), .A2(n421), .ZN(n294) );
  NAND2_X1 U313 ( .A1(n295), .A2(n294), .ZN(n397) );
  MUX2_X1 U314 ( .A(product[0]), .B(n545), .S(n325), .Z(n433) );
  MUX2_X1 U315 ( .A(n545), .B(n546), .S(n325), .Z(n435) );
  AND2_X1 U316 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n296) );
  MUX2_X1 U317 ( .A(n546), .B(n296), .S(n325), .Z(n437) );
  MUX2_X1 U318 ( .A(product[1]), .B(n548), .S(n325), .Z(n439) );
  MUX2_X1 U319 ( .A(n548), .B(n549), .S(n325), .Z(n441) );
  OR2_X1 U320 ( .A1(n298), .A2(n297), .ZN(n299) );
  AND2_X1 U321 ( .A1(n299), .A2(n304), .ZN(n300) );
  MUX2_X1 U322 ( .A(n549), .B(n300), .S(n325), .Z(n443) );
  MUX2_X1 U323 ( .A(product[2]), .B(n551), .S(n325), .Z(n445) );
  MUX2_X1 U324 ( .A(n551), .B(n552), .S(n325), .Z(n447) );
  INV_X1 U325 ( .A(n301), .ZN(n303) );
  NAND2_X1 U326 ( .A1(n303), .A2(n302), .ZN(n305) );
  XOR2_X1 U327 ( .A(n305), .B(n304), .Z(n306) );
  MUX2_X1 U328 ( .A(n552), .B(n306), .S(n325), .Z(n449) );
  MUX2_X1 U329 ( .A(product[3]), .B(n554), .S(n325), .Z(n451) );
  MUX2_X1 U330 ( .A(n554), .B(n555), .S(n325), .Z(n453) );
  NAND2_X1 U331 ( .A1(n308), .A2(n307), .ZN(n310) );
  XNOR2_X1 U332 ( .A(n310), .B(n309), .ZN(n311) );
  MUX2_X1 U333 ( .A(n555), .B(n311), .S(n325), .Z(n455) );
  MUX2_X1 U334 ( .A(product[4]), .B(n557), .S(n325), .Z(n457) );
  MUX2_X1 U335 ( .A(n557), .B(n558), .S(n325), .Z(n459) );
  INV_X1 U336 ( .A(n312), .ZN(n314) );
  NAND2_X1 U337 ( .A1(n314), .A2(n313), .ZN(n316) );
  XOR2_X1 U338 ( .A(n316), .B(n315), .Z(n317) );
  MUX2_X1 U339 ( .A(n558), .B(n317), .S(n325), .Z(n461) );
  MUX2_X1 U340 ( .A(product[5]), .B(n560), .S(n325), .Z(n463) );
  MUX2_X1 U341 ( .A(n560), .B(n561), .S(n325), .Z(n465) );
  NAND2_X1 U342 ( .A1(n319), .A2(n318), .ZN(n321) );
  XNOR2_X1 U343 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U344 ( .A(n561), .B(n322), .S(n325), .Z(n467) );
  MUX2_X1 U345 ( .A(product[6]), .B(n563), .S(n325), .Z(n469) );
  MUX2_X1 U346 ( .A(n563), .B(n564), .S(n325), .Z(n471) );
  MUX2_X1 U347 ( .A(product[7]), .B(n566), .S(n325), .Z(n475) );
  NAND2_X1 U348 ( .A1(n367), .A2(n377), .ZN(n323) );
  XNOR2_X1 U349 ( .A(n382), .B(n323), .ZN(n324) );
  MUX2_X1 U350 ( .A(n566), .B(n324), .S(n325), .Z(n477) );
  MUX2_X1 U351 ( .A(product[8]), .B(n568), .S(n325), .Z(n479) );
  AOI21_X1 U352 ( .B1(n382), .B2(n367), .A(n422), .ZN(n328) );
  NAND2_X1 U353 ( .A1(n423), .A2(n376), .ZN(n326) );
  XOR2_X1 U354 ( .A(n328), .B(n326), .Z(n327) );
  BUF_X4 U355 ( .A(en), .Z(n363) );
  MUX2_X1 U356 ( .A(n568), .B(n327), .S(n363), .Z(n481) );
  MUX2_X1 U357 ( .A(product[9]), .B(n570), .S(n363), .Z(n483) );
  OAI21_X1 U358 ( .B1(n328), .B2(n375), .A(n376), .ZN(n336) );
  INV_X1 U359 ( .A(n336), .ZN(n331) );
  NAND2_X1 U360 ( .A1(n424), .A2(n374), .ZN(n329) );
  XOR2_X1 U361 ( .A(n331), .B(n329), .Z(n330) );
  MUX2_X1 U362 ( .A(n570), .B(n330), .S(n363), .Z(n485) );
  MUX2_X1 U363 ( .A(product[10]), .B(n572), .S(n363), .Z(n487) );
  OAI21_X1 U364 ( .B1(n331), .B2(n373), .A(n374), .ZN(n333) );
  NAND2_X1 U365 ( .A1(n425), .A2(n379), .ZN(n332) );
  XNOR2_X1 U366 ( .A(n333), .B(n332), .ZN(n334) );
  MUX2_X1 U367 ( .A(n572), .B(n334), .S(n363), .Z(n489) );
  MUX2_X1 U368 ( .A(product[11]), .B(n574), .S(n363), .Z(n491) );
  NOR2_X1 U369 ( .A1(n378), .A2(n373), .ZN(n337) );
  OAI21_X1 U370 ( .B1(n378), .B2(n374), .A(n379), .ZN(n335) );
  AOI21_X1 U371 ( .B1(n337), .B2(n336), .A(n335), .ZN(n359) );
  NAND2_X1 U372 ( .A1(n364), .A2(n372), .ZN(n338) );
  XOR2_X1 U373 ( .A(n359), .B(n338), .Z(n339) );
  MUX2_X1 U374 ( .A(n574), .B(n339), .S(n363), .Z(n493) );
  MUX2_X1 U375 ( .A(product[12]), .B(n576), .S(n363), .Z(n495) );
  OAI21_X1 U376 ( .B1(n359), .B2(n371), .A(n372), .ZN(n341) );
  NAND2_X1 U377 ( .A1(n366), .A2(n380), .ZN(n340) );
  XNOR2_X1 U378 ( .A(n341), .B(n340), .ZN(n342) );
  MUX2_X1 U379 ( .A(n576), .B(n342), .S(n363), .Z(n497) );
  MUX2_X1 U380 ( .A(product[13]), .B(n578), .S(n363), .Z(n499) );
  NAND2_X1 U381 ( .A1(n364), .A2(n366), .ZN(n344) );
  AOI21_X1 U382 ( .B1(n421), .B2(n366), .A(n426), .ZN(n343) );
  OAI21_X1 U383 ( .B1(n359), .B2(n344), .A(n343), .ZN(n346) );
  NAND2_X1 U384 ( .A1(n368), .A2(n381), .ZN(n345) );
  XNOR2_X1 U385 ( .A(n346), .B(n345), .ZN(n347) );
  MUX2_X1 U386 ( .A(n578), .B(n347), .S(n363), .Z(n501) );
  MUX2_X1 U387 ( .A(product[14]), .B(n580), .S(n363), .Z(n503) );
  NAND2_X1 U388 ( .A1(n366), .A2(n368), .ZN(n349) );
  NOR2_X1 U389 ( .A1(n371), .A2(n349), .ZN(n355) );
  INV_X1 U390 ( .A(n355), .ZN(n351) );
  AOI21_X1 U391 ( .B1(n426), .B2(n368), .A(n420), .ZN(n348) );
  OAI21_X1 U392 ( .B1(n349), .B2(n372), .A(n348), .ZN(n356) );
  INV_X1 U393 ( .A(n356), .ZN(n350) );
  OAI21_X1 U394 ( .B1(n359), .B2(n351), .A(n350), .ZN(n353) );
  NAND2_X1 U395 ( .A1(n365), .A2(n370), .ZN(n352) );
  XNOR2_X1 U396 ( .A(n353), .B(n352), .ZN(n354) );
  MUX2_X1 U397 ( .A(n580), .B(n354), .S(n363), .Z(n505) );
  MUX2_X1 U398 ( .A(product[15]), .B(n582), .S(n363), .Z(n507) );
  NAND2_X1 U399 ( .A1(n355), .A2(n365), .ZN(n358) );
  AOI21_X1 U400 ( .B1(n356), .B2(n365), .A(n419), .ZN(n357) );
  OAI21_X1 U401 ( .B1(n359), .B2(n358), .A(n357), .ZN(n360) );
  XNOR2_X1 U402 ( .A(n360), .B(n369), .ZN(n361) );
  MUX2_X1 U403 ( .A(n582), .B(n361), .S(n363), .Z(n509) );
  MUX2_X1 U404 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n363), .Z(n511) );
  MUX2_X1 U405 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n363), .Z(n513) );
  MUX2_X1 U406 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n363), .Z(n515) );
  MUX2_X1 U407 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n363), .Z(n517) );
  MUX2_X1 U408 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n363), .Z(n519) );
  MUX2_X1 U409 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n363), .Z(n521) );
  MUX2_X1 U410 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n363), .Z(n523) );
  MUX2_X1 U411 ( .A(n7), .B(B_extended[7]), .S(n363), .Z(n525) );
  MUX2_X1 U412 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n363), .Z(n527) );
  MUX2_X1 U413 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n363), .Z(n529) );
  MUX2_X1 U414 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n363), .Z(n531) );
  MUX2_X1 U415 ( .A(n93), .B(A_extended[3]), .S(n363), .Z(n533) );
  MUX2_X1 U416 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n363), .Z(n535) );
  MUX2_X1 U417 ( .A(n362), .B(A_extended[5]), .S(n363), .Z(n537) );
  MUX2_X1 U418 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n363), .Z(n539) );
  MUX2_X1 U419 ( .A(n8), .B(A_extended[7]), .S(n363), .Z(n541) );
  OR2_X1 U420 ( .A1(n363), .A2(n584), .ZN(n543) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_11 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n364, n366, n368, n370, n372, n374, n376,
         n378, n380, n382, n384, n386, n388, n390, n392, n394, n396, n398,
         n400, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n505, n507, n509, n511, n513, n515, n517, n519,
         n521, n523, n525, n526, n528, n529, n531, n532, n534, n535, n537,
         n538, n540, n541, n543, n545, n547, n549, n551, n553, n555, n557,
         n559, n561, n562, n563, n564;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n413), .SE(n523), .CK(clk), .Q(n563), 
        .QN(n20) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n413), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n26) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n413), .SE(n517), .CK(clk), .Q(n562), 
        .QN(n25) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n413), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n27) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n413), .SE(n511), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n24) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n413), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n12) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n413), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n14) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n413), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n19) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n412), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n15) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n412), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n13) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n412), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n16) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n412), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n18) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n412), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n17) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n412), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n412), .SE(n489), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n412), .SE(n487), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n412), .SE(n485), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n412), .SE(n483), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n412), .SE(n481), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n413), .SE(n479), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n413), .SE(n477), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n412), .SE(n475), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n413), .SE(n473), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n412), .SE(n471), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n413), .SE(n469), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n412), .SE(n467), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n413), .SE(n465), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n413), .SE(n463), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n413), .SE(n461), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n412), .SE(n459), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n413), .SE(n457), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n412), .SE(n455), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n412), .SE(n453), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n413), .SE(n451), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n413), .SE(n449), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n413), .SE(n447), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n412), .SE(n445), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n413), .SE(n443), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n413), .SE(n441), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n413), .SE(n439), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n413), .SE(n437), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n413), .SE(n435), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n412), .SE(n433), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n413), .SE(n431), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n413), .SE(n429), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n412), .SE(n427), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n413), .SE(n425), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n413), .SE(n423), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n412), .SE(n421), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n413), .SE(n419), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n413), .SE(n417), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n412), .SE(n415), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n413), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n30) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n564), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n564), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n564), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n359), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n564), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n358), .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n564), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n357), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n564), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n356), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n564), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n355), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n564), .SE(n386), .CK(
        clk), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n564), .SE(n384), .CK(
        clk), .Q(n410), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n564), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n564), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n351), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n564), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n350), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n564), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n349), .QN(n29) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n564), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n348), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n564), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n564), .SE(n370), .CK(
        clk), .Q(n403), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n564), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n345), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n564), .SE(n366), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n564), .SE(n364), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n564), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n342) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n413), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n22) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n413), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n21) );
  BUF_X1 U2 ( .A(en), .Z(n341) );
  BUF_X2 U3 ( .A(n341), .Z(n8) );
  BUF_X2 U4 ( .A(n341), .Z(n9) );
  CLKBUF_X2 U5 ( .A(rst_n), .Z(n413) );
  INV_X1 U6 ( .A(n22), .ZN(n10) );
  BUF_X1 U7 ( .A(n562), .Z(n5) );
  NOR2_X1 U8 ( .A1(n13), .A2(n90), .ZN(n260) );
  NAND2_X1 U9 ( .A1(n51), .A2(n50), .ZN(n263) );
  NAND2_X1 U10 ( .A1(n175), .A2(n174), .ZN(n50) );
  OR2_X1 U11 ( .A1(n175), .A2(n174), .ZN(n49) );
  XNOR2_X1 U12 ( .A(n23), .B(n150), .ZN(n180) );
  NAND2_X1 U13 ( .A1(n156), .A2(n155), .ZN(n179) );
  NAND2_X1 U14 ( .A1(n154), .A2(n153), .ZN(n155) );
  NAND2_X1 U15 ( .A1(n152), .A2(n151), .ZN(n156) );
  OR2_X1 U16 ( .A1(n154), .A2(n153), .ZN(n151) );
  XNOR2_X1 U17 ( .A(n152), .B(n97), .ZN(n239) );
  XNOR2_X1 U18 ( .A(n154), .B(n153), .ZN(n97) );
  NAND2_X1 U19 ( .A1(n131), .A2(n130), .ZN(n184) );
  NAND2_X1 U20 ( .A1(n23), .A2(n129), .ZN(n131) );
  NAND2_X1 U21 ( .A1(n54), .A2(n53), .ZN(n255) );
  NAND2_X1 U22 ( .A1(n52), .A2(n261), .ZN(n54) );
  OAI21_X1 U23 ( .B1(n52), .B2(n261), .A(n263), .ZN(n53) );
  OAI21_X1 U24 ( .B1(n164), .B2(n31), .A(n163), .ZN(n190) );
  NAND2_X1 U25 ( .A1(n162), .A2(n161), .ZN(n163) );
  NOR2_X1 U26 ( .A1(n162), .A2(n161), .ZN(n164) );
  OR2_X1 U27 ( .A1(n62), .A2(n61), .ZN(n275) );
  NAND2_X1 U28 ( .A1(n62), .A2(n61), .ZN(n272) );
  NAND2_X1 U29 ( .A1(n302), .A2(n157), .ZN(n159) );
  INV_X1 U30 ( .A(n179), .ZN(n157) );
  NAND2_X1 U31 ( .A1(n56), .A2(n55), .ZN(n394) );
  OR2_X1 U32 ( .A1(n302), .A2(n28), .ZN(n55) );
  OAI21_X1 U33 ( .B1(n256), .B2(n255), .A(n302), .ZN(n56) );
  INV_X1 U34 ( .A(n21), .ZN(n6) );
  NAND2_X1 U35 ( .A1(n20), .A2(\mult_x_1/n310 ), .ZN(n90) );
  OAI22_X1 U36 ( .A1(n116), .A2(n113), .B1(n44), .B2(n114), .ZN(n7) );
  OAI22_X1 U37 ( .A1(n116), .A2(n113), .B1(n44), .B2(n114), .ZN(n172) );
  XNOR2_X1 U38 ( .A(n25), .B(n26), .ZN(n33) );
  XNOR2_X1 U39 ( .A(n128), .B(n140), .ZN(n149) );
  OAI22_X1 U40 ( .A1(n212), .A2(n38), .B1(n214), .B2(n47), .ZN(n11) );
  BUF_X1 U41 ( .A(rst_n), .Z(n412) );
  INV_X1 U42 ( .A(rst_n), .ZN(n564) );
  XOR2_X1 U43 ( .A(n134), .B(n133), .Z(n23) );
  BUF_X1 U44 ( .A(n341), .Z(n253) );
  INV_X1 U45 ( .A(n31), .ZN(n160) );
  NAND2_X1 U46 ( .A1(n133), .A2(n134), .ZN(n31) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(n26), .ZN(n32) );
  NAND2_X2 U48 ( .A1(n32), .A2(n33), .ZN(n223) );
  XNOR2_X1 U49 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n40) );
  CLKBUF_X2 U50 ( .A(n33), .Z(n224) );
  XNOR2_X1 U51 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n37) );
  OAI22_X1 U52 ( .A1(n223), .A2(n40), .B1(n224), .B2(n37), .ZN(n259) );
  XNOR2_X1 U53 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n36) );
  INV_X1 U54 ( .A(n36), .ZN(n34) );
  INV_X2 U55 ( .A(n34), .ZN(n212) );
  AND2_X1 U56 ( .A1(n563), .A2(\mult_x_1/n281 ), .ZN(n198) );
  XNOR2_X1 U57 ( .A(n198), .B(n5), .ZN(n38) );
  XNOR2_X1 U58 ( .A(n562), .B(n27), .ZN(n35) );
  NAND2_X1 U59 ( .A1(n35), .A2(n36), .ZN(n214) );
  XNOR2_X1 U60 ( .A(n5), .B(\mult_x_1/n281 ), .ZN(n47) );
  OAI22_X1 U61 ( .A1(n212), .A2(n38), .B1(n214), .B2(n47), .ZN(n200) );
  INV_X1 U62 ( .A(n200), .ZN(n258) );
  NOR2_X1 U63 ( .A1(n15), .A2(n90), .ZN(n196) );
  XNOR2_X1 U64 ( .A(n6), .B(\mult_x_1/n281 ), .ZN(n199) );
  OAI22_X1 U65 ( .A1(n223), .A2(n37), .B1(n224), .B2(n199), .ZN(n202) );
  AOI21_X1 U66 ( .B1(n212), .B2(n214), .A(n38), .ZN(n39) );
  INV_X1 U67 ( .A(n39), .ZN(n201) );
  FA_X1 U68 ( .A(n260), .B(n259), .CI(n258), .S(n52) );
  XNOR2_X1 U69 ( .A(n6), .B(\mult_x_1/n284 ), .ZN(n46) );
  OAI22_X1 U70 ( .A1(n223), .A2(n46), .B1(n224), .B2(n40), .ZN(n173) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n312 ), .B(n24), .ZN(n41) );
  XNOR2_X1 U72 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n42) );
  NAND2_X1 U73 ( .A1(n41), .A2(n42), .ZN(n116) );
  XNOR2_X1 U74 ( .A(n10), .B(\mult_x_1/n281 ), .ZN(n113) );
  XNOR2_X1 U75 ( .A(n198), .B(\mult_x_1/n312 ), .ZN(n44) );
  INV_X1 U76 ( .A(n42), .ZN(n43) );
  INV_X2 U77 ( .A(n43), .ZN(n114) );
  AOI21_X1 U78 ( .B1(n114), .B2(n116), .A(n44), .ZN(n45) );
  INV_X1 U79 ( .A(n45), .ZN(n171) );
  XNOR2_X1 U80 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n123) );
  OAI22_X1 U81 ( .A1(n223), .A2(n123), .B1(n224), .B2(n46), .ZN(n137) );
  XNOR2_X1 U82 ( .A(n5), .B(\mult_x_1/n283 ), .ZN(n111) );
  XNOR2_X1 U83 ( .A(n5), .B(\mult_x_1/n282 ), .ZN(n48) );
  OAI22_X1 U84 ( .A1(n214), .A2(n111), .B1(n212), .B2(n48), .ZN(n136) );
  INV_X1 U85 ( .A(n172), .ZN(n135) );
  NOR2_X1 U86 ( .A1(n16), .A2(n90), .ZN(n175) );
  OAI22_X1 U87 ( .A1(n214), .A2(n48), .B1(n212), .B2(n47), .ZN(n174) );
  NAND2_X1 U88 ( .A1(n177), .A2(n49), .ZN(n51) );
  BUF_X4 U89 ( .A(en), .Z(n302) );
  XNOR2_X1 U90 ( .A(n10), .B(\mult_x_1/n286 ), .ZN(n60) );
  XNOR2_X1 U91 ( .A(n10), .B(\mult_x_1/n285 ), .ZN(n102) );
  OAI22_X1 U92 ( .A1(n116), .A2(n60), .B1(n114), .B2(n102), .ZN(n249) );
  NAND2_X1 U93 ( .A1(n12), .A2(\mult_x_1/n313 ), .ZN(n126) );
  BUF_X2 U94 ( .A(\mult_x_1/n313 ), .Z(n94) );
  XNOR2_X1 U95 ( .A(n94), .B(\mult_x_1/n284 ), .ZN(n59) );
  XNOR2_X1 U96 ( .A(n94), .B(\mult_x_1/n283 ), .ZN(n99) );
  OAI22_X1 U97 ( .A1(n126), .A2(n59), .B1(n99), .B2(n12), .ZN(n248) );
  OR2_X1 U98 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n57) );
  OAI22_X1 U99 ( .A1(n214), .A2(n25), .B1(n57), .B2(n212), .ZN(n210) );
  XNOR2_X1 U100 ( .A(n5), .B(\mult_x_1/n288 ), .ZN(n58) );
  XNOR2_X1 U101 ( .A(n5), .B(\mult_x_1/n287 ), .ZN(n213) );
  OAI22_X1 U102 ( .A1(n214), .A2(n58), .B1(n212), .B2(n213), .ZN(n209) );
  XNOR2_X1 U103 ( .A(n94), .B(\mult_x_1/n285 ), .ZN(n68) );
  OAI22_X1 U104 ( .A1(n126), .A2(n68), .B1(n59), .B2(n12), .ZN(n65) );
  AND2_X1 U105 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n64) );
  XNOR2_X1 U106 ( .A(n10), .B(\mult_x_1/n287 ), .ZN(n66) );
  OAI22_X1 U107 ( .A1(n116), .A2(n66), .B1(n114), .B2(n60), .ZN(n63) );
  NAND2_X1 U108 ( .A1(n275), .A2(n272), .ZN(n84) );
  FA_X1 U109 ( .A(n65), .B(n64), .CI(n63), .CO(n61), .S(n82) );
  XNOR2_X1 U110 ( .A(n10), .B(\mult_x_1/n288 ), .ZN(n67) );
  OAI22_X1 U111 ( .A1(n116), .A2(n67), .B1(n114), .B2(n66), .ZN(n70) );
  XNOR2_X1 U112 ( .A(n94), .B(\mult_x_1/n286 ), .ZN(n72) );
  OAI22_X1 U113 ( .A1(n126), .A2(n72), .B1(n68), .B2(n12), .ZN(n69) );
  NOR2_X1 U114 ( .A1(n82), .A2(n81), .ZN(n293) );
  HA_X1 U115 ( .A(n70), .B(n69), .CO(n81), .S(n79) );
  OR2_X1 U116 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n71) );
  OAI22_X1 U117 ( .A1(n116), .A2(n22), .B1(n71), .B2(n114), .ZN(n78) );
  OR2_X1 U118 ( .A1(n79), .A2(n78), .ZN(n289) );
  XNOR2_X1 U119 ( .A(n94), .B(\mult_x_1/n287 ), .ZN(n74) );
  OAI22_X1 U120 ( .A1(n126), .A2(n74), .B1(n72), .B2(n12), .ZN(n77) );
  INV_X1 U121 ( .A(n114), .ZN(n73) );
  AND2_X1 U122 ( .A1(\mult_x_1/n288 ), .A2(n73), .ZN(n76) );
  NOR2_X1 U123 ( .A1(n77), .A2(n76), .ZN(n282) );
  OAI22_X1 U124 ( .A1(n126), .A2(\mult_x_1/n288 ), .B1(n74), .B2(n12), .ZN(
        n279) );
  OR2_X1 U125 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n75) );
  NAND2_X1 U126 ( .A1(n75), .A2(n126), .ZN(n278) );
  NAND2_X1 U127 ( .A1(n279), .A2(n278), .ZN(n285) );
  NAND2_X1 U128 ( .A1(n77), .A2(n76), .ZN(n283) );
  OAI21_X1 U129 ( .B1(n282), .B2(n285), .A(n283), .ZN(n290) );
  NAND2_X1 U130 ( .A1(n79), .A2(n78), .ZN(n288) );
  INV_X1 U131 ( .A(n288), .ZN(n80) );
  AOI21_X1 U132 ( .B1(n289), .B2(n290), .A(n80), .ZN(n296) );
  NAND2_X1 U133 ( .A1(n82), .A2(n81), .ZN(n294) );
  OAI21_X1 U134 ( .B1(n293), .B2(n296), .A(n294), .ZN(n274) );
  INV_X1 U135 ( .A(n274), .ZN(n83) );
  XNOR2_X1 U136 ( .A(n84), .B(n83), .ZN(n87) );
  INV_X1 U137 ( .A(n302), .ZN(n86) );
  NAND2_X1 U138 ( .A1(n86), .A2(n541), .ZN(n85) );
  OAI21_X1 U139 ( .B1(n87), .B2(n86), .A(n85), .ZN(n449) );
  XNOR2_X1 U140 ( .A(n5), .B(\mult_x_1/n285 ), .ZN(n93) );
  XNOR2_X1 U141 ( .A(n5), .B(\mult_x_1/n284 ), .ZN(n112) );
  OAI22_X1 U142 ( .A1(n214), .A2(n93), .B1(n212), .B2(n112), .ZN(n122) );
  XNOR2_X1 U143 ( .A(n10), .B(\mult_x_1/n283 ), .ZN(n96) );
  XNOR2_X1 U144 ( .A(n10), .B(\mult_x_1/n282 ), .ZN(n115) );
  OAI22_X1 U145 ( .A1(n116), .A2(n96), .B1(n114), .B2(n115), .ZN(n121) );
  OR2_X1 U146 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n88) );
  OAI22_X1 U147 ( .A1(n223), .A2(n21), .B1(n88), .B2(n224), .ZN(n104) );
  XNOR2_X1 U148 ( .A(n6), .B(\mult_x_1/n288 ), .ZN(n89) );
  XNOR2_X1 U149 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n92) );
  OAI22_X1 U150 ( .A1(n223), .A2(n89), .B1(n224), .B2(n92), .ZN(n103) );
  INV_X1 U151 ( .A(n90), .ZN(n91) );
  AND2_X1 U152 ( .A1(\mult_x_1/n288 ), .A2(n91), .ZN(n119) );
  XNOR2_X1 U153 ( .A(n94), .B(\mult_x_1/n281 ), .ZN(n95) );
  XNOR2_X1 U154 ( .A(n198), .B(n94), .ZN(n125) );
  OAI22_X1 U155 ( .A1(n126), .A2(n95), .B1(n125), .B2(n12), .ZN(n118) );
  XNOR2_X1 U156 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n124) );
  OAI22_X1 U157 ( .A1(n223), .A2(n92), .B1(n224), .B2(n124), .ZN(n117) );
  XNOR2_X1 U158 ( .A(n5), .B(\mult_x_1/n286 ), .ZN(n211) );
  OAI22_X1 U159 ( .A1(n214), .A2(n211), .B1(n212), .B2(n93), .ZN(n107) );
  XNOR2_X1 U160 ( .A(n94), .B(\mult_x_1/n282 ), .ZN(n98) );
  OAI22_X1 U161 ( .A1(n126), .A2(n98), .B1(n95), .B2(n12), .ZN(n106) );
  XNOR2_X1 U162 ( .A(n10), .B(\mult_x_1/n284 ), .ZN(n101) );
  OAI22_X1 U163 ( .A1(n116), .A2(n101), .B1(n114), .B2(n96), .ZN(n105) );
  OAI22_X1 U164 ( .A1(n126), .A2(n99), .B1(n98), .B2(n12), .ZN(n217) );
  INV_X1 U165 ( .A(n224), .ZN(n100) );
  AND2_X1 U166 ( .A1(\mult_x_1/n288 ), .A2(n100), .ZN(n216) );
  OAI22_X1 U167 ( .A1(n116), .A2(n102), .B1(n114), .B2(n101), .ZN(n215) );
  HA_X1 U168 ( .A(n104), .B(n103), .CO(n120), .S(n207) );
  FA_X1 U169 ( .A(n107), .B(n106), .CI(n105), .CO(n153), .S(n206) );
  NAND2_X1 U170 ( .A1(n239), .A2(n238), .ZN(n108) );
  NAND2_X1 U171 ( .A1(n108), .A2(n253), .ZN(n110) );
  OR2_X1 U172 ( .A1(n253), .A2(n29), .ZN(n109) );
  NAND2_X1 U173 ( .A1(n110), .A2(n109), .ZN(n376) );
  OAI22_X1 U174 ( .A1(n214), .A2(n112), .B1(n212), .B2(n111), .ZN(n139) );
  OAI22_X1 U175 ( .A1(n116), .A2(n115), .B1(n114), .B2(n113), .ZN(n138) );
  XNOR2_X1 U176 ( .A(n139), .B(n138), .ZN(n134) );
  FA_X1 U177 ( .A(n119), .B(n118), .CI(n117), .CO(n133), .S(n154) );
  FA_X1 U178 ( .A(n122), .B(n121), .CI(n120), .CO(n148), .S(n152) );
  OAI22_X1 U179 ( .A1(n223), .A2(n124), .B1(n224), .B2(n123), .ZN(n142) );
  AOI21_X1 U180 ( .B1(n126), .B2(n12), .A(n125), .ZN(n127) );
  INV_X1 U181 ( .A(n127), .ZN(n141) );
  XNOR2_X1 U182 ( .A(n142), .B(n141), .ZN(n128) );
  NOR2_X1 U183 ( .A1(n17), .A2(n90), .ZN(n140) );
  OR2_X1 U184 ( .A1(n148), .A2(n149), .ZN(n129) );
  NAND2_X1 U185 ( .A1(n149), .A2(n148), .ZN(n130) );
  INV_X1 U186 ( .A(n184), .ZN(n132) );
  NAND2_X1 U187 ( .A1(n132), .A2(n302), .ZN(n147) );
  FA_X1 U188 ( .A(n137), .B(n136), .CI(n135), .CO(n177), .S(n161) );
  XNOR2_X1 U189 ( .A(n160), .B(n161), .ZN(n146) );
  OR2_X1 U190 ( .A1(n139), .A2(n138), .ZN(n168) );
  NOR2_X1 U191 ( .A1(n18), .A2(n90), .ZN(n167) );
  XNOR2_X1 U192 ( .A(n168), .B(n167), .ZN(n145) );
  OAI21_X1 U193 ( .B1(n142), .B2(n141), .A(n140), .ZN(n144) );
  NAND2_X1 U194 ( .A1(n142), .A2(n141), .ZN(n143) );
  NAND2_X1 U195 ( .A1(n144), .A2(n143), .ZN(n166) );
  XNOR2_X1 U196 ( .A(n145), .B(n166), .ZN(n162) );
  XNOR2_X1 U197 ( .A(n146), .B(n162), .ZN(n185) );
  OAI22_X1 U198 ( .A1(n147), .A2(n185), .B1(n302), .B2(n410), .ZN(n384) );
  XNOR2_X1 U199 ( .A(n149), .B(n148), .ZN(n150) );
  INV_X1 U200 ( .A(n302), .ZN(n187) );
  NAND2_X1 U201 ( .A1(n187), .A2(n357), .ZN(n158) );
  OAI21_X1 U202 ( .B1(n180), .B2(n159), .A(n158), .ZN(n392) );
  INV_X1 U203 ( .A(n190), .ZN(n165) );
  NAND2_X1 U204 ( .A1(n253), .A2(n165), .ZN(n178) );
  OAI21_X1 U205 ( .B1(n167), .B2(n168), .A(n166), .ZN(n170) );
  NAND2_X1 U206 ( .A1(n168), .A2(n167), .ZN(n169) );
  NAND2_X1 U207 ( .A1(n170), .A2(n169), .ZN(n267) );
  FA_X1 U208 ( .A(n173), .B(n7), .CI(n171), .CO(n261), .S(n266) );
  XNOR2_X1 U209 ( .A(n175), .B(n174), .ZN(n176) );
  XNOR2_X1 U210 ( .A(n177), .B(n176), .ZN(n265) );
  OAI22_X1 U211 ( .A1(n178), .A2(n191), .B1(n341), .B2(n403), .ZN(n370) );
  NAND2_X1 U212 ( .A1(n180), .A2(n179), .ZN(n181) );
  NAND2_X1 U213 ( .A1(n181), .A2(n253), .ZN(n183) );
  NAND2_X1 U214 ( .A1(n86), .A2(n347), .ZN(n182) );
  NAND2_X1 U215 ( .A1(n183), .A2(n182), .ZN(n372) );
  NAND2_X1 U216 ( .A1(n185), .A2(n184), .ZN(n186) );
  NAND2_X1 U217 ( .A1(n186), .A2(n302), .ZN(n189) );
  NAND2_X1 U218 ( .A1(n187), .A2(n354), .ZN(n188) );
  NAND2_X1 U219 ( .A1(n189), .A2(n188), .ZN(n386) );
  NAND2_X1 U220 ( .A1(n191), .A2(n190), .ZN(n192) );
  NAND2_X1 U221 ( .A1(n192), .A2(n302), .ZN(n194) );
  OR2_X1 U222 ( .A1(n302), .A2(n404), .ZN(n193) );
  NAND2_X1 U223 ( .A1(n194), .A2(n193), .ZN(n396) );
  FA_X1 U244 ( .A(n197), .B(n196), .CI(n195), .CO(n235), .S(n256) );
  INV_X1 U245 ( .A(n235), .ZN(n204) );
  NOR2_X1 U246 ( .A1(n19), .A2(n90), .ZN(n221) );
  XNOR2_X1 U247 ( .A(n198), .B(n6), .ZN(n222) );
  OAI22_X1 U248 ( .A1(n223), .A2(n199), .B1(n222), .B2(n224), .ZN(n229) );
  INV_X1 U249 ( .A(n229), .ZN(n220) );
  FA_X1 U250 ( .A(n202), .B(n201), .CI(n11), .CO(n219), .S(n195) );
  INV_X1 U251 ( .A(n236), .ZN(n203) );
  NAND2_X1 U252 ( .A1(n204), .A2(n203), .ZN(n205) );
  MUX2_X1 U253 ( .A(n342), .B(n205), .S(n253), .Z(n362) );
  FA_X1 U254 ( .A(n208), .B(n207), .CI(n206), .CO(n238), .S(n242) );
  HA_X1 U255 ( .A(n210), .B(n209), .CO(n246), .S(n247) );
  OAI22_X1 U256 ( .A1(n214), .A2(n213), .B1(n212), .B2(n211), .ZN(n245) );
  FA_X1 U257 ( .A(n217), .B(n216), .CI(n215), .CO(n208), .S(n244) );
  OR2_X1 U258 ( .A1(n242), .A2(n241), .ZN(n218) );
  MUX2_X1 U259 ( .A(n343), .B(n218), .S(n302), .Z(n364) );
  FA_X1 U260 ( .A(n221), .B(n220), .CI(n219), .CO(n231), .S(n236) );
  AOI21_X1 U261 ( .B1(n224), .B2(n223), .A(n222), .ZN(n225) );
  INV_X1 U262 ( .A(n225), .ZN(n227) );
  NOR2_X1 U263 ( .A1(n14), .A2(n90), .ZN(n226) );
  XOR2_X1 U264 ( .A(n227), .B(n226), .Z(n228) );
  XOR2_X1 U265 ( .A(n229), .B(n228), .Z(n230) );
  OR2_X1 U266 ( .A1(n231), .A2(n230), .ZN(n233) );
  NAND2_X1 U267 ( .A1(n231), .A2(n230), .ZN(n232) );
  NAND2_X1 U268 ( .A1(n233), .A2(n232), .ZN(n234) );
  MUX2_X1 U269 ( .A(n344), .B(n234), .S(n302), .Z(n366) );
  NAND2_X1 U270 ( .A1(n236), .A2(n235), .ZN(n237) );
  MUX2_X1 U271 ( .A(n345), .B(n237), .S(n341), .Z(n368) );
  NOR2_X1 U272 ( .A1(n239), .A2(n238), .ZN(n240) );
  MUX2_X1 U273 ( .A(n348), .B(n240), .S(n302), .Z(n374) );
  NAND2_X1 U274 ( .A1(n242), .A2(n241), .ZN(n243) );
  MUX2_X1 U275 ( .A(n350), .B(n243), .S(n8), .Z(n378) );
  FA_X1 U276 ( .A(n246), .B(n245), .CI(n244), .CO(n241), .S(n252) );
  FA_X1 U277 ( .A(n249), .B(n248), .CI(n247), .CO(n251), .S(n62) );
  NOR2_X1 U278 ( .A1(n252), .A2(n251), .ZN(n250) );
  MUX2_X1 U279 ( .A(n351), .B(n250), .S(n302), .Z(n380) );
  NAND2_X1 U280 ( .A1(n252), .A2(n251), .ZN(n254) );
  MUX2_X1 U281 ( .A(n352), .B(n254), .S(n253), .Z(n382) );
  NAND2_X1 U282 ( .A1(n256), .A2(n255), .ZN(n257) );
  MUX2_X1 U283 ( .A(n355), .B(n257), .S(n302), .Z(n388) );
  FA_X1 U284 ( .A(n260), .B(n259), .CI(n258), .CO(n197), .S(n262) );
  XNOR2_X1 U285 ( .A(n262), .B(n261), .ZN(n264) );
  XNOR2_X1 U286 ( .A(n264), .B(n263), .ZN(n270) );
  FA_X1 U287 ( .A(n267), .B(n266), .CI(n265), .CO(n269), .S(n191) );
  NAND2_X1 U288 ( .A1(n270), .A2(n269), .ZN(n268) );
  MUX2_X1 U289 ( .A(n356), .B(n268), .S(n302), .Z(n390) );
  OR2_X1 U290 ( .A1(n270), .A2(n269), .ZN(n271) );
  MUX2_X1 U291 ( .A(n360), .B(n271), .S(n302), .Z(n398) );
  INV_X1 U292 ( .A(n272), .ZN(n273) );
  AOI21_X1 U293 ( .B1(n275), .B2(n274), .A(n273), .ZN(n276) );
  MUX2_X1 U294 ( .A(n361), .B(n276), .S(n302), .Z(n400) );
  MUX2_X1 U295 ( .A(product[0]), .B(n525), .S(n302), .Z(n415) );
  MUX2_X1 U296 ( .A(n525), .B(n526), .S(n302), .Z(n417) );
  AND2_X1 U297 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n277) );
  MUX2_X1 U298 ( .A(n526), .B(n277), .S(n302), .Z(n419) );
  MUX2_X1 U299 ( .A(product[1]), .B(n528), .S(n302), .Z(n421) );
  MUX2_X1 U300 ( .A(n528), .B(n529), .S(n302), .Z(n423) );
  OR2_X1 U301 ( .A1(n279), .A2(n278), .ZN(n280) );
  AND2_X1 U302 ( .A1(n280), .A2(n285), .ZN(n281) );
  MUX2_X1 U303 ( .A(n529), .B(n281), .S(n302), .Z(n425) );
  MUX2_X1 U304 ( .A(product[2]), .B(n531), .S(n302), .Z(n427) );
  MUX2_X1 U305 ( .A(n531), .B(n532), .S(n302), .Z(n429) );
  INV_X1 U306 ( .A(n282), .ZN(n284) );
  NAND2_X1 U307 ( .A1(n284), .A2(n283), .ZN(n286) );
  XOR2_X1 U308 ( .A(n286), .B(n285), .Z(n287) );
  MUX2_X1 U309 ( .A(n532), .B(n287), .S(n302), .Z(n431) );
  MUX2_X1 U310 ( .A(product[3]), .B(n534), .S(n302), .Z(n433) );
  MUX2_X1 U311 ( .A(n534), .B(n535), .S(n302), .Z(n435) );
  NAND2_X1 U312 ( .A1(n289), .A2(n288), .ZN(n291) );
  XNOR2_X1 U313 ( .A(n291), .B(n290), .ZN(n292) );
  MUX2_X1 U314 ( .A(n535), .B(n292), .S(n302), .Z(n437) );
  MUX2_X1 U315 ( .A(product[4]), .B(n537), .S(n302), .Z(n439) );
  MUX2_X1 U316 ( .A(n537), .B(n538), .S(n302), .Z(n441) );
  INV_X1 U317 ( .A(n293), .ZN(n295) );
  NAND2_X1 U318 ( .A1(n295), .A2(n294), .ZN(n297) );
  XOR2_X1 U319 ( .A(n297), .B(n296), .Z(n298) );
  MUX2_X1 U320 ( .A(n538), .B(n298), .S(n302), .Z(n443) );
  MUX2_X1 U321 ( .A(product[5]), .B(n540), .S(n302), .Z(n445) );
  MUX2_X1 U322 ( .A(n540), .B(n541), .S(n302), .Z(n447) );
  MUX2_X1 U323 ( .A(product[6]), .B(n543), .S(n302), .Z(n451) );
  NAND2_X1 U324 ( .A1(n405), .A2(n352), .ZN(n299) );
  XOR2_X1 U325 ( .A(n299), .B(n361), .Z(n300) );
  MUX2_X1 U326 ( .A(n543), .B(n300), .S(n302), .Z(n453) );
  MUX2_X1 U327 ( .A(product[7]), .B(n545), .S(n302), .Z(n455) );
  OAI21_X1 U328 ( .B1(n351), .B2(n361), .A(n352), .ZN(n304) );
  NAND2_X1 U329 ( .A1(n343), .A2(n350), .ZN(n301) );
  XNOR2_X1 U330 ( .A(n304), .B(n301), .ZN(n303) );
  MUX2_X1 U331 ( .A(n545), .B(n303), .S(n302), .Z(n457) );
  MUX2_X1 U332 ( .A(product[8]), .B(n547), .S(n9), .Z(n459) );
  AOI21_X1 U333 ( .B1(n304), .B2(n343), .A(n407), .ZN(n307) );
  NAND2_X1 U334 ( .A1(n408), .A2(n349), .ZN(n305) );
  XOR2_X1 U335 ( .A(n307), .B(n305), .Z(n306) );
  MUX2_X1 U336 ( .A(n547), .B(n306), .S(n9), .Z(n461) );
  MUX2_X1 U337 ( .A(product[9]), .B(n549), .S(n9), .Z(n463) );
  OAI21_X1 U338 ( .B1(n307), .B2(n348), .A(n349), .ZN(n315) );
  INV_X1 U339 ( .A(n315), .ZN(n310) );
  NAND2_X1 U340 ( .A1(n409), .A2(n347), .ZN(n308) );
  XOR2_X1 U341 ( .A(n310), .B(n308), .Z(n309) );
  MUX2_X1 U342 ( .A(n549), .B(n309), .S(n9), .Z(n465) );
  MUX2_X1 U343 ( .A(product[10]), .B(n551), .S(n8), .Z(n467) );
  OAI21_X1 U344 ( .B1(n310), .B2(n357), .A(n347), .ZN(n312) );
  NAND2_X1 U345 ( .A1(n410), .A2(n354), .ZN(n311) );
  XNOR2_X1 U346 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U347 ( .A(n551), .B(n313), .S(n9), .Z(n469) );
  MUX2_X1 U348 ( .A(product[11]), .B(n553), .S(n8), .Z(n471) );
  NOR2_X1 U349 ( .A1(n353), .A2(n357), .ZN(n316) );
  OAI21_X1 U350 ( .B1(n353), .B2(n347), .A(n354), .ZN(n314) );
  AOI21_X1 U351 ( .B1(n316), .B2(n315), .A(n314), .ZN(n338) );
  NAND2_X1 U352 ( .A1(n403), .A2(n359), .ZN(n317) );
  XOR2_X1 U353 ( .A(n338), .B(n317), .Z(n318) );
  MUX2_X1 U354 ( .A(n553), .B(n318), .S(n9), .Z(n473) );
  MUX2_X1 U355 ( .A(product[12]), .B(n555), .S(n8), .Z(n475) );
  OAI21_X1 U356 ( .B1(n338), .B2(n346), .A(n359), .ZN(n320) );
  NAND2_X1 U357 ( .A1(n360), .A2(n356), .ZN(n319) );
  XNOR2_X1 U358 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U359 ( .A(n555), .B(n321), .S(n9), .Z(n477) );
  MUX2_X1 U360 ( .A(product[13]), .B(n557), .S(n8), .Z(n479) );
  NAND2_X1 U361 ( .A1(n403), .A2(n360), .ZN(n323) );
  AOI21_X1 U362 ( .B1(n404), .B2(n360), .A(n411), .ZN(n322) );
  OAI21_X1 U363 ( .B1(n338), .B2(n323), .A(n322), .ZN(n325) );
  NAND2_X1 U364 ( .A1(n358), .A2(n355), .ZN(n324) );
  XNOR2_X1 U365 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U366 ( .A(n557), .B(n326), .S(n9), .Z(n481) );
  MUX2_X1 U367 ( .A(product[14]), .B(n559), .S(n8), .Z(n483) );
  NAND2_X1 U368 ( .A1(n360), .A2(n358), .ZN(n328) );
  NOR2_X1 U369 ( .A1(n346), .A2(n328), .ZN(n334) );
  INV_X1 U370 ( .A(n334), .ZN(n330) );
  AOI21_X1 U371 ( .B1(n411), .B2(n358), .A(n402), .ZN(n327) );
  OAI21_X1 U372 ( .B1(n328), .B2(n359), .A(n327), .ZN(n335) );
  INV_X1 U373 ( .A(n335), .ZN(n329) );
  OAI21_X1 U374 ( .B1(n338), .B2(n330), .A(n329), .ZN(n332) );
  NAND2_X1 U375 ( .A1(n342), .A2(n345), .ZN(n331) );
  XNOR2_X1 U376 ( .A(n332), .B(n331), .ZN(n333) );
  MUX2_X1 U377 ( .A(n559), .B(n333), .S(n9), .Z(n485) );
  MUX2_X1 U378 ( .A(product[15]), .B(n561), .S(n8), .Z(n487) );
  NAND2_X1 U379 ( .A1(n334), .A2(n342), .ZN(n337) );
  AOI21_X1 U380 ( .B1(n335), .B2(n342), .A(n406), .ZN(n336) );
  OAI21_X1 U381 ( .B1(n338), .B2(n337), .A(n336), .ZN(n339) );
  XNOR2_X1 U382 ( .A(n339), .B(n344), .ZN(n340) );
  MUX2_X1 U383 ( .A(n561), .B(n340), .S(n9), .Z(n489) );
  MUX2_X1 U384 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n9), .Z(n491) );
  MUX2_X1 U385 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n9), .Z(n493) );
  MUX2_X1 U386 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n8), .Z(n495) );
  MUX2_X1 U387 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n9), .Z(n497) );
  MUX2_X1 U388 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n8), .Z(n499) );
  MUX2_X1 U389 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n9), .Z(n501) );
  MUX2_X1 U390 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n8), .Z(n503) );
  MUX2_X1 U391 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n8), .Z(n505) );
  MUX2_X1 U392 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n8), .Z(n507) );
  MUX2_X1 U393 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n8), .Z(n509) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n9), .Z(n511) );
  MUX2_X1 U395 ( .A(n10), .B(A_extended[3]), .S(n8), .Z(n513) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n8), .Z(n515) );
  MUX2_X1 U397 ( .A(n5), .B(A_extended[5]), .S(n8), .Z(n517) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n8), .Z(n519) );
  MUX2_X1 U399 ( .A(n6), .B(A_extended[7]), .S(n9), .Z(n521) );
  OR2_X1 U400 ( .A1(n9), .A2(n563), .ZN(n523) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_12 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n356,
         n358, n360, n362, n364, n366, n368, n370, n372, n374, n376, n378,
         n380, n382, n384, n386, n388, n390, n392, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n409,
         n411, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n505, n507, n509, n511, n513, n515, n517, n519,
         n520, n522, n523, n525, n526, n528, n529, n531, n532, n534, n535,
         n537, n539, n541, n543, n545, n547, n549, n551, n553, n555, n556,
         n557, n558, n559, n560, n561;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n407), .SE(n517), .CK(clk), .Q(n560), 
        .QN(n20) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n407), .SE(n513), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n28) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n407), .SE(n511), .CK(clk), .Q(n558), 
        .QN(n25) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n407), .SE(n509), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n30) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n407), .SE(n507), .CK(clk), .Q(n557), 
        .QN(n23) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n407), .SE(n505), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n29) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n407), .SE(n503), .CK(clk), .Q(n556), 
        .QN(n32) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n407), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n21) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n407), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n17) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n406), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n19) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n406), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n18) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n406), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n16) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n406), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n15) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n406), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n26) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n406), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n406), .SE(n483), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n406), .SE(n481), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n406), .SE(n479), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n406), .SE(n477), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n406), .SE(n475), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n406), .SE(n473), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n406), .SE(n471), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n407), .SE(n469), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n406), .SE(n467), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n406), .SE(n465), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n406), .SE(n463), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n406), .SE(n461), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n407), .SE(n459), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n407), .SE(n457), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n406), .SE(n455), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n407), .SE(n453), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n406), .SE(n451), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n406), .SE(n449), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n406), .SE(n447), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n406), .SE(n445), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n406), .SE(n443), .CK(clk), .Q(n535), 
        .QN(n333) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n407), .SE(n441), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n406), .SE(n439), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n406), .SE(n437), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n407), .SE(n435), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n407), .SE(n433), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n406), .SE(n431), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n406), .SE(n429), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n406), .SE(n427), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n407), .SE(n425), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n406), .SE(n423), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n406), .SE(n421), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n407), .SE(n419), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n406), .SE(n417), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n415), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n413), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n411), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n409), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n407), .SE(n515), .CK(clk), .Q(n559), 
        .QN(n27) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n561), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n561), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n352), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n561), .SE(n388), .CK(
        clk), .Q(n404), .QN(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n561), .SE(n386), .CK(
        clk), .Q(n398), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n561), .SE(n384), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n561), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n348), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n561), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n561), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n346), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n561), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n345), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n561), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n561), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n343), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n561), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n561), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n341), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n561), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n340), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n561), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n339), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n561), .SE(n362), .CK(
        clk), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n561), .SE(n360), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n561), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n336), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n561), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n561), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n334), .QN(n397) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n407), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n14) );
  BUF_X2 U2 ( .A(en), .Z(n290) );
  CLKBUF_X2 U3 ( .A(n556), .Z(n329) );
  XNOR2_X1 U4 ( .A(n24), .B(n5), .ZN(n251) );
  XNOR2_X1 U5 ( .A(n232), .B(n231), .ZN(n5) );
  INV_X1 U6 ( .A(n9), .ZN(n162) );
  INV_X1 U7 ( .A(n38), .ZN(n179) );
  XNOR2_X1 U8 ( .A(n130), .B(n82), .ZN(n241) );
  NAND2_X1 U9 ( .A1(n71), .A2(n70), .ZN(n243) );
  XNOR2_X1 U10 ( .A(n131), .B(n132), .ZN(n82) );
  NAND2_X1 U11 ( .A1(n99), .A2(n98), .ZN(n102) );
  NAND2_X1 U12 ( .A1(n22), .A2(n228), .ZN(n98) );
  OAI21_X1 U13 ( .B1(n22), .B2(n228), .A(n229), .ZN(n99) );
  NAND2_X1 U14 ( .A1(n192), .A2(n191), .ZN(n89) );
  NAND2_X1 U15 ( .A1(n132), .A2(n131), .ZN(n133) );
  NAND2_X1 U16 ( .A1(n97), .A2(n31), .ZN(n71) );
  NAND2_X1 U17 ( .A1(n94), .A2(n95), .ZN(n70) );
  CLKBUF_X1 U18 ( .A(n125), .Z(n13) );
  XNOR2_X1 U19 ( .A(n194), .B(n193), .ZN(n204) );
  XNOR2_X1 U20 ( .A(n192), .B(n191), .ZN(n194) );
  NAND2_X1 U21 ( .A1(n136), .A2(n135), .ZN(n225) );
  NAND2_X1 U22 ( .A1(n240), .A2(n237), .ZN(n135) );
  OAI21_X1 U23 ( .B1(n240), .B2(n237), .A(n238), .ZN(n136) );
  BUF_X4 U24 ( .A(en), .Z(n332) );
  OAI211_X1 U25 ( .C1(n106), .C2(n6), .A(n101), .B(n100), .ZN(n366) );
  OR2_X1 U26 ( .A1(n102), .A2(n6), .ZN(n100) );
  NAND2_X1 U27 ( .A1(n6), .A2(n351), .ZN(n104) );
  NAND2_X1 U28 ( .A1(n103), .A2(n262), .ZN(n105) );
  INV_X1 U29 ( .A(n102), .ZN(n103) );
  NAND2_X1 U30 ( .A1(n352), .A2(n6), .ZN(n7) );
  NAND2_X1 U31 ( .A1(n244), .A2(n262), .ZN(n8) );
  NAND2_X1 U32 ( .A1(n7), .A2(n8), .ZN(n390) );
  INV_X1 U33 ( .A(n262), .ZN(n6) );
  BUF_X4 U34 ( .A(en), .Z(n262) );
  XOR2_X1 U35 ( .A(n27), .B(n28), .Z(n68) );
  XOR2_X1 U36 ( .A(\mult_x_1/a[6] ), .B(n558), .Z(n9) );
  NAND2_X1 U37 ( .A1(n68), .A2(n69), .ZN(n12) );
  XNOR2_X1 U38 ( .A(n108), .B(n330), .ZN(n10) );
  OR2_X1 U39 ( .A1(n75), .A2(n74), .ZN(n11) );
  NAND2_X1 U40 ( .A1(n11), .A2(n73), .ZN(n125) );
  AND2_X1 U41 ( .A1(n560), .A2(\mult_x_1/n281 ), .ZN(n108) );
  XNOR2_X1 U42 ( .A(\mult_x_1/a[2] ), .B(n23), .ZN(n34) );
  NAND2_X1 U43 ( .A1(n68), .A2(n69), .ZN(n161) );
  BUF_X1 U44 ( .A(rst_n), .Z(n407) );
  INV_X1 U45 ( .A(rst_n), .ZN(n561) );
  AND2_X1 U46 ( .A1(n177), .A2(n176), .ZN(n22) );
  XOR2_X1 U47 ( .A(n177), .B(n176), .Z(n24) );
  OR2_X1 U48 ( .A1(n94), .A2(n95), .ZN(n31) );
  OR2_X1 U49 ( .A1(n290), .A2(n333), .ZN(n33) );
  BUF_X2 U50 ( .A(n557), .Z(n330) );
  XNOR2_X1 U51 ( .A(n29), .B(n556), .ZN(n35) );
  INV_X1 U52 ( .A(n35), .ZN(n72) );
  NAND2_X1 U53 ( .A1(n34), .A2(n72), .ZN(n75) );
  BUF_X1 U54 ( .A(n75), .Z(n185) );
  XNOR2_X1 U55 ( .A(n330), .B(\mult_x_1/n286 ), .ZN(n42) );
  INV_X1 U56 ( .A(n35), .ZN(n183) );
  XNOR2_X1 U57 ( .A(n330), .B(\mult_x_1/n285 ), .ZN(n140) );
  OAI22_X1 U58 ( .A1(n185), .A2(n42), .B1(n183), .B2(n140), .ZN(n220) );
  NAND2_X1 U59 ( .A1(n329), .A2(n21), .ZN(n146) );
  XNOR2_X1 U60 ( .A(n329), .B(\mult_x_1/n284 ), .ZN(n41) );
  XNOR2_X1 U61 ( .A(n329), .B(\mult_x_1/n283 ), .ZN(n138) );
  OAI22_X1 U62 ( .A1(n146), .A2(n41), .B1(n138), .B2(n21), .ZN(n219) );
  XNOR2_X1 U63 ( .A(n558), .B(n30), .ZN(n36) );
  XNOR2_X1 U64 ( .A(\mult_x_1/a[4] ), .B(n557), .ZN(n37) );
  NAND2_X1 U65 ( .A1(n36), .A2(n37), .ZN(n181) );
  BUF_X2 U66 ( .A(n558), .Z(n331) );
  OR2_X1 U67 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n39) );
  INV_X1 U68 ( .A(n37), .ZN(n38) );
  OAI22_X1 U69 ( .A1(n181), .A2(n25), .B1(n39), .B2(n179), .ZN(n150) );
  XNOR2_X1 U70 ( .A(n331), .B(\mult_x_1/n288 ), .ZN(n40) );
  XNOR2_X1 U71 ( .A(n331), .B(\mult_x_1/n287 ), .ZN(n152) );
  OAI22_X1 U72 ( .A1(n181), .A2(n40), .B1(n179), .B2(n152), .ZN(n149) );
  XNOR2_X1 U73 ( .A(n329), .B(\mult_x_1/n285 ), .ZN(n50) );
  OAI22_X1 U74 ( .A1(n146), .A2(n50), .B1(n41), .B2(n21), .ZN(n47) );
  AND2_X1 U75 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n46) );
  BUF_X1 U76 ( .A(n75), .Z(n148) );
  XNOR2_X1 U77 ( .A(n330), .B(\mult_x_1/n287 ), .ZN(n48) );
  OAI22_X1 U78 ( .A1(n148), .A2(n48), .B1(n183), .B2(n42), .ZN(n45) );
  OR2_X1 U79 ( .A1(n44), .A2(n43), .ZN(n248) );
  NAND2_X1 U80 ( .A1(n44), .A2(n43), .ZN(n245) );
  NAND2_X1 U81 ( .A1(n248), .A2(n245), .ZN(n65) );
  FA_X1 U82 ( .A(n47), .B(n46), .CI(n45), .CO(n43), .S(n63) );
  XNOR2_X1 U83 ( .A(n330), .B(\mult_x_1/n288 ), .ZN(n49) );
  OAI22_X1 U84 ( .A1(n185), .A2(n49), .B1(n183), .B2(n48), .ZN(n52) );
  XNOR2_X1 U85 ( .A(n329), .B(\mult_x_1/n286 ), .ZN(n54) );
  OAI22_X1 U86 ( .A1(n146), .A2(n54), .B1(n50), .B2(n21), .ZN(n51) );
  NOR2_X1 U87 ( .A1(n63), .A2(n62), .ZN(n281) );
  HA_X1 U88 ( .A(n52), .B(n51), .CO(n62), .S(n60) );
  OR2_X1 U89 ( .A1(\mult_x_1/n288 ), .A2(n23), .ZN(n53) );
  OAI22_X1 U90 ( .A1(n148), .A2(n23), .B1(n53), .B2(n183), .ZN(n59) );
  OR2_X1 U91 ( .A1(n60), .A2(n59), .ZN(n277) );
  XNOR2_X1 U92 ( .A(n329), .B(\mult_x_1/n287 ), .ZN(n55) );
  OAI22_X1 U93 ( .A1(n146), .A2(n55), .B1(n54), .B2(n21), .ZN(n58) );
  AND2_X1 U94 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n57) );
  NOR2_X1 U95 ( .A1(n58), .A2(n57), .ZN(n270) );
  OAI22_X1 U96 ( .A1(n146), .A2(\mult_x_1/n288 ), .B1(n55), .B2(n21), .ZN(n267) );
  OR2_X1 U97 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n56) );
  NAND2_X1 U98 ( .A1(n56), .A2(n146), .ZN(n266) );
  NAND2_X1 U99 ( .A1(n267), .A2(n266), .ZN(n273) );
  NAND2_X1 U100 ( .A1(n58), .A2(n57), .ZN(n271) );
  OAI21_X1 U101 ( .B1(n270), .B2(n273), .A(n271), .ZN(n278) );
  NAND2_X1 U102 ( .A1(n60), .A2(n59), .ZN(n276) );
  INV_X1 U103 ( .A(n276), .ZN(n61) );
  AOI21_X1 U104 ( .B1(n277), .B2(n278), .A(n61), .ZN(n284) );
  NAND2_X1 U105 ( .A1(n63), .A2(n62), .ZN(n282) );
  OAI21_X1 U106 ( .B1(n284), .B2(n281), .A(n282), .ZN(n247) );
  INV_X1 U107 ( .A(n247), .ZN(n64) );
  XNOR2_X1 U108 ( .A(n65), .B(n64), .ZN(n66) );
  OAI21_X1 U109 ( .B1(n66), .B2(n6), .A(n33), .ZN(n443) );
  XNOR2_X1 U110 ( .A(n108), .B(n329), .ZN(n85) );
  AOI21_X1 U111 ( .B1(n146), .B2(n21), .A(n85), .ZN(n67) );
  INV_X1 U112 ( .A(n67), .ZN(n190) );
  XNOR2_X1 U113 ( .A(\mult_x_1/a[6] ), .B(n558), .ZN(n69) );
  XNOR2_X1 U114 ( .A(n559), .B(\mult_x_1/n286 ), .ZN(n88) );
  XNOR2_X1 U115 ( .A(n559), .B(\mult_x_1/n285 ), .ZN(n79) );
  OAI22_X1 U116 ( .A1(n12), .A2(n88), .B1(n162), .B2(n79), .ZN(n189) );
  NAND2_X1 U117 ( .A1(n559), .A2(n20), .ZN(n86) );
  NOR2_X1 U118 ( .A1(n26), .A2(n86), .ZN(n188) );
  XNOR2_X1 U119 ( .A(n331), .B(\mult_x_1/n284 ), .ZN(n178) );
  XNOR2_X1 U120 ( .A(n331), .B(\mult_x_1/n283 ), .ZN(n80) );
  OAI22_X1 U121 ( .A1(n181), .A2(n178), .B1(n179), .B2(n80), .ZN(n84) );
  XNOR2_X1 U122 ( .A(n330), .B(\mult_x_1/n282 ), .ZN(n182) );
  XNOR2_X1 U123 ( .A(n330), .B(\mult_x_1/n281 ), .ZN(n74) );
  OAI22_X1 U124 ( .A1(n75), .A2(n182), .B1(n183), .B2(n74), .ZN(n83) );
  OR2_X1 U125 ( .A1(n84), .A2(n83), .ZN(n94) );
  NOR2_X1 U126 ( .A1(n15), .A2(n86), .ZN(n95) );
  XNOR2_X1 U127 ( .A(n559), .B(\mult_x_1/n284 ), .ZN(n78) );
  XNOR2_X1 U128 ( .A(n559), .B(\mult_x_1/n283 ), .ZN(n113) );
  OAI22_X1 U129 ( .A1(n12), .A2(n78), .B1(n162), .B2(n113), .ZN(n126) );
  XNOR2_X1 U130 ( .A(n108), .B(n330), .ZN(n76) );
  OR2_X1 U131 ( .A1(n76), .A2(n72), .ZN(n73) );
  AOI21_X1 U132 ( .B1(n183), .B2(n185), .A(n10), .ZN(n77) );
  INV_X1 U133 ( .A(n77), .ZN(n124) );
  OAI22_X1 U134 ( .A1(n161), .A2(n79), .B1(n162), .B2(n78), .ZN(n93) );
  XNOR2_X1 U135 ( .A(n331), .B(\mult_x_1/n282 ), .ZN(n81) );
  OAI22_X1 U136 ( .A1(n181), .A2(n80), .B1(n179), .B2(n81), .ZN(n92) );
  INV_X1 U137 ( .A(n125), .ZN(n91) );
  NOR2_X1 U138 ( .A1(n16), .A2(n86), .ZN(n131) );
  XNOR2_X1 U139 ( .A(n331), .B(\mult_x_1/n281 ), .ZN(n109) );
  OAI22_X1 U140 ( .A1(n181), .A2(n81), .B1(n179), .B2(n109), .ZN(n132) );
  NAND2_X1 U141 ( .A1(n6), .A2(n340), .ZN(n101) );
  XNOR2_X1 U142 ( .A(n84), .B(n83), .ZN(n177) );
  XNOR2_X1 U143 ( .A(n329), .B(\mult_x_1/n281 ), .ZN(n144) );
  OAI22_X1 U144 ( .A1(n146), .A2(n144), .B1(n85), .B2(n21), .ZN(n191) );
  INV_X1 U145 ( .A(n86), .ZN(n87) );
  AND2_X1 U146 ( .A1(\mult_x_1/n288 ), .A2(n87), .ZN(n192) );
  XNOR2_X1 U147 ( .A(n559), .B(\mult_x_1/n287 ), .ZN(n142) );
  OAI22_X1 U148 ( .A1(n12), .A2(n142), .B1(n162), .B2(n88), .ZN(n193) );
  OAI21_X1 U149 ( .B1(n191), .B2(n192), .A(n193), .ZN(n90) );
  NAND2_X1 U150 ( .A1(n90), .A2(n89), .ZN(n176) );
  FA_X1 U151 ( .A(n93), .B(n92), .CI(n91), .CO(n130), .S(n228) );
  XNOR2_X1 U152 ( .A(n95), .B(n94), .ZN(n96) );
  XNOR2_X1 U153 ( .A(n97), .B(n96), .ZN(n229) );
  OAI21_X1 U154 ( .B1(n106), .B2(n105), .A(n104), .ZN(n388) );
  NOR2_X1 U175 ( .A1(n17), .A2(n86), .ZN(n159) );
  XNOR2_X1 U176 ( .A(n559), .B(\mult_x_1/n281 ), .ZN(n107) );
  XNOR2_X1 U177 ( .A(n108), .B(n559), .ZN(n160) );
  OAI22_X1 U178 ( .A1(n12), .A2(n107), .B1(n160), .B2(n162), .ZN(n167) );
  INV_X1 U179 ( .A(n167), .ZN(n158) );
  XNOR2_X1 U180 ( .A(n559), .B(\mult_x_1/n282 ), .ZN(n112) );
  OAI22_X1 U181 ( .A1(n12), .A2(n112), .B1(n162), .B2(n107), .ZN(n116) );
  XNOR2_X1 U182 ( .A(n108), .B(n331), .ZN(n110) );
  OAI22_X1 U183 ( .A1(n181), .A2(n109), .B1(n110), .B2(n179), .ZN(n115) );
  AOI21_X1 U184 ( .B1(n179), .B2(n181), .A(n110), .ZN(n111) );
  INV_X1 U185 ( .A(n111), .ZN(n114) );
  INV_X1 U186 ( .A(n115), .ZN(n123) );
  OAI22_X1 U187 ( .A1(n12), .A2(n113), .B1(n162), .B2(n112), .ZN(n122) );
  NOR2_X1 U188 ( .A1(n18), .A2(n86), .ZN(n121) );
  NOR2_X1 U189 ( .A1(n19), .A2(n86), .ZN(n119) );
  FA_X1 U190 ( .A(n116), .B(n115), .CI(n114), .CO(n157), .S(n118) );
  OR2_X1 U191 ( .A1(n174), .A2(n173), .ZN(n117) );
  MUX2_X1 U192 ( .A(n334), .B(n117), .S(n290), .Z(n354) );
  FA_X1 U193 ( .A(n120), .B(n119), .CI(n118), .CO(n173), .S(n226) );
  FA_X1 U194 ( .A(n123), .B(n122), .CI(n121), .CO(n120), .S(n240) );
  FA_X1 U195 ( .A(n126), .B(n13), .CI(n124), .CO(n237), .S(n242) );
  INV_X1 U196 ( .A(n132), .ZN(n128) );
  INV_X1 U197 ( .A(n131), .ZN(n127) );
  NAND2_X1 U198 ( .A1(n128), .A2(n127), .ZN(n129) );
  NAND2_X1 U199 ( .A1(n130), .A2(n129), .ZN(n134) );
  NAND2_X1 U200 ( .A1(n134), .A2(n133), .ZN(n238) );
  OR2_X1 U201 ( .A1(n226), .A2(n225), .ZN(n137) );
  MUX2_X1 U202 ( .A(n335), .B(n137), .S(n262), .Z(n356) );
  XNOR2_X1 U203 ( .A(n329), .B(\mult_x_1/n282 ), .ZN(n145) );
  OAI22_X1 U204 ( .A1(n146), .A2(n138), .B1(n145), .B2(n21), .ZN(n155) );
  INV_X1 U205 ( .A(n162), .ZN(n139) );
  AND2_X1 U206 ( .A1(\mult_x_1/n288 ), .A2(n139), .ZN(n154) );
  XNOR2_X1 U207 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n147) );
  OAI22_X1 U208 ( .A1(n148), .A2(n140), .B1(n183), .B2(n147), .ZN(n153) );
  OR2_X1 U209 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n141) );
  OAI22_X1 U210 ( .A1(n161), .A2(n27), .B1(n141), .B2(n162), .ZN(n187) );
  XNOR2_X1 U211 ( .A(n559), .B(\mult_x_1/n288 ), .ZN(n143) );
  OAI22_X1 U212 ( .A1(n161), .A2(n143), .B1(n162), .B2(n142), .ZN(n186) );
  XNOR2_X1 U213 ( .A(n331), .B(\mult_x_1/n286 ), .ZN(n151) );
  XNOR2_X1 U214 ( .A(n331), .B(\mult_x_1/n285 ), .ZN(n180) );
  OAI22_X1 U215 ( .A1(n181), .A2(n151), .B1(n179), .B2(n180), .ZN(n197) );
  OAI22_X1 U216 ( .A1(n146), .A2(n145), .B1(n144), .B2(n21), .ZN(n196) );
  XNOR2_X1 U217 ( .A(n330), .B(\mult_x_1/n283 ), .ZN(n184) );
  OAI22_X1 U218 ( .A1(n148), .A2(n147), .B1(n183), .B2(n184), .ZN(n195) );
  HA_X1 U219 ( .A(n150), .B(n149), .CO(n217), .S(n218) );
  OAI22_X1 U220 ( .A1(n181), .A2(n152), .B1(n179), .B2(n151), .ZN(n216) );
  FA_X1 U221 ( .A(n155), .B(n154), .CI(n153), .CO(n207), .S(n215) );
  OR2_X1 U222 ( .A1(n213), .A2(n212), .ZN(n156) );
  MUX2_X1 U223 ( .A(n337), .B(n156), .S(n262), .Z(n360) );
  FA_X1 U224 ( .A(n159), .B(n158), .CI(n157), .CO(n169), .S(n174) );
  AOI21_X1 U225 ( .B1(n162), .B2(n12), .A(n160), .ZN(n163) );
  INV_X1 U226 ( .A(n163), .ZN(n165) );
  NOR2_X1 U227 ( .A1(n14), .A2(n86), .ZN(n164) );
  XOR2_X1 U228 ( .A(n165), .B(n164), .Z(n166) );
  XOR2_X1 U229 ( .A(n167), .B(n166), .Z(n168) );
  OR2_X1 U230 ( .A1(n169), .A2(n168), .ZN(n171) );
  NAND2_X1 U231 ( .A1(n169), .A2(n168), .ZN(n170) );
  NAND2_X1 U232 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U233 ( .A(n338), .B(n172), .S(n262), .Z(n362) );
  NAND2_X1 U234 ( .A1(n174), .A2(n173), .ZN(n175) );
  MUX2_X1 U235 ( .A(n339), .B(n175), .S(n262), .Z(n364) );
  OAI22_X1 U236 ( .A1(n181), .A2(n180), .B1(n179), .B2(n178), .ZN(n200) );
  OAI22_X1 U237 ( .A1(n185), .A2(n184), .B1(n183), .B2(n182), .ZN(n199) );
  HA_X1 U238 ( .A(n187), .B(n186), .CO(n198), .S(n206) );
  FA_X1 U239 ( .A(n190), .B(n188), .CI(n189), .CO(n97), .S(n231) );
  FA_X1 U240 ( .A(n197), .B(n196), .CI(n195), .CO(n203), .S(n205) );
  FA_X1 U241 ( .A(n200), .B(n199), .CI(n198), .CO(n232), .S(n202) );
  NOR2_X1 U242 ( .A1(n251), .A2(n250), .ZN(n201) );
  MUX2_X1 U243 ( .A(n341), .B(n201), .S(n262), .Z(n368) );
  FA_X1 U244 ( .A(n204), .B(n203), .CI(n202), .CO(n250), .S(n210) );
  FA_X1 U245 ( .A(n207), .B(n206), .CI(n205), .CO(n209), .S(n213) );
  NOR2_X1 U246 ( .A1(n210), .A2(n209), .ZN(n208) );
  MUX2_X1 U247 ( .A(n343), .B(n208), .S(n262), .Z(n372) );
  NAND2_X1 U248 ( .A1(n210), .A2(n209), .ZN(n211) );
  MUX2_X1 U249 ( .A(n344), .B(n211), .S(n262), .Z(n374) );
  NAND2_X1 U250 ( .A1(n213), .A2(n212), .ZN(n214) );
  MUX2_X1 U251 ( .A(n345), .B(n214), .S(n290), .Z(n376) );
  FA_X1 U252 ( .A(n217), .B(n216), .CI(n215), .CO(n212), .S(n223) );
  FA_X1 U253 ( .A(n220), .B(n219), .CI(n218), .CO(n222), .S(n44) );
  NOR2_X1 U254 ( .A1(n223), .A2(n222), .ZN(n221) );
  MUX2_X1 U255 ( .A(n346), .B(n221), .S(n262), .Z(n378) );
  NAND2_X1 U256 ( .A1(n223), .A2(n222), .ZN(n224) );
  MUX2_X1 U257 ( .A(n347), .B(n224), .S(n262), .Z(n380) );
  NAND2_X1 U258 ( .A1(n226), .A2(n225), .ZN(n227) );
  MUX2_X1 U259 ( .A(n348), .B(n227), .S(n262), .Z(n382) );
  XNOR2_X1 U260 ( .A(n22), .B(n228), .ZN(n230) );
  XNOR2_X1 U261 ( .A(n230), .B(n229), .ZN(n260) );
  NAND2_X1 U262 ( .A1(n24), .A2(n232), .ZN(n235) );
  NAND2_X1 U263 ( .A1(n24), .A2(n231), .ZN(n234) );
  NAND2_X1 U264 ( .A1(n232), .A2(n231), .ZN(n233) );
  NAND3_X1 U265 ( .A1(n235), .A2(n234), .A3(n233), .ZN(n259) );
  NOR2_X1 U266 ( .A1(n260), .A2(n259), .ZN(n236) );
  MUX2_X1 U267 ( .A(n350), .B(n236), .S(n262), .Z(n386) );
  XNOR2_X1 U268 ( .A(n238), .B(n237), .ZN(n239) );
  XNOR2_X1 U269 ( .A(n240), .B(n239), .ZN(n256) );
  FA_X1 U270 ( .A(n243), .B(n242), .CI(n241), .CO(n255), .S(n106) );
  NAND2_X1 U271 ( .A1(n256), .A2(n255), .ZN(n244) );
  INV_X1 U272 ( .A(n245), .ZN(n246) );
  AOI21_X1 U273 ( .B1(n248), .B2(n247), .A(n246), .ZN(n249) );
  MUX2_X1 U274 ( .A(n353), .B(n249), .S(n262), .Z(n392) );
  NAND2_X1 U275 ( .A1(n342), .A2(n6), .ZN(n254) );
  NAND2_X1 U276 ( .A1(n251), .A2(n250), .ZN(n252) );
  NAND2_X1 U277 ( .A1(n252), .A2(n290), .ZN(n253) );
  NAND2_X1 U278 ( .A1(n254), .A2(n253), .ZN(n370) );
  OR2_X1 U279 ( .A1(n290), .A2(n396), .ZN(n258) );
  OAI21_X1 U280 ( .B1(n255), .B2(n256), .A(n290), .ZN(n257) );
  NAND2_X1 U281 ( .A1(n258), .A2(n257), .ZN(n358) );
  NAND2_X1 U282 ( .A1(n260), .A2(n259), .ZN(n261) );
  NAND2_X1 U283 ( .A1(n261), .A2(n262), .ZN(n264) );
  NAND2_X1 U284 ( .A1(n6), .A2(n349), .ZN(n263) );
  NAND2_X1 U285 ( .A1(n264), .A2(n263), .ZN(n384) );
  BUF_X2 U286 ( .A(rst_n), .Z(n406) );
  MUX2_X1 U287 ( .A(product[0]), .B(n519), .S(n290), .Z(n409) );
  MUX2_X1 U288 ( .A(n519), .B(n520), .S(n290), .Z(n411) );
  AND2_X1 U289 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n265) );
  MUX2_X1 U290 ( .A(n520), .B(n265), .S(n290), .Z(n413) );
  MUX2_X1 U291 ( .A(product[1]), .B(n522), .S(n290), .Z(n415) );
  MUX2_X1 U292 ( .A(n522), .B(n523), .S(n290), .Z(n417) );
  OR2_X1 U293 ( .A1(n267), .A2(n266), .ZN(n268) );
  AND2_X1 U294 ( .A1(n268), .A2(n273), .ZN(n269) );
  MUX2_X1 U295 ( .A(n523), .B(n269), .S(n290), .Z(n419) );
  MUX2_X1 U296 ( .A(product[2]), .B(n525), .S(n290), .Z(n421) );
  MUX2_X1 U297 ( .A(n525), .B(n526), .S(n290), .Z(n423) );
  INV_X1 U298 ( .A(n270), .ZN(n272) );
  NAND2_X1 U299 ( .A1(n272), .A2(n271), .ZN(n274) );
  XOR2_X1 U300 ( .A(n274), .B(n273), .Z(n275) );
  MUX2_X1 U301 ( .A(n526), .B(n275), .S(n290), .Z(n425) );
  MUX2_X1 U302 ( .A(product[3]), .B(n528), .S(n290), .Z(n427) );
  MUX2_X1 U303 ( .A(n528), .B(n529), .S(n290), .Z(n429) );
  NAND2_X1 U304 ( .A1(n277), .A2(n276), .ZN(n279) );
  XNOR2_X1 U305 ( .A(n279), .B(n278), .ZN(n280) );
  MUX2_X1 U306 ( .A(n529), .B(n280), .S(n290), .Z(n431) );
  MUX2_X1 U307 ( .A(product[4]), .B(n531), .S(n290), .Z(n433) );
  MUX2_X1 U308 ( .A(n531), .B(n532), .S(n290), .Z(n435) );
  INV_X1 U309 ( .A(n281), .ZN(n283) );
  NAND2_X1 U310 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U311 ( .A(n285), .B(n284), .Z(n286) );
  MUX2_X1 U312 ( .A(n532), .B(n286), .S(n290), .Z(n437) );
  MUX2_X1 U313 ( .A(product[5]), .B(n534), .S(n290), .Z(n439) );
  MUX2_X1 U314 ( .A(n534), .B(n535), .S(n290), .Z(n441) );
  MUX2_X1 U315 ( .A(product[6]), .B(n537), .S(n290), .Z(n445) );
  NAND2_X1 U316 ( .A1(n399), .A2(n347), .ZN(n287) );
  XOR2_X1 U317 ( .A(n287), .B(n353), .Z(n288) );
  MUX2_X1 U318 ( .A(n537), .B(n288), .S(n290), .Z(n447) );
  MUX2_X1 U319 ( .A(product[7]), .B(n539), .S(n290), .Z(n449) );
  OAI21_X1 U320 ( .B1(n346), .B2(n353), .A(n347), .ZN(n292) );
  NAND2_X1 U321 ( .A1(n337), .A2(n345), .ZN(n289) );
  XNOR2_X1 U322 ( .A(n292), .B(n289), .ZN(n291) );
  MUX2_X1 U323 ( .A(n539), .B(n291), .S(n290), .Z(n451) );
  MUX2_X1 U324 ( .A(product[8]), .B(n541), .S(n332), .Z(n453) );
  AOI21_X1 U325 ( .B1(n292), .B2(n337), .A(n401), .ZN(n295) );
  NAND2_X1 U326 ( .A1(n402), .A2(n344), .ZN(n293) );
  XOR2_X1 U327 ( .A(n295), .B(n293), .Z(n294) );
  MUX2_X1 U328 ( .A(n541), .B(n294), .S(n332), .Z(n455) );
  MUX2_X1 U329 ( .A(product[9]), .B(n543), .S(n332), .Z(n457) );
  OAI21_X1 U330 ( .B1(n295), .B2(n343), .A(n344), .ZN(n303) );
  INV_X1 U331 ( .A(n303), .ZN(n298) );
  NAND2_X1 U332 ( .A1(n403), .A2(n342), .ZN(n296) );
  XOR2_X1 U333 ( .A(n298), .B(n296), .Z(n297) );
  MUX2_X1 U334 ( .A(n543), .B(n297), .S(n332), .Z(n459) );
  MUX2_X1 U335 ( .A(product[10]), .B(n545), .S(n332), .Z(n461) );
  OAI21_X1 U336 ( .B1(n298), .B2(n341), .A(n342), .ZN(n300) );
  NAND2_X1 U337 ( .A1(n398), .A2(n349), .ZN(n299) );
  XNOR2_X1 U338 ( .A(n300), .B(n299), .ZN(n301) );
  MUX2_X1 U339 ( .A(n545), .B(n301), .S(n332), .Z(n463) );
  MUX2_X1 U340 ( .A(product[11]), .B(n547), .S(n332), .Z(n465) );
  NOR2_X1 U341 ( .A1(n350), .A2(n341), .ZN(n304) );
  OAI21_X1 U342 ( .B1(n350), .B2(n342), .A(n349), .ZN(n302) );
  AOI21_X1 U343 ( .B1(n304), .B2(n303), .A(n302), .ZN(n326) );
  NAND2_X1 U344 ( .A1(n404), .A2(n340), .ZN(n305) );
  XOR2_X1 U345 ( .A(n326), .B(n305), .Z(n306) );
  MUX2_X1 U346 ( .A(n547), .B(n306), .S(n332), .Z(n467) );
  MUX2_X1 U347 ( .A(product[12]), .B(n549), .S(n332), .Z(n469) );
  OAI21_X1 U348 ( .B1(n326), .B2(n351), .A(n340), .ZN(n308) );
  NAND2_X1 U349 ( .A1(n336), .A2(n352), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U351 ( .A(n549), .B(n309), .S(n332), .Z(n471) );
  MUX2_X1 U352 ( .A(product[13]), .B(n551), .S(n332), .Z(n473) );
  NAND2_X1 U353 ( .A1(n404), .A2(n336), .ZN(n311) );
  AOI21_X1 U354 ( .B1(n395), .B2(n336), .A(n405), .ZN(n310) );
  OAI21_X1 U355 ( .B1(n326), .B2(n311), .A(n310), .ZN(n313) );
  NAND2_X1 U356 ( .A1(n335), .A2(n348), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  MUX2_X1 U358 ( .A(n551), .B(n314), .S(n332), .Z(n475) );
  MUX2_X1 U359 ( .A(product[14]), .B(n553), .S(n332), .Z(n477) );
  NAND2_X1 U360 ( .A1(n336), .A2(n335), .ZN(n321) );
  OR2_X1 U361 ( .A1(n351), .A2(n321), .ZN(n317) );
  AOI21_X1 U362 ( .B1(n405), .B2(n335), .A(n400), .ZN(n315) );
  OAI21_X1 U363 ( .B1(n321), .B2(n340), .A(n315), .ZN(n323) );
  INV_X1 U364 ( .A(n323), .ZN(n316) );
  OAI21_X1 U365 ( .B1(n326), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U366 ( .A1(n334), .A2(n339), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U368 ( .A(n553), .B(n320), .S(n332), .Z(n479) );
  MUX2_X1 U369 ( .A(product[15]), .B(n555), .S(n332), .Z(n481) );
  NOR2_X1 U370 ( .A1(n321), .A2(n397), .ZN(n322) );
  NAND2_X1 U371 ( .A1(n404), .A2(n322), .ZN(n325) );
  AOI21_X1 U372 ( .B1(n323), .B2(n334), .A(n394), .ZN(n324) );
  OAI21_X1 U373 ( .B1(n326), .B2(n325), .A(n324), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n327), .B(n338), .ZN(n328) );
  MUX2_X1 U375 ( .A(n555), .B(n328), .S(n332), .Z(n483) );
  MUX2_X1 U376 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n332), .Z(n485) );
  MUX2_X1 U377 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n332), .Z(n487) );
  MUX2_X1 U378 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n332), .Z(n489) );
  MUX2_X1 U379 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n332), .Z(n491) );
  MUX2_X1 U380 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n332), .Z(n493) );
  MUX2_X1 U381 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n332), .Z(n495) );
  MUX2_X1 U382 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n332), .Z(n497) );
  MUX2_X1 U383 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n332), .Z(n499) );
  MUX2_X1 U384 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n332), .Z(n501) );
  MUX2_X1 U385 ( .A(n329), .B(A_extended[1]), .S(n332), .Z(n503) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n332), .Z(n505) );
  MUX2_X1 U387 ( .A(n330), .B(A_extended[3]), .S(n332), .Z(n507) );
  MUX2_X1 U388 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n332), .Z(n509) );
  MUX2_X1 U389 ( .A(n331), .B(A_extended[5]), .S(n332), .Z(n511) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n332), .Z(n513) );
  MUX2_X1 U391 ( .A(n559), .B(A_extended[7]), .S(n332), .Z(n515) );
  OR2_X1 U392 ( .A1(n332), .A2(n560), .ZN(n517) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_13 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n362,
         n364, n366, n368, n370, n372, n374, n376, n378, n380, n382, n384,
         n386, n388, n390, n392, n394, n396, n398, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n411, n413, n415, n417, n419,
         n421, n423, n425, n427, n429, n431, n433, n435, n437, n439, n441,
         n443, n445, n447, n449, n451, n453, n455, n457, n459, n461, n463,
         n465, n467, n469, n471, n473, n475, n477, n479, n481, n483, n485,
         n487, n489, n491, n493, n495, n497, n499, n501, n503, n505, n507,
         n509, n511, n513, n515, n517, n519, n521, n522, n524, n525, n527,
         n528, n530, n531, n533, n534, n536, n537, n539, n541, n543, n545,
         n547, n549, n551, n553, n555, n557, n558, n559, n560, n561;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n409), .SE(n519), .CK(clk), .Q(n560), 
        .QN(n27) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n409), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n409), .SE(n513), .CK(clk), .Q(n559), 
        .QN(n338) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n409), .SE(n511), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n409), .SE(n509), .CK(clk), .Q(n558), 
        .QN(n29) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n409), .SE(n507), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n409), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n409), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n408), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n26) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n408), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n20) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n408), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n22) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n408), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n408), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n23) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n408), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n408), .SE(n485), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n408), .SE(n483), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n408), .SE(n481), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n408), .SE(n479), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n408), .SE(n477), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n408), .SE(n475), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n408), .SE(n473), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n409), .SE(n471), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n409), .SE(n469), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n409), .SE(n467), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n409), .SE(n465), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n409), .SE(n463), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n408), .SE(n461), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n409), .SE(n459), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n408), .SE(n457), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n409), .SE(n455), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n408), .SE(n453), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n408), .SE(n451), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n409), .SE(n449), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n409), .SE(n447), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n409), .SE(n445), .CK(clk), .Q(n537), 
        .QN(n30) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n409), .SE(n443), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n409), .SE(n441), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n409), .SE(n439), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n409), .SE(n437), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n409), .SE(n435), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n408), .SE(n433), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n408), .SE(n431), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n429), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n409), .SE(n427), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n425), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n409), .SE(n423), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n421), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n408), .SE(n419), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n417), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n409), .SE(n415), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n409), .SE(n413), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n409), .SE(n411), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n409), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n31) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n561), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n561), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n561), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n561), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n356), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n561), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n355), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n561), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n561), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n353), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n561), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n352), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n561), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n561), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n350), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n561), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n561), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n348), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n561), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n347), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n561), .SE(n372), .CK(
        clk), .Q(n339), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n561), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n345), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n561), .SE(n368), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n561), .SE(n366), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n561), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n561), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n561), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n340) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n409), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n337) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n409), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n21) );
  BUF_X1 U2 ( .A(n559), .Z(n334) );
  XNOR2_X1 U3 ( .A(n112), .B(n154), .ZN(n6) );
  INV_X1 U4 ( .A(n19), .ZN(n7) );
  XNOR2_X1 U5 ( .A(n112), .B(n333), .ZN(n8) );
  NAND2_X1 U6 ( .A1(n33), .A2(n34), .ZN(n114) );
  NAND2_X1 U7 ( .A1(n154), .A2(n5), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n154), .A2(n5), .ZN(n163) );
  NAND2_X1 U9 ( .A1(n121), .A2(n120), .ZN(n122) );
  INV_X1 U10 ( .A(n17), .ZN(n120) );
  NAND2_X1 U11 ( .A1(n119), .A2(n131), .ZN(n121) );
  XNOR2_X1 U12 ( .A(n98), .B(n97), .ZN(n99) );
  INV_X1 U13 ( .A(n239), .ZN(n235) );
  INV_X1 U14 ( .A(n238), .ZN(n234) );
  NAND2_X1 U15 ( .A1(n139), .A2(n138), .ZN(n140) );
  INV_X1 U16 ( .A(n143), .ZN(n139) );
  NAND2_X1 U17 ( .A1(n102), .A2(n101), .ZN(n105) );
  NAND2_X1 U18 ( .A1(n28), .A2(n258), .ZN(n101) );
  NAND2_X1 U19 ( .A1(n241), .A2(n240), .ZN(n243) );
  NAND2_X1 U20 ( .A1(n239), .A2(n238), .ZN(n240) );
  NAND2_X1 U21 ( .A1(n237), .A2(n236), .ZN(n241) );
  NAND2_X1 U22 ( .A1(n235), .A2(n234), .ZN(n236) );
  NAND2_X1 U23 ( .A1(n123), .A2(n122), .ZN(n129) );
  CLKBUF_X1 U24 ( .A(n249), .Z(n16) );
  XNOR2_X1 U25 ( .A(n259), .B(n28), .ZN(n260) );
  INV_X1 U26 ( .A(n19), .ZN(n18) );
  XOR2_X1 U27 ( .A(n220), .B(n219), .Z(n10) );
  XOR2_X1 U28 ( .A(n218), .B(n10), .Z(n226) );
  NAND2_X1 U29 ( .A1(n218), .A2(n220), .ZN(n11) );
  NAND2_X1 U30 ( .A1(n218), .A2(n219), .ZN(n12) );
  NAND2_X1 U31 ( .A1(n220), .A2(n219), .ZN(n13) );
  NAND3_X1 U32 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n215) );
  NAND2_X2 U33 ( .A1(n37), .A2(n38), .ZN(n14) );
  NAND2_X1 U34 ( .A1(n37), .A2(n38), .ZN(n83) );
  CLKBUF_X1 U35 ( .A(\mult_x_1/n281 ), .Z(n15) );
  MUX2_X1 U36 ( .A(n153), .B(n342), .S(n69), .Z(n364) );
  OAI22_X1 U37 ( .A1(n114), .A2(n113), .B1(n115), .B2(n196), .ZN(n17) );
  NAND2_X1 U38 ( .A1(n143), .A2(n142), .ZN(n144) );
  INV_X1 U39 ( .A(n142), .ZN(n138) );
  XNOR2_X1 U40 ( .A(n143), .B(n142), .ZN(n75) );
  OAI21_X1 U41 ( .B1(n28), .B2(n258), .A(n257), .ZN(n102) );
  XNOR2_X1 U42 ( .A(n258), .B(n257), .ZN(n259) );
  XNOR2_X1 U43 ( .A(n100), .B(n99), .ZN(n257) );
  OR2_X2 U44 ( .A1(n93), .A2(n92), .ZN(n98) );
  XOR2_X1 U45 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .Z(n19) );
  XNOR2_X1 U46 ( .A(n141), .B(n75), .ZN(n152) );
  BUF_X1 U47 ( .A(en), .Z(n107) );
  BUF_X1 U48 ( .A(rst_n), .Z(n408) );
  AND2_X1 U49 ( .A1(n203), .A2(n202), .ZN(n28) );
  INV_X1 U50 ( .A(rst_n), .ZN(n561) );
  OR2_X1 U51 ( .A1(n288), .A2(n30), .ZN(n32) );
  BUF_X4 U52 ( .A(en), .Z(n336) );
  INV_X1 U53 ( .A(n132), .ZN(n119) );
  XNOR2_X1 U54 ( .A(n338), .B(\mult_x_1/a[4] ), .ZN(n33) );
  XNOR2_X1 U55 ( .A(n558), .B(\mult_x_1/a[4] ), .ZN(n34) );
  OR2_X1 U56 ( .A1(\mult_x_1/n288 ), .A2(n338), .ZN(n35) );
  INV_X1 U57 ( .A(n34), .ZN(n41) );
  INV_X2 U58 ( .A(n41), .ZN(n196) );
  OAI22_X1 U59 ( .A1(n114), .A2(n338), .B1(n35), .B2(n196), .ZN(n166) );
  XNOR2_X1 U60 ( .A(n334), .B(\mult_x_1/n288 ), .ZN(n36) );
  XNOR2_X1 U61 ( .A(n334), .B(\mult_x_1/n287 ), .ZN(n168) );
  OAI22_X1 U62 ( .A1(n114), .A2(n36), .B1(n196), .B2(n168), .ZN(n165) );
  XOR2_X1 U63 ( .A(\mult_x_1/a[2] ), .B(n558), .Z(n37) );
  XNOR2_X1 U64 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n38) );
  BUF_X2 U65 ( .A(n558), .Z(n333) );
  XNOR2_X1 U66 ( .A(n333), .B(\mult_x_1/n286 ), .ZN(n42) );
  XNOR2_X1 U67 ( .A(n333), .B(\mult_x_1/n285 ), .ZN(n157) );
  OAI22_X1 U68 ( .A1(n14), .A2(n42), .B1(n18), .B2(n157), .ZN(n239) );
  BUF_X2 U69 ( .A(\mult_x_1/n313 ), .Z(n154) );
  XNOR2_X1 U70 ( .A(n154), .B(\mult_x_1/n284 ), .ZN(n40) );
  XNOR2_X1 U71 ( .A(n154), .B(\mult_x_1/n283 ), .ZN(n155) );
  OAI22_X1 U72 ( .A1(n9), .A2(n40), .B1(n155), .B2(n5), .ZN(n238) );
  XNOR2_X1 U73 ( .A(n239), .B(n238), .ZN(n39) );
  XNOR2_X1 U74 ( .A(n237), .B(n39), .ZN(n46) );
  INV_X1 U75 ( .A(n46), .ZN(n44) );
  XNOR2_X1 U76 ( .A(n154), .B(\mult_x_1/n285 ), .ZN(n52) );
  OAI22_X1 U77 ( .A1(n9), .A2(n52), .B1(n40), .B2(n5), .ZN(n49) );
  AND2_X1 U78 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n48) );
  XNOR2_X1 U79 ( .A(n333), .B(\mult_x_1/n287 ), .ZN(n50) );
  OAI22_X1 U80 ( .A1(n14), .A2(n50), .B1(n18), .B2(n42), .ZN(n47) );
  INV_X1 U81 ( .A(n45), .ZN(n43) );
  NAND2_X1 U82 ( .A1(n44), .A2(n43), .ZN(n255) );
  NAND2_X1 U83 ( .A1(n46), .A2(n45), .ZN(n252) );
  NAND2_X1 U84 ( .A1(n255), .A2(n252), .ZN(n68) );
  FA_X1 U85 ( .A(n49), .B(n48), .CI(n47), .CO(n45), .S(n66) );
  XNOR2_X1 U86 ( .A(n333), .B(\mult_x_1/n288 ), .ZN(n51) );
  OAI22_X1 U87 ( .A1(n14), .A2(n51), .B1(n18), .B2(n50), .ZN(n54) );
  XNOR2_X1 U88 ( .A(n154), .B(\mult_x_1/n286 ), .ZN(n56) );
  OAI22_X1 U89 ( .A1(n9), .A2(n56), .B1(n52), .B2(n5), .ZN(n53) );
  NOR2_X1 U90 ( .A1(n66), .A2(n65), .ZN(n281) );
  HA_X1 U91 ( .A(n54), .B(n53), .CO(n65), .S(n63) );
  OR2_X1 U92 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n55) );
  OAI22_X1 U93 ( .A1(n14), .A2(n29), .B1(n55), .B2(n18), .ZN(n62) );
  OR2_X1 U94 ( .A1(n63), .A2(n62), .ZN(n277) );
  XNOR2_X1 U95 ( .A(n154), .B(\mult_x_1/n287 ), .ZN(n58) );
  OAI22_X1 U96 ( .A1(n9), .A2(n58), .B1(n56), .B2(n5), .ZN(n61) );
  INV_X1 U97 ( .A(n18), .ZN(n57) );
  AND2_X1 U98 ( .A1(\mult_x_1/n288 ), .A2(n57), .ZN(n60) );
  NOR2_X1 U99 ( .A1(n61), .A2(n60), .ZN(n270) );
  OAI22_X1 U100 ( .A1(n9), .A2(\mult_x_1/n288 ), .B1(n58), .B2(n5), .ZN(n267)
         );
  OR2_X1 U101 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n59) );
  NAND2_X1 U102 ( .A1(n59), .A2(n9), .ZN(n266) );
  NAND2_X1 U103 ( .A1(n267), .A2(n266), .ZN(n273) );
  NAND2_X1 U104 ( .A1(n61), .A2(n60), .ZN(n271) );
  OAI21_X1 U105 ( .B1(n270), .B2(n273), .A(n271), .ZN(n278) );
  NAND2_X1 U106 ( .A1(n63), .A2(n62), .ZN(n276) );
  INV_X1 U107 ( .A(n276), .ZN(n64) );
  AOI21_X1 U108 ( .B1(n277), .B2(n278), .A(n64), .ZN(n284) );
  NAND2_X1 U109 ( .A1(n66), .A2(n65), .ZN(n282) );
  OAI21_X1 U110 ( .B1(n281), .B2(n284), .A(n282), .ZN(n254) );
  INV_X1 U111 ( .A(n254), .ZN(n67) );
  XNOR2_X1 U112 ( .A(n68), .B(n67), .ZN(n70) );
  BUF_X2 U113 ( .A(n107), .Z(n288) );
  INV_X1 U114 ( .A(n288), .ZN(n69) );
  OAI21_X1 U115 ( .B1(n70), .B2(n69), .A(n32), .ZN(n445) );
  XOR2_X1 U116 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n71) );
  XNOR2_X1 U117 ( .A(n559), .B(\mult_x_1/a[6] ), .ZN(n72) );
  NAND2_X1 U118 ( .A1(n71), .A2(n72), .ZN(n177) );
  INV_X2 U119 ( .A(n337), .ZN(n335) );
  XNOR2_X1 U120 ( .A(n335), .B(\mult_x_1/n285 ), .ZN(n80) );
  INV_X1 U121 ( .A(n72), .ZN(n73) );
  INV_X2 U122 ( .A(n73), .ZN(n178) );
  XNOR2_X1 U123 ( .A(n335), .B(\mult_x_1/n284 ), .ZN(n76) );
  OAI22_X1 U124 ( .A1(n177), .A2(n80), .B1(n178), .B2(n76), .ZN(n96) );
  XNOR2_X1 U125 ( .A(n334), .B(\mult_x_1/n283 ), .ZN(n81) );
  XNOR2_X1 U126 ( .A(n334), .B(\mult_x_1/n282 ), .ZN(n74) );
  OAI22_X1 U127 ( .A1(n114), .A2(n81), .B1(n196), .B2(n74), .ZN(n95) );
  XNOR2_X1 U128 ( .A(n333), .B(n15), .ZN(n82) );
  AND2_X1 U129 ( .A1(n560), .A2(\mult_x_1/n281 ), .ZN(n112) );
  XNOR2_X1 U130 ( .A(n112), .B(n333), .ZN(n77) );
  OAI22_X1 U131 ( .A1(n83), .A2(n82), .B1(n8), .B2(n7), .ZN(n136) );
  INV_X1 U132 ( .A(n136), .ZN(n94) );
  NAND2_X1 U133 ( .A1(n27), .A2(\mult_x_1/n310 ), .ZN(n90) );
  NOR2_X1 U134 ( .A1(n22), .A2(n90), .ZN(n143) );
  XNOR2_X1 U135 ( .A(n334), .B(n15), .ZN(n113) );
  OAI22_X1 U136 ( .A1(n114), .A2(n74), .B1(n196), .B2(n113), .ZN(n142) );
  XNOR2_X1 U137 ( .A(n335), .B(\mult_x_1/n283 ), .ZN(n118) );
  OAI22_X1 U138 ( .A1(n177), .A2(n76), .B1(n178), .B2(n118), .ZN(n137) );
  AOI21_X1 U139 ( .B1(n18), .B2(n14), .A(n77), .ZN(n78) );
  INV_X1 U140 ( .A(n78), .ZN(n135) );
  XNOR2_X1 U141 ( .A(n112), .B(n154), .ZN(n89) );
  AOI21_X1 U142 ( .B1(n163), .B2(n5), .A(n6), .ZN(n79) );
  INV_X1 U143 ( .A(n79), .ZN(n194) );
  XNOR2_X1 U144 ( .A(n335), .B(\mult_x_1/n286 ), .ZN(n88) );
  OAI22_X1 U145 ( .A1(n177), .A2(n88), .B1(n178), .B2(n80), .ZN(n193) );
  NOR2_X1 U146 ( .A1(n23), .A2(n90), .ZN(n192) );
  XNOR2_X1 U147 ( .A(n334), .B(\mult_x_1/n284 ), .ZN(n195) );
  OAI22_X1 U148 ( .A1(n114), .A2(n195), .B1(n196), .B2(n81), .ZN(n93) );
  XNOR2_X1 U149 ( .A(n333), .B(\mult_x_1/n282 ), .ZN(n198) );
  OAI22_X1 U150 ( .A1(n14), .A2(n198), .B1(n7), .B2(n82), .ZN(n92) );
  INV_X1 U151 ( .A(n98), .ZN(n85) );
  NOR2_X1 U152 ( .A1(n24), .A2(n90), .ZN(n97) );
  INV_X1 U153 ( .A(n97), .ZN(n84) );
  NAND2_X1 U154 ( .A1(n85), .A2(n84), .ZN(n86) );
  AOI22_X1 U155 ( .A1(n100), .A2(n86), .B1(n97), .B2(n98), .ZN(n87) );
  INV_X1 U156 ( .A(n87), .ZN(n150) );
  XNOR2_X1 U157 ( .A(n335), .B(\mult_x_1/n287 ), .ZN(n159) );
  OAI22_X1 U158 ( .A1(n177), .A2(n159), .B1(n178), .B2(n88), .ZN(n207) );
  XNOR2_X1 U159 ( .A(n154), .B(n15), .ZN(n161) );
  OAI22_X1 U160 ( .A1(n9), .A2(n161), .B1(n89), .B2(n5), .ZN(n206) );
  INV_X1 U161 ( .A(n90), .ZN(n91) );
  AND2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n91), .ZN(n205) );
  XNOR2_X1 U163 ( .A(n93), .B(n92), .ZN(n202) );
  FA_X1 U164 ( .A(n96), .B(n95), .CI(n94), .CO(n141), .S(n258) );
  INV_X1 U165 ( .A(n105), .ZN(n103) );
  NAND2_X1 U166 ( .A1(n288), .A2(n103), .ZN(n104) );
  OAI22_X1 U167 ( .A1(n104), .A2(n106), .B1(n336), .B2(n339), .ZN(n372) );
  NAND2_X1 U168 ( .A1(n106), .A2(n105), .ZN(n108) );
  BUF_X2 U169 ( .A(n107), .Z(n291) );
  NAND2_X1 U170 ( .A1(n108), .A2(n291), .ZN(n110) );
  NAND2_X1 U171 ( .A1(n69), .A2(n347), .ZN(n109) );
  NAND2_X1 U172 ( .A1(n110), .A2(n109), .ZN(n374) );
  NOR2_X1 U193 ( .A1(n25), .A2(n90), .ZN(n175) );
  XNOR2_X1 U194 ( .A(n335), .B(n15), .ZN(n111) );
  XNOR2_X1 U195 ( .A(n112), .B(n335), .ZN(n176) );
  OAI22_X1 U196 ( .A1(n177), .A2(n111), .B1(n176), .B2(n178), .ZN(n183) );
  INV_X1 U197 ( .A(n183), .ZN(n174) );
  XNOR2_X1 U198 ( .A(n335), .B(\mult_x_1/n282 ), .ZN(n117) );
  OAI22_X1 U199 ( .A1(n177), .A2(n117), .B1(n178), .B2(n111), .ZN(n125) );
  XNOR2_X1 U200 ( .A(n112), .B(n334), .ZN(n115) );
  OAI22_X1 U201 ( .A1(n114), .A2(n113), .B1(n115), .B2(n196), .ZN(n133) );
  AOI21_X1 U202 ( .B1(n196), .B2(n114), .A(n115), .ZN(n116) );
  INV_X1 U203 ( .A(n116), .ZN(n124) );
  OAI22_X1 U204 ( .A1(n177), .A2(n118), .B1(n178), .B2(n117), .ZN(n132) );
  NOR2_X1 U205 ( .A1(n20), .A2(n90), .ZN(n130) );
  NAND2_X1 U206 ( .A1(n132), .A2(n130), .ZN(n123) );
  NOR2_X1 U207 ( .A1(n26), .A2(n90), .ZN(n128) );
  FA_X1 U208 ( .A(n125), .B(n133), .CI(n124), .CO(n173), .S(n127) );
  OR2_X1 U209 ( .A1(n190), .A2(n189), .ZN(n126) );
  MUX2_X1 U210 ( .A(n340), .B(n126), .S(n336), .Z(n360) );
  FA_X1 U211 ( .A(n129), .B(n128), .CI(n127), .CO(n189), .S(n247) );
  INV_X1 U212 ( .A(n130), .ZN(n131) );
  XNOR2_X1 U213 ( .A(n132), .B(n131), .ZN(n134) );
  XNOR2_X1 U214 ( .A(n134), .B(n17), .ZN(n149) );
  FA_X1 U215 ( .A(n137), .B(n136), .CI(n135), .CO(n148), .S(n151) );
  NAND2_X1 U216 ( .A1(n141), .A2(n140), .ZN(n145) );
  NAND2_X1 U217 ( .A1(n145), .A2(n144), .ZN(n147) );
  OR2_X1 U218 ( .A1(n247), .A2(n246), .ZN(n146) );
  MUX2_X1 U219 ( .A(n341), .B(n146), .S(n291), .Z(n362) );
  FA_X1 U220 ( .A(n149), .B(n148), .CI(n147), .CO(n246), .S(n250) );
  FA_X1 U221 ( .A(n152), .B(n151), .CI(n150), .CO(n249), .S(n106) );
  OR2_X1 U222 ( .A1(n250), .A2(n249), .ZN(n153) );
  XNOR2_X1 U223 ( .A(n154), .B(\mult_x_1/n282 ), .ZN(n162) );
  OAI22_X1 U224 ( .A1(n9), .A2(n155), .B1(n162), .B2(n5), .ZN(n171) );
  INV_X1 U225 ( .A(n178), .ZN(n156) );
  AND2_X1 U226 ( .A1(\mult_x_1/n288 ), .A2(n156), .ZN(n170) );
  XNOR2_X1 U227 ( .A(n333), .B(\mult_x_1/n284 ), .ZN(n164) );
  OAI22_X1 U228 ( .A1(n14), .A2(n157), .B1(n18), .B2(n164), .ZN(n169) );
  OR2_X1 U229 ( .A1(\mult_x_1/n288 ), .A2(n337), .ZN(n158) );
  OAI22_X1 U230 ( .A1(n177), .A2(n337), .B1(n158), .B2(n178), .ZN(n201) );
  XNOR2_X1 U231 ( .A(n335), .B(\mult_x_1/n288 ), .ZN(n160) );
  OAI22_X1 U232 ( .A1(n177), .A2(n160), .B1(n178), .B2(n159), .ZN(n200) );
  XNOR2_X1 U233 ( .A(n334), .B(\mult_x_1/n286 ), .ZN(n167) );
  XNOR2_X1 U234 ( .A(n334), .B(\mult_x_1/n285 ), .ZN(n197) );
  OAI22_X1 U235 ( .A1(n114), .A2(n167), .B1(n196), .B2(n197), .ZN(n210) );
  OAI22_X1 U236 ( .A1(n9), .A2(n162), .B1(n161), .B2(n5), .ZN(n209) );
  XNOR2_X1 U237 ( .A(n333), .B(\mult_x_1/n283 ), .ZN(n199) );
  OAI22_X1 U238 ( .A1(n14), .A2(n164), .B1(n18), .B2(n199), .ZN(n208) );
  HA_X1 U239 ( .A(n166), .B(n165), .CO(n233), .S(n237) );
  OAI22_X1 U240 ( .A1(n114), .A2(n168), .B1(n196), .B2(n167), .ZN(n232) );
  FA_X1 U241 ( .A(n171), .B(n170), .CI(n169), .CO(n223), .S(n231) );
  OR2_X1 U242 ( .A1(n229), .A2(n228), .ZN(n172) );
  MUX2_X1 U243 ( .A(n343), .B(n172), .S(n291), .Z(n366) );
  FA_X1 U244 ( .A(n175), .B(n174), .CI(n173), .CO(n185), .S(n190) );
  AOI21_X1 U245 ( .B1(n178), .B2(n177), .A(n176), .ZN(n179) );
  INV_X1 U246 ( .A(n179), .ZN(n181) );
  NOR2_X1 U247 ( .A1(n21), .A2(n90), .ZN(n180) );
  XOR2_X1 U248 ( .A(n181), .B(n180), .Z(n182) );
  XOR2_X1 U249 ( .A(n183), .B(n182), .Z(n184) );
  OR2_X1 U250 ( .A1(n185), .A2(n184), .ZN(n187) );
  NAND2_X1 U251 ( .A1(n185), .A2(n184), .ZN(n186) );
  NAND2_X1 U252 ( .A1(n187), .A2(n186), .ZN(n188) );
  MUX2_X1 U253 ( .A(n344), .B(n188), .S(n336), .Z(n368) );
  NAND2_X1 U254 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U255 ( .A(n345), .B(n191), .S(n291), .Z(n370) );
  FA_X1 U256 ( .A(n194), .B(n193), .CI(n192), .CO(n100), .S(n263) );
  OAI22_X1 U257 ( .A1(n114), .A2(n197), .B1(n196), .B2(n195), .ZN(n213) );
  OAI22_X1 U258 ( .A1(n14), .A2(n199), .B1(n18), .B2(n198), .ZN(n212) );
  HA_X1 U259 ( .A(n201), .B(n200), .CO(n211), .S(n222) );
  INV_X1 U260 ( .A(n202), .ZN(n204) );
  XNOR2_X1 U261 ( .A(n204), .B(n203), .ZN(n261) );
  FA_X1 U262 ( .A(n207), .B(n206), .CI(n205), .CO(n203), .S(n220) );
  FA_X1 U263 ( .A(n210), .B(n209), .CI(n208), .CO(n219), .S(n221) );
  FA_X1 U264 ( .A(n213), .B(n212), .CI(n211), .CO(n262), .S(n218) );
  NOR2_X1 U265 ( .A1(n216), .A2(n215), .ZN(n214) );
  MUX2_X1 U266 ( .A(n348), .B(n214), .S(n336), .Z(n376) );
  NAND2_X1 U267 ( .A1(n216), .A2(n215), .ZN(n217) );
  MUX2_X1 U268 ( .A(n349), .B(n217), .S(n291), .Z(n378) );
  FA_X1 U269 ( .A(n223), .B(n222), .CI(n221), .CO(n225), .S(n229) );
  NOR2_X1 U270 ( .A1(n226), .A2(n225), .ZN(n224) );
  MUX2_X1 U271 ( .A(n350), .B(n224), .S(n291), .Z(n380) );
  NAND2_X1 U272 ( .A1(n226), .A2(n225), .ZN(n227) );
  MUX2_X1 U273 ( .A(n351), .B(n227), .S(n336), .Z(n382) );
  NAND2_X1 U274 ( .A1(n229), .A2(n228), .ZN(n230) );
  MUX2_X1 U275 ( .A(n352), .B(n230), .S(n288), .Z(n384) );
  FA_X1 U276 ( .A(n233), .B(n232), .CI(n231), .CO(n228), .S(n244) );
  NOR2_X1 U277 ( .A1(n244), .A2(n243), .ZN(n242) );
  MUX2_X1 U278 ( .A(n353), .B(n242), .S(n291), .Z(n386) );
  NAND2_X1 U279 ( .A1(n244), .A2(n243), .ZN(n245) );
  MUX2_X1 U280 ( .A(n354), .B(n245), .S(n336), .Z(n388) );
  NAND2_X1 U281 ( .A1(n247), .A2(n246), .ZN(n248) );
  MUX2_X1 U282 ( .A(n355), .B(n248), .S(n291), .Z(n390) );
  NAND2_X1 U283 ( .A1(n250), .A2(n16), .ZN(n251) );
  MUX2_X1 U284 ( .A(n356), .B(n251), .S(n336), .Z(n392) );
  INV_X1 U285 ( .A(n252), .ZN(n253) );
  AOI21_X1 U286 ( .B1(n255), .B2(n254), .A(n253), .ZN(n256) );
  MUX2_X1 U287 ( .A(n357), .B(n256), .S(n291), .Z(n394) );
  MUX2_X1 U288 ( .A(n358), .B(n260), .S(n336), .Z(n396) );
  FA_X1 U289 ( .A(n263), .B(n262), .CI(n261), .CO(n264), .S(n216) );
  MUX2_X1 U290 ( .A(n359), .B(n264), .S(n291), .Z(n398) );
  BUF_X2 U291 ( .A(rst_n), .Z(n409) );
  MUX2_X1 U292 ( .A(product[0]), .B(n521), .S(n288), .Z(n411) );
  MUX2_X1 U293 ( .A(n521), .B(n522), .S(n291), .Z(n413) );
  AND2_X1 U294 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n265) );
  MUX2_X1 U295 ( .A(n522), .B(n265), .S(n288), .Z(n415) );
  MUX2_X1 U296 ( .A(product[1]), .B(n524), .S(n291), .Z(n417) );
  MUX2_X1 U297 ( .A(n524), .B(n525), .S(n288), .Z(n419) );
  OR2_X1 U298 ( .A1(n267), .A2(n266), .ZN(n268) );
  AND2_X1 U299 ( .A1(n268), .A2(n273), .ZN(n269) );
  MUX2_X1 U300 ( .A(n525), .B(n269), .S(n291), .Z(n421) );
  MUX2_X1 U301 ( .A(product[2]), .B(n527), .S(n288), .Z(n423) );
  MUX2_X1 U302 ( .A(n527), .B(n528), .S(n291), .Z(n425) );
  INV_X1 U303 ( .A(n270), .ZN(n272) );
  NAND2_X1 U304 ( .A1(n272), .A2(n271), .ZN(n274) );
  XOR2_X1 U305 ( .A(n274), .B(n273), .Z(n275) );
  MUX2_X1 U306 ( .A(n528), .B(n275), .S(n288), .Z(n427) );
  MUX2_X1 U307 ( .A(product[3]), .B(n530), .S(n291), .Z(n429) );
  MUX2_X1 U308 ( .A(n530), .B(n531), .S(n288), .Z(n431) );
  NAND2_X1 U309 ( .A1(n277), .A2(n276), .ZN(n279) );
  XNOR2_X1 U310 ( .A(n279), .B(n278), .ZN(n280) );
  MUX2_X1 U311 ( .A(n531), .B(n280), .S(n291), .Z(n433) );
  MUX2_X1 U312 ( .A(product[4]), .B(n533), .S(n288), .Z(n435) );
  MUX2_X1 U313 ( .A(n533), .B(n534), .S(n291), .Z(n437) );
  INV_X1 U314 ( .A(n281), .ZN(n283) );
  NAND2_X1 U315 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U316 ( .A(n285), .B(n284), .Z(n286) );
  MUX2_X1 U317 ( .A(n534), .B(n286), .S(n288), .Z(n439) );
  MUX2_X1 U318 ( .A(product[5]), .B(n536), .S(n291), .Z(n441) );
  MUX2_X1 U319 ( .A(n536), .B(n537), .S(n288), .Z(n443) );
  MUX2_X1 U320 ( .A(product[6]), .B(n539), .S(n288), .Z(n447) );
  NAND2_X1 U321 ( .A1(n402), .A2(n354), .ZN(n287) );
  XOR2_X1 U322 ( .A(n287), .B(n357), .Z(n289) );
  MUX2_X1 U323 ( .A(n539), .B(n289), .S(n288), .Z(n449) );
  MUX2_X1 U324 ( .A(product[7]), .B(n541), .S(n291), .Z(n451) );
  OAI21_X1 U325 ( .B1(n353), .B2(n357), .A(n354), .ZN(n293) );
  NAND2_X1 U326 ( .A1(n343), .A2(n352), .ZN(n290) );
  XNOR2_X1 U327 ( .A(n293), .B(n290), .ZN(n292) );
  MUX2_X1 U328 ( .A(n541), .B(n292), .S(n291), .Z(n453) );
  MUX2_X1 U329 ( .A(product[8]), .B(n543), .S(n336), .Z(n455) );
  AOI21_X1 U330 ( .B1(n293), .B2(n343), .A(n404), .ZN(n296) );
  NAND2_X1 U331 ( .A1(n405), .A2(n351), .ZN(n294) );
  XOR2_X1 U332 ( .A(n296), .B(n294), .Z(n295) );
  MUX2_X1 U333 ( .A(n543), .B(n295), .S(n336), .Z(n457) );
  MUX2_X1 U334 ( .A(product[9]), .B(n545), .S(n336), .Z(n459) );
  OAI21_X1 U335 ( .B1(n296), .B2(n350), .A(n351), .ZN(n307) );
  INV_X1 U336 ( .A(n307), .ZN(n299) );
  NAND2_X1 U337 ( .A1(n406), .A2(n349), .ZN(n297) );
  XOR2_X1 U338 ( .A(n299), .B(n297), .Z(n298) );
  MUX2_X1 U339 ( .A(n545), .B(n298), .S(n336), .Z(n461) );
  MUX2_X1 U340 ( .A(product[10]), .B(n547), .S(n336), .Z(n463) );
  OAI21_X1 U341 ( .B1(n299), .B2(n348), .A(n349), .ZN(n302) );
  NOR2_X1 U342 ( .A1(n358), .A2(n359), .ZN(n305) );
  INV_X1 U343 ( .A(n305), .ZN(n300) );
  NAND2_X1 U344 ( .A1(n358), .A2(n359), .ZN(n304) );
  NAND2_X1 U345 ( .A1(n300), .A2(n304), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n303) );
  MUX2_X1 U347 ( .A(n547), .B(n303), .S(n336), .Z(n465) );
  MUX2_X1 U348 ( .A(product[11]), .B(n549), .S(n336), .Z(n467) );
  NOR2_X1 U349 ( .A1(n305), .A2(n348), .ZN(n308) );
  OAI21_X1 U350 ( .B1(n305), .B2(n349), .A(n304), .ZN(n306) );
  AOI21_X1 U351 ( .B1(n308), .B2(n307), .A(n306), .ZN(n330) );
  NAND2_X1 U352 ( .A1(n339), .A2(n347), .ZN(n309) );
  XOR2_X1 U353 ( .A(n330), .B(n309), .Z(n310) );
  MUX2_X1 U354 ( .A(n549), .B(n310), .S(n336), .Z(n469) );
  MUX2_X1 U355 ( .A(product[12]), .B(n551), .S(n336), .Z(n471) );
  OAI21_X1 U356 ( .B1(n330), .B2(n346), .A(n347), .ZN(n312) );
  NAND2_X1 U357 ( .A1(n342), .A2(n356), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U359 ( .A(n551), .B(n313), .S(n336), .Z(n473) );
  MUX2_X1 U360 ( .A(product[13]), .B(n553), .S(n336), .Z(n475) );
  NAND2_X1 U361 ( .A1(n339), .A2(n342), .ZN(n315) );
  AOI21_X1 U362 ( .B1(n401), .B2(n342), .A(n407), .ZN(n314) );
  OAI21_X1 U363 ( .B1(n330), .B2(n315), .A(n314), .ZN(n317) );
  NAND2_X1 U364 ( .A1(n341), .A2(n355), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U366 ( .A(n553), .B(n318), .S(n336), .Z(n477) );
  MUX2_X1 U367 ( .A(product[14]), .B(n555), .S(n336), .Z(n479) );
  NAND2_X1 U368 ( .A1(n342), .A2(n341), .ZN(n320) );
  NOR2_X1 U369 ( .A1(n346), .A2(n320), .ZN(n326) );
  INV_X1 U370 ( .A(n326), .ZN(n322) );
  AOI21_X1 U371 ( .B1(n407), .B2(n341), .A(n403), .ZN(n319) );
  OAI21_X1 U372 ( .B1(n320), .B2(n347), .A(n319), .ZN(n327) );
  INV_X1 U373 ( .A(n327), .ZN(n321) );
  OAI21_X1 U374 ( .B1(n330), .B2(n322), .A(n321), .ZN(n324) );
  NAND2_X1 U375 ( .A1(n340), .A2(n345), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  MUX2_X1 U377 ( .A(n555), .B(n325), .S(n336), .Z(n481) );
  MUX2_X1 U378 ( .A(product[15]), .B(n557), .S(n336), .Z(n483) );
  NAND2_X1 U379 ( .A1(n326), .A2(n340), .ZN(n329) );
  AOI21_X1 U380 ( .B1(n327), .B2(n340), .A(n400), .ZN(n328) );
  OAI21_X1 U381 ( .B1(n330), .B2(n329), .A(n328), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n331), .B(n344), .ZN(n332) );
  MUX2_X1 U383 ( .A(n557), .B(n332), .S(n336), .Z(n485) );
  MUX2_X1 U384 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n336), .Z(n487) );
  MUX2_X1 U385 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n336), .Z(n489) );
  MUX2_X1 U386 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n336), .Z(n491) );
  MUX2_X1 U387 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n336), .Z(n493) );
  MUX2_X1 U388 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n336), .Z(n495) );
  MUX2_X1 U389 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n336), .Z(n497) );
  MUX2_X1 U390 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n336), .Z(n499) );
  MUX2_X1 U391 ( .A(n15), .B(B_extended[7]), .S(n336), .Z(n501) );
  MUX2_X1 U392 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n336), .Z(n503) );
  MUX2_X1 U393 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n336), .Z(n505) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n336), .Z(n507) );
  MUX2_X1 U395 ( .A(n333), .B(A_extended[3]), .S(n336), .Z(n509) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n336), .Z(n511) );
  MUX2_X1 U397 ( .A(n334), .B(A_extended[5]), .S(n336), .Z(n513) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n336), .Z(n515) );
  MUX2_X1 U399 ( .A(n335), .B(A_extended[7]), .S(n336), .Z(n517) );
  OR2_X1 U400 ( .A1(n336), .A2(n560), .ZN(n519) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_14 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n9, n10, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n373, n375, n377,
         n379, n381, n383, n385, n387, n389, n391, n393, n395, n397, n399,
         n401, n403, n405, n407, n409, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n422, n424, n426, n428, n430, n432, n434,
         n436, n438, n440, n442, n444, n446, n448, n450, n452, n454, n456,
         n458, n460, n462, n464, n466, n468, n470, n472, n474, n476, n478,
         n480, n482, n484, n486, n488, n490, n492, n494, n496, n498, n500,
         n502, n504, n506, n508, n510, n512, n514, n516, n518, n520, n522,
         n524, n526, n528, n530, n532, n533, n535, n536, n538, n539, n541,
         n542, n544, n545, n547, n548, n550, n552, n554, n556, n558, n560,
         n562, n564, n566, n568, n569, n570, n571, n572;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n530), .CK(clk), .Q(n571), 
        .QN(n32) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n526), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n31) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(rst_n), .SE(n518), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n27) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n29) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n28) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n26) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n25) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n21) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(rst_n), .SE(n496), .CK(clk), .Q(n568)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(rst_n), .SE(n492), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(rst_n), .SE(n490), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(rst_n), .SE(n488), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(rst_n), .SE(n486), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(n562)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(rst_n), .SE(n482), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(rst_n), .SE(n480), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(rst_n), .SE(n478), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(rst_n), .SE(n476), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(rst_n), .SE(n474), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n470), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n468), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n466), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n464), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n462), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n460), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n458), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n456), .CK(clk), .Q(n548), 
        .QN(n35) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n454), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n450), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n448), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n442), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n440), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n438), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n434), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n430), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n428), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n426), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(
        product[0]) );
  SDFF_X2 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n528), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n20) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(rst_n), .SE(n516), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n34) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n572), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n370) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n572), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n369), .QN(n420) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n572), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n368), .QN(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n572), .SE(n403), .CK(
        clk), .Q(n419), .QN(n367) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n572), .SE(n401), .CK(
        clk), .QN(n366) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n572), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n365) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n572), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n364), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n572), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n363), .QN(n415) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n572), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n572), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n361), .QN(n416) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n572), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n360), .QN(n33) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n572), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n359), .QN(n418) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n572), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n358), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n572), .SE(n383), .CK(
        clk), .Q(n417), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n572), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n356), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n572), .SE(n379), .CK(
        clk), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n572), .SE(n377), .CK(
        clk), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n572), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n572), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n572), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n351) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n522), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n350) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n524), .CK(clk), .Q(n570), 
        .QN(n30) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n520), .CK(clk), .Q(n569), 
        .QN(n349) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n23) );
  CLKBUF_X1 U2 ( .A(n10), .Z(n6) );
  BUF_X2 U3 ( .A(n10), .Z(n7) );
  BUF_X2 U4 ( .A(en), .Z(n308) );
  CLKBUF_X2 U5 ( .A(en), .Z(n279) );
  BUF_X1 U6 ( .A(n37), .Z(n10) );
  CLKBUF_X2 U7 ( .A(n15), .Z(n16) );
  BUF_X1 U8 ( .A(\mult_x_1/n281 ), .Z(n9) );
  NAND2_X1 U9 ( .A1(n101), .A2(n100), .ZN(n78) );
  XNOR2_X1 U10 ( .A(n190), .B(n189), .ZN(n89) );
  CLKBUF_X2 U11 ( .A(n569), .Z(n14) );
  XNOR2_X1 U12 ( .A(n110), .B(n109), .ZN(n162) );
  NAND2_X1 U13 ( .A1(n258), .A2(n254), .ZN(n195) );
  NAND2_X1 U14 ( .A1(n46), .A2(n45), .ZN(n266) );
  NAND2_X1 U15 ( .A1(n274), .A2(n367), .ZN(n154) );
  CLKBUF_X1 U16 ( .A(n96), .Z(n12) );
  OAI22_X1 U17 ( .A1(n169), .A2(n168), .B1(n170), .B2(n16), .ZN(n13) );
  NAND2_X1 U18 ( .A1(n32), .A2(\mult_x_1/n310 ), .ZN(n217) );
  XNOR2_X1 U19 ( .A(\mult_x_1/n310 ), .B(n31), .ZN(n74) );
  XNOR2_X1 U20 ( .A(n349), .B(n350), .ZN(n15) );
  XNOR2_X1 U21 ( .A(n349), .B(n350), .ZN(n39) );
  BUF_X1 U22 ( .A(n570), .Z(n347) );
  AOI21_X1 U23 ( .B1(n193), .B2(n192), .A(n191), .ZN(n17) );
  CLKBUF_X1 U24 ( .A(n185), .Z(n18) );
  XNOR2_X1 U25 ( .A(n350), .B(n570), .ZN(n38) );
  AND2_X1 U26 ( .A1(n202), .A2(n201), .ZN(n19) );
  INV_X1 U27 ( .A(rst_n), .ZN(n572) );
  AND2_X1 U28 ( .A1(n138), .A2(n136), .ZN(n22) );
  XOR2_X1 U29 ( .A(\mult_x_1/a[2] ), .B(n569), .Z(n36) );
  XNOR2_X1 U30 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n37) );
  NAND2_X1 U31 ( .A1(n36), .A2(n37), .ZN(n81) );
  BUF_X2 U32 ( .A(n81), .Z(n127) );
  XNOR2_X1 U33 ( .A(n14), .B(\mult_x_1/n286 ), .ZN(n44) );
  XNOR2_X1 U34 ( .A(n14), .B(\mult_x_1/n285 ), .ZN(n126) );
  OAI22_X1 U35 ( .A1(n127), .A2(n44), .B1(n7), .B2(n126), .ZN(n246) );
  BUF_X2 U36 ( .A(\mult_x_1/n313 ), .Z(n111) );
  NAND2_X1 U37 ( .A1(n111), .A2(n5), .ZN(n123) );
  XNOR2_X1 U38 ( .A(n111), .B(\mult_x_1/n284 ), .ZN(n43) );
  XNOR2_X1 U39 ( .A(n111), .B(\mult_x_1/n283 ), .ZN(n122) );
  OAI22_X1 U40 ( .A1(n123), .A2(n43), .B1(n122), .B2(n5), .ZN(n245) );
  NAND2_X1 U41 ( .A1(n38), .A2(n39), .ZN(n84) );
  BUF_X2 U42 ( .A(n84), .Z(n169) );
  OR2_X1 U43 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n41) );
  INV_X1 U44 ( .A(n15), .ZN(n40) );
  OAI22_X1 U45 ( .A1(n169), .A2(n30), .B1(n41), .B2(n16), .ZN(n202) );
  XNOR2_X1 U46 ( .A(n347), .B(\mult_x_1/n288 ), .ZN(n42) );
  XNOR2_X1 U47 ( .A(n347), .B(\mult_x_1/n287 ), .ZN(n204) );
  OAI22_X1 U48 ( .A1(n169), .A2(n42), .B1(n16), .B2(n204), .ZN(n201) );
  XOR2_X1 U49 ( .A(n202), .B(n201), .Z(n244) );
  XNOR2_X1 U50 ( .A(n111), .B(\mult_x_1/n285 ), .ZN(n52) );
  OAI22_X1 U51 ( .A1(n123), .A2(n52), .B1(n43), .B2(n5), .ZN(n49) );
  AND2_X1 U52 ( .A1(\mult_x_1/n288 ), .A2(n40), .ZN(n48) );
  XNOR2_X1 U53 ( .A(n14), .B(\mult_x_1/n287 ), .ZN(n50) );
  OAI22_X1 U54 ( .A1(n127), .A2(n50), .B1(n7), .B2(n44), .ZN(n47) );
  OR2_X1 U55 ( .A1(n46), .A2(n45), .ZN(n269) );
  NAND2_X1 U56 ( .A1(n269), .A2(n266), .ZN(n68) );
  FA_X1 U57 ( .A(n49), .B(n48), .CI(n47), .CO(n45), .S(n66) );
  XNOR2_X1 U58 ( .A(n14), .B(\mult_x_1/n288 ), .ZN(n51) );
  OAI22_X1 U59 ( .A1(n127), .A2(n51), .B1(n7), .B2(n50), .ZN(n54) );
  XNOR2_X1 U60 ( .A(n111), .B(\mult_x_1/n286 ), .ZN(n56) );
  OAI22_X1 U61 ( .A1(n123), .A2(n56), .B1(n52), .B2(n5), .ZN(n53) );
  NOR2_X1 U62 ( .A1(n66), .A2(n65), .ZN(n298) );
  HA_X1 U63 ( .A(n54), .B(n53), .CO(n65), .S(n63) );
  OR2_X1 U64 ( .A1(\mult_x_1/n288 ), .A2(n349), .ZN(n55) );
  OAI22_X1 U65 ( .A1(n127), .A2(n349), .B1(n55), .B2(n7), .ZN(n62) );
  OR2_X1 U66 ( .A1(n63), .A2(n62), .ZN(n294) );
  XNOR2_X1 U67 ( .A(n111), .B(\mult_x_1/n287 ), .ZN(n58) );
  OAI22_X1 U68 ( .A1(n123), .A2(n58), .B1(n56), .B2(n5), .ZN(n61) );
  INV_X1 U69 ( .A(n7), .ZN(n57) );
  AND2_X1 U70 ( .A1(\mult_x_1/n288 ), .A2(n57), .ZN(n60) );
  NOR2_X1 U71 ( .A1(n61), .A2(n60), .ZN(n287) );
  OAI22_X1 U72 ( .A1(n123), .A2(\mult_x_1/n288 ), .B1(n58), .B2(n5), .ZN(n284)
         );
  OR2_X1 U73 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n59) );
  NAND2_X1 U74 ( .A1(n59), .A2(n123), .ZN(n283) );
  NAND2_X1 U75 ( .A1(n284), .A2(n283), .ZN(n290) );
  NAND2_X1 U76 ( .A1(n61), .A2(n60), .ZN(n288) );
  OAI21_X1 U77 ( .B1(n287), .B2(n290), .A(n288), .ZN(n295) );
  NAND2_X1 U78 ( .A1(n63), .A2(n62), .ZN(n293) );
  INV_X1 U79 ( .A(n293), .ZN(n64) );
  AOI21_X1 U80 ( .B1(n294), .B2(n295), .A(n64), .ZN(n301) );
  NAND2_X1 U81 ( .A1(n66), .A2(n65), .ZN(n300) );
  OAI21_X1 U82 ( .B1(n298), .B2(n301), .A(n300), .ZN(n268) );
  INV_X1 U83 ( .A(n268), .ZN(n67) );
  XNOR2_X1 U84 ( .A(n68), .B(n67), .ZN(n70) );
  OR2_X1 U85 ( .A1(n308), .A2(n35), .ZN(n69) );
  OAI21_X1 U86 ( .B1(n70), .B2(n274), .A(n69), .ZN(n456) );
  NAND2_X1 U87 ( .A1(n358), .A2(n274), .ZN(n106) );
  XNOR2_X1 U88 ( .A(n347), .B(\mult_x_1/n284 ), .ZN(n115) );
  XNOR2_X1 U89 ( .A(n570), .B(\mult_x_1/n283 ), .ZN(n85) );
  OAI22_X1 U90 ( .A1(n169), .A2(n115), .B1(n16), .B2(n85), .ZN(n96) );
  XNOR2_X1 U91 ( .A(n14), .B(\mult_x_1/n282 ), .ZN(n113) );
  XNOR2_X1 U92 ( .A(n569), .B(n9), .ZN(n80) );
  OAI22_X1 U93 ( .A1(n81), .A2(n113), .B1(n7), .B2(n80), .ZN(n95) );
  OR2_X2 U94 ( .A1(n96), .A2(n95), .ZN(n101) );
  INV_X1 U95 ( .A(n101), .ZN(n72) );
  NOR2_X1 U96 ( .A1(n24), .A2(n217), .ZN(n100) );
  INV_X1 U97 ( .A(n100), .ZN(n71) );
  NAND2_X1 U98 ( .A1(n72), .A2(n71), .ZN(n77) );
  AND2_X1 U99 ( .A1(n571), .A2(\mult_x_1/n281 ), .ZN(n167) );
  XNOR2_X1 U100 ( .A(n167), .B(n111), .ZN(n91) );
  AOI21_X1 U101 ( .B1(n123), .B2(n5), .A(n91), .ZN(n73) );
  INV_X1 U102 ( .A(n73), .ZN(n149) );
  XNOR2_X1 U103 ( .A(n570), .B(\mult_x_1/a[6] ), .ZN(n75) );
  NAND2_X2 U104 ( .A1(n75), .A2(n74), .ZN(n214) );
  XNOR2_X1 U105 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n92) );
  INV_X1 U106 ( .A(n75), .ZN(n76) );
  INV_X2 U107 ( .A(n76), .ZN(n215) );
  XNOR2_X1 U108 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n87) );
  OAI22_X1 U109 ( .A1(n214), .A2(n92), .B1(n215), .B2(n87), .ZN(n148) );
  NOR2_X1 U110 ( .A1(n25), .A2(n217), .ZN(n147) );
  NAND2_X1 U111 ( .A1(n77), .A2(n102), .ZN(n79) );
  NAND2_X1 U112 ( .A1(n79), .A2(n78), .ZN(n261) );
  XNOR2_X1 U113 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n86) );
  XNOR2_X1 U114 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n173) );
  OAI22_X1 U115 ( .A1(n214), .A2(n86), .B1(n215), .B2(n173), .ZN(n186) );
  XNOR2_X1 U116 ( .A(n167), .B(n569), .ZN(n82) );
  OAI22_X1 U117 ( .A1(n81), .A2(n80), .B1(n82), .B2(n6), .ZN(n185) );
  AOI21_X1 U118 ( .B1(n7), .B2(n127), .A(n82), .ZN(n83) );
  INV_X1 U119 ( .A(n83), .ZN(n184) );
  XNOR2_X1 U120 ( .A(n261), .B(n260), .ZN(n90) );
  INV_X1 U121 ( .A(n185), .ZN(n99) );
  BUF_X1 U122 ( .A(n84), .Z(n205) );
  XNOR2_X1 U123 ( .A(n347), .B(\mult_x_1/n282 ), .ZN(n88) );
  OAI22_X1 U124 ( .A1(n205), .A2(n85), .B1(n16), .B2(n88), .ZN(n98) );
  OAI22_X1 U125 ( .A1(n214), .A2(n87), .B1(n215), .B2(n86), .ZN(n97) );
  NOR2_X1 U126 ( .A1(n26), .A2(n217), .ZN(n190) );
  XNOR2_X1 U127 ( .A(n570), .B(n9), .ZN(n168) );
  OAI22_X1 U128 ( .A1(n205), .A2(n88), .B1(n16), .B2(n168), .ZN(n189) );
  XNOR2_X1 U129 ( .A(n193), .B(n89), .ZN(n259) );
  XNOR2_X1 U130 ( .A(n90), .B(n259), .ZN(n231) );
  XNOR2_X1 U131 ( .A(n111), .B(n9), .ZN(n112) );
  OAI22_X1 U132 ( .A1(n123), .A2(n112), .B1(n91), .B2(n5), .ZN(n107) );
  XNOR2_X1 U133 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n118) );
  OAI22_X1 U134 ( .A1(n214), .A2(n118), .B1(n215), .B2(n92), .ZN(n108) );
  NOR2_X1 U135 ( .A1(n217), .A2(n21), .ZN(n109) );
  OAI21_X1 U136 ( .B1(n107), .B2(n108), .A(n109), .ZN(n94) );
  NAND2_X1 U137 ( .A1(n108), .A2(n107), .ZN(n93) );
  NAND2_X1 U138 ( .A1(n94), .A2(n93), .ZN(n138) );
  XNOR2_X1 U139 ( .A(n12), .B(n95), .ZN(n136) );
  FA_X1 U140 ( .A(n99), .B(n98), .CI(n97), .CO(n193), .S(n135) );
  XNOR2_X1 U141 ( .A(n101), .B(n100), .ZN(n103) );
  XNOR2_X1 U142 ( .A(n103), .B(n102), .ZN(n134) );
  NAND2_X1 U143 ( .A1(n231), .A2(n230), .ZN(n104) );
  NAND2_X1 U144 ( .A1(n104), .A2(n279), .ZN(n105) );
  NAND2_X1 U145 ( .A1(n106), .A2(n105), .ZN(n385) );
  XNOR2_X1 U146 ( .A(n108), .B(n107), .ZN(n110) );
  XNOR2_X1 U147 ( .A(n347), .B(\mult_x_1/n286 ), .ZN(n203) );
  XNOR2_X1 U148 ( .A(n347), .B(\mult_x_1/n285 ), .ZN(n116) );
  OAI22_X1 U149 ( .A1(n169), .A2(n203), .B1(n16), .B2(n116), .ZN(n132) );
  XNOR2_X1 U150 ( .A(n111), .B(\mult_x_1/n282 ), .ZN(n121) );
  OAI22_X1 U151 ( .A1(n123), .A2(n121), .B1(n112), .B2(n5), .ZN(n131) );
  XNOR2_X1 U152 ( .A(n14), .B(\mult_x_1/n284 ), .ZN(n125) );
  XNOR2_X1 U153 ( .A(n14), .B(\mult_x_1/n283 ), .ZN(n114) );
  OAI22_X1 U154 ( .A1(n127), .A2(n125), .B1(n7), .B2(n114), .ZN(n130) );
  OAI22_X1 U155 ( .A1(n127), .A2(n114), .B1(n7), .B2(n113), .ZN(n144) );
  OAI22_X1 U156 ( .A1(n169), .A2(n116), .B1(n16), .B2(n115), .ZN(n143) );
  XNOR2_X1 U157 ( .A(n144), .B(n143), .ZN(n120) );
  OR2_X1 U158 ( .A1(\mult_x_1/n288 ), .A2(n20), .ZN(n117) );
  OAI22_X1 U159 ( .A1(n214), .A2(n20), .B1(n117), .B2(n215), .ZN(n129) );
  XNOR2_X1 U160 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n119) );
  OAI22_X1 U161 ( .A1(n214), .A2(n119), .B1(n215), .B2(n118), .ZN(n128) );
  XNOR2_X1 U162 ( .A(n120), .B(n141), .ZN(n160) );
  OAI22_X1 U163 ( .A1(n123), .A2(n122), .B1(n121), .B2(n5), .ZN(n208) );
  INV_X1 U164 ( .A(n215), .ZN(n124) );
  AND2_X1 U165 ( .A1(\mult_x_1/n288 ), .A2(n124), .ZN(n207) );
  OAI22_X1 U166 ( .A1(n127), .A2(n126), .B1(n7), .B2(n125), .ZN(n206) );
  HA_X1 U167 ( .A(n129), .B(n128), .CO(n141), .S(n199) );
  FA_X1 U168 ( .A(n132), .B(n131), .CI(n130), .CO(n161), .S(n198) );
  NAND2_X1 U169 ( .A1(n237), .A2(n236), .ZN(n133) );
  MUX2_X1 U170 ( .A(n362), .B(n133), .S(n279), .Z(n393) );
  FA_X1 U171 ( .A(n22), .B(n135), .CI(n134), .CO(n230), .S(n272) );
  INV_X1 U172 ( .A(n136), .ZN(n137) );
  XNOR2_X1 U173 ( .A(n138), .B(n137), .ZN(n158) );
  INV_X1 U174 ( .A(n144), .ZN(n140) );
  INV_X1 U175 ( .A(n143), .ZN(n139) );
  NAND2_X1 U176 ( .A1(n140), .A2(n139), .ZN(n142) );
  NAND2_X1 U177 ( .A1(n142), .A2(n141), .ZN(n146) );
  NAND2_X1 U178 ( .A1(n144), .A2(n143), .ZN(n145) );
  NAND2_X1 U179 ( .A1(n146), .A2(n145), .ZN(n156) );
  NAND2_X1 U180 ( .A1(n158), .A2(n156), .ZN(n152) );
  FA_X1 U181 ( .A(n149), .B(n147), .CI(n148), .CO(n102), .S(n157) );
  NAND2_X1 U182 ( .A1(n158), .A2(n157), .ZN(n151) );
  NAND2_X1 U183 ( .A1(n156), .A2(n157), .ZN(n150) );
  NAND3_X1 U184 ( .A1(n152), .A2(n151), .A3(n150), .ZN(n271) );
  INV_X1 U185 ( .A(n271), .ZN(n153) );
  NAND2_X1 U186 ( .A1(n153), .A2(n279), .ZN(n155) );
  OAI21_X1 U187 ( .B1(n272), .B2(n155), .A(n154), .ZN(n403) );
  XNOR2_X1 U188 ( .A(n157), .B(n156), .ZN(n159) );
  XNOR2_X1 U189 ( .A(n159), .B(n158), .ZN(n234) );
  FA_X1 U190 ( .A(n162), .B(n161), .CI(n160), .CO(n233), .S(n237) );
  NAND2_X1 U191 ( .A1(n234), .A2(n233), .ZN(n163) );
  NAND2_X1 U192 ( .A1(n163), .A2(n279), .ZN(n165) );
  OR2_X1 U193 ( .A1(n279), .A2(n33), .ZN(n164) );
  NAND2_X1 U194 ( .A1(n165), .A2(n164), .ZN(n389) );
  NOR2_X1 U215 ( .A1(n27), .A2(n217), .ZN(n212) );
  XNOR2_X1 U216 ( .A(\mult_x_1/n310 ), .B(n9), .ZN(n166) );
  XNOR2_X1 U217 ( .A(n167), .B(\mult_x_1/n310 ), .ZN(n213) );
  OAI22_X1 U218 ( .A1(n214), .A2(n166), .B1(n213), .B2(n215), .ZN(n221) );
  INV_X1 U219 ( .A(n221), .ZN(n211) );
  XNOR2_X1 U220 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n172) );
  OAI22_X1 U221 ( .A1(n214), .A2(n172), .B1(n215), .B2(n166), .ZN(n176) );
  XNOR2_X1 U222 ( .A(n167), .B(n570), .ZN(n170) );
  OAI22_X1 U223 ( .A1(n169), .A2(n168), .B1(n170), .B2(n16), .ZN(n175) );
  AOI21_X1 U224 ( .B1(n16), .B2(n205), .A(n170), .ZN(n171) );
  INV_X1 U225 ( .A(n171), .ZN(n174) );
  INV_X1 U226 ( .A(n175), .ZN(n183) );
  OAI22_X1 U227 ( .A1(n214), .A2(n173), .B1(n215), .B2(n172), .ZN(n182) );
  NOR2_X1 U228 ( .A1(n28), .A2(n217), .ZN(n181) );
  NOR2_X1 U229 ( .A1(n29), .A2(n217), .ZN(n179) );
  FA_X1 U230 ( .A(n176), .B(n13), .CI(n174), .CO(n210), .S(n178) );
  OR2_X1 U231 ( .A1(n228), .A2(n227), .ZN(n177) );
  MUX2_X1 U232 ( .A(n351), .B(n177), .S(n279), .Z(n371) );
  FA_X1 U233 ( .A(n180), .B(n179), .CI(n178), .CO(n227), .S(n252) );
  FA_X1 U234 ( .A(n183), .B(n182), .CI(n181), .CO(n180), .S(n258) );
  FA_X1 U235 ( .A(n186), .B(n18), .CI(n184), .CO(n254), .S(n260) );
  INV_X1 U236 ( .A(n190), .ZN(n188) );
  INV_X1 U237 ( .A(n189), .ZN(n187) );
  NAND2_X1 U238 ( .A1(n188), .A2(n187), .ZN(n192) );
  AND2_X1 U239 ( .A1(n190), .A2(n189), .ZN(n191) );
  AOI21_X1 U240 ( .B1(n193), .B2(n192), .A(n191), .ZN(n256) );
  INV_X1 U241 ( .A(n17), .ZN(n194) );
  OAI21_X1 U242 ( .B1(n258), .B2(n254), .A(n194), .ZN(n196) );
  NAND2_X1 U243 ( .A1(n196), .A2(n195), .ZN(n251) );
  OR2_X1 U244 ( .A1(n252), .A2(n251), .ZN(n197) );
  MUX2_X1 U245 ( .A(n352), .B(n197), .S(n279), .Z(n373) );
  FA_X1 U246 ( .A(n200), .B(n199), .CI(n198), .CO(n236), .S(n240) );
  OAI22_X1 U247 ( .A1(n205), .A2(n204), .B1(n16), .B2(n203), .ZN(n243) );
  FA_X1 U248 ( .A(n208), .B(n207), .CI(n206), .CO(n200), .S(n242) );
  OR2_X1 U249 ( .A1(n240), .A2(n239), .ZN(n209) );
  MUX2_X1 U250 ( .A(n354), .B(n209), .S(n279), .Z(n377) );
  FA_X1 U251 ( .A(n212), .B(n211), .CI(n210), .CO(n223), .S(n228) );
  AOI21_X1 U252 ( .B1(n215), .B2(n214), .A(n213), .ZN(n216) );
  INV_X1 U253 ( .A(n216), .ZN(n219) );
  NOR2_X1 U254 ( .A1(n23), .A2(n217), .ZN(n218) );
  XOR2_X1 U255 ( .A(n219), .B(n218), .Z(n220) );
  XOR2_X1 U256 ( .A(n221), .B(n220), .Z(n222) );
  OR2_X1 U257 ( .A1(n223), .A2(n222), .ZN(n225) );
  NAND2_X1 U258 ( .A1(n223), .A2(n222), .ZN(n224) );
  NAND2_X1 U259 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U260 ( .A(n355), .B(n226), .S(n279), .Z(n379) );
  NAND2_X1 U261 ( .A1(n228), .A2(n227), .ZN(n229) );
  MUX2_X1 U262 ( .A(n356), .B(n229), .S(n279), .Z(n381) );
  NOR2_X1 U263 ( .A1(n231), .A2(n230), .ZN(n232) );
  MUX2_X1 U264 ( .A(n357), .B(n232), .S(n279), .Z(n383) );
  NOR2_X1 U265 ( .A1(n234), .A2(n233), .ZN(n235) );
  MUX2_X1 U266 ( .A(n359), .B(n235), .S(n279), .Z(n387) );
  NOR2_X1 U267 ( .A1(n237), .A2(n236), .ZN(n238) );
  MUX2_X1 U268 ( .A(n361), .B(n238), .S(n279), .Z(n391) );
  NAND2_X1 U269 ( .A1(n240), .A2(n239), .ZN(n241) );
  MUX2_X1 U270 ( .A(n363), .B(n241), .S(n279), .Z(n395) );
  FA_X1 U271 ( .A(n19), .B(n243), .CI(n242), .CO(n239), .S(n249) );
  FA_X1 U272 ( .A(n246), .B(n245), .CI(n244), .CO(n248), .S(n46) );
  NOR2_X1 U273 ( .A1(n249), .A2(n248), .ZN(n247) );
  MUX2_X1 U274 ( .A(n364), .B(n247), .S(n279), .Z(n397) );
  NAND2_X1 U275 ( .A1(n249), .A2(n248), .ZN(n250) );
  MUX2_X1 U276 ( .A(n365), .B(n250), .S(n348), .Z(n399) );
  NAND2_X1 U277 ( .A1(n252), .A2(n251), .ZN(n253) );
  MUX2_X1 U278 ( .A(n368), .B(n253), .S(n348), .Z(n405) );
  INV_X1 U279 ( .A(n254), .ZN(n255) );
  XNOR2_X1 U280 ( .A(n256), .B(n255), .ZN(n257) );
  XNOR2_X1 U281 ( .A(n258), .B(n257), .ZN(n278) );
  NAND2_X1 U282 ( .A1(n259), .A2(n260), .ZN(n264) );
  NAND2_X1 U283 ( .A1(n259), .A2(n261), .ZN(n263) );
  NAND2_X1 U284 ( .A1(n261), .A2(n260), .ZN(n262) );
  NAND3_X1 U285 ( .A1(n264), .A2(n263), .A3(n262), .ZN(n277) );
  NAND2_X1 U286 ( .A1(n278), .A2(n277), .ZN(n265) );
  MUX2_X1 U287 ( .A(n369), .B(n265), .S(n279), .Z(n407) );
  INV_X1 U288 ( .A(n266), .ZN(n267) );
  AOI21_X1 U289 ( .B1(n269), .B2(n268), .A(n267), .ZN(n270) );
  MUX2_X1 U290 ( .A(n370), .B(n270), .S(n348), .Z(n409) );
  NAND2_X1 U291 ( .A1(n272), .A2(n271), .ZN(n273) );
  NAND2_X1 U292 ( .A1(n273), .A2(n348), .ZN(n276) );
  INV_X1 U293 ( .A(n279), .ZN(n274) );
  NAND2_X1 U294 ( .A1(n274), .A2(n366), .ZN(n275) );
  NAND2_X1 U295 ( .A1(n276), .A2(n275), .ZN(n401) );
  OAI21_X1 U296 ( .B1(n277), .B2(n278), .A(n279), .ZN(n281) );
  NAND2_X1 U297 ( .A1(n274), .A2(n353), .ZN(n280) );
  NAND2_X1 U298 ( .A1(n281), .A2(n280), .ZN(n375) );
  MUX2_X1 U299 ( .A(product[0]), .B(n532), .S(n308), .Z(n422) );
  MUX2_X1 U300 ( .A(n532), .B(n533), .S(n308), .Z(n424) );
  AND2_X1 U301 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n282) );
  MUX2_X1 U302 ( .A(n533), .B(n282), .S(n308), .Z(n426) );
  MUX2_X1 U303 ( .A(product[1]), .B(n535), .S(n308), .Z(n428) );
  MUX2_X1 U304 ( .A(n535), .B(n536), .S(n308), .Z(n430) );
  OR2_X1 U305 ( .A1(n284), .A2(n283), .ZN(n285) );
  AND2_X1 U306 ( .A1(n285), .A2(n290), .ZN(n286) );
  MUX2_X1 U307 ( .A(n536), .B(n286), .S(n308), .Z(n432) );
  MUX2_X1 U308 ( .A(product[2]), .B(n538), .S(n308), .Z(n434) );
  MUX2_X1 U309 ( .A(n538), .B(n539), .S(n308), .Z(n436) );
  INV_X1 U310 ( .A(n287), .ZN(n289) );
  NAND2_X1 U311 ( .A1(n289), .A2(n288), .ZN(n291) );
  XOR2_X1 U312 ( .A(n291), .B(n290), .Z(n292) );
  MUX2_X1 U313 ( .A(n539), .B(n292), .S(n308), .Z(n438) );
  MUX2_X1 U314 ( .A(product[3]), .B(n541), .S(n308), .Z(n440) );
  MUX2_X1 U315 ( .A(n541), .B(n542), .S(n308), .Z(n442) );
  NAND2_X1 U316 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U317 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U318 ( .A(n542), .B(n297), .S(n308), .Z(n444) );
  MUX2_X1 U319 ( .A(product[4]), .B(n544), .S(n308), .Z(n446) );
  MUX2_X1 U320 ( .A(n544), .B(n545), .S(n308), .Z(n448) );
  INV_X1 U321 ( .A(n298), .ZN(n299) );
  NAND2_X1 U322 ( .A1(n300), .A2(n299), .ZN(n303) );
  INV_X1 U323 ( .A(n301), .ZN(n302) );
  XNOR2_X1 U324 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U325 ( .A(n545), .B(n304), .S(n308), .Z(n450) );
  MUX2_X1 U326 ( .A(product[5]), .B(n547), .S(n308), .Z(n452) );
  MUX2_X1 U327 ( .A(n547), .B(n548), .S(n308), .Z(n454) );
  MUX2_X1 U328 ( .A(product[6]), .B(n550), .S(n308), .Z(n458) );
  NAND2_X1 U329 ( .A1(n413), .A2(n365), .ZN(n305) );
  XOR2_X1 U330 ( .A(n305), .B(n370), .Z(n306) );
  MUX2_X1 U331 ( .A(n550), .B(n306), .S(n308), .Z(n460) );
  MUX2_X1 U332 ( .A(product[7]), .B(n552), .S(n308), .Z(n462) );
  OAI21_X1 U333 ( .B1(n364), .B2(n370), .A(n365), .ZN(n310) );
  NAND2_X1 U334 ( .A1(n354), .A2(n363), .ZN(n307) );
  XNOR2_X1 U335 ( .A(n310), .B(n307), .ZN(n309) );
  MUX2_X1 U336 ( .A(n552), .B(n309), .S(n308), .Z(n464) );
  BUF_X4 U337 ( .A(en), .Z(n348) );
  MUX2_X1 U338 ( .A(product[8]), .B(n554), .S(n348), .Z(n466) );
  AOI21_X1 U339 ( .B1(n310), .B2(n354), .A(n415), .ZN(n313) );
  NAND2_X1 U340 ( .A1(n416), .A2(n362), .ZN(n311) );
  XOR2_X1 U341 ( .A(n313), .B(n311), .Z(n312) );
  MUX2_X1 U342 ( .A(n554), .B(n312), .S(n348), .Z(n468) );
  MUX2_X1 U343 ( .A(product[9]), .B(n556), .S(n348), .Z(n470) );
  OAI21_X1 U344 ( .B1(n313), .B2(n361), .A(n362), .ZN(n321) );
  INV_X1 U345 ( .A(n321), .ZN(n316) );
  NAND2_X1 U346 ( .A1(n418), .A2(n360), .ZN(n314) );
  XOR2_X1 U347 ( .A(n316), .B(n314), .Z(n315) );
  MUX2_X1 U348 ( .A(n556), .B(n315), .S(n348), .Z(n472) );
  MUX2_X1 U349 ( .A(product[10]), .B(n558), .S(n348), .Z(n474) );
  OAI21_X1 U350 ( .B1(n316), .B2(n359), .A(n360), .ZN(n318) );
  NAND2_X1 U351 ( .A1(n419), .A2(n366), .ZN(n317) );
  XNOR2_X1 U352 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U353 ( .A(n558), .B(n319), .S(n348), .Z(n476) );
  MUX2_X1 U354 ( .A(product[11]), .B(n560), .S(n348), .Z(n478) );
  NOR2_X1 U355 ( .A1(n367), .A2(n359), .ZN(n322) );
  OAI21_X1 U356 ( .B1(n367), .B2(n360), .A(n366), .ZN(n320) );
  AOI21_X1 U357 ( .B1(n322), .B2(n321), .A(n320), .ZN(n344) );
  NAND2_X1 U358 ( .A1(n417), .A2(n358), .ZN(n323) );
  XOR2_X1 U359 ( .A(n344), .B(n323), .Z(n324) );
  MUX2_X1 U360 ( .A(n560), .B(n324), .S(n348), .Z(n480) );
  MUX2_X1 U361 ( .A(product[12]), .B(n562), .S(n348), .Z(n482) );
  OAI21_X1 U362 ( .B1(n344), .B2(n357), .A(n358), .ZN(n326) );
  NAND2_X1 U363 ( .A1(n353), .A2(n369), .ZN(n325) );
  XNOR2_X1 U364 ( .A(n326), .B(n325), .ZN(n327) );
  MUX2_X1 U365 ( .A(n562), .B(n327), .S(n348), .Z(n484) );
  MUX2_X1 U366 ( .A(product[13]), .B(n564), .S(n348), .Z(n486) );
  NAND2_X1 U367 ( .A1(n417), .A2(n353), .ZN(n329) );
  AOI21_X1 U368 ( .B1(n412), .B2(n353), .A(n420), .ZN(n328) );
  OAI21_X1 U369 ( .B1(n344), .B2(n329), .A(n328), .ZN(n331) );
  NAND2_X1 U370 ( .A1(n352), .A2(n368), .ZN(n330) );
  XNOR2_X1 U371 ( .A(n331), .B(n330), .ZN(n332) );
  MUX2_X1 U372 ( .A(n564), .B(n332), .S(n348), .Z(n488) );
  MUX2_X1 U373 ( .A(product[14]), .B(n566), .S(n348), .Z(n490) );
  NAND2_X1 U374 ( .A1(n353), .A2(n352), .ZN(n334) );
  NOR2_X1 U375 ( .A1(n357), .A2(n334), .ZN(n340) );
  INV_X1 U376 ( .A(n340), .ZN(n336) );
  AOI21_X1 U377 ( .B1(n420), .B2(n352), .A(n414), .ZN(n333) );
  OAI21_X1 U378 ( .B1(n334), .B2(n358), .A(n333), .ZN(n341) );
  INV_X1 U379 ( .A(n341), .ZN(n335) );
  OAI21_X1 U380 ( .B1(n344), .B2(n336), .A(n335), .ZN(n338) );
  NAND2_X1 U381 ( .A1(n351), .A2(n356), .ZN(n337) );
  XNOR2_X1 U382 ( .A(n338), .B(n337), .ZN(n339) );
  MUX2_X1 U383 ( .A(n566), .B(n339), .S(n348), .Z(n492) );
  MUX2_X1 U384 ( .A(product[15]), .B(n568), .S(n348), .Z(n494) );
  NAND2_X1 U385 ( .A1(n340), .A2(n351), .ZN(n343) );
  AOI21_X1 U386 ( .B1(n341), .B2(n351), .A(n411), .ZN(n342) );
  OAI21_X1 U387 ( .B1(n344), .B2(n343), .A(n342), .ZN(n345) );
  XNOR2_X1 U388 ( .A(n345), .B(n355), .ZN(n346) );
  MUX2_X1 U389 ( .A(n568), .B(n346), .S(n348), .Z(n496) );
  MUX2_X1 U390 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n348), .Z(n498) );
  MUX2_X1 U391 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n348), .Z(n500) );
  MUX2_X1 U392 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n348), .Z(n502) );
  MUX2_X1 U393 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n348), .Z(n504) );
  MUX2_X1 U394 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n348), .Z(n506) );
  MUX2_X1 U395 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n348), .Z(n508) );
  MUX2_X1 U396 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n348), .Z(n510) );
  MUX2_X1 U397 ( .A(n9), .B(B_extended[7]), .S(n348), .Z(n512) );
  MUX2_X1 U398 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n348), .Z(n514) );
  MUX2_X1 U399 ( .A(n111), .B(A_extended[1]), .S(n348), .Z(n516) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n348), .Z(n518) );
  MUX2_X1 U401 ( .A(n14), .B(A_extended[3]), .S(n348), .Z(n520) );
  MUX2_X1 U402 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n348), .Z(n522) );
  MUX2_X1 U403 ( .A(n347), .B(A_extended[5]), .S(n348), .Z(n524) );
  MUX2_X1 U404 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n348), .Z(n526) );
  MUX2_X1 U405 ( .A(\mult_x_1/n310 ), .B(A_extended[7]), .S(n348), .Z(n528) );
  OR2_X1 U406 ( .A1(n348), .A2(n571), .ZN(n530) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_15 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n352,
         n354, n356, n358, n360, n362, n364, n366, n368, n370, n372, n374,
         n376, n378, n380, n382, n384, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n397, n399, n401, n403, n405, n407, n409,
         n411, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n505, n507, n509, n510, n512, n513, n515, n516,
         n518, n519, n521, n522, n524, n525, n527, n528, n530, n532, n534,
         n536, n538, n540, n542, n544, n546, n547, n548, n549, n550;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n259), .SE(n507), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n395), .SE(n503), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n395), .SE(n499), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n11) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n395), .SE(n495), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n28) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n395), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n395), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n26) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n395), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n259), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n24) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n259), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n23) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n259), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n21) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n259), .SE(n477), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n22) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n259), .SE(n475), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n259), .SE(n473), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n259), .SE(n471), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n259), .SE(n469), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n259), .SE(n467), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n259), .SE(n465), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n259), .SE(n463), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n395), .SE(n461), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n395), .SE(n459), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n395), .SE(n457), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n395), .SE(n455), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n395), .SE(n453), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n395), .SE(n451), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n259), .SE(n449), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n395), .SE(n447), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n395), .SE(n445), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n259), .SE(n443), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n395), .SE(n441), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n259), .SE(n439), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n395), .SE(n437), .CK(clk), .Q(n528), 
        .QN(n331) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n395), .SE(n435), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n395), .SE(n433), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n395), .SE(n431), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n395), .SE(n429), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n259), .SE(n427), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n259), .SE(n425), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n395), .SE(n423), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n395), .SE(n421), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n395), .SE(n419), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n395), .SE(n417), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n395), .SE(n415), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n395), .SE(n413), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n395), .SE(n411), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n395), .SE(n409), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n395), .SE(n407), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n395), .SE(n405), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n395), .SE(n403), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n395), .SE(n401), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n395), .SE(n399), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n395), .SE(n397), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n395), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n30) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n395), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n20) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n395), .SE(n501), .CK(clk), .Q(n547), 
        .QN(n27) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n395), .SE(n505), .CK(clk), .Q(n548), 
        .QN(n18) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n550), .SE(n384), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n550), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n348), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n550), .SE(n380), .CK(
        clk), .Q(n393), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n550), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n346), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n550), .SE(n376), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n550), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n344), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n550), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n550), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n342), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n550), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n550), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n340), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n550), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n339), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n550), .SE(n362), .CK(
        clk), .Q(n392), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n550), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n337), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n550), .SE(n358), .CK(
        clk), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n550), .SE(n356), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n550), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n550), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n550), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n332) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n395), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n19) );
  AOI21_X1 U2 ( .B1(n182), .B2(n181), .A(n61), .ZN(n60) );
  XNOR2_X1 U3 ( .A(n59), .B(n77), .ZN(n182) );
  CLKBUF_X2 U4 ( .A(n260), .Z(n256) );
  OAI21_X1 U5 ( .B1(n50), .B2(n49), .A(n48), .ZN(n79) );
  INV_X2 U6 ( .A(n34), .ZN(n191) );
  BUF_X4 U7 ( .A(\mult_x_1/n313 ), .Z(n113) );
  BUF_X1 U8 ( .A(n67), .Z(n6) );
  INV_X1 U9 ( .A(n7), .ZN(n168) );
  XNOR2_X1 U10 ( .A(n155), .B(n121), .ZN(n126) );
  XNOR2_X1 U11 ( .A(n157), .B(n156), .ZN(n121) );
  XNOR2_X1 U12 ( .A(n227), .B(n196), .ZN(n208) );
  OR2_X1 U13 ( .A1(n126), .A2(n125), .ZN(n249) );
  INV_X1 U14 ( .A(n10), .ZN(n16) );
  CLKBUF_X1 U15 ( .A(n139), .Z(n15) );
  NAND2_X1 U16 ( .A1(n47), .A2(n46), .ZN(n48) );
  NOR2_X1 U17 ( .A1(n47), .A2(n46), .ZN(n49) );
  XNOR2_X1 U18 ( .A(n71), .B(n72), .ZN(n58) );
  NAND2_X1 U19 ( .A1(n159), .A2(n158), .ZN(n220) );
  NAND2_X1 U20 ( .A1(n157), .A2(n156), .ZN(n158) );
  NAND2_X1 U21 ( .A1(n155), .A2(n154), .ZN(n159) );
  OR2_X1 U22 ( .A1(n157), .A2(n156), .ZN(n154) );
  NAND2_X1 U23 ( .A1(n241), .A2(n240), .ZN(n254) );
  NAND2_X1 U24 ( .A1(n239), .A2(n238), .ZN(n240) );
  NAND2_X1 U25 ( .A1(n237), .A2(n236), .ZN(n241) );
  OR2_X1 U26 ( .A1(n239), .A2(n238), .ZN(n236) );
  INV_X1 U27 ( .A(n184), .ZN(n35) );
  NAND2_X1 U28 ( .A1(n231), .A2(n230), .ZN(n243) );
  NAND2_X1 U29 ( .A1(n227), .A2(n226), .ZN(n231) );
  NAND2_X1 U30 ( .A1(n208), .A2(n207), .ZN(n209) );
  INV_X1 U31 ( .A(n249), .ZN(n252) );
  OAI21_X1 U32 ( .B1(n129), .B2(n61), .A(n128), .ZN(n437) );
  OR2_X1 U33 ( .A1(n291), .A2(n331), .ZN(n128) );
  XNOR2_X1 U34 ( .A(n8), .B(n548), .ZN(n7) );
  NAND2_X1 U35 ( .A1(n549), .A2(n548), .ZN(n8) );
  XNOR2_X1 U36 ( .A(n229), .B(n228), .ZN(n196) );
  OR2_X1 U37 ( .A1(n229), .A2(n228), .ZN(n226) );
  NAND2_X1 U38 ( .A1(n229), .A2(n228), .ZN(n230) );
  OR2_X2 U39 ( .A1(n34), .A2(n9), .ZN(n193) );
  XOR2_X1 U40 ( .A(n28), .B(\mult_x_1/n312 ), .Z(n9) );
  XNOR2_X2 U41 ( .A(n11), .B(n20), .ZN(n10) );
  NAND2_X2 U42 ( .A1(n32), .A2(n33), .ZN(n85) );
  XNOR2_X1 U43 ( .A(n136), .B(n113), .ZN(n12) );
  CLKBUF_X1 U44 ( .A(\mult_x_1/n281 ), .Z(n13) );
  OAI22_X1 U45 ( .A1(n193), .A2(n190), .B1(n191), .B2(n37), .ZN(n14) );
  NAND2_X2 U46 ( .A1(n113), .A2(n5), .ZN(n152) );
  AOI21_X1 U47 ( .B1(n284), .B2(n285), .A(n112), .ZN(n17) );
  XNOR2_X1 U48 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n33) );
  OR2_X1 U49 ( .A1(n39), .A2(n14), .ZN(n47) );
  BUF_X2 U50 ( .A(n548), .Z(n330) );
  INV_X1 U51 ( .A(rst_n), .ZN(n550) );
  BUF_X2 U52 ( .A(n547), .Z(n329) );
  XOR2_X1 U53 ( .A(n39), .B(n38), .Z(n29) );
  XNOR2_X1 U54 ( .A(n547), .B(\mult_x_1/a[6] ), .ZN(n115) );
  AND2_X1 U55 ( .A1(\mult_x_1/n288 ), .A2(n7), .ZN(n199) );
  XNOR2_X1 U56 ( .A(n113), .B(n13), .ZN(n150) );
  AND2_X1 U57 ( .A1(n549), .A2(\mult_x_1/n281 ), .ZN(n136) );
  XNOR2_X1 U58 ( .A(n136), .B(n113), .ZN(n40) );
  OAI22_X1 U59 ( .A1(n152), .A2(n150), .B1(n40), .B2(n5), .ZN(n198) );
  XOR2_X1 U60 ( .A(\mult_x_1/a[6] ), .B(n548), .Z(n31) );
  NAND2_X2 U61 ( .A1(n31), .A2(n115), .ZN(n165) );
  XNOR2_X1 U62 ( .A(n330), .B(\mult_x_1/n287 ), .ZN(n146) );
  BUF_X2 U63 ( .A(n115), .Z(n166) );
  XNOR2_X1 U64 ( .A(n330), .B(\mult_x_1/n286 ), .ZN(n43) );
  OAI22_X1 U65 ( .A1(n165), .A2(n146), .B1(n166), .B2(n43), .ZN(n197) );
  XOR2_X1 U66 ( .A(\mult_x_1/a[4] ), .B(n547), .Z(n32) );
  XNOR2_X1 U67 ( .A(n329), .B(\mult_x_1/n284 ), .ZN(n188) );
  XNOR2_X1 U68 ( .A(n329), .B(\mult_x_1/n283 ), .ZN(n36) );
  OAI22_X1 U69 ( .A1(n85), .A2(n188), .B1(n10), .B2(n36), .ZN(n39) );
  XNOR2_X1 U70 ( .A(n28), .B(\mult_x_1/n313 ), .ZN(n34) );
  BUF_X2 U71 ( .A(\mult_x_1/n312 ), .Z(n328) );
  XNOR2_X1 U72 ( .A(n328), .B(\mult_x_1/n282 ), .ZN(n190) );
  XNOR2_X1 U73 ( .A(n328), .B(n13), .ZN(n37) );
  OAI22_X1 U74 ( .A1(n193), .A2(n190), .B1(n191), .B2(n37), .ZN(n38) );
  NOR2_X1 U75 ( .A1(n35), .A2(n29), .ZN(n225) );
  XNOR2_X1 U76 ( .A(n330), .B(\mult_x_1/n285 ), .ZN(n42) );
  XNOR2_X1 U77 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n51) );
  OAI22_X1 U78 ( .A1(n165), .A2(n42), .B1(n166), .B2(n51), .ZN(n56) );
  XNOR2_X1 U79 ( .A(n329), .B(\mult_x_1/n282 ), .ZN(n57) );
  OAI22_X1 U80 ( .A1(n85), .A2(n36), .B1(n10), .B2(n57), .ZN(n55) );
  XNOR2_X1 U81 ( .A(n136), .B(n328), .ZN(n52) );
  OAI22_X1 U82 ( .A1(n52), .A2(n191), .B1(n37), .B2(n193), .ZN(n67) );
  INV_X1 U83 ( .A(n67), .ZN(n54) );
  NOR2_X1 U84 ( .A1(n21), .A2(n168), .ZN(n46) );
  XNOR2_X1 U85 ( .A(n47), .B(n46), .ZN(n44) );
  AOI21_X1 U86 ( .B1(n152), .B2(n5), .A(n12), .ZN(n41) );
  INV_X1 U87 ( .A(n41), .ZN(n187) );
  OAI22_X1 U88 ( .A1(n165), .A2(n43), .B1(n166), .B2(n42), .ZN(n186) );
  NOR2_X1 U89 ( .A1(n22), .A2(n168), .ZN(n185) );
  XNOR2_X1 U90 ( .A(n44), .B(n45), .ZN(n223) );
  INV_X1 U91 ( .A(n45), .ZN(n50) );
  XNOR2_X1 U92 ( .A(n330), .B(\mult_x_1/n283 ), .ZN(n65) );
  OAI22_X1 U93 ( .A1(n165), .A2(n51), .B1(n166), .B2(n65), .ZN(n68) );
  AOI21_X1 U94 ( .B1(n191), .B2(n193), .A(n52), .ZN(n53) );
  INV_X1 U95 ( .A(n53), .ZN(n66) );
  XNOR2_X1 U96 ( .A(n79), .B(n78), .ZN(n59) );
  FA_X1 U97 ( .A(n56), .B(n55), .CI(n54), .CO(n74), .S(n224) );
  NOR2_X1 U98 ( .A1(n23), .A2(n168), .ZN(n71) );
  XNOR2_X1 U99 ( .A(n329), .B(n13), .ZN(n64) );
  OAI22_X1 U100 ( .A1(n85), .A2(n57), .B1(n10), .B2(n64), .ZN(n72) );
  XNOR2_X1 U101 ( .A(n74), .B(n58), .ZN(n77) );
  CLKBUF_X1 U102 ( .A(en), .Z(n260) );
  INV_X1 U103 ( .A(n256), .ZN(n61) );
  INV_X1 U104 ( .A(n60), .ZN(n63) );
  NAND2_X1 U105 ( .A1(n61), .A2(n339), .ZN(n62) );
  NAND2_X1 U106 ( .A1(n63), .A2(n62), .ZN(n364) );
  XNOR2_X1 U107 ( .A(n136), .B(n329), .ZN(n134) );
  OAI22_X1 U108 ( .A1(n85), .A2(n64), .B1(n134), .B2(n10), .ZN(n139) );
  INV_X1 U109 ( .A(n139), .ZN(n132) );
  XNOR2_X1 U110 ( .A(n330), .B(\mult_x_1/n282 ), .ZN(n133) );
  OAI22_X1 U111 ( .A1(n165), .A2(n65), .B1(n166), .B2(n133), .ZN(n131) );
  NOR2_X1 U112 ( .A1(n24), .A2(n168), .ZN(n130) );
  FA_X1 U113 ( .A(n68), .B(n66), .CI(n6), .CO(n238), .S(n78) );
  XNOR2_X1 U114 ( .A(n239), .B(n238), .ZN(n76) );
  INV_X1 U115 ( .A(n72), .ZN(n70) );
  INV_X1 U116 ( .A(n71), .ZN(n69) );
  NAND2_X1 U117 ( .A1(n70), .A2(n69), .ZN(n73) );
  AOI22_X1 U118 ( .A1(n74), .A2(n73), .B1(n72), .B2(n71), .ZN(n75) );
  INV_X1 U119 ( .A(n75), .ZN(n237) );
  XNOR2_X1 U120 ( .A(n76), .B(n237), .ZN(n247) );
  NAND2_X1 U121 ( .A1(n77), .A2(n79), .ZN(n82) );
  NAND2_X1 U122 ( .A1(n77), .A2(n78), .ZN(n81) );
  NAND2_X1 U123 ( .A1(n79), .A2(n78), .ZN(n80) );
  NAND3_X1 U124 ( .A1(n82), .A2(n81), .A3(n80), .ZN(n246) );
  OAI21_X1 U125 ( .B1(n247), .B2(n246), .A(n256), .ZN(n84) );
  NAND2_X1 U126 ( .A1(n61), .A2(n334), .ZN(n83) );
  NAND2_X1 U127 ( .A1(n84), .A2(n83), .ZN(n354) );
  XNOR2_X1 U128 ( .A(n328), .B(\mult_x_1/n286 ), .ZN(n89) );
  XNOR2_X1 U129 ( .A(n328), .B(\mult_x_1/n285 ), .ZN(n117) );
  OAI22_X1 U130 ( .A1(n193), .A2(n89), .B1(n191), .B2(n117), .ZN(n124) );
  XNOR2_X1 U131 ( .A(n113), .B(\mult_x_1/n284 ), .ZN(n88) );
  XNOR2_X1 U132 ( .A(n113), .B(\mult_x_1/n283 ), .ZN(n114) );
  OAI22_X1 U133 ( .A1(n152), .A2(n88), .B1(n114), .B2(n5), .ZN(n123) );
  OR2_X1 U134 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n86) );
  OAI22_X1 U135 ( .A1(n85), .A2(n27), .B1(n86), .B2(n10), .ZN(n119) );
  XNOR2_X1 U136 ( .A(n329), .B(\mult_x_1/n288 ), .ZN(n87) );
  XNOR2_X1 U137 ( .A(n329), .B(\mult_x_1/n287 ), .ZN(n120) );
  OAI22_X1 U138 ( .A1(n85), .A2(n87), .B1(n10), .B2(n120), .ZN(n118) );
  XOR2_X1 U139 ( .A(n119), .B(n118), .Z(n122) );
  XNOR2_X1 U140 ( .A(n113), .B(\mult_x_1/n285 ), .ZN(n95) );
  OAI22_X1 U141 ( .A1(n152), .A2(n95), .B1(n88), .B2(n5), .ZN(n92) );
  AND2_X1 U142 ( .A1(\mult_x_1/n288 ), .A2(n16), .ZN(n91) );
  XNOR2_X1 U143 ( .A(n328), .B(\mult_x_1/n287 ), .ZN(n93) );
  OAI22_X1 U144 ( .A1(n193), .A2(n93), .B1(n191), .B2(n89), .ZN(n90) );
  OR2_X1 U145 ( .A1(n111), .A2(n110), .ZN(n284) );
  FA_X1 U146 ( .A(n92), .B(n91), .CI(n90), .CO(n110), .S(n109) );
  XNOR2_X1 U147 ( .A(n328), .B(\mult_x_1/n288 ), .ZN(n94) );
  OAI22_X1 U148 ( .A1(n193), .A2(n94), .B1(n191), .B2(n93), .ZN(n97) );
  XNOR2_X1 U149 ( .A(n113), .B(\mult_x_1/n286 ), .ZN(n99) );
  OAI22_X1 U150 ( .A1(n152), .A2(n99), .B1(n95), .B2(n5), .ZN(n96) );
  NOR2_X1 U151 ( .A1(n109), .A2(n108), .ZN(n277) );
  HA_X1 U152 ( .A(n97), .B(n96), .CO(n108), .S(n106) );
  OR2_X1 U153 ( .A1(\mult_x_1/n288 ), .A2(n20), .ZN(n98) );
  OAI22_X1 U154 ( .A1(n193), .A2(n20), .B1(n98), .B2(n191), .ZN(n105) );
  OR2_X1 U155 ( .A1(n106), .A2(n105), .ZN(n273) );
  XNOR2_X1 U156 ( .A(n113), .B(\mult_x_1/n287 ), .ZN(n101) );
  OAI22_X1 U157 ( .A1(n152), .A2(n101), .B1(n99), .B2(n5), .ZN(n104) );
  INV_X1 U158 ( .A(n191), .ZN(n100) );
  AND2_X1 U159 ( .A1(\mult_x_1/n288 ), .A2(n100), .ZN(n103) );
  NOR2_X1 U160 ( .A1(n104), .A2(n103), .ZN(n266) );
  OAI22_X1 U161 ( .A1(n152), .A2(\mult_x_1/n288 ), .B1(n101), .B2(n5), .ZN(
        n263) );
  OR2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n102) );
  NAND2_X1 U163 ( .A1(n102), .A2(n152), .ZN(n262) );
  NAND2_X1 U164 ( .A1(n263), .A2(n262), .ZN(n269) );
  NAND2_X1 U165 ( .A1(n104), .A2(n103), .ZN(n267) );
  OAI21_X1 U166 ( .B1(n266), .B2(n269), .A(n267), .ZN(n274) );
  NAND2_X1 U167 ( .A1(n106), .A2(n105), .ZN(n272) );
  INV_X1 U168 ( .A(n272), .ZN(n107) );
  AOI21_X1 U169 ( .B1(n273), .B2(n274), .A(n107), .ZN(n280) );
  NAND2_X1 U170 ( .A1(n109), .A2(n108), .ZN(n278) );
  OAI21_X1 U171 ( .B1(n277), .B2(n280), .A(n278), .ZN(n285) );
  NAND2_X1 U172 ( .A1(n111), .A2(n110), .ZN(n283) );
  INV_X1 U173 ( .A(n283), .ZN(n112) );
  AOI21_X1 U174 ( .B1(n284), .B2(n285), .A(n112), .ZN(n251) );
  XNOR2_X1 U175 ( .A(n113), .B(\mult_x_1/n282 ), .ZN(n151) );
  OAI22_X1 U176 ( .A1(n152), .A2(n114), .B1(n151), .B2(n5), .ZN(n144) );
  INV_X1 U177 ( .A(n166), .ZN(n116) );
  AND2_X1 U178 ( .A1(\mult_x_1/n288 ), .A2(n116), .ZN(n143) );
  XNOR2_X1 U179 ( .A(n328), .B(\mult_x_1/n284 ), .ZN(n153) );
  OAI22_X1 U180 ( .A1(n193), .A2(n117), .B1(n191), .B2(n153), .ZN(n142) );
  AND2_X1 U181 ( .A1(n119), .A2(n118), .ZN(n157) );
  XNOR2_X1 U182 ( .A(n329), .B(\mult_x_1/n286 ), .ZN(n148) );
  OAI22_X1 U183 ( .A1(n85), .A2(n120), .B1(n10), .B2(n148), .ZN(n156) );
  FA_X1 U184 ( .A(n124), .B(n123), .CI(n122), .CO(n125), .S(n111) );
  NAND2_X1 U185 ( .A1(n126), .A2(n125), .ZN(n250) );
  NAND2_X1 U186 ( .A1(n249), .A2(n250), .ZN(n127) );
  XNOR2_X1 U187 ( .A(n251), .B(n127), .ZN(n129) );
  BUF_X2 U188 ( .A(n260), .Z(n291) );
  FA_X1 U207 ( .A(n132), .B(n131), .CI(n130), .CO(n235), .S(n239) );
  NOR2_X1 U208 ( .A1(n25), .A2(n168), .ZN(n234) );
  XNOR2_X1 U209 ( .A(n330), .B(n13), .ZN(n137) );
  OAI22_X1 U210 ( .A1(n165), .A2(n133), .B1(n166), .B2(n137), .ZN(n140) );
  AOI21_X1 U211 ( .B1(n10), .B2(n85), .A(n134), .ZN(n135) );
  INV_X1 U212 ( .A(n135), .ZN(n138) );
  NOR2_X1 U213 ( .A1(n26), .A2(n168), .ZN(n163) );
  XNOR2_X1 U214 ( .A(n136), .B(n330), .ZN(n164) );
  OAI22_X1 U215 ( .A1(n165), .A2(n137), .B1(n164), .B2(n166), .ZN(n172) );
  INV_X1 U216 ( .A(n172), .ZN(n162) );
  FA_X1 U217 ( .A(n140), .B(n15), .CI(n138), .CO(n161), .S(n233) );
  OR2_X1 U218 ( .A1(n178), .A2(n179), .ZN(n141) );
  MUX2_X1 U219 ( .A(n332), .B(n141), .S(n256), .Z(n350) );
  FA_X1 U220 ( .A(n144), .B(n143), .CI(n142), .CO(n215), .S(n155) );
  OR2_X1 U221 ( .A1(\mult_x_1/n288 ), .A2(n18), .ZN(n145) );
  OAI22_X1 U222 ( .A1(n165), .A2(n18), .B1(n145), .B2(n166), .ZN(n195) );
  XNOR2_X1 U223 ( .A(n330), .B(\mult_x_1/n288 ), .ZN(n147) );
  OAI22_X1 U224 ( .A1(n165), .A2(n147), .B1(n166), .B2(n146), .ZN(n194) );
  XNOR2_X1 U225 ( .A(n329), .B(\mult_x_1/n285 ), .ZN(n189) );
  OAI22_X1 U226 ( .A1(n85), .A2(n148), .B1(n10), .B2(n189), .ZN(n202) );
  OAI22_X1 U227 ( .A1(n152), .A2(n151), .B1(n150), .B2(n5), .ZN(n201) );
  XNOR2_X1 U228 ( .A(n328), .B(\mult_x_1/n283 ), .ZN(n192) );
  OAI22_X1 U229 ( .A1(n193), .A2(n153), .B1(n191), .B2(n192), .ZN(n200) );
  OR2_X1 U230 ( .A1(n221), .A2(n220), .ZN(n160) );
  MUX2_X1 U231 ( .A(n335), .B(n160), .S(n256), .Z(n356) );
  FA_X1 U232 ( .A(n163), .B(n162), .CI(n161), .CO(n174), .S(n179) );
  AOI21_X1 U233 ( .B1(n166), .B2(n165), .A(n164), .ZN(n167) );
  INV_X1 U234 ( .A(n167), .ZN(n170) );
  NOR2_X1 U235 ( .A1(n19), .A2(n168), .ZN(n169) );
  XOR2_X1 U236 ( .A(n170), .B(n169), .Z(n171) );
  XOR2_X1 U237 ( .A(n172), .B(n171), .Z(n173) );
  OR2_X1 U238 ( .A1(n174), .A2(n173), .ZN(n176) );
  NAND2_X1 U239 ( .A1(n174), .A2(n173), .ZN(n175) );
  NAND2_X1 U240 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U241 ( .A(n336), .B(n177), .S(n256), .Z(n358) );
  NAND2_X1 U242 ( .A1(n179), .A2(n178), .ZN(n180) );
  MUX2_X1 U243 ( .A(n337), .B(n180), .S(n256), .Z(n360) );
  NOR2_X1 U244 ( .A1(n182), .A2(n181), .ZN(n183) );
  MUX2_X1 U245 ( .A(n338), .B(n183), .S(n256), .Z(n362) );
  XNOR2_X1 U246 ( .A(n184), .B(n29), .ZN(n227) );
  FA_X1 U247 ( .A(n187), .B(n186), .CI(n185), .CO(n45), .S(n229) );
  OAI22_X1 U248 ( .A1(n85), .A2(n189), .B1(n10), .B2(n188), .ZN(n205) );
  OAI22_X1 U249 ( .A1(n193), .A2(n192), .B1(n191), .B2(n190), .ZN(n204) );
  HA_X1 U250 ( .A(n195), .B(n194), .CO(n203), .S(n214) );
  FA_X1 U251 ( .A(n199), .B(n198), .CI(n197), .CO(n184), .S(n212) );
  FA_X1 U252 ( .A(n202), .B(n201), .CI(n200), .CO(n211), .S(n213) );
  FA_X1 U253 ( .A(n205), .B(n204), .CI(n203), .CO(n228), .S(n210) );
  NOR2_X1 U254 ( .A1(n208), .A2(n207), .ZN(n206) );
  MUX2_X1 U255 ( .A(n340), .B(n206), .S(n256), .Z(n366) );
  MUX2_X1 U256 ( .A(n341), .B(n209), .S(n256), .Z(n368) );
  FA_X1 U257 ( .A(n212), .B(n211), .CI(n210), .CO(n207), .S(n218) );
  FA_X1 U258 ( .A(n215), .B(n214), .CI(n213), .CO(n217), .S(n221) );
  NOR2_X1 U259 ( .A1(n218), .A2(n217), .ZN(n216) );
  MUX2_X1 U260 ( .A(n342), .B(n216), .S(n256), .Z(n370) );
  NAND2_X1 U261 ( .A1(n218), .A2(n217), .ZN(n219) );
  MUX2_X1 U262 ( .A(n343), .B(n219), .S(n256), .Z(n372) );
  NAND2_X1 U263 ( .A1(n221), .A2(n220), .ZN(n222) );
  MUX2_X1 U264 ( .A(n344), .B(n222), .S(n288), .Z(n374) );
  FA_X1 U265 ( .A(n225), .B(n224), .CI(n223), .CO(n181), .S(n244) );
  NAND2_X1 U266 ( .A1(n244), .A2(n243), .ZN(n232) );
  MUX2_X1 U267 ( .A(n345), .B(n232), .S(n291), .Z(n376) );
  FA_X1 U268 ( .A(n235), .B(n234), .CI(n233), .CO(n178), .S(n255) );
  NAND2_X1 U269 ( .A1(n255), .A2(n254), .ZN(n242) );
  MUX2_X1 U270 ( .A(n346), .B(n242), .S(n288), .Z(n378) );
  NOR2_X1 U271 ( .A1(n244), .A2(n243), .ZN(n245) );
  MUX2_X1 U272 ( .A(n347), .B(n245), .S(n291), .Z(n380) );
  NAND2_X1 U273 ( .A1(n247), .A2(n246), .ZN(n248) );
  MUX2_X1 U274 ( .A(n348), .B(n248), .S(n288), .Z(n382) );
  OAI21_X1 U275 ( .B1(n252), .B2(n17), .A(n250), .ZN(n253) );
  MUX2_X1 U276 ( .A(n349), .B(n253), .S(n291), .Z(n384) );
  OAI21_X1 U277 ( .B1(n255), .B2(n254), .A(n256), .ZN(n258) );
  NAND2_X1 U278 ( .A1(n61), .A2(n333), .ZN(n257) );
  NAND2_X1 U279 ( .A1(n258), .A2(n257), .ZN(n352) );
  BUF_X2 U280 ( .A(rst_n), .Z(n395) );
  BUF_X1 U281 ( .A(rst_n), .Z(n259) );
  MUX2_X1 U282 ( .A(product[0]), .B(n509), .S(n291), .Z(n397) );
  BUF_X2 U283 ( .A(n260), .Z(n288) );
  MUX2_X1 U284 ( .A(n509), .B(n510), .S(n288), .Z(n399) );
  AND2_X1 U285 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n261) );
  MUX2_X1 U286 ( .A(n510), .B(n261), .S(n291), .Z(n401) );
  MUX2_X1 U287 ( .A(product[1]), .B(n512), .S(n288), .Z(n403) );
  MUX2_X1 U288 ( .A(n512), .B(n513), .S(n291), .Z(n405) );
  OR2_X1 U289 ( .A1(n263), .A2(n262), .ZN(n264) );
  AND2_X1 U290 ( .A1(n264), .A2(n269), .ZN(n265) );
  MUX2_X1 U291 ( .A(n513), .B(n265), .S(n288), .Z(n407) );
  MUX2_X1 U292 ( .A(product[2]), .B(n515), .S(n288), .Z(n409) );
  MUX2_X1 U293 ( .A(n515), .B(n516), .S(n291), .Z(n411) );
  INV_X1 U294 ( .A(n266), .ZN(n268) );
  NAND2_X1 U295 ( .A1(n268), .A2(n267), .ZN(n270) );
  XOR2_X1 U296 ( .A(n270), .B(n269), .Z(n271) );
  MUX2_X1 U297 ( .A(n516), .B(n271), .S(n288), .Z(n413) );
  MUX2_X1 U298 ( .A(product[3]), .B(n518), .S(n288), .Z(n415) );
  MUX2_X1 U299 ( .A(n518), .B(n519), .S(n291), .Z(n417) );
  NAND2_X1 U300 ( .A1(n273), .A2(n272), .ZN(n275) );
  XNOR2_X1 U301 ( .A(n275), .B(n274), .ZN(n276) );
  MUX2_X1 U302 ( .A(n519), .B(n276), .S(n288), .Z(n419) );
  MUX2_X1 U303 ( .A(product[4]), .B(n521), .S(n288), .Z(n421) );
  MUX2_X1 U304 ( .A(n521), .B(n522), .S(n291), .Z(n423) );
  INV_X1 U305 ( .A(n277), .ZN(n279) );
  NAND2_X1 U306 ( .A1(n279), .A2(n278), .ZN(n281) );
  XOR2_X1 U307 ( .A(n281), .B(n280), .Z(n282) );
  MUX2_X1 U308 ( .A(n522), .B(n282), .S(n288), .Z(n425) );
  MUX2_X1 U309 ( .A(product[5]), .B(n524), .S(n288), .Z(n427) );
  MUX2_X1 U310 ( .A(n524), .B(n525), .S(n291), .Z(n429) );
  NAND2_X1 U311 ( .A1(n284), .A2(n283), .ZN(n286) );
  XNOR2_X1 U312 ( .A(n286), .B(n285), .ZN(n287) );
  MUX2_X1 U313 ( .A(n525), .B(n287), .S(n288), .Z(n431) );
  MUX2_X1 U314 ( .A(product[6]), .B(n527), .S(n291), .Z(n433) );
  MUX2_X1 U315 ( .A(n527), .B(n528), .S(n288), .Z(n435) );
  MUX2_X1 U316 ( .A(product[7]), .B(n530), .S(n291), .Z(n439) );
  NAND2_X1 U317 ( .A1(n335), .A2(n344), .ZN(n289) );
  XNOR2_X1 U318 ( .A(n349), .B(n289), .ZN(n290) );
  MUX2_X1 U319 ( .A(n530), .B(n290), .S(n291), .Z(n441) );
  MUX2_X1 U320 ( .A(product[8]), .B(n532), .S(n291), .Z(n443) );
  AOI21_X1 U321 ( .B1(n349), .B2(n335), .A(n389), .ZN(n294) );
  NAND2_X1 U322 ( .A1(n390), .A2(n343), .ZN(n292) );
  XOR2_X1 U323 ( .A(n294), .B(n292), .Z(n293) );
  MUX2_X1 U324 ( .A(n532), .B(n293), .S(n288), .Z(n445) );
  MUX2_X1 U325 ( .A(product[9]), .B(n534), .S(n288), .Z(n447) );
  OAI21_X1 U326 ( .B1(n294), .B2(n342), .A(n343), .ZN(n302) );
  INV_X1 U327 ( .A(n302), .ZN(n297) );
  NAND2_X1 U328 ( .A1(n391), .A2(n341), .ZN(n295) );
  XOR2_X1 U329 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U330 ( .A(n534), .B(n296), .S(n291), .Z(n449) );
  MUX2_X1 U331 ( .A(product[10]), .B(n536), .S(n288), .Z(n451) );
  OAI21_X1 U332 ( .B1(n297), .B2(n340), .A(n341), .ZN(n299) );
  NAND2_X1 U333 ( .A1(n393), .A2(n345), .ZN(n298) );
  XNOR2_X1 U334 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U335 ( .A(n536), .B(n300), .S(n291), .Z(n453) );
  MUX2_X1 U336 ( .A(product[11]), .B(n538), .S(n291), .Z(n455) );
  NOR2_X1 U337 ( .A1(n347), .A2(n340), .ZN(n303) );
  OAI21_X1 U338 ( .B1(n347), .B2(n341), .A(n345), .ZN(n301) );
  AOI21_X1 U339 ( .B1(n303), .B2(n302), .A(n301), .ZN(n325) );
  NAND2_X1 U340 ( .A1(n392), .A2(n339), .ZN(n304) );
  XOR2_X1 U341 ( .A(n325), .B(n304), .Z(n305) );
  MUX2_X1 U342 ( .A(n538), .B(n305), .S(n288), .Z(n457) );
  MUX2_X1 U343 ( .A(product[12]), .B(n540), .S(n291), .Z(n459) );
  OAI21_X1 U344 ( .B1(n325), .B2(n338), .A(n339), .ZN(n307) );
  NAND2_X1 U345 ( .A1(n334), .A2(n348), .ZN(n306) );
  XNOR2_X1 U346 ( .A(n307), .B(n306), .ZN(n308) );
  MUX2_X1 U347 ( .A(n540), .B(n308), .S(n288), .Z(n461) );
  MUX2_X1 U348 ( .A(product[13]), .B(n542), .S(n291), .Z(n463) );
  NAND2_X1 U349 ( .A1(n392), .A2(n334), .ZN(n310) );
  AOI21_X1 U350 ( .B1(n388), .B2(n334), .A(n394), .ZN(n309) );
  OAI21_X1 U351 ( .B1(n325), .B2(n310), .A(n309), .ZN(n312) );
  NAND2_X1 U352 ( .A1(n333), .A2(n346), .ZN(n311) );
  XNOR2_X1 U353 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U354 ( .A(n542), .B(n313), .S(n291), .Z(n465) );
  MUX2_X1 U355 ( .A(product[14]), .B(n544), .S(n288), .Z(n467) );
  NAND2_X1 U356 ( .A1(n334), .A2(n333), .ZN(n315) );
  NOR2_X1 U357 ( .A1(n338), .A2(n315), .ZN(n321) );
  INV_X1 U358 ( .A(n321), .ZN(n317) );
  AOI21_X1 U359 ( .B1(n394), .B2(n333), .A(n387), .ZN(n314) );
  OAI21_X1 U360 ( .B1(n315), .B2(n339), .A(n314), .ZN(n322) );
  INV_X1 U361 ( .A(n322), .ZN(n316) );
  OAI21_X1 U362 ( .B1(n325), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U363 ( .A1(n332), .A2(n337), .ZN(n318) );
  XNOR2_X1 U364 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U365 ( .A(n544), .B(n320), .S(n291), .Z(n469) );
  MUX2_X1 U366 ( .A(product[15]), .B(n546), .S(n288), .Z(n471) );
  NAND2_X1 U367 ( .A1(n321), .A2(n332), .ZN(n324) );
  AOI21_X1 U368 ( .B1(n322), .B2(n332), .A(n386), .ZN(n323) );
  OAI21_X1 U369 ( .B1(n325), .B2(n324), .A(n323), .ZN(n326) );
  XNOR2_X1 U370 ( .A(n326), .B(n336), .ZN(n327) );
  MUX2_X1 U371 ( .A(n546), .B(n327), .S(n291), .Z(n473) );
  MUX2_X1 U372 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n288), .Z(n475) );
  MUX2_X1 U373 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n291), .Z(n477) );
  MUX2_X1 U374 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n288), .Z(n479) );
  MUX2_X1 U375 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n291), .Z(n481) );
  MUX2_X1 U376 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n288), .Z(n483) );
  MUX2_X1 U377 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n291), .Z(n485) );
  MUX2_X1 U378 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n288), .Z(n487) );
  MUX2_X1 U379 ( .A(n13), .B(B_extended[7]), .S(n291), .Z(n489) );
  MUX2_X1 U380 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n288), .Z(n491) );
  MUX2_X1 U381 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n291), .Z(n493) );
  MUX2_X1 U382 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n288), .Z(n495) );
  MUX2_X1 U383 ( .A(n328), .B(A_extended[3]), .S(n291), .Z(n497) );
  MUX2_X1 U384 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n288), .Z(n499) );
  MUX2_X1 U385 ( .A(n329), .B(A_extended[5]), .S(n291), .Z(n501) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n288), .Z(n503) );
  MUX2_X1 U387 ( .A(n330), .B(A_extended[7]), .S(n291), .Z(n505) );
  OR2_X1 U388 ( .A1(n288), .A2(n549), .ZN(n507) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_16 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n385, n387, n389, n391, n393, n395, n397, n399, n401, n403, n405,
         n407, n409, n411, n413, n415, n417, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n429, n431, n433, n435, n437, n439, n441,
         n443, n445, n447, n449, n451, n453, n455, n457, n459, n461, n463,
         n465, n467, n469, n471, n473, n475, n477, n479, n481, n483, n485,
         n487, n489, n491, n493, n495, n497, n499, n501, n503, n505, n507,
         n509, n511, n513, n515, n517, n519, n521, n523, n525, n527, n529,
         n531, n533, n535, n537, n539, n541, n542, n544, n545, n547, n548,
         n550, n551, n553, n554, n556, n557, n559, n560, n562, n564, n566,
         n568, n570, n572, n574, n576, n578, n579, n580, n581, n582;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n291), .SE(n539), .CK(clk), .Q(n581), 
        .QN(n27) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n427), .SE(n535), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n39) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n427), .SE(n533), .CK(clk), .Q(n580), 
        .QN(n31) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n427), .SE(n531), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n24) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n427), .SE(n529), .CK(clk), .Q(n579), 
        .QN(n29) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n427), .SE(n527), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n10) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n427), .SE(n523), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n9) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n427), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n30) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n427), .SE(n519), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n37) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n427), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n36) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n291), .SE(n515), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n35) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n291), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n34) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n291), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n33) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n291), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n32) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n291), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n291), .SE(n505), .CK(clk), .Q(n578)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n291), .SE(n503), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n291), .SE(n501), .CK(clk), .Q(n576)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n291), .SE(n499), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n291), .SE(n497), .CK(clk), .Q(n574)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n291), .SE(n495), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n427), .SE(n493), .CK(clk), .Q(n572)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n427), .SE(n491), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n427), .SE(n489), .CK(clk), .Q(n570)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n427), .SE(n487), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n427), .SE(n485), .CK(clk), .Q(n568)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n427), .SE(n483), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n291), .SE(n481), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n427), .SE(n479), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n427), .SE(n477), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n291), .SE(n475), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n427), .SE(n473), .CK(clk), .Q(n562)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n427), .SE(n471), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n427), .SE(n469), .CK(clk), .Q(n560), 
        .QN(n364) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n291), .SE(n467), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n427), .SE(n465), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n427), .SE(n463), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n291), .SE(n461), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n427), .SE(n459), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n427), .SE(n457), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n427), .SE(n455), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n291), .SE(n453), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n427), .SE(n451), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n427), .SE(n449), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n427), .SE(n447), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n427), .SE(n445), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n427), .SE(n443), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n427), .SE(n441), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n427), .SE(n439), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n427), .SE(n437), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n427), .SE(n435), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n427), .SE(n433), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n427), .SE(n431), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n427), .SE(n429), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n427), .SE(n525), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n42) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n582), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n382) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n582), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n381) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n582), .SE(n413), .CK(
        clk), .QN(n380) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n582), .SI(1'b1), .SE(n411), .CK(clk), 
        .Q(n379), .QN(n421) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n582), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n378), .QN(n426) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n582), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n377), .QN(n422) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n582), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n376) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n582), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n375), .QN(n423) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n582), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n374), .QN(n41) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n582), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n373), .QN(n425) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n582), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n372), .QN(n420) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n582), .SE(n395), .CK(
        clk), .Q(n424), .QN(n371) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n582), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n370), .QN(n419) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n582), .SE(n391), .CK(
        clk), .QN(n369) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n582), .SE(n389), .CK(
        clk), .QN(n368) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n582), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n367) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n582), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n366) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n582), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n365) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n427), .SE(n537), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n28) );
  BUF_X1 U2 ( .A(n267), .Z(n22) );
  AOI21_X1 U3 ( .B1(n304), .B2(n305), .A(n115), .ZN(n314) );
  NAND2_X1 U4 ( .A1(n7), .A2(n5), .ZN(n413) );
  OR2_X1 U5 ( .A1(n322), .A2(n6), .ZN(n5) );
  INV_X1 U6 ( .A(n380), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n279), .A2(n322), .ZN(n7) );
  XNOR2_X1 U8 ( .A(n89), .B(n88), .ZN(n90) );
  OAI21_X1 U9 ( .B1(n17), .B2(n93), .A(n8), .ZN(n88) );
  OR2_X1 U10 ( .A1(n82), .A2(n9), .ZN(n8) );
  INV_X1 U11 ( .A(en), .ZN(n21) );
  INV_X1 U12 ( .A(n46), .ZN(n148) );
  BUF_X2 U13 ( .A(n45), .Z(n14) );
  INV_X1 U14 ( .A(n10), .ZN(n11) );
  NAND2_X1 U15 ( .A1(n144), .A2(n26), .ZN(n12) );
  NAND2_X1 U16 ( .A1(n144), .A2(n26), .ZN(n13) );
  NAND2_X1 U17 ( .A1(n144), .A2(n26), .ZN(n147) );
  AND2_X2 U18 ( .A1(n581), .A2(\mult_x_1/n281 ), .ZN(n184) );
  MUX2_X1 U19 ( .A(n218), .B(n367), .S(n21), .Z(n387) );
  BUF_X1 U20 ( .A(n45), .Z(n180) );
  NAND2_X1 U21 ( .A1(n45), .A2(n44), .ZN(n15) );
  NAND2_X1 U22 ( .A1(n45), .A2(n44), .ZN(n179) );
  CLKBUF_X1 U23 ( .A(n15), .Z(n16) );
  CLKBUF_X1 U24 ( .A(n109), .Z(n17) );
  NAND2_X1 U25 ( .A1(n108), .A2(n9), .ZN(n109) );
  NAND2_X1 U26 ( .A1(n204), .A2(n203), .ZN(n205) );
  CLKBUF_X1 U27 ( .A(n197), .Z(n20) );
  NAND2_X1 U28 ( .A1(n284), .A2(n283), .ZN(n285) );
  INV_X1 U29 ( .A(n287), .ZN(n284) );
  INV_X1 U30 ( .A(n286), .ZN(n283) );
  NAND2_X1 U31 ( .A1(n161), .A2(n160), .ZN(n139) );
  NAND2_X1 U32 ( .A1(n99), .A2(n98), .ZN(n125) );
  NAND2_X1 U33 ( .A1(n97), .A2(n96), .ZN(n98) );
  NAND2_X1 U34 ( .A1(n118), .A2(n95), .ZN(n99) );
  NAND2_X1 U35 ( .A1(n85), .A2(n84), .ZN(n86) );
  NAND2_X1 U36 ( .A1(n89), .A2(n88), .ZN(n84) );
  NAND2_X1 U37 ( .A1(n91), .A2(n83), .ZN(n85) );
  OR2_X1 U38 ( .A1(n89), .A2(n88), .ZN(n83) );
  NAND2_X1 U39 ( .A1(n223), .A2(n222), .ZN(n260) );
  NAND2_X1 U40 ( .A1(n215), .A2(n213), .ZN(n207) );
  CLKBUF_X1 U41 ( .A(n214), .Z(n18) );
  XNOR2_X1 U42 ( .A(n161), .B(n160), .ZN(n162) );
  NAND2_X1 U43 ( .A1(n167), .A2(n166), .ZN(n168) );
  NAND2_X1 U44 ( .A1(n289), .A2(n288), .ZN(n290) );
  NAND2_X1 U45 ( .A1(n287), .A2(n286), .ZN(n288) );
  NAND2_X1 U46 ( .A1(n38), .A2(n285), .ZN(n289) );
  XNOR2_X1 U47 ( .A(n29), .B(\mult_x_1/a[2] ), .ZN(n144) );
  XOR2_X1 U48 ( .A(n216), .B(n215), .Z(n19) );
  INV_X2 U49 ( .A(n28), .ZN(n23) );
  XNOR2_X1 U50 ( .A(n29), .B(n24), .ZN(n45) );
  OAI22_X1 U51 ( .A1(n13), .A2(n101), .B1(n148), .B2(n92), .ZN(n118) );
  OAI22_X1 U52 ( .A1(n12), .A2(n29), .B1(n148), .B2(n105), .ZN(n113) );
  OAI22_X1 U53 ( .A1(n13), .A2(n81), .B1(n148), .B2(n73), .ZN(n221) );
  OAI22_X1 U54 ( .A1(n13), .A2(n65), .B1(n148), .B2(n51), .ZN(n67) );
  OAI22_X1 U55 ( .A1(n12), .A2(n73), .B1(n148), .B2(n65), .ZN(n226) );
  OAI22_X1 U56 ( .A1(n13), .A2(n92), .B1(n148), .B2(n81), .ZN(n89) );
  AOI21_X1 U57 ( .B1(n148), .B2(n12), .A(n146), .ZN(n149) );
  XOR2_X1 U58 ( .A(n91), .B(n90), .Z(n25) );
  CLKBUF_X1 U59 ( .A(n143), .Z(n26) );
  NAND2_X1 U60 ( .A1(n208), .A2(n207), .ZN(n272) );
  NAND2_X1 U61 ( .A1(n117), .A2(n116), .ZN(n95) );
  INV_X1 U62 ( .A(n116), .ZN(n97) );
  AND2_X1 U63 ( .A1(n121), .A2(n120), .ZN(n122) );
  OAI22_X1 U64 ( .A1(n147), .A2(n102), .B1(n148), .B2(n101), .ZN(n121) );
  OAI21_X1 U65 ( .B1(n221), .B2(n220), .A(n219), .ZN(n223) );
  NAND2_X1 U66 ( .A1(n221), .A2(n220), .ZN(n222) );
  INV_X1 U67 ( .A(rst_n), .ZN(n582) );
  XOR2_X1 U68 ( .A(n156), .B(n155), .Z(n38) );
  AND2_X1 U69 ( .A1(n156), .A2(n155), .ZN(n40) );
  OR2_X1 U70 ( .A1(n166), .A2(n21), .ZN(n43) );
  XOR2_X1 U71 ( .A(\mult_x_1/a[4] ), .B(n580), .Z(n44) );
  CLKBUF_X2 U72 ( .A(n580), .Z(n362) );
  XNOR2_X1 U73 ( .A(n362), .B(\mult_x_1/n284 ), .ZN(n50) );
  XNOR2_X1 U74 ( .A(n362), .B(\mult_x_1/n283 ), .ZN(n152) );
  OAI22_X1 U75 ( .A1(n179), .A2(n50), .B1(n14), .B2(n152), .ZN(n131) );
  XNOR2_X1 U76 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n143) );
  XNOR2_X1 U77 ( .A(n579), .B(\mult_x_1/n282 ), .ZN(n51) );
  INV_X1 U78 ( .A(n143), .ZN(n46) );
  XNOR2_X1 U79 ( .A(n579), .B(\mult_x_1/n281 ), .ZN(n141) );
  OAI22_X1 U80 ( .A1(n12), .A2(n51), .B1(n148), .B2(n141), .ZN(n132) );
  XNOR2_X1 U81 ( .A(n131), .B(n132), .ZN(n156) );
  XNOR2_X1 U82 ( .A(\mult_x_1/a[6] ), .B(n580), .ZN(n48) );
  XNOR2_X1 U83 ( .A(\mult_x_1/n310 ), .B(n39), .ZN(n47) );
  NAND2_X2 U84 ( .A1(n48), .A2(n47), .ZN(n240) );
  XNOR2_X1 U85 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n53) );
  BUF_X2 U86 ( .A(n48), .Z(n241) );
  XNOR2_X1 U87 ( .A(n23), .B(\mult_x_1/n286 ), .ZN(n57) );
  OAI22_X1 U88 ( .A1(n240), .A2(n53), .B1(n241), .B2(n57), .ZN(n62) );
  BUF_X2 U89 ( .A(\mult_x_1/n313 ), .Z(n108) );
  XNOR2_X1 U90 ( .A(n108), .B(\mult_x_1/n281 ), .ZN(n64) );
  XNOR2_X1 U91 ( .A(n184), .B(n108), .ZN(n55) );
  OAI22_X1 U92 ( .A1(n17), .A2(n64), .B1(n55), .B2(n9), .ZN(n61) );
  NAND2_X1 U93 ( .A1(n27), .A2(n23), .ZN(n58) );
  INV_X1 U94 ( .A(n58), .ZN(n49) );
  AND2_X1 U95 ( .A1(\mult_x_1/n288 ), .A2(n49), .ZN(n60) );
  XNOR2_X1 U96 ( .A(n362), .B(\mult_x_1/n285 ), .ZN(n63) );
  OAI22_X1 U97 ( .A1(n15), .A2(n63), .B1(n14), .B2(n50), .ZN(n68) );
  XNOR2_X1 U98 ( .A(n579), .B(\mult_x_1/n283 ), .ZN(n65) );
  OR2_X1 U99 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n52) );
  OAI22_X1 U100 ( .A1(n240), .A2(n28), .B1(n52), .B2(n241), .ZN(n225) );
  XNOR2_X1 U101 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n54) );
  OAI22_X1 U102 ( .A1(n240), .A2(n54), .B1(n241), .B2(n53), .ZN(n224) );
  AOI21_X1 U103 ( .B1(n109), .B2(n9), .A(n55), .ZN(n56) );
  INV_X1 U104 ( .A(n56), .ZN(n137) );
  XNOR2_X1 U105 ( .A(n23), .B(\mult_x_1/n285 ), .ZN(n151) );
  OAI22_X1 U106 ( .A1(n240), .A2(n57), .B1(n241), .B2(n151), .ZN(n136) );
  NOR2_X1 U107 ( .A1(n32), .A2(n58), .ZN(n135) );
  XNOR2_X1 U108 ( .A(n287), .B(n286), .ZN(n59) );
  XNOR2_X1 U109 ( .A(n38), .B(n59), .ZN(n167) );
  FA_X1 U110 ( .A(n62), .B(n61), .CI(n60), .CO(n155), .S(n257) );
  XNOR2_X1 U111 ( .A(n362), .B(\mult_x_1/n286 ), .ZN(n71) );
  OAI22_X1 U112 ( .A1(n15), .A2(n71), .B1(n14), .B2(n63), .ZN(n228) );
  XNOR2_X1 U113 ( .A(n108), .B(\mult_x_1/n282 ), .ZN(n74) );
  OAI22_X1 U114 ( .A1(n17), .A2(n74), .B1(n64), .B2(n9), .ZN(n227) );
  XNOR2_X1 U115 ( .A(n579), .B(\mult_x_1/n284 ), .ZN(n73) );
  FA_X1 U116 ( .A(n68), .B(n67), .CI(n66), .CO(n287), .S(n255) );
  BUF_X1 U117 ( .A(en), .Z(n267) );
  OAI22_X1 U118 ( .A1(n167), .A2(n43), .B1(n22), .B2(n425), .ZN(n399) );
  OR2_X1 U119 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n69) );
  OAI22_X1 U120 ( .A1(n15), .A2(n31), .B1(n69), .B2(n180), .ZN(n80) );
  XNOR2_X1 U121 ( .A(n362), .B(\mult_x_1/n288 ), .ZN(n70) );
  XNOR2_X1 U122 ( .A(n362), .B(\mult_x_1/n287 ), .ZN(n72) );
  OAI22_X1 U123 ( .A1(n15), .A2(n70), .B1(n180), .B2(n72), .ZN(n79) );
  OAI22_X1 U124 ( .A1(n16), .A2(n72), .B1(n14), .B2(n71), .ZN(n230) );
  XOR2_X1 U125 ( .A(n231), .B(n230), .Z(n78) );
  XNOR2_X1 U126 ( .A(n579), .B(\mult_x_1/n285 ), .ZN(n81) );
  XNOR2_X1 U127 ( .A(n108), .B(\mult_x_1/n283 ), .ZN(n82) );
  OAI22_X1 U128 ( .A1(n109), .A2(n82), .B1(n74), .B2(n9), .ZN(n220) );
  INV_X1 U129 ( .A(n241), .ZN(n75) );
  AND2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n75), .ZN(n219) );
  XNOR2_X1 U131 ( .A(n220), .B(n219), .ZN(n76) );
  XNOR2_X1 U132 ( .A(n221), .B(n76), .ZN(n229) );
  INV_X1 U133 ( .A(n229), .ZN(n77) );
  XNOR2_X1 U134 ( .A(n78), .B(n77), .ZN(n87) );
  HA_X1 U135 ( .A(n80), .B(n79), .CO(n231), .S(n91) );
  XNOR2_X1 U136 ( .A(n579), .B(\mult_x_1/n286 ), .ZN(n92) );
  XNOR2_X1 U137 ( .A(n108), .B(\mult_x_1/n284 ), .ZN(n93) );
  OR2_X1 U138 ( .A1(n87), .A2(n86), .ZN(n275) );
  NAND2_X1 U139 ( .A1(n87), .A2(n86), .ZN(n276) );
  NAND2_X1 U140 ( .A1(n275), .A2(n276), .ZN(n128) );
  XNOR2_X1 U141 ( .A(n91), .B(n90), .ZN(n126) );
  XNOR2_X1 U142 ( .A(n579), .B(\mult_x_1/n287 ), .ZN(n101) );
  XNOR2_X1 U143 ( .A(n108), .B(\mult_x_1/n285 ), .ZN(n103) );
  OAI22_X1 U144 ( .A1(n109), .A2(n103), .B1(n93), .B2(n9), .ZN(n96) );
  INV_X1 U145 ( .A(n96), .ZN(n117) );
  INV_X1 U146 ( .A(n180), .ZN(n94) );
  NAND2_X1 U147 ( .A1(n94), .A2(\mult_x_1/n288 ), .ZN(n116) );
  INV_X1 U148 ( .A(n125), .ZN(n100) );
  NAND2_X1 U149 ( .A1(n25), .A2(n100), .ZN(n316) );
  XNOR2_X1 U150 ( .A(n579), .B(\mult_x_1/n288 ), .ZN(n102) );
  XNOR2_X1 U151 ( .A(n108), .B(\mult_x_1/n286 ), .ZN(n106) );
  OAI22_X1 U152 ( .A1(n109), .A2(n106), .B1(n103), .B2(n9), .ZN(n120) );
  INV_X1 U153 ( .A(n120), .ZN(n104) );
  XNOR2_X1 U154 ( .A(n121), .B(n104), .ZN(n114) );
  OR2_X1 U155 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n105) );
  OR2_X1 U156 ( .A1(n114), .A2(n113), .ZN(n304) );
  XNOR2_X1 U157 ( .A(n108), .B(\mult_x_1/n287 ), .ZN(n107) );
  OAI22_X1 U158 ( .A1(n17), .A2(n107), .B1(n106), .B2(n9), .ZN(n112) );
  AND2_X1 U159 ( .A1(\mult_x_1/n288 ), .A2(n46), .ZN(n111) );
  NOR2_X1 U160 ( .A1(n112), .A2(n111), .ZN(n297) );
  OAI22_X1 U161 ( .A1(n109), .A2(\mult_x_1/n288 ), .B1(n107), .B2(n9), .ZN(
        n294) );
  OR2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n42), .ZN(n110) );
  NAND2_X1 U163 ( .A1(n110), .A2(n17), .ZN(n293) );
  NAND2_X1 U164 ( .A1(n294), .A2(n293), .ZN(n300) );
  NAND2_X1 U165 ( .A1(n112), .A2(n111), .ZN(n298) );
  OAI21_X1 U166 ( .B1(n297), .B2(n300), .A(n298), .ZN(n305) );
  NAND2_X1 U167 ( .A1(n114), .A2(n113), .ZN(n303) );
  INV_X1 U168 ( .A(n303), .ZN(n115) );
  XNOR2_X1 U169 ( .A(n117), .B(n116), .ZN(n119) );
  XNOR2_X1 U170 ( .A(n119), .B(n118), .ZN(n123) );
  NOR2_X1 U171 ( .A1(n123), .A2(n122), .ZN(n308) );
  NAND2_X1 U172 ( .A1(n123), .A2(n122), .ZN(n312) );
  OAI21_X1 U173 ( .B1(n314), .B2(n308), .A(n312), .ZN(n124) );
  NAND2_X1 U174 ( .A1(n316), .A2(n124), .ZN(n127) );
  NAND2_X1 U175 ( .A1(n126), .A2(n125), .ZN(n315) );
  AND2_X1 U176 ( .A1(n127), .A2(n315), .ZN(n278) );
  XNOR2_X1 U177 ( .A(n128), .B(n278), .ZN(n130) );
  BUF_X4 U178 ( .A(n267), .Z(n322) );
  OR2_X1 U179 ( .A1(n322), .A2(n364), .ZN(n129) );
  OAI21_X1 U180 ( .B1(n130), .B2(n21), .A(n129), .ZN(n469) );
  OR2_X2 U181 ( .A1(n132), .A2(n131), .ZN(n161) );
  INV_X1 U182 ( .A(n161), .ZN(n134) );
  NOR2_X1 U183 ( .A1(n33), .A2(n58), .ZN(n160) );
  INV_X1 U184 ( .A(n160), .ZN(n133) );
  NAND2_X1 U185 ( .A1(n134), .A2(n133), .ZN(n138) );
  FA_X1 U186 ( .A(n137), .B(n136), .CI(n135), .CO(n163), .S(n286) );
  NAND2_X1 U187 ( .A1(n138), .A2(n163), .ZN(n140) );
  NAND2_X1 U188 ( .A1(n140), .A2(n139), .ZN(n212) );
  XNOR2_X1 U189 ( .A(n23), .B(\mult_x_1/n284 ), .ZN(n150) );
  XNOR2_X1 U190 ( .A(n23), .B(\mult_x_1/n283 ), .ZN(n177) );
  OAI22_X1 U191 ( .A1(n240), .A2(n150), .B1(n241), .B2(n177), .ZN(n198) );
  XNOR2_X1 U192 ( .A(n579), .B(n184), .ZN(n146) );
  INV_X1 U193 ( .A(n141), .ZN(n142) );
  NAND3_X1 U194 ( .A1(n142), .A2(n26), .A3(n144), .ZN(n145) );
  OAI21_X1 U195 ( .B1(n146), .B2(n148), .A(n145), .ZN(n197) );
  INV_X1 U196 ( .A(n149), .ZN(n196) );
  OAI22_X1 U197 ( .A1(n240), .A2(n151), .B1(n241), .B2(n150), .ZN(n159) );
  XNOR2_X1 U198 ( .A(n362), .B(\mult_x_1/n282 ), .ZN(n153) );
  OAI22_X1 U199 ( .A1(n179), .A2(n152), .B1(n180), .B2(n153), .ZN(n158) );
  INV_X1 U200 ( .A(n197), .ZN(n157) );
  NOR2_X1 U201 ( .A1(n34), .A2(n58), .ZN(n204) );
  XNOR2_X1 U202 ( .A(n362), .B(\mult_x_1/n281 ), .ZN(n176) );
  OAI22_X1 U203 ( .A1(n15), .A2(n153), .B1(n14), .B2(n176), .ZN(n203) );
  XNOR2_X1 U204 ( .A(n204), .B(n203), .ZN(n154) );
  XNOR2_X1 U205 ( .A(n202), .B(n154), .ZN(n210) );
  FA_X1 U206 ( .A(n158), .B(n159), .CI(n157), .CO(n202), .S(n281) );
  XNOR2_X1 U207 ( .A(n163), .B(n162), .ZN(n280) );
  INV_X1 U208 ( .A(n171), .ZN(n164) );
  NAND2_X1 U209 ( .A1(n164), .A2(n22), .ZN(n165) );
  OAI22_X1 U210 ( .A1(n172), .A2(n165), .B1(n22), .B2(n424), .ZN(n395) );
  NAND2_X1 U211 ( .A1(n168), .A2(n22), .ZN(n170) );
  OR2_X1 U212 ( .A1(n22), .A2(n41), .ZN(n169) );
  NAND2_X1 U213 ( .A1(n170), .A2(n169), .ZN(n401) );
  NAND2_X1 U214 ( .A1(n172), .A2(n171), .ZN(n173) );
  NAND2_X1 U215 ( .A1(n173), .A2(n22), .ZN(n175) );
  OR2_X1 U216 ( .A1(n22), .A2(n420), .ZN(n174) );
  NAND2_X1 U217 ( .A1(n175), .A2(n174), .ZN(n397) );
  XNOR2_X1 U236 ( .A(n184), .B(n362), .ZN(n181) );
  OAI22_X1 U237 ( .A1(n179), .A2(n176), .B1(n181), .B2(n180), .ZN(n186) );
  INV_X1 U238 ( .A(n186), .ZN(n195) );
  XNOR2_X1 U239 ( .A(n23), .B(\mult_x_1/n282 ), .ZN(n178) );
  OAI22_X1 U240 ( .A1(n240), .A2(n177), .B1(n241), .B2(n178), .ZN(n194) );
  NOR2_X1 U241 ( .A1(n35), .A2(n58), .ZN(n193) );
  NOR2_X1 U242 ( .A1(n36), .A2(n58), .ZN(n191) );
  XNOR2_X1 U243 ( .A(n23), .B(\mult_x_1/n281 ), .ZN(n185) );
  OAI22_X1 U244 ( .A1(n240), .A2(n178), .B1(n241), .B2(n185), .ZN(n188) );
  NAND2_X1 U245 ( .A1(n14), .A2(n179), .ZN(n183) );
  INV_X1 U246 ( .A(n181), .ZN(n182) );
  NAND2_X1 U247 ( .A1(n183), .A2(n182), .ZN(n187) );
  NOR2_X1 U248 ( .A1(n37), .A2(n58), .ZN(n238) );
  XNOR2_X1 U249 ( .A(n184), .B(n23), .ZN(n239) );
  OAI22_X1 U250 ( .A1(n240), .A2(n185), .B1(n239), .B2(n241), .ZN(n246) );
  INV_X1 U251 ( .A(n246), .ZN(n237) );
  FA_X1 U252 ( .A(n188), .B(n187), .CI(n186), .CO(n236), .S(n190) );
  OR2_X1 U253 ( .A1(n252), .A2(n253), .ZN(n189) );
  MUX2_X1 U254 ( .A(n365), .B(n189), .S(n22), .Z(n383) );
  FA_X1 U255 ( .A(n192), .B(n191), .CI(n190), .CO(n252), .S(n273) );
  FA_X1 U256 ( .A(n195), .B(n194), .CI(n193), .CO(n192), .S(n215) );
  FA_X1 U257 ( .A(n198), .B(n196), .CI(n20), .CO(n213), .S(n211) );
  INV_X1 U258 ( .A(n204), .ZN(n200) );
  INV_X1 U259 ( .A(n203), .ZN(n199) );
  NAND2_X1 U260 ( .A1(n200), .A2(n199), .ZN(n201) );
  NAND2_X1 U261 ( .A1(n202), .A2(n201), .ZN(n206) );
  NAND2_X1 U262 ( .A1(n206), .A2(n205), .ZN(n214) );
  OAI21_X1 U263 ( .B1(n215), .B2(n213), .A(n18), .ZN(n208) );
  OR2_X1 U264 ( .A1(n273), .A2(n272), .ZN(n209) );
  MUX2_X1 U265 ( .A(n366), .B(n209), .S(n22), .Z(n385) );
  FA_X1 U266 ( .A(n212), .B(n211), .CI(n210), .CO(n269), .S(n172) );
  INV_X1 U267 ( .A(n269), .ZN(n217) );
  XNOR2_X1 U268 ( .A(n214), .B(n213), .ZN(n216) );
  XNOR2_X1 U269 ( .A(n216), .B(n215), .ZN(n270) );
  NAND2_X1 U270 ( .A1(n19), .A2(n217), .ZN(n218) );
  HA_X1 U271 ( .A(n225), .B(n224), .CO(n66), .S(n259) );
  FA_X1 U272 ( .A(n228), .B(n227), .CI(n226), .CO(n256), .S(n258) );
  NAND2_X1 U273 ( .A1(n229), .A2(n231), .ZN(n234) );
  NAND2_X1 U274 ( .A1(n229), .A2(n230), .ZN(n233) );
  NAND2_X1 U275 ( .A1(n231), .A2(n230), .ZN(n232) );
  NAND3_X1 U276 ( .A1(n234), .A2(n233), .A3(n232), .ZN(n265) );
  OR2_X1 U277 ( .A1(n266), .A2(n265), .ZN(n235) );
  MUX2_X1 U278 ( .A(n368), .B(n235), .S(n22), .Z(n389) );
  FA_X1 U279 ( .A(n238), .B(n237), .CI(n236), .CO(n248), .S(n253) );
  AOI21_X1 U280 ( .B1(n241), .B2(n240), .A(n239), .ZN(n242) );
  INV_X1 U281 ( .A(n242), .ZN(n244) );
  NOR2_X1 U282 ( .A1(n30), .A2(n58), .ZN(n243) );
  XOR2_X1 U283 ( .A(n244), .B(n243), .Z(n245) );
  XOR2_X1 U284 ( .A(n246), .B(n245), .Z(n247) );
  OR2_X1 U285 ( .A1(n248), .A2(n247), .ZN(n250) );
  NAND2_X1 U286 ( .A1(n248), .A2(n247), .ZN(n249) );
  NAND2_X1 U287 ( .A1(n250), .A2(n249), .ZN(n251) );
  MUX2_X1 U288 ( .A(n369), .B(n251), .S(n22), .Z(n391) );
  NAND2_X1 U289 ( .A1(n253), .A2(n252), .ZN(n254) );
  MUX2_X1 U290 ( .A(n370), .B(n254), .S(n22), .Z(n393) );
  FA_X1 U291 ( .A(n257), .B(n256), .CI(n255), .CO(n166), .S(n263) );
  FA_X1 U292 ( .A(n260), .B(n259), .CI(n258), .CO(n262), .S(n266) );
  NOR2_X1 U293 ( .A1(n263), .A2(n262), .ZN(n261) );
  MUX2_X1 U294 ( .A(n375), .B(n261), .S(n22), .Z(n403) );
  NAND2_X1 U295 ( .A1(n263), .A2(n262), .ZN(n264) );
  MUX2_X1 U296 ( .A(n376), .B(n264), .S(n22), .Z(n405) );
  NAND2_X1 U297 ( .A1(n266), .A2(n265), .ZN(n268) );
  MUX2_X1 U298 ( .A(n377), .B(n268), .S(n322), .Z(n407) );
  NAND2_X1 U299 ( .A1(n270), .A2(n269), .ZN(n271) );
  MUX2_X1 U300 ( .A(n378), .B(n271), .S(n322), .Z(n409) );
  NAND2_X1 U301 ( .A1(n273), .A2(n272), .ZN(n274) );
  MUX2_X1 U302 ( .A(n379), .B(n274), .S(n322), .Z(n411) );
  INV_X1 U303 ( .A(n275), .ZN(n277) );
  OAI21_X1 U304 ( .B1(n278), .B2(n277), .A(n276), .ZN(n279) );
  FA_X1 U305 ( .A(n40), .B(n281), .CI(n280), .CO(n171), .S(n282) );
  MUX2_X1 U306 ( .A(n381), .B(n282), .S(n322), .Z(n415) );
  MUX2_X1 U307 ( .A(n382), .B(n290), .S(n322), .Z(n417) );
  BUF_X2 U308 ( .A(rst_n), .Z(n427) );
  BUF_X1 U309 ( .A(rst_n), .Z(n291) );
  MUX2_X1 U310 ( .A(product[0]), .B(n541), .S(n322), .Z(n429) );
  MUX2_X1 U311 ( .A(n541), .B(n542), .S(n322), .Z(n431) );
  AND2_X1 U312 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n292) );
  MUX2_X1 U313 ( .A(n542), .B(n292), .S(n322), .Z(n433) );
  MUX2_X1 U314 ( .A(product[1]), .B(n544), .S(n322), .Z(n435) );
  MUX2_X1 U315 ( .A(n544), .B(n545), .S(n322), .Z(n437) );
  OR2_X1 U316 ( .A1(n294), .A2(n293), .ZN(n295) );
  AND2_X1 U317 ( .A1(n295), .A2(n300), .ZN(n296) );
  MUX2_X1 U318 ( .A(n545), .B(n296), .S(n322), .Z(n439) );
  MUX2_X1 U319 ( .A(product[2]), .B(n547), .S(n322), .Z(n441) );
  MUX2_X1 U320 ( .A(n547), .B(n548), .S(n322), .Z(n443) );
  INV_X1 U321 ( .A(n297), .ZN(n299) );
  NAND2_X1 U322 ( .A1(n299), .A2(n298), .ZN(n301) );
  XOR2_X1 U323 ( .A(n301), .B(n300), .Z(n302) );
  MUX2_X1 U324 ( .A(n548), .B(n302), .S(n322), .Z(n445) );
  MUX2_X1 U325 ( .A(product[3]), .B(n550), .S(n322), .Z(n447) );
  MUX2_X1 U326 ( .A(n550), .B(n551), .S(n322), .Z(n449) );
  NAND2_X1 U327 ( .A1(n304), .A2(n303), .ZN(n306) );
  XNOR2_X1 U328 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U329 ( .A(n551), .B(n307), .S(n322), .Z(n451) );
  MUX2_X1 U330 ( .A(product[4]), .B(n553), .S(n322), .Z(n453) );
  MUX2_X1 U331 ( .A(n553), .B(n554), .S(n322), .Z(n455) );
  INV_X1 U332 ( .A(n308), .ZN(n311) );
  NAND2_X1 U333 ( .A1(n311), .A2(n312), .ZN(n309) );
  XOR2_X1 U334 ( .A(n314), .B(n309), .Z(n310) );
  MUX2_X1 U335 ( .A(n554), .B(n310), .S(n322), .Z(n457) );
  MUX2_X1 U336 ( .A(product[5]), .B(n556), .S(n322), .Z(n459) );
  MUX2_X1 U337 ( .A(n556), .B(n557), .S(n322), .Z(n461) );
  INV_X1 U338 ( .A(n311), .ZN(n313) );
  OAI21_X1 U339 ( .B1(n314), .B2(n313), .A(n312), .ZN(n318) );
  NAND2_X1 U340 ( .A1(n316), .A2(n315), .ZN(n317) );
  XNOR2_X1 U341 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U342 ( .A(n557), .B(n319), .S(n322), .Z(n463) );
  MUX2_X1 U343 ( .A(product[6]), .B(n559), .S(n322), .Z(n465) );
  MUX2_X1 U344 ( .A(n559), .B(n560), .S(n322), .Z(n467) );
  MUX2_X1 U345 ( .A(product[7]), .B(n562), .S(n322), .Z(n471) );
  NAND2_X1 U346 ( .A1(n368), .A2(n377), .ZN(n320) );
  XNOR2_X1 U347 ( .A(n380), .B(n320), .ZN(n321) );
  MUX2_X1 U348 ( .A(n562), .B(n321), .S(n322), .Z(n473) );
  MUX2_X1 U349 ( .A(product[8]), .B(n564), .S(n322), .Z(n475) );
  AOI21_X1 U350 ( .B1(n380), .B2(n368), .A(n422), .ZN(n325) );
  NAND2_X1 U351 ( .A1(n423), .A2(n376), .ZN(n323) );
  XOR2_X1 U352 ( .A(n325), .B(n323), .Z(n324) );
  BUF_X2 U353 ( .A(en), .Z(n363) );
  MUX2_X1 U354 ( .A(n564), .B(n324), .S(n363), .Z(n477) );
  MUX2_X1 U355 ( .A(product[9]), .B(n566), .S(n363), .Z(n479) );
  OAI21_X1 U356 ( .B1(n325), .B2(n375), .A(n376), .ZN(n336) );
  INV_X1 U357 ( .A(n336), .ZN(n328) );
  NAND2_X1 U358 ( .A1(n425), .A2(n374), .ZN(n326) );
  XOR2_X1 U359 ( .A(n328), .B(n326), .Z(n327) );
  MUX2_X1 U360 ( .A(n566), .B(n327), .S(n363), .Z(n481) );
  MUX2_X1 U361 ( .A(product[10]), .B(n568), .S(n363), .Z(n483) );
  OAI21_X1 U362 ( .B1(n328), .B2(n373), .A(n374), .ZN(n331) );
  NOR2_X1 U363 ( .A1(n381), .A2(n382), .ZN(n334) );
  INV_X1 U364 ( .A(n334), .ZN(n329) );
  NAND2_X1 U365 ( .A1(n381), .A2(n382), .ZN(n333) );
  NAND2_X1 U366 ( .A1(n329), .A2(n333), .ZN(n330) );
  XNOR2_X1 U367 ( .A(n331), .B(n330), .ZN(n332) );
  MUX2_X1 U368 ( .A(n568), .B(n332), .S(n363), .Z(n485) );
  MUX2_X1 U369 ( .A(product[11]), .B(n570), .S(n363), .Z(n487) );
  NOR2_X1 U370 ( .A1(n334), .A2(n373), .ZN(n337) );
  OAI21_X1 U371 ( .B1(n334), .B2(n374), .A(n333), .ZN(n335) );
  AOI21_X1 U372 ( .B1(n337), .B2(n336), .A(n335), .ZN(n359) );
  NAND2_X1 U373 ( .A1(n424), .A2(n372), .ZN(n338) );
  XOR2_X1 U374 ( .A(n359), .B(n338), .Z(n339) );
  MUX2_X1 U375 ( .A(n570), .B(n339), .S(n363), .Z(n489) );
  MUX2_X1 U376 ( .A(product[12]), .B(n572), .S(n363), .Z(n491) );
  OAI21_X1 U377 ( .B1(n359), .B2(n371), .A(n372), .ZN(n341) );
  NAND2_X1 U378 ( .A1(n367), .A2(n378), .ZN(n340) );
  XNOR2_X1 U379 ( .A(n341), .B(n340), .ZN(n342) );
  MUX2_X1 U380 ( .A(n572), .B(n342), .S(n363), .Z(n493) );
  MUX2_X1 U381 ( .A(product[13]), .B(n574), .S(n363), .Z(n495) );
  NAND2_X1 U382 ( .A1(n424), .A2(n367), .ZN(n344) );
  AOI21_X1 U383 ( .B1(n420), .B2(n367), .A(n426), .ZN(n343) );
  OAI21_X1 U384 ( .B1(n359), .B2(n344), .A(n343), .ZN(n346) );
  NAND2_X1 U385 ( .A1(n366), .A2(n379), .ZN(n345) );
  XNOR2_X1 U386 ( .A(n346), .B(n345), .ZN(n347) );
  MUX2_X1 U387 ( .A(n574), .B(n347), .S(n363), .Z(n497) );
  MUX2_X1 U388 ( .A(product[14]), .B(n576), .S(n363), .Z(n499) );
  NAND2_X1 U389 ( .A1(n367), .A2(n366), .ZN(n349) );
  NOR2_X1 U390 ( .A1(n371), .A2(n349), .ZN(n355) );
  INV_X1 U391 ( .A(n355), .ZN(n351) );
  AOI21_X1 U392 ( .B1(n426), .B2(n366), .A(n421), .ZN(n348) );
  OAI21_X1 U393 ( .B1(n349), .B2(n372), .A(n348), .ZN(n356) );
  INV_X1 U394 ( .A(n356), .ZN(n350) );
  OAI21_X1 U395 ( .B1(n359), .B2(n351), .A(n350), .ZN(n353) );
  NAND2_X1 U396 ( .A1(n365), .A2(n370), .ZN(n352) );
  XNOR2_X1 U397 ( .A(n353), .B(n352), .ZN(n354) );
  MUX2_X1 U398 ( .A(n576), .B(n354), .S(n363), .Z(n501) );
  MUX2_X1 U399 ( .A(product[15]), .B(n578), .S(n363), .Z(n503) );
  NAND2_X1 U400 ( .A1(n355), .A2(n365), .ZN(n358) );
  AOI21_X1 U401 ( .B1(n356), .B2(n365), .A(n419), .ZN(n357) );
  OAI21_X1 U402 ( .B1(n359), .B2(n358), .A(n357), .ZN(n360) );
  XNOR2_X1 U403 ( .A(n360), .B(n369), .ZN(n361) );
  MUX2_X1 U404 ( .A(n578), .B(n361), .S(n363), .Z(n505) );
  MUX2_X1 U405 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n363), .Z(n507) );
  MUX2_X1 U406 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n363), .Z(n509) );
  MUX2_X1 U407 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n363), .Z(n511) );
  MUX2_X1 U408 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n363), .Z(n513) );
  MUX2_X1 U409 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n363), .Z(n515) );
  MUX2_X1 U410 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n363), .Z(n517) );
  MUX2_X1 U411 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n363), .Z(n519) );
  MUX2_X1 U412 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n363), .Z(n521) );
  MUX2_X1 U413 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n363), .Z(n523) );
  MUX2_X1 U414 ( .A(n108), .B(A_extended[1]), .S(n363), .Z(n525) );
  MUX2_X1 U415 ( .A(n11), .B(A_extended[2]), .S(n363), .Z(n527) );
  MUX2_X1 U416 ( .A(n579), .B(A_extended[3]), .S(n363), .Z(n529) );
  MUX2_X1 U417 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n363), .Z(n531) );
  MUX2_X1 U418 ( .A(n362), .B(A_extended[5]), .S(n363), .Z(n533) );
  MUX2_X1 U419 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n363), .Z(n535) );
  MUX2_X1 U420 ( .A(n23), .B(A_extended[7]), .S(n363), .Z(n537) );
  OR2_X1 U421 ( .A1(n363), .A2(n581), .ZN(n539) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_17 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n374, n376,
         n378, n380, n382, n384, n386, n388, n390, n392, n394, n396, n398,
         n400, n402, n404, n406, n408, n409, n410, n411, n412, n413, n414,
         n415, n417, n419, n421, n423, n425, n427, n429, n431, n433, n435,
         n437, n439, n441, n443, n445, n447, n449, n451, n453, n455, n457,
         n459, n461, n463, n465, n467, n469, n471, n473, n475, n477, n479,
         n481, n483, n485, n487, n489, n491, n493, n495, n497, n499, n501,
         n503, n505, n507, n509, n511, n513, n515, n517, n519, n521, n523,
         n525, n527, n529, n530, n532, n533, n535, n536, n538, n539, n541,
         n542, n544, n545, n547, n548, n550, n552, n554, n556, n558, n560,
         n562, n564, n566, n567, n568, n569, n570;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n281), .SE(n527), .CK(clk), .Q(n569)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n415), .SE(n523), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n22) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n415), .SE(n521), .CK(clk), .Q(n568), 
        .QN(n31) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n415), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n20) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n415), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n18) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n415), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n9) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n415), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n23) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n415), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n28) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n415), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n281), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n27) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n281), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n281), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n25) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n281), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n281), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n281), .SE(n493), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n281), .SE(n491), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n281), .SE(n489), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n281), .SE(n487), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n281), .SE(n485), .CK(clk), .Q(n562)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n281), .SE(n483), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n415), .SE(n481), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n415), .SE(n479), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n415), .SE(n477), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n415), .SE(n475), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n415), .SE(n473), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n415), .SE(n471), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n281), .SE(n469), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n415), .SE(n467), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n415), .SE(n465), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n281), .SE(n463), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n415), .SE(n461), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n415), .SE(n459), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n415), .SE(n457), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n415), .SE(n455), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n415), .SE(n453), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n415), .SE(n451), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n415), .SE(n449), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n415), .SE(n447), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n415), .SE(n445), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n415), .SE(n443), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n415), .SE(n441), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n415), .SE(n439), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n415), .SE(n437), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n415), .SE(n435), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n415), .SE(n433), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n415), .SE(n431), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n281), .SE(n429), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n415), .SE(n427), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n281), .SE(n425), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n415), .SE(n423), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n415), .SE(n421), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n281), .SE(n419), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n415), .SE(n417), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n415), .SE(n517), .CK(clk), .Q(n567), 
        .QN(n32) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n415), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n36) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n570), .SE(n406), .CK(
        clk), .QN(n371) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n570), .SI(1'b1), .SE(n404), .CK(clk), 
        .Q(n370), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n570), .SE(n402), .CK(
        clk), .Q(n353), .QN(n369) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n570), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n368), .QN(n33) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n570), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n367), .QN(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n570), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n366), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n570), .SE(n394), .CK(
        clk), .Q(n37), .QN(n365) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n570), .SE(n392), .CK(
        clk), .Q(n352), .QN(n364) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n570), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n363), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n570), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n362) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n570), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n361), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n570), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n360), .QN(n35) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n570), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n358), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n570), .SE(n378), .CK(
        clk), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n570), .SE(n376), .CK(
        clk), .QN(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n570), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n570), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n354) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n415), .SE(n525), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n21) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n570), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n359), .QN(n413) );
  BUF_X1 U2 ( .A(n173), .Z(n246) );
  NAND2_X1 U3 ( .A1(n41), .A2(n12), .ZN(n245) );
  NAND2_X1 U4 ( .A1(n7), .A2(n5), .ZN(n388) );
  OR2_X1 U5 ( .A1(n311), .A2(n6), .ZN(n5) );
  INV_X1 U6 ( .A(n362), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n8), .A2(n311), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n268), .A2(n267), .ZN(n8) );
  BUF_X4 U9 ( .A(en), .Z(n311) );
  OR2_X1 U10 ( .A1(n188), .A2(n187), .ZN(n11) );
  XNOR2_X1 U11 ( .A(\mult_x_1/a[6] ), .B(n568), .ZN(n12) );
  XNOR2_X1 U12 ( .A(n32), .B(n27), .ZN(n175) );
  INV_X1 U13 ( .A(n184), .ZN(n180) );
  INV_X1 U14 ( .A(n86), .ZN(n83) );
  INV_X1 U15 ( .A(n85), .ZN(n82) );
  XNOR2_X1 U16 ( .A(n30), .B(n53), .ZN(n199) );
  XNOR2_X1 U17 ( .A(n86), .B(n85), .ZN(n53) );
  XNOR2_X1 U18 ( .A(n57), .B(n56), .ZN(n262) );
  XNOR2_X1 U19 ( .A(n55), .B(n54), .ZN(n57) );
  NAND2_X1 U20 ( .A1(n103), .A2(n102), .ZN(n126) );
  XNOR2_X1 U21 ( .A(\mult_x_1/n310 ), .B(n22), .ZN(n41) );
  BUF_X1 U22 ( .A(n153), .Z(n19) );
  CLKBUF_X1 U23 ( .A(n176), .Z(n15) );
  INV_X1 U24 ( .A(n101), .ZN(n97) );
  NAND2_X1 U25 ( .A1(n186), .A2(n185), .ZN(n187) );
  NAND2_X1 U26 ( .A1(n182), .A2(n181), .ZN(n186) );
  NAND2_X1 U27 ( .A1(n180), .A2(n179), .ZN(n181) );
  NAND2_X1 U28 ( .A1(n88), .A2(n87), .ZN(n193) );
  NAND2_X1 U29 ( .A1(n86), .A2(n85), .ZN(n87) );
  INV_X1 U30 ( .A(n198), .ZN(n66) );
  OR2_X1 U31 ( .A1(n311), .A2(n33), .ZN(n132) );
  OAI21_X1 U32 ( .B1(n131), .B2(n130), .A(n351), .ZN(n133) );
  INV_X1 U33 ( .A(n203), .ZN(n95) );
  INV_X1 U34 ( .A(n23), .ZN(n13) );
  XNOR2_X1 U35 ( .A(n40), .B(n21), .ZN(n14) );
  INV_X1 U36 ( .A(n14), .ZN(n47) );
  BUF_X2 U37 ( .A(\mult_x_1/n310 ), .Z(n350) );
  INV_X1 U38 ( .A(n39), .ZN(n176) );
  INV_X1 U39 ( .A(n172), .ZN(n16) );
  INV_X1 U40 ( .A(n16), .ZN(n17) );
  NAND2_X1 U41 ( .A1(n153), .A2(n9), .ZN(n172) );
  NAND2_X1 U42 ( .A1(n184), .A2(n183), .ZN(n185) );
  INV_X1 U43 ( .A(n183), .ZN(n179) );
  XNOR2_X1 U44 ( .A(n184), .B(n183), .ZN(n137) );
  XNOR2_X1 U45 ( .A(n18), .B(\mult_x_1/n313 ), .ZN(n39) );
  XOR2_X1 U46 ( .A(n20), .B(n31), .Z(n59) );
  BUF_X2 U47 ( .A(n568), .Z(n349) );
  XNOR2_X1 U48 ( .A(n182), .B(n137), .ZN(n163) );
  INV_X1 U49 ( .A(rst_n), .ZN(n570) );
  XOR2_X1 U50 ( .A(n71), .B(n70), .Z(n30) );
  BUF_X2 U51 ( .A(n567), .Z(n348) );
  AND2_X1 U52 ( .A1(n70), .A2(n71), .ZN(n34) );
  NAND2_X1 U53 ( .A1(n191), .A2(n359), .ZN(n69) );
  XNOR2_X1 U54 ( .A(n567), .B(\mult_x_1/a[4] ), .ZN(n58) );
  NAND2_X1 U55 ( .A1(n59), .A2(n58), .ZN(n212) );
  XNOR2_X1 U56 ( .A(n349), .B(\mult_x_1/n284 ), .ZN(n48) );
  BUF_X2 U57 ( .A(n58), .Z(n213) );
  XNOR2_X1 U58 ( .A(n349), .B(\mult_x_1/n283 ), .ZN(n73) );
  OAI22_X1 U59 ( .A1(n212), .A2(n48), .B1(n213), .B2(n73), .ZN(n76) );
  XNOR2_X1 U60 ( .A(n567), .B(\mult_x_1/a[2] ), .ZN(n38) );
  OR2_X2 U61 ( .A1(n39), .A2(n38), .ZN(n178) );
  XNOR2_X1 U62 ( .A(n348), .B(\mult_x_1/n282 ), .ZN(n49) );
  XNOR2_X1 U63 ( .A(n348), .B(\mult_x_1/n281 ), .ZN(n74) );
  OAI22_X1 U64 ( .A1(n178), .A2(n49), .B1(n176), .B2(n74), .ZN(n75) );
  XNOR2_X1 U65 ( .A(n76), .B(n75), .ZN(n71) );
  AND2_X1 U66 ( .A1(\mult_x_1/n310 ), .A2(n569), .ZN(n40) );
  AND2_X1 U67 ( .A1(\mult_x_1/n288 ), .A2(n14), .ZN(n56) );
  BUF_X2 U68 ( .A(\mult_x_1/n313 ), .Z(n153) );
  XNOR2_X1 U69 ( .A(n19), .B(\mult_x_1/n281 ), .ZN(n61) );
  AND2_X1 U70 ( .A1(n569), .A2(\mult_x_1/n281 ), .ZN(n208) );
  XNOR2_X1 U71 ( .A(n208), .B(n153), .ZN(n44) );
  OAI22_X1 U72 ( .A1(n172), .A2(n61), .B1(n44), .B2(n9), .ZN(n55) );
  XNOR2_X1 U73 ( .A(\mult_x_1/a[6] ), .B(n568), .ZN(n173) );
  XNOR2_X1 U74 ( .A(n350), .B(\mult_x_1/n287 ), .ZN(n51) );
  XNOR2_X1 U75 ( .A(n350), .B(\mult_x_1/n286 ), .ZN(n46) );
  OAI22_X1 U76 ( .A1(n245), .A2(n51), .B1(n246), .B2(n46), .ZN(n54) );
  OAI21_X1 U77 ( .B1(n56), .B2(n55), .A(n54), .ZN(n43) );
  NAND2_X1 U78 ( .A1(n56), .A2(n55), .ZN(n42) );
  NAND2_X1 U79 ( .A1(n43), .A2(n42), .ZN(n70) );
  AOI21_X1 U80 ( .B1(n172), .B2(n9), .A(n44), .ZN(n45) );
  INV_X1 U81 ( .A(n45), .ZN(n79) );
  XNOR2_X1 U82 ( .A(n350), .B(\mult_x_1/n285 ), .ZN(n72) );
  OAI22_X1 U83 ( .A1(n245), .A2(n46), .B1(n246), .B2(n72), .ZN(n78) );
  NOR2_X1 U84 ( .A1(n24), .A2(n47), .ZN(n77) );
  NAND2_X1 U85 ( .A1(n59), .A2(n58), .ZN(n169) );
  XNOR2_X1 U86 ( .A(n349), .B(\mult_x_1/n285 ), .ZN(n60) );
  OAI22_X1 U87 ( .A1(n169), .A2(n60), .B1(n213), .B2(n48), .ZN(n65) );
  XNOR2_X1 U88 ( .A(n348), .B(\mult_x_1/n283 ), .ZN(n62) );
  OAI22_X1 U89 ( .A1(n178), .A2(n62), .B1(n15), .B2(n49), .ZN(n64) );
  OR2_X1 U90 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n50) );
  OAI22_X1 U91 ( .A1(n245), .A2(n21), .B1(n50), .B2(n246), .ZN(n233) );
  XNOR2_X1 U92 ( .A(n350), .B(\mult_x_1/n288 ), .ZN(n52) );
  OAI22_X1 U93 ( .A1(n245), .A2(n52), .B1(n246), .B2(n51), .ZN(n232) );
  INV_X1 U94 ( .A(n199), .ZN(n67) );
  NAND2_X1 U95 ( .A1(n59), .A2(n58), .ZN(n136) );
  XNOR2_X1 U96 ( .A(n349), .B(\mult_x_1/n286 ), .ZN(n167) );
  OAI22_X1 U97 ( .A1(n136), .A2(n167), .B1(n213), .B2(n60), .ZN(n236) );
  XNOR2_X1 U98 ( .A(n153), .B(\mult_x_1/n282 ), .ZN(n170) );
  OAI22_X1 U99 ( .A1(n17), .A2(n170), .B1(n61), .B2(n9), .ZN(n235) );
  OAI22_X1 U100 ( .A1(n178), .A2(n175), .B1(n15), .B2(n62), .ZN(n234) );
  FA_X1 U101 ( .A(n65), .B(n64), .CI(n63), .CO(n85), .S(n260) );
  NAND3_X1 U102 ( .A1(n67), .A2(n66), .A3(n311), .ZN(n68) );
  NAND2_X1 U103 ( .A1(n69), .A2(n68), .ZN(n382) );
  XNOR2_X1 U104 ( .A(n350), .B(\mult_x_1/n284 ), .ZN(n104) );
  OAI22_X1 U105 ( .A1(n245), .A2(n72), .B1(n246), .B2(n104), .ZN(n109) );
  XNOR2_X1 U106 ( .A(n349), .B(\mult_x_1/n282 ), .ZN(n110) );
  OAI22_X1 U107 ( .A1(n169), .A2(n73), .B1(n213), .B2(n110), .ZN(n108) );
  XNOR2_X1 U108 ( .A(n348), .B(n208), .ZN(n105) );
  OAI22_X1 U109 ( .A1(n178), .A2(n74), .B1(n105), .B2(n176), .ZN(n116) );
  INV_X1 U110 ( .A(n116), .ZN(n107) );
  OR2_X1 U111 ( .A1(n76), .A2(n75), .ZN(n101) );
  NOR2_X1 U112 ( .A1(n25), .A2(n47), .ZN(n100) );
  XNOR2_X1 U113 ( .A(n101), .B(n100), .ZN(n80) );
  FA_X1 U114 ( .A(n79), .B(n78), .CI(n77), .CO(n99), .S(n86) );
  XNOR2_X1 U115 ( .A(n80), .B(n99), .ZN(n93) );
  INV_X1 U116 ( .A(n351), .ZN(n81) );
  NOR2_X1 U117 ( .A1(n194), .A2(n81), .ZN(n90) );
  NAND2_X1 U118 ( .A1(n83), .A2(n82), .ZN(n84) );
  NAND2_X1 U119 ( .A1(n30), .A2(n84), .ZN(n88) );
  INV_X1 U120 ( .A(n193), .ZN(n89) );
  NAND2_X1 U121 ( .A1(n90), .A2(n89), .ZN(n92) );
  OR2_X1 U122 ( .A1(n311), .A2(n352), .ZN(n91) );
  NAND2_X1 U123 ( .A1(n92), .A2(n91), .ZN(n392) );
  FA_X1 U124 ( .A(n34), .B(n94), .CI(n93), .CO(n203), .S(n194) );
  NAND2_X1 U125 ( .A1(n95), .A2(n351), .ZN(n112) );
  INV_X1 U126 ( .A(n100), .ZN(n96) );
  NAND2_X1 U127 ( .A1(n97), .A2(n96), .ZN(n98) );
  NAND2_X1 U128 ( .A1(n99), .A2(n98), .ZN(n103) );
  NAND2_X1 U129 ( .A1(n101), .A2(n100), .ZN(n102) );
  XNOR2_X1 U130 ( .A(n350), .B(\mult_x_1/n283 ), .ZN(n113) );
  OAI22_X1 U131 ( .A1(n245), .A2(n104), .B1(n246), .B2(n113), .ZN(n117) );
  AOI21_X1 U132 ( .B1(n15), .B2(n178), .A(n105), .ZN(n106) );
  INV_X1 U133 ( .A(n106), .ZN(n115) );
  FA_X1 U134 ( .A(n109), .B(n108), .CI(n107), .CO(n119), .S(n94) );
  XNOR2_X1 U135 ( .A(n349), .B(\mult_x_1/n281 ), .ZN(n114) );
  OAI22_X1 U136 ( .A1(n136), .A2(n110), .B1(n213), .B2(n114), .ZN(n121) );
  NOR2_X1 U137 ( .A1(n26), .A2(n47), .ZN(n120) );
  XNOR2_X1 U138 ( .A(n121), .B(n120), .ZN(n111) );
  XNOR2_X1 U139 ( .A(n119), .B(n111), .ZN(n124) );
  OAI22_X1 U140 ( .A1(n112), .A2(n204), .B1(n311), .B2(n353), .ZN(n402) );
  NOR2_X1 U141 ( .A1(n27), .A2(n47), .ZN(n217) );
  XNOR2_X1 U142 ( .A(n350), .B(\mult_x_1/n282 ), .ZN(n210) );
  OAI22_X1 U143 ( .A1(n245), .A2(n113), .B1(n246), .B2(n210), .ZN(n216) );
  XNOR2_X1 U144 ( .A(n208), .B(n349), .ZN(n211) );
  OAI22_X1 U145 ( .A1(n136), .A2(n114), .B1(n211), .B2(n213), .ZN(n218) );
  INV_X1 U146 ( .A(n218), .ZN(n215) );
  FA_X1 U147 ( .A(n117), .B(n116), .CI(n115), .CO(n226), .S(n125) );
  OR2_X1 U148 ( .A1(n121), .A2(n120), .ZN(n118) );
  NAND2_X1 U149 ( .A1(n119), .A2(n118), .ZN(n123) );
  NAND2_X1 U150 ( .A1(n121), .A2(n120), .ZN(n122) );
  NAND2_X1 U151 ( .A1(n123), .A2(n122), .ZN(n225) );
  FA_X1 U152 ( .A(n126), .B(n125), .CI(n124), .CO(n130), .S(n204) );
  NAND2_X1 U153 ( .A1(n131), .A2(n130), .ZN(n127) );
  NAND2_X1 U154 ( .A1(n127), .A2(n311), .ZN(n129) );
  OR2_X1 U155 ( .A1(n351), .A2(n414), .ZN(n128) );
  NAND2_X1 U156 ( .A1(n129), .A2(n128), .ZN(n398) );
  NAND2_X1 U157 ( .A1(n133), .A2(n132), .ZN(n400) );
  OR2_X1 U158 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n134) );
  OAI22_X1 U159 ( .A1(n169), .A2(n31), .B1(n134), .B2(n213), .ZN(n166) );
  XNOR2_X1 U160 ( .A(n349), .B(\mult_x_1/n288 ), .ZN(n135) );
  XNOR2_X1 U161 ( .A(n349), .B(\mult_x_1/n287 ), .ZN(n168) );
  OAI22_X1 U162 ( .A1(n136), .A2(n135), .B1(n213), .B2(n168), .ZN(n165) );
  XNOR2_X1 U163 ( .A(n348), .B(\mult_x_1/n286 ), .ZN(n140) );
  XNOR2_X1 U164 ( .A(n348), .B(\mult_x_1/n285 ), .ZN(n177) );
  OAI22_X1 U165 ( .A1(n178), .A2(n140), .B1(n176), .B2(n177), .ZN(n184) );
  XNOR2_X1 U166 ( .A(n19), .B(\mult_x_1/n284 ), .ZN(n138) );
  XNOR2_X1 U167 ( .A(n153), .B(\mult_x_1/n283 ), .ZN(n171) );
  OAI22_X1 U168 ( .A1(n17), .A2(n138), .B1(n171), .B2(n9), .ZN(n183) );
  XNOR2_X1 U169 ( .A(n153), .B(\mult_x_1/n285 ), .ZN(n146) );
  OAI22_X1 U170 ( .A1(n172), .A2(n146), .B1(n138), .B2(n9), .ZN(n143) );
  INV_X1 U171 ( .A(n213), .ZN(n139) );
  AND2_X1 U172 ( .A1(\mult_x_1/n288 ), .A2(n139), .ZN(n142) );
  XNOR2_X1 U173 ( .A(n348), .B(\mult_x_1/n287 ), .ZN(n144) );
  OAI22_X1 U174 ( .A1(n178), .A2(n144), .B1(n176), .B2(n140), .ZN(n141) );
  OR2_X1 U175 ( .A1(n163), .A2(n162), .ZN(n305) );
  FA_X1 U176 ( .A(n143), .B(n142), .CI(n141), .CO(n162), .S(n161) );
  XNOR2_X1 U177 ( .A(n348), .B(\mult_x_1/n288 ), .ZN(n145) );
  OAI22_X1 U178 ( .A1(n178), .A2(n145), .B1(n176), .B2(n144), .ZN(n148) );
  XNOR2_X1 U179 ( .A(n153), .B(\mult_x_1/n286 ), .ZN(n150) );
  OAI22_X1 U180 ( .A1(n172), .A2(n150), .B1(n146), .B2(n9), .ZN(n147) );
  NOR2_X1 U181 ( .A1(n161), .A2(n160), .ZN(n298) );
  HA_X1 U182 ( .A(n148), .B(n147), .CO(n160), .S(n158) );
  OR2_X1 U183 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n149) );
  OAI22_X1 U184 ( .A1(n178), .A2(n32), .B1(n149), .B2(n15), .ZN(n157) );
  OR2_X1 U185 ( .A1(n158), .A2(n157), .ZN(n294) );
  XNOR2_X1 U186 ( .A(n19), .B(\mult_x_1/n287 ), .ZN(n152) );
  OAI22_X1 U187 ( .A1(n17), .A2(n152), .B1(n150), .B2(n9), .ZN(n156) );
  INV_X1 U188 ( .A(n176), .ZN(n151) );
  AND2_X1 U189 ( .A1(\mult_x_1/n288 ), .A2(n151), .ZN(n155) );
  NOR2_X1 U190 ( .A1(n156), .A2(n155), .ZN(n287) );
  OAI22_X1 U191 ( .A1(n17), .A2(\mult_x_1/n288 ), .B1(n152), .B2(n9), .ZN(n284) );
  OR2_X1 U192 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n154) );
  NAND2_X1 U193 ( .A1(n154), .A2(n17), .ZN(n283) );
  NAND2_X1 U194 ( .A1(n284), .A2(n283), .ZN(n290) );
  NAND2_X1 U195 ( .A1(n156), .A2(n155), .ZN(n288) );
  OAI21_X1 U196 ( .B1(n287), .B2(n290), .A(n288), .ZN(n295) );
  NAND2_X1 U197 ( .A1(n158), .A2(n157), .ZN(n293) );
  INV_X1 U198 ( .A(n293), .ZN(n159) );
  AOI21_X1 U199 ( .B1(n294), .B2(n295), .A(n159), .ZN(n301) );
  NAND2_X1 U200 ( .A1(n161), .A2(n160), .ZN(n299) );
  OAI21_X1 U201 ( .B1(n298), .B2(n301), .A(n299), .ZN(n306) );
  NAND2_X1 U202 ( .A1(n163), .A2(n162), .ZN(n304) );
  INV_X1 U203 ( .A(n304), .ZN(n164) );
  AOI21_X1 U204 ( .B1(n305), .B2(n306), .A(n164), .ZN(n278) );
  HA_X1 U205 ( .A(n166), .B(n165), .CO(n239), .S(n182) );
  OAI22_X1 U206 ( .A1(n169), .A2(n168), .B1(n213), .B2(n167), .ZN(n238) );
  OAI22_X1 U207 ( .A1(n172), .A2(n171), .B1(n170), .B2(n9), .ZN(n231) );
  INV_X1 U208 ( .A(n173), .ZN(n174) );
  AND2_X1 U209 ( .A1(\mult_x_1/n288 ), .A2(n174), .ZN(n230) );
  OAI22_X1 U210 ( .A1(n178), .A2(n177), .B1(n176), .B2(n175), .ZN(n229) );
  OR2_X1 U211 ( .A1(n188), .A2(n187), .ZN(n276) );
  NAND2_X1 U212 ( .A1(n188), .A2(n187), .ZN(n277) );
  NAND2_X1 U213 ( .A1(n11), .A2(n277), .ZN(n189) );
  XNOR2_X1 U214 ( .A(n278), .B(n189), .ZN(n192) );
  INV_X1 U215 ( .A(n351), .ZN(n191) );
  NAND2_X1 U216 ( .A1(n191), .A2(n548), .ZN(n190) );
  OAI21_X1 U217 ( .B1(n192), .B2(n191), .A(n190), .ZN(n457) );
  NAND2_X1 U218 ( .A1(n194), .A2(n193), .ZN(n195) );
  NAND2_X1 U219 ( .A1(n195), .A2(n311), .ZN(n197) );
  OR2_X1 U220 ( .A1(n311), .A2(n37), .ZN(n196) );
  NAND2_X1 U221 ( .A1(n197), .A2(n196), .ZN(n394) );
  NAND2_X1 U222 ( .A1(n199), .A2(n198), .ZN(n200) );
  NAND2_X1 U223 ( .A1(n200), .A2(n311), .ZN(n202) );
  OR2_X1 U224 ( .A1(n311), .A2(n35), .ZN(n201) );
  NAND2_X1 U225 ( .A1(n202), .A2(n201), .ZN(n384) );
  NAND2_X1 U226 ( .A1(n204), .A2(n203), .ZN(n205) );
  NAND2_X1 U227 ( .A1(n205), .A2(n311), .ZN(n207) );
  OR2_X1 U228 ( .A1(n351), .A2(n409), .ZN(n206) );
  NAND2_X1 U229 ( .A1(n207), .A2(n206), .ZN(n404) );
  NOR2_X1 U248 ( .A1(n28), .A2(n47), .ZN(n243) );
  XNOR2_X1 U249 ( .A(n350), .B(n13), .ZN(n209) );
  XNOR2_X1 U250 ( .A(n208), .B(n350), .ZN(n244) );
  OAI22_X1 U251 ( .A1(n245), .A2(n209), .B1(n244), .B2(n246), .ZN(n251) );
  INV_X1 U252 ( .A(n251), .ZN(n242) );
  OAI22_X1 U253 ( .A1(n245), .A2(n210), .B1(n246), .B2(n209), .ZN(n220) );
  AOI21_X1 U254 ( .B1(n213), .B2(n212), .A(n211), .ZN(n214) );
  INV_X1 U255 ( .A(n214), .ZN(n219) );
  FA_X1 U256 ( .A(n217), .B(n216), .CI(n215), .CO(n224), .S(n227) );
  NOR2_X1 U257 ( .A1(n29), .A2(n47), .ZN(n223) );
  FA_X1 U258 ( .A(n220), .B(n219), .CI(n218), .CO(n241), .S(n222) );
  OR2_X1 U259 ( .A1(n258), .A2(n257), .ZN(n221) );
  MUX2_X1 U260 ( .A(n354), .B(n221), .S(n311), .Z(n372) );
  FA_X1 U261 ( .A(n224), .B(n223), .CI(n222), .CO(n257), .S(n274) );
  FA_X1 U262 ( .A(n227), .B(n226), .CI(n225), .CO(n273), .S(n131) );
  OR2_X1 U263 ( .A1(n274), .A2(n273), .ZN(n228) );
  MUX2_X1 U264 ( .A(n355), .B(n228), .S(n311), .Z(n374) );
  FA_X1 U265 ( .A(n231), .B(n230), .CI(n229), .CO(n265), .S(n237) );
  HA_X1 U266 ( .A(n233), .B(n232), .CO(n63), .S(n264) );
  FA_X1 U267 ( .A(n236), .B(n235), .CI(n234), .CO(n261), .S(n263) );
  FA_X1 U268 ( .A(n239), .B(n238), .CI(n237), .CO(n270), .S(n188) );
  OR2_X1 U269 ( .A1(n271), .A2(n270), .ZN(n240) );
  MUX2_X1 U270 ( .A(n356), .B(n240), .S(n311), .Z(n376) );
  FA_X1 U271 ( .A(n243), .B(n242), .CI(n241), .CO(n253), .S(n258) );
  AOI21_X1 U272 ( .B1(n246), .B2(n245), .A(n244), .ZN(n247) );
  INV_X1 U273 ( .A(n247), .ZN(n249) );
  NOR2_X1 U274 ( .A1(n23), .A2(n47), .ZN(n248) );
  XOR2_X1 U275 ( .A(n249), .B(n248), .Z(n250) );
  XOR2_X1 U276 ( .A(n251), .B(n250), .Z(n252) );
  OR2_X1 U277 ( .A1(n253), .A2(n252), .ZN(n255) );
  NAND2_X1 U278 ( .A1(n253), .A2(n252), .ZN(n254) );
  NAND2_X1 U279 ( .A1(n255), .A2(n254), .ZN(n256) );
  MUX2_X1 U280 ( .A(n357), .B(n256), .S(n311), .Z(n378) );
  NAND2_X1 U281 ( .A1(n258), .A2(n257), .ZN(n259) );
  MUX2_X1 U282 ( .A(n358), .B(n259), .S(n351), .Z(n380) );
  FA_X1 U283 ( .A(n262), .B(n261), .CI(n260), .CO(n198), .S(n268) );
  FA_X1 U284 ( .A(n265), .B(n264), .CI(n263), .CO(n267), .S(n271) );
  NOR2_X1 U285 ( .A1(n268), .A2(n267), .ZN(n266) );
  MUX2_X1 U286 ( .A(n361), .B(n266), .S(n311), .Z(n386) );
  NAND2_X1 U287 ( .A1(n271), .A2(n270), .ZN(n272) );
  MUX2_X1 U288 ( .A(n363), .B(n272), .S(n311), .Z(n390) );
  NAND2_X1 U289 ( .A1(n274), .A2(n273), .ZN(n275) );
  MUX2_X1 U290 ( .A(n366), .B(n275), .S(n311), .Z(n396) );
  INV_X1 U291 ( .A(n276), .ZN(n279) );
  OAI21_X1 U292 ( .B1(n279), .B2(n278), .A(n277), .ZN(n280) );
  MUX2_X1 U293 ( .A(n371), .B(n280), .S(n351), .Z(n406) );
  BUF_X2 U294 ( .A(rst_n), .Z(n415) );
  BUF_X1 U295 ( .A(rst_n), .Z(n281) );
  MUX2_X1 U296 ( .A(product[0]), .B(n529), .S(n311), .Z(n417) );
  MUX2_X1 U297 ( .A(n529), .B(n530), .S(n311), .Z(n419) );
  AND2_X1 U298 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n282) );
  MUX2_X1 U299 ( .A(n530), .B(n282), .S(n311), .Z(n421) );
  MUX2_X1 U300 ( .A(product[1]), .B(n532), .S(n311), .Z(n423) );
  MUX2_X1 U301 ( .A(n532), .B(n533), .S(n351), .Z(n425) );
  OR2_X1 U302 ( .A1(n284), .A2(n283), .ZN(n285) );
  AND2_X1 U303 ( .A1(n285), .A2(n290), .ZN(n286) );
  MUX2_X1 U304 ( .A(n533), .B(n286), .S(n311), .Z(n427) );
  MUX2_X1 U305 ( .A(product[2]), .B(n535), .S(n311), .Z(n429) );
  MUX2_X1 U306 ( .A(n535), .B(n536), .S(n311), .Z(n431) );
  INV_X1 U307 ( .A(n287), .ZN(n289) );
  NAND2_X1 U308 ( .A1(n289), .A2(n288), .ZN(n291) );
  XOR2_X1 U309 ( .A(n291), .B(n290), .Z(n292) );
  MUX2_X1 U310 ( .A(n536), .B(n292), .S(n311), .Z(n433) );
  MUX2_X1 U311 ( .A(product[3]), .B(n538), .S(n351), .Z(n435) );
  MUX2_X1 U312 ( .A(n538), .B(n539), .S(n311), .Z(n437) );
  NAND2_X1 U313 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U314 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U315 ( .A(n539), .B(n297), .S(n311), .Z(n439) );
  MUX2_X1 U316 ( .A(product[4]), .B(n541), .S(n311), .Z(n441) );
  MUX2_X1 U317 ( .A(n541), .B(n542), .S(n311), .Z(n443) );
  INV_X1 U318 ( .A(n298), .ZN(n300) );
  NAND2_X1 U319 ( .A1(n300), .A2(n299), .ZN(n302) );
  XOR2_X1 U320 ( .A(n302), .B(n301), .Z(n303) );
  MUX2_X1 U321 ( .A(n542), .B(n303), .S(n351), .Z(n445) );
  MUX2_X1 U322 ( .A(product[5]), .B(n544), .S(n311), .Z(n447) );
  MUX2_X1 U323 ( .A(n544), .B(n545), .S(n311), .Z(n449) );
  NAND2_X1 U324 ( .A1(n305), .A2(n304), .ZN(n307) );
  XNOR2_X1 U325 ( .A(n307), .B(n306), .ZN(n308) );
  MUX2_X1 U326 ( .A(n545), .B(n308), .S(n311), .Z(n451) );
  MUX2_X1 U327 ( .A(product[6]), .B(n547), .S(n311), .Z(n453) );
  MUX2_X1 U328 ( .A(n547), .B(n548), .S(n351), .Z(n455) );
  MUX2_X1 U329 ( .A(product[7]), .B(n550), .S(n311), .Z(n459) );
  NAND2_X1 U330 ( .A1(n356), .A2(n363), .ZN(n309) );
  XNOR2_X1 U331 ( .A(n371), .B(n309), .ZN(n310) );
  MUX2_X1 U332 ( .A(n550), .B(n310), .S(n311), .Z(n461) );
  MUX2_X1 U333 ( .A(product[8]), .B(n552), .S(n311), .Z(n463) );
  AOI21_X1 U334 ( .B1(n371), .B2(n356), .A(n411), .ZN(n314) );
  NAND2_X1 U335 ( .A1(n412), .A2(n362), .ZN(n312) );
  XOR2_X1 U336 ( .A(n314), .B(n312), .Z(n313) );
  BUF_X2 U337 ( .A(en), .Z(n351) );
  MUX2_X1 U338 ( .A(n552), .B(n313), .S(n311), .Z(n465) );
  MUX2_X1 U339 ( .A(product[9]), .B(n554), .S(n351), .Z(n467) );
  OAI21_X1 U340 ( .B1(n314), .B2(n361), .A(n362), .ZN(n322) );
  INV_X1 U341 ( .A(n322), .ZN(n317) );
  NAND2_X1 U342 ( .A1(n413), .A2(n360), .ZN(n315) );
  XOR2_X1 U343 ( .A(n317), .B(n315), .Z(n316) );
  MUX2_X1 U344 ( .A(n554), .B(n316), .S(n311), .Z(n469) );
  MUX2_X1 U345 ( .A(product[10]), .B(n556), .S(n351), .Z(n471) );
  OAI21_X1 U346 ( .B1(n317), .B2(n359), .A(n360), .ZN(n319) );
  NAND2_X1 U347 ( .A1(n352), .A2(n365), .ZN(n318) );
  XNOR2_X1 U348 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U349 ( .A(n556), .B(n320), .S(n311), .Z(n473) );
  MUX2_X1 U350 ( .A(product[11]), .B(n558), .S(n311), .Z(n475) );
  NOR2_X1 U351 ( .A1(n364), .A2(n359), .ZN(n323) );
  OAI21_X1 U352 ( .B1(n364), .B2(n360), .A(n365), .ZN(n321) );
  AOI21_X1 U353 ( .B1(n323), .B2(n322), .A(n321), .ZN(n345) );
  NAND2_X1 U354 ( .A1(n353), .A2(n370), .ZN(n324) );
  XOR2_X1 U355 ( .A(n345), .B(n324), .Z(n325) );
  MUX2_X1 U356 ( .A(n558), .B(n325), .S(n311), .Z(n477) );
  MUX2_X1 U357 ( .A(product[12]), .B(n560), .S(n311), .Z(n479) );
  OAI21_X1 U358 ( .B1(n345), .B2(n369), .A(n370), .ZN(n327) );
  NAND2_X1 U359 ( .A1(n368), .A2(n367), .ZN(n326) );
  XNOR2_X1 U360 ( .A(n327), .B(n326), .ZN(n328) );
  MUX2_X1 U361 ( .A(n560), .B(n328), .S(n311), .Z(n481) );
  MUX2_X1 U362 ( .A(product[13]), .B(n562), .S(n311), .Z(n483) );
  NAND2_X1 U363 ( .A1(n353), .A2(n368), .ZN(n330) );
  AOI21_X1 U364 ( .B1(n409), .B2(n368), .A(n414), .ZN(n329) );
  OAI21_X1 U365 ( .B1(n345), .B2(n330), .A(n329), .ZN(n332) );
  NAND2_X1 U366 ( .A1(n355), .A2(n366), .ZN(n331) );
  XNOR2_X1 U367 ( .A(n332), .B(n331), .ZN(n333) );
  MUX2_X1 U368 ( .A(n562), .B(n333), .S(n351), .Z(n485) );
  MUX2_X1 U369 ( .A(product[14]), .B(n564), .S(n311), .Z(n487) );
  NAND2_X1 U370 ( .A1(n368), .A2(n355), .ZN(n335) );
  NOR2_X1 U371 ( .A1(n369), .A2(n335), .ZN(n341) );
  INV_X1 U372 ( .A(n341), .ZN(n337) );
  AOI21_X1 U373 ( .B1(n414), .B2(n355), .A(n410), .ZN(n334) );
  OAI21_X1 U374 ( .B1(n335), .B2(n370), .A(n334), .ZN(n342) );
  INV_X1 U375 ( .A(n342), .ZN(n336) );
  OAI21_X1 U376 ( .B1(n345), .B2(n337), .A(n336), .ZN(n339) );
  NAND2_X1 U377 ( .A1(n354), .A2(n358), .ZN(n338) );
  XNOR2_X1 U378 ( .A(n339), .B(n338), .ZN(n340) );
  MUX2_X1 U379 ( .A(n564), .B(n340), .S(n311), .Z(n489) );
  MUX2_X1 U380 ( .A(product[15]), .B(n566), .S(n311), .Z(n491) );
  NAND2_X1 U381 ( .A1(n341), .A2(n354), .ZN(n344) );
  AOI21_X1 U382 ( .B1(n342), .B2(n354), .A(n408), .ZN(n343) );
  OAI21_X1 U383 ( .B1(n345), .B2(n344), .A(n343), .ZN(n346) );
  XNOR2_X1 U384 ( .A(n346), .B(n357), .ZN(n347) );
  MUX2_X1 U385 ( .A(n566), .B(n347), .S(n351), .Z(n493) );
  MUX2_X1 U386 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n311), .Z(n495) );
  MUX2_X1 U387 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n351), .Z(n497) );
  MUX2_X1 U388 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n351), .Z(n499) );
  MUX2_X1 U389 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n311), .Z(n501) );
  MUX2_X1 U390 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n351), .Z(n503) );
  MUX2_X1 U391 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n311), .Z(n505) );
  MUX2_X1 U392 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n311), .Z(n507) );
  MUX2_X1 U393 ( .A(n13), .B(B_extended[7]), .S(n311), .Z(n509) );
  MUX2_X1 U394 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n351), .Z(n511) );
  MUX2_X1 U395 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n311), .Z(n513) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n311), .Z(n515) );
  MUX2_X1 U397 ( .A(n348), .B(A_extended[3]), .S(n311), .Z(n517) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n351), .Z(n519) );
  MUX2_X1 U399 ( .A(n349), .B(A_extended[5]), .S(n311), .Z(n521) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n311), .Z(n523) );
  MUX2_X1 U401 ( .A(n350), .B(A_extended[7]), .S(n311), .Z(n525) );
  OR2_X1 U402 ( .A1(n311), .A2(n569), .ZN(n527) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_18 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n355, n357, n359, n361, n363, n365, n367, n369, n371,
         n373, n375, n377, n379, n381, n383, n385, n387, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n399, n401, n403, n405, n407,
         n409, n411, n413, n415, n417, n419, n421, n423, n425, n427, n429,
         n431, n433, n435, n437, n439, n441, n443, n445, n447, n449, n451,
         n453, n455, n457, n459, n461, n463, n465, n467, n469, n471, n473,
         n475, n477, n479, n481, n483, n485, n487, n489, n491, n493, n495,
         n497, n499, n501, n503, n505, n507, n509, n511, n512, n514, n515,
         n517, n518, n520, n521, n523, n524, n526, n527, n529, n530, n532,
         n534, n536, n538, n540, n542, n544, n546, n548, n549, n550, n551,
         n552;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n260), .SE(n509), .CK(clk), .Q(n551), 
        .QN(n36) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n397), .SE(n507), .CK(clk), .Q(n550), 
        .QN(n24) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n397), .SE(n505), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n397), .SE(n503), .CK(clk), .Q(n549), 
        .QN(n27) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n397), .SE(n501), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n34) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n397), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n26) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n397), .SE(n497), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n397), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n397), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n29) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n397), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n31) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n260), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n260), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n32) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n260), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n33) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n260), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n28) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n260), .SE(n477), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n22) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n260), .SE(n475), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n260), .SE(n473), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n260), .SE(n471), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n260), .SE(n469), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n260), .SE(n467), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n260), .SE(n465), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n397), .SE(n463), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n397), .SE(n461), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n397), .SE(n459), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n397), .SE(n457), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n397), .SE(n455), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n397), .SE(n453), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n260), .SE(n451), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n397), .SE(n449), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n397), .SE(n447), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n260), .SE(n445), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n397), .SE(n443), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n397), .SE(n441), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n397), .SE(n439), .CK(clk), .Q(n530), 
        .QN(n334) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n397), .SE(n437), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n397), .SE(n435), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n397), .SE(n433), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n397), .SE(n431), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n397), .SE(n429), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n397), .SE(n427), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n397), .SE(n425), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n397), .SE(n423), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n397), .SE(n421), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n397), .SE(n419), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n397), .SE(n417), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n397), .SE(n415), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n397), .SE(n413), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n260), .SE(n411), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n397), .SE(n409), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n260), .SE(n407), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n397), .SE(n405), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n397), .SE(n403), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n260), .SE(n401), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n397), .SE(n399), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n397), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n38) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n552), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n552), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n552), .SE(n383), .CK(
        clk), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n552), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n349), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n552), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n348), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n552), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n552), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n346), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n552), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n345), .QN(n37) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n552), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n344), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n552), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n343), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n552), .SE(n367), .CK(
        clk), .Q(n395), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n552), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n341), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n552), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n340), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n552), .SE(n361), .CK(
        clk), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n552), .SE(n359), .CK(
        clk), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n552), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n552), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n552), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n335) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n397), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n25) );
  BUF_X4 U2 ( .A(en), .Z(n69) );
  OR2_X1 U3 ( .A1(n38), .A2(\mult_x_1/n180 ), .ZN(n104) );
  OR2_X1 U4 ( .A1(n18), .A2(n21), .ZN(n40) );
  CLKBUF_X2 U5 ( .A(n550), .Z(n332) );
  BUF_X1 U6 ( .A(n549), .Z(n331) );
  CLKBUF_X1 U7 ( .A(n207), .Z(n6) );
  INV_X1 U8 ( .A(n47), .ZN(n20) );
  INV_X1 U9 ( .A(n115), .ZN(n111) );
  INV_X1 U10 ( .A(n114), .ZN(n110) );
  OAI22_X1 U11 ( .A1(n148), .A2(n88), .B1(n20), .B2(n109), .ZN(n115) );
  NAND2_X1 U12 ( .A1(n117), .A2(n116), .ZN(n118) );
  NAND2_X1 U13 ( .A1(n115), .A2(n114), .ZN(n116) );
  NAND2_X1 U14 ( .A1(n113), .A2(n112), .ZN(n117) );
  NAND2_X1 U15 ( .A1(n111), .A2(n110), .ZN(n112) );
  AND2_X1 U16 ( .A1(n169), .A2(n167), .ZN(n56) );
  XNOR2_X1 U17 ( .A(n113), .B(n91), .ZN(n96) );
  XNOR2_X1 U18 ( .A(n115), .B(n114), .ZN(n91) );
  NAND2_X1 U19 ( .A1(n209), .A2(n208), .ZN(n256) );
  NAND2_X1 U20 ( .A1(n67), .A2(n66), .ZN(n123) );
  NAND2_X1 U21 ( .A1(n228), .A2(n227), .ZN(n66) );
  NAND2_X1 U22 ( .A1(n230), .A2(n65), .ZN(n67) );
  OR2_X1 U23 ( .A1(n228), .A2(n227), .ZN(n65) );
  XNOR2_X1 U24 ( .A(n230), .B(n229), .ZN(n236) );
  XNOR2_X1 U25 ( .A(n228), .B(n227), .ZN(n229) );
  INV_X1 U26 ( .A(n167), .ZN(n168) );
  OR2_X1 U27 ( .A1(n119), .A2(n118), .ZN(n244) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(n245) );
  XNOR2_X1 U29 ( .A(n198), .B(n199), .ZN(n211) );
  AOI21_X1 U30 ( .B1(n11), .B2(n284), .A(n97), .ZN(n7) );
  CLKBUF_X1 U31 ( .A(n144), .Z(n8) );
  CLKBUF_X1 U32 ( .A(n144), .Z(n9) );
  CLKBUF_X1 U33 ( .A(n144), .Z(n10) );
  XNOR2_X1 U34 ( .A(n26), .B(n32), .ZN(n109) );
  OAI21_X1 U35 ( .B1(n277), .B2(n280), .A(n278), .ZN(n11) );
  XOR2_X1 U36 ( .A(n141), .B(n140), .Z(n12) );
  XOR2_X1 U37 ( .A(n142), .B(n12), .Z(n197) );
  NAND2_X1 U38 ( .A1(n142), .A2(n141), .ZN(n13) );
  NAND2_X1 U39 ( .A1(n142), .A2(n140), .ZN(n14) );
  NAND2_X1 U40 ( .A1(n141), .A2(n140), .ZN(n15) );
  NAND3_X1 U41 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n139) );
  XNOR2_X1 U42 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n16) );
  BUF_X2 U43 ( .A(n89), .Z(n17) );
  AOI21_X2 U44 ( .B1(n273), .B2(n274), .A(n83), .ZN(n280) );
  AND2_X1 U45 ( .A1(n104), .A2(n5), .ZN(n18) );
  CLKBUF_X1 U46 ( .A(\mult_x_1/n281 ), .Z(n19) );
  OAI21_X1 U47 ( .B1(n220), .B2(n219), .A(n221), .ZN(n209) );
  NAND2_X1 U48 ( .A1(n220), .A2(n219), .ZN(n208) );
  INV_X1 U49 ( .A(n47), .ZN(n149) );
  XNOR2_X1 U50 ( .A(n145), .B(n89), .ZN(n21) );
  AND2_X1 U51 ( .A1(n551), .A2(\mult_x_1/n281 ), .ZN(n145) );
  XNOR2_X1 U52 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n46) );
  AND2_X1 U53 ( .A1(n212), .A2(n211), .ZN(n23) );
  INV_X1 U54 ( .A(rst_n), .ZN(n552) );
  XNOR2_X1 U55 ( .A(n206), .B(n205), .ZN(n35) );
  INV_X1 U56 ( .A(n46), .ZN(n47) );
  OR2_X1 U57 ( .A1(n123), .A2(n68), .ZN(n39) );
  BUF_X2 U58 ( .A(\mult_x_1/n313 ), .Z(n89) );
  XNOR2_X1 U59 ( .A(n145), .B(n17), .ZN(n52) );
  XOR2_X1 U60 ( .A(\mult_x_1/a[6] ), .B(n550), .Z(n41) );
  XNOR2_X1 U61 ( .A(n549), .B(\mult_x_1/a[6] ), .ZN(n105) );
  NAND2_X1 U62 ( .A1(n41), .A2(n105), .ZN(n144) );
  XNOR2_X1 U63 ( .A(n332), .B(\mult_x_1/n286 ), .ZN(n50) );
  BUF_X2 U64 ( .A(n105), .Z(n181) );
  XNOR2_X1 U65 ( .A(n332), .B(\mult_x_1/n285 ), .ZN(n152) );
  OAI22_X1 U66 ( .A1(n8), .A2(n50), .B1(n181), .B2(n152), .ZN(n201) );
  NAND2_X1 U67 ( .A1(n332), .A2(n36), .ZN(n128) );
  NOR2_X1 U68 ( .A1(n28), .A2(n128), .ZN(n200) );
  XNOR2_X1 U69 ( .A(n549), .B(n34), .ZN(n42) );
  XNOR2_X1 U70 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n43) );
  NAND2_X1 U71 ( .A1(n42), .A2(n43), .ZN(n157) );
  XNOR2_X1 U72 ( .A(n331), .B(\mult_x_1/n285 ), .ZN(n62) );
  INV_X1 U73 ( .A(n43), .ZN(n44) );
  INV_X2 U74 ( .A(n44), .ZN(n155) );
  XNOR2_X1 U75 ( .A(n331), .B(\mult_x_1/n284 ), .ZN(n54) );
  OAI22_X1 U76 ( .A1(n157), .A2(n62), .B1(n155), .B2(n54), .ZN(n58) );
  XOR2_X1 U77 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[2] ), .Z(n45) );
  NAND2_X1 U78 ( .A1(n45), .A2(n46), .ZN(n107) );
  BUF_X2 U79 ( .A(n107), .Z(n148) );
  BUF_X2 U80 ( .A(\mult_x_1/n312 ), .Z(n330) );
  XNOR2_X1 U81 ( .A(n330), .B(\mult_x_1/n283 ), .ZN(n64) );
  XNOR2_X1 U82 ( .A(n330), .B(\mult_x_1/n282 ), .ZN(n53) );
  OAI22_X1 U83 ( .A1(n148), .A2(n64), .B1(n20), .B2(n53), .ZN(n57) );
  XNOR2_X1 U84 ( .A(n332), .B(\mult_x_1/n288 ), .ZN(n48) );
  XNOR2_X1 U85 ( .A(n332), .B(\mult_x_1/n287 ), .ZN(n51) );
  OAI22_X1 U86 ( .A1(n10), .A2(n48), .B1(n181), .B2(n51), .ZN(n169) );
  OR2_X1 U87 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n49) );
  OAI22_X1 U88 ( .A1(n10), .A2(n24), .B1(n49), .B2(n181), .ZN(n167) );
  OAI22_X1 U89 ( .A1(n8), .A2(n51), .B1(n181), .B2(n50), .ZN(n61) );
  NOR2_X1 U90 ( .A1(n128), .A2(n22), .ZN(n60) );
  XNOR2_X1 U91 ( .A(n17), .B(n19), .ZN(n63) );
  OAI22_X1 U92 ( .A1(n104), .A2(n63), .B1(n52), .B2(n5), .ZN(n59) );
  INV_X1 U93 ( .A(n212), .ZN(n55) );
  XNOR2_X1 U94 ( .A(n330), .B(n19), .ZN(n146) );
  OAI22_X1 U95 ( .A1(n148), .A2(n53), .B1(n20), .B2(n146), .ZN(n198) );
  XNOR2_X1 U96 ( .A(n331), .B(\mult_x_1/n283 ), .ZN(n153) );
  OAI22_X1 U97 ( .A1(n157), .A2(n54), .B1(n155), .B2(n153), .ZN(n199) );
  XNOR2_X1 U98 ( .A(n55), .B(n211), .ZN(n252) );
  FA_X1 U99 ( .A(n58), .B(n57), .CI(n56), .CO(n253), .S(n230) );
  FA_X1 U100 ( .A(n61), .B(n60), .CI(n59), .CO(n212), .S(n228) );
  XNOR2_X1 U101 ( .A(n331), .B(\mult_x_1/n286 ), .ZN(n100) );
  OAI22_X1 U102 ( .A1(n157), .A2(n100), .B1(n155), .B2(n62), .ZN(n172) );
  XNOR2_X1 U103 ( .A(n89), .B(\mult_x_1/n282 ), .ZN(n102) );
  OAI22_X1 U104 ( .A1(n104), .A2(n102), .B1(n63), .B2(n5), .ZN(n171) );
  XNOR2_X1 U105 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n108) );
  OAI22_X1 U106 ( .A1(n148), .A2(n108), .B1(n20), .B2(n64), .ZN(n170) );
  INV_X1 U107 ( .A(en), .ZN(n68) );
  OAI22_X1 U108 ( .A1(n124), .A2(n39), .B1(n69), .B2(n394), .ZN(n371) );
  XNOR2_X1 U109 ( .A(n89), .B(\mult_x_1/n285 ), .ZN(n72) );
  XNOR2_X1 U110 ( .A(n89), .B(\mult_x_1/n284 ), .ZN(n90) );
  OAI22_X1 U111 ( .A1(n104), .A2(n72), .B1(n90), .B2(n5), .ZN(n94) );
  AND2_X1 U112 ( .A1(\mult_x_1/n288 ), .A2(n44), .ZN(n93) );
  XNOR2_X1 U113 ( .A(n330), .B(\mult_x_1/n287 ), .ZN(n70) );
  XNOR2_X1 U114 ( .A(n330), .B(\mult_x_1/n286 ), .ZN(n88) );
  OAI22_X1 U115 ( .A1(n148), .A2(n70), .B1(n20), .B2(n88), .ZN(n92) );
  XNOR2_X1 U116 ( .A(n330), .B(\mult_x_1/n288 ), .ZN(n71) );
  OAI22_X1 U117 ( .A1(n148), .A2(n71), .B1(n20), .B2(n70), .ZN(n74) );
  XNOR2_X1 U118 ( .A(n17), .B(\mult_x_1/n286 ), .ZN(n76) );
  OAI22_X1 U119 ( .A1(n104), .A2(n76), .B1(n72), .B2(n5), .ZN(n73) );
  NOR2_X1 U120 ( .A1(n85), .A2(n84), .ZN(n277) );
  HA_X1 U121 ( .A(n74), .B(n73), .CO(n84), .S(n82) );
  OR2_X1 U122 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n75) );
  OAI22_X1 U123 ( .A1(n148), .A2(n26), .B1(n75), .B2(n20), .ZN(n81) );
  OR2_X1 U124 ( .A1(n82), .A2(n81), .ZN(n273) );
  XNOR2_X1 U125 ( .A(n17), .B(\mult_x_1/n287 ), .ZN(n77) );
  OAI22_X1 U126 ( .A1(n104), .A2(n77), .B1(n76), .B2(n5), .ZN(n80) );
  AND2_X1 U127 ( .A1(\mult_x_1/n288 ), .A2(n47), .ZN(n79) );
  NOR2_X1 U128 ( .A1(n80), .A2(n79), .ZN(n266) );
  OAI22_X1 U129 ( .A1(n104), .A2(\mult_x_1/n288 ), .B1(n77), .B2(n5), .ZN(n263) );
  OR2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n78) );
  NAND2_X1 U131 ( .A1(n78), .A2(n104), .ZN(n262) );
  NAND2_X1 U132 ( .A1(n263), .A2(n262), .ZN(n269) );
  NAND2_X1 U133 ( .A1(n80), .A2(n79), .ZN(n267) );
  OAI21_X1 U134 ( .B1(n266), .B2(n269), .A(n267), .ZN(n274) );
  NAND2_X1 U135 ( .A1(n82), .A2(n81), .ZN(n272) );
  INV_X1 U136 ( .A(n272), .ZN(n83) );
  NAND2_X1 U137 ( .A1(n85), .A2(n84), .ZN(n278) );
  OAI21_X1 U138 ( .B1(n277), .B2(n280), .A(n278), .ZN(n285) );
  OR2_X1 U139 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n86) );
  OAI22_X1 U140 ( .A1(n157), .A2(n27), .B1(n86), .B2(n155), .ZN(n99) );
  XNOR2_X1 U141 ( .A(n331), .B(\mult_x_1/n288 ), .ZN(n87) );
  XNOR2_X1 U142 ( .A(n331), .B(\mult_x_1/n287 ), .ZN(n101) );
  OAI22_X1 U143 ( .A1(n157), .A2(n87), .B1(n155), .B2(n101), .ZN(n98) );
  XNOR2_X1 U144 ( .A(n89), .B(\mult_x_1/n283 ), .ZN(n103) );
  OAI22_X1 U145 ( .A1(n104), .A2(n90), .B1(n103), .B2(n5), .ZN(n114) );
  FA_X1 U146 ( .A(n94), .B(n93), .CI(n92), .CO(n95), .S(n85) );
  OR2_X1 U147 ( .A1(n96), .A2(n95), .ZN(n284) );
  NAND2_X1 U148 ( .A1(n96), .A2(n95), .ZN(n283) );
  INV_X1 U149 ( .A(n283), .ZN(n97) );
  AOI21_X1 U150 ( .B1(n11), .B2(n284), .A(n97), .ZN(n246) );
  HA_X1 U151 ( .A(n99), .B(n98), .CO(n175), .S(n113) );
  OAI22_X1 U152 ( .A1(n157), .A2(n101), .B1(n155), .B2(n100), .ZN(n174) );
  OAI22_X1 U153 ( .A1(n104), .A2(n103), .B1(n102), .B2(n5), .ZN(n166) );
  INV_X1 U154 ( .A(n105), .ZN(n106) );
  AND2_X1 U155 ( .A1(\mult_x_1/n288 ), .A2(n106), .ZN(n165) );
  OAI22_X1 U156 ( .A1(n107), .A2(n109), .B1(n149), .B2(n16), .ZN(n164) );
  NAND2_X1 U157 ( .A1(n244), .A2(n245), .ZN(n120) );
  XNOR2_X1 U158 ( .A(n7), .B(n120), .ZN(n122) );
  OR2_X1 U159 ( .A1(n69), .A2(n334), .ZN(n121) );
  OAI21_X1 U160 ( .B1(n122), .B2(n68), .A(n121), .ZN(n439) );
  NAND2_X1 U161 ( .A1(n124), .A2(n123), .ZN(n125) );
  NAND2_X1 U162 ( .A1(n125), .A2(n69), .ZN(n127) );
  OR2_X1 U163 ( .A1(n69), .A2(n37), .ZN(n126) );
  NAND2_X1 U164 ( .A1(n127), .A2(n126), .ZN(n373) );
  NOR2_X1 U183 ( .A1(n29), .A2(n128), .ZN(n179) );
  XNOR2_X1 U184 ( .A(n332), .B(n19), .ZN(n129) );
  XNOR2_X1 U185 ( .A(n145), .B(n332), .ZN(n180) );
  OAI22_X1 U186 ( .A1(n10), .A2(n129), .B1(n180), .B2(n181), .ZN(n186) );
  INV_X1 U187 ( .A(n186), .ZN(n178) );
  XNOR2_X1 U188 ( .A(n332), .B(\mult_x_1/n282 ), .ZN(n132) );
  OAI22_X1 U189 ( .A1(n9), .A2(n132), .B1(n181), .B2(n129), .ZN(n135) );
  XNOR2_X1 U190 ( .A(n331), .B(n19), .ZN(n154) );
  XNOR2_X1 U191 ( .A(n145), .B(n331), .ZN(n130) );
  OAI22_X1 U192 ( .A1(n157), .A2(n154), .B1(n130), .B2(n155), .ZN(n134) );
  AOI21_X1 U193 ( .B1(n155), .B2(n157), .A(n130), .ZN(n131) );
  INV_X1 U194 ( .A(n131), .ZN(n133) );
  INV_X1 U195 ( .A(n134), .ZN(n142) );
  XNOR2_X1 U196 ( .A(n332), .B(\mult_x_1/n283 ), .ZN(n143) );
  OAI22_X1 U197 ( .A1(n10), .A2(n143), .B1(n181), .B2(n132), .ZN(n141) );
  NOR2_X1 U198 ( .A1(n30), .A2(n128), .ZN(n140) );
  NOR2_X1 U199 ( .A1(n31), .A2(n128), .ZN(n138) );
  FA_X1 U200 ( .A(n135), .B(n134), .CI(n133), .CO(n177), .S(n137) );
  OR2_X1 U201 ( .A1(n193), .A2(n192), .ZN(n136) );
  MUX2_X1 U202 ( .A(n335), .B(n136), .S(n69), .Z(n353) );
  FA_X1 U203 ( .A(n139), .B(n138), .CI(n137), .CO(n192), .S(n242) );
  XNOR2_X1 U204 ( .A(n332), .B(\mult_x_1/n284 ), .ZN(n151) );
  OAI22_X1 U205 ( .A1(n9), .A2(n151), .B1(n181), .B2(n143), .ZN(n204) );
  XNOR2_X1 U206 ( .A(n330), .B(n145), .ZN(n147) );
  OAI22_X1 U207 ( .A1(n107), .A2(n146), .B1(n147), .B2(n149), .ZN(n203) );
  AOI21_X1 U208 ( .B1(n20), .B2(n148), .A(n147), .ZN(n150) );
  INV_X1 U209 ( .A(n150), .ZN(n202) );
  OAI22_X1 U210 ( .A1(n9), .A2(n152), .B1(n181), .B2(n151), .ZN(n215) );
  XNOR2_X1 U211 ( .A(n331), .B(\mult_x_1/n282 ), .ZN(n156) );
  OAI22_X1 U212 ( .A1(n157), .A2(n153), .B1(n155), .B2(n156), .ZN(n214) );
  INV_X1 U213 ( .A(n203), .ZN(n213) );
  NOR2_X1 U214 ( .A1(n32), .A2(n128), .ZN(n206) );
  INV_X1 U215 ( .A(n206), .ZN(n159) );
  OAI22_X1 U216 ( .A1(n157), .A2(n156), .B1(n155), .B2(n154), .ZN(n205) );
  INV_X1 U217 ( .A(n205), .ZN(n158) );
  NAND2_X1 U218 ( .A1(n159), .A2(n158), .ZN(n160) );
  NAND2_X1 U219 ( .A1(n207), .A2(n160), .ZN(n162) );
  NAND2_X1 U220 ( .A1(n206), .A2(n205), .ZN(n161) );
  NAND2_X1 U221 ( .A1(n162), .A2(n161), .ZN(n195) );
  OR2_X1 U222 ( .A1(n242), .A2(n241), .ZN(n163) );
  MUX2_X1 U223 ( .A(n336), .B(n163), .S(n69), .Z(n355) );
  FA_X1 U224 ( .A(n166), .B(n165), .CI(n164), .CO(n233), .S(n173) );
  XNOR2_X1 U225 ( .A(n169), .B(n168), .ZN(n232) );
  FA_X1 U226 ( .A(n172), .B(n171), .CI(n170), .CO(n227), .S(n231) );
  FA_X1 U227 ( .A(n175), .B(n174), .CI(n173), .CO(n238), .S(n119) );
  OR2_X1 U228 ( .A1(n239), .A2(n238), .ZN(n176) );
  MUX2_X1 U229 ( .A(n338), .B(n176), .S(n69), .Z(n359) );
  FA_X1 U230 ( .A(n179), .B(n178), .CI(n177), .CO(n188), .S(n193) );
  AOI21_X1 U231 ( .B1(n181), .B2(n9), .A(n180), .ZN(n182) );
  INV_X1 U232 ( .A(n182), .ZN(n184) );
  NOR2_X1 U233 ( .A1(n25), .A2(n128), .ZN(n183) );
  XOR2_X1 U234 ( .A(n184), .B(n183), .Z(n185) );
  XOR2_X1 U235 ( .A(n186), .B(n185), .Z(n187) );
  OR2_X1 U236 ( .A1(n188), .A2(n187), .ZN(n190) );
  NAND2_X1 U237 ( .A1(n188), .A2(n187), .ZN(n189) );
  NAND2_X1 U238 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U239 ( .A(n339), .B(n191), .S(n69), .Z(n361) );
  NAND2_X1 U240 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U241 ( .A(n340), .B(n194), .S(n69), .Z(n363) );
  FA_X1 U242 ( .A(n197), .B(n196), .CI(n195), .CO(n241), .S(n257) );
  OR2_X1 U243 ( .A1(n198), .A2(n199), .ZN(n218) );
  NOR2_X1 U244 ( .A1(n33), .A2(n128), .ZN(n217) );
  FA_X1 U245 ( .A(n40), .B(n201), .CI(n200), .CO(n216), .S(n254) );
  FA_X1 U246 ( .A(n204), .B(n203), .CI(n202), .CO(n196), .S(n219) );
  XNOR2_X1 U247 ( .A(n6), .B(n35), .ZN(n221) );
  NAND2_X1 U248 ( .A1(n257), .A2(n256), .ZN(n210) );
  MUX2_X1 U249 ( .A(n341), .B(n210), .S(n69), .Z(n365) );
  FA_X1 U250 ( .A(n215), .B(n214), .CI(n213), .CO(n207), .S(n250) );
  FA_X1 U251 ( .A(n218), .B(n217), .CI(n216), .CO(n220), .S(n249) );
  XNOR2_X1 U252 ( .A(n220), .B(n219), .ZN(n222) );
  XNOR2_X1 U253 ( .A(n222), .B(n221), .ZN(n225) );
  NOR2_X1 U254 ( .A1(n224), .A2(n225), .ZN(n223) );
  MUX2_X1 U255 ( .A(n342), .B(n223), .S(n69), .Z(n367) );
  NAND2_X1 U256 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U257 ( .A(n343), .B(n226), .S(n69), .Z(n369) );
  FA_X1 U258 ( .A(n233), .B(n232), .CI(n231), .CO(n235), .S(n239) );
  NOR2_X1 U259 ( .A1(n236), .A2(n235), .ZN(n234) );
  MUX2_X1 U260 ( .A(n346), .B(n234), .S(n69), .Z(n375) );
  NAND2_X1 U261 ( .A1(n236), .A2(n235), .ZN(n237) );
  MUX2_X1 U262 ( .A(n347), .B(n237), .S(n333), .Z(n377) );
  NAND2_X1 U263 ( .A1(n239), .A2(n238), .ZN(n240) );
  MUX2_X1 U264 ( .A(n348), .B(n240), .S(n333), .Z(n379) );
  NAND2_X1 U265 ( .A1(n242), .A2(n241), .ZN(n243) );
  MUX2_X1 U266 ( .A(n349), .B(n243), .S(n333), .Z(n381) );
  INV_X1 U267 ( .A(n244), .ZN(n247) );
  OAI21_X1 U268 ( .B1(n247), .B2(n246), .A(n245), .ZN(n248) );
  MUX2_X1 U269 ( .A(n350), .B(n248), .S(n333), .Z(n383) );
  FA_X1 U270 ( .A(n23), .B(n250), .CI(n249), .CO(n224), .S(n251) );
  MUX2_X1 U271 ( .A(n351), .B(n251), .S(n333), .Z(n385) );
  FA_X1 U272 ( .A(n254), .B(n253), .CI(n252), .CO(n255), .S(n124) );
  MUX2_X1 U273 ( .A(n352), .B(n255), .S(n333), .Z(n387) );
  OAI21_X1 U274 ( .B1(n257), .B2(n256), .A(n69), .ZN(n259) );
  NAND2_X1 U275 ( .A1(n68), .A2(n337), .ZN(n258) );
  NAND2_X1 U276 ( .A1(n259), .A2(n258), .ZN(n357) );
  BUF_X2 U277 ( .A(rst_n), .Z(n397) );
  BUF_X1 U278 ( .A(rst_n), .Z(n260) );
  MUX2_X1 U279 ( .A(product[0]), .B(n511), .S(n69), .Z(n399) );
  MUX2_X1 U280 ( .A(n511), .B(n512), .S(n69), .Z(n401) );
  AND2_X1 U281 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n261) );
  MUX2_X1 U282 ( .A(n512), .B(n261), .S(n69), .Z(n403) );
  MUX2_X1 U283 ( .A(product[1]), .B(n514), .S(n69), .Z(n405) );
  MUX2_X1 U284 ( .A(n514), .B(n515), .S(n69), .Z(n407) );
  OR2_X1 U285 ( .A1(n263), .A2(n262), .ZN(n264) );
  AND2_X1 U286 ( .A1(n264), .A2(n269), .ZN(n265) );
  MUX2_X1 U287 ( .A(n515), .B(n265), .S(n69), .Z(n409) );
  MUX2_X1 U288 ( .A(product[2]), .B(n517), .S(n69), .Z(n411) );
  MUX2_X1 U289 ( .A(n517), .B(n518), .S(n69), .Z(n413) );
  INV_X1 U290 ( .A(n266), .ZN(n268) );
  NAND2_X1 U291 ( .A1(n268), .A2(n267), .ZN(n270) );
  XOR2_X1 U292 ( .A(n270), .B(n269), .Z(n271) );
  MUX2_X1 U293 ( .A(n518), .B(n271), .S(n69), .Z(n415) );
  MUX2_X1 U294 ( .A(product[3]), .B(n520), .S(n69), .Z(n417) );
  MUX2_X1 U295 ( .A(n520), .B(n521), .S(n69), .Z(n419) );
  NAND2_X1 U296 ( .A1(n273), .A2(n272), .ZN(n275) );
  XNOR2_X1 U297 ( .A(n275), .B(n274), .ZN(n276) );
  MUX2_X1 U298 ( .A(n521), .B(n276), .S(n69), .Z(n421) );
  MUX2_X1 U299 ( .A(product[4]), .B(n523), .S(n69), .Z(n423) );
  MUX2_X1 U300 ( .A(n523), .B(n524), .S(n69), .Z(n425) );
  INV_X1 U301 ( .A(n277), .ZN(n279) );
  NAND2_X1 U302 ( .A1(n279), .A2(n278), .ZN(n281) );
  XOR2_X1 U303 ( .A(n281), .B(n280), .Z(n282) );
  MUX2_X1 U304 ( .A(n524), .B(n282), .S(n69), .Z(n427) );
  MUX2_X1 U305 ( .A(product[5]), .B(n526), .S(n69), .Z(n429) );
  MUX2_X1 U306 ( .A(n526), .B(n527), .S(n69), .Z(n431) );
  NAND2_X1 U307 ( .A1(n284), .A2(n283), .ZN(n286) );
  XNOR2_X1 U308 ( .A(n286), .B(n285), .ZN(n287) );
  MUX2_X1 U309 ( .A(n527), .B(n287), .S(n69), .Z(n433) );
  MUX2_X1 U310 ( .A(product[6]), .B(n529), .S(n69), .Z(n435) );
  MUX2_X1 U311 ( .A(n529), .B(n530), .S(n69), .Z(n437) );
  MUX2_X1 U312 ( .A(product[7]), .B(n532), .S(n69), .Z(n441) );
  NAND2_X1 U313 ( .A1(n338), .A2(n348), .ZN(n288) );
  XNOR2_X1 U314 ( .A(n350), .B(n288), .ZN(n289) );
  MUX2_X1 U315 ( .A(n532), .B(n289), .S(n69), .Z(n443) );
  MUX2_X1 U316 ( .A(product[8]), .B(n534), .S(n69), .Z(n445) );
  AOI21_X1 U317 ( .B1(n350), .B2(n338), .A(n392), .ZN(n293) );
  NAND2_X1 U318 ( .A1(n393), .A2(n347), .ZN(n291) );
  XOR2_X1 U319 ( .A(n293), .B(n291), .Z(n292) );
  BUF_X4 U320 ( .A(en), .Z(n333) );
  MUX2_X1 U321 ( .A(n534), .B(n292), .S(n333), .Z(n447) );
  MUX2_X1 U322 ( .A(product[9]), .B(n536), .S(n333), .Z(n449) );
  OAI21_X1 U323 ( .B1(n293), .B2(n346), .A(n347), .ZN(n304) );
  INV_X1 U324 ( .A(n304), .ZN(n296) );
  NAND2_X1 U325 ( .A1(n394), .A2(n345), .ZN(n294) );
  XOR2_X1 U326 ( .A(n296), .B(n294), .Z(n295) );
  MUX2_X1 U327 ( .A(n536), .B(n295), .S(n333), .Z(n451) );
  MUX2_X1 U328 ( .A(product[10]), .B(n538), .S(n333), .Z(n453) );
  OAI21_X1 U329 ( .B1(n296), .B2(n344), .A(n345), .ZN(n299) );
  NOR2_X1 U330 ( .A1(n351), .A2(n352), .ZN(n302) );
  INV_X1 U331 ( .A(n302), .ZN(n297) );
  NAND2_X1 U332 ( .A1(n351), .A2(n352), .ZN(n301) );
  NAND2_X1 U333 ( .A1(n297), .A2(n301), .ZN(n298) );
  XNOR2_X1 U334 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U335 ( .A(n538), .B(n300), .S(n333), .Z(n455) );
  MUX2_X1 U336 ( .A(product[11]), .B(n540), .S(n333), .Z(n457) );
  NOR2_X1 U337 ( .A1(n302), .A2(n344), .ZN(n305) );
  OAI21_X1 U338 ( .B1(n302), .B2(n345), .A(n301), .ZN(n303) );
  AOI21_X1 U339 ( .B1(n305), .B2(n304), .A(n303), .ZN(n327) );
  NAND2_X1 U340 ( .A1(n395), .A2(n343), .ZN(n306) );
  XOR2_X1 U341 ( .A(n327), .B(n306), .Z(n307) );
  MUX2_X1 U342 ( .A(n540), .B(n307), .S(n333), .Z(n459) );
  MUX2_X1 U343 ( .A(product[12]), .B(n542), .S(n333), .Z(n461) );
  OAI21_X1 U344 ( .B1(n327), .B2(n342), .A(n343), .ZN(n309) );
  NAND2_X1 U345 ( .A1(n337), .A2(n341), .ZN(n308) );
  XNOR2_X1 U346 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U347 ( .A(n542), .B(n310), .S(n333), .Z(n463) );
  MUX2_X1 U348 ( .A(product[13]), .B(n544), .S(n333), .Z(n465) );
  NAND2_X1 U349 ( .A1(n395), .A2(n337), .ZN(n312) );
  AOI21_X1 U350 ( .B1(n390), .B2(n337), .A(n396), .ZN(n311) );
  OAI21_X1 U351 ( .B1(n327), .B2(n312), .A(n311), .ZN(n314) );
  NAND2_X1 U352 ( .A1(n336), .A2(n349), .ZN(n313) );
  XNOR2_X1 U353 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U354 ( .A(n544), .B(n315), .S(n333), .Z(n467) );
  MUX2_X1 U355 ( .A(product[14]), .B(n546), .S(n333), .Z(n469) );
  NAND2_X1 U356 ( .A1(n337), .A2(n336), .ZN(n317) );
  NOR2_X1 U357 ( .A1(n342), .A2(n317), .ZN(n323) );
  INV_X1 U358 ( .A(n323), .ZN(n319) );
  AOI21_X1 U359 ( .B1(n396), .B2(n336), .A(n391), .ZN(n316) );
  OAI21_X1 U360 ( .B1(n317), .B2(n343), .A(n316), .ZN(n324) );
  INV_X1 U361 ( .A(n324), .ZN(n318) );
  OAI21_X1 U362 ( .B1(n327), .B2(n319), .A(n318), .ZN(n321) );
  NAND2_X1 U363 ( .A1(n335), .A2(n340), .ZN(n320) );
  XNOR2_X1 U364 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U365 ( .A(n546), .B(n322), .S(n333), .Z(n471) );
  MUX2_X1 U366 ( .A(product[15]), .B(n548), .S(n333), .Z(n473) );
  NAND2_X1 U367 ( .A1(n323), .A2(n335), .ZN(n326) );
  AOI21_X1 U368 ( .B1(n324), .B2(n335), .A(n389), .ZN(n325) );
  OAI21_X1 U369 ( .B1(n327), .B2(n326), .A(n325), .ZN(n328) );
  XNOR2_X1 U370 ( .A(n328), .B(n339), .ZN(n329) );
  MUX2_X1 U371 ( .A(n548), .B(n329), .S(n333), .Z(n475) );
  MUX2_X1 U372 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n333), .Z(n477) );
  MUX2_X1 U373 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n333), .Z(n479) );
  MUX2_X1 U374 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n333), .Z(n481) );
  MUX2_X1 U375 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n333), .Z(n483) );
  MUX2_X1 U376 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n333), .Z(n485) );
  MUX2_X1 U377 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n333), .Z(n487) );
  MUX2_X1 U378 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n333), .Z(n489) );
  MUX2_X1 U379 ( .A(n19), .B(B_extended[7]), .S(n333), .Z(n491) );
  MUX2_X1 U380 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n333), .Z(n493) );
  MUX2_X1 U381 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n333), .Z(n495) );
  MUX2_X1 U382 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n333), .Z(n497) );
  MUX2_X1 U383 ( .A(n330), .B(A_extended[3]), .S(n333), .Z(n499) );
  MUX2_X1 U384 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n333), .Z(n501) );
  MUX2_X1 U385 ( .A(n331), .B(A_extended[5]), .S(n333), .Z(n503) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n333), .Z(n505) );
  MUX2_X1 U387 ( .A(n332), .B(A_extended[7]), .S(n333), .Z(n507) );
  OR2_X1 U388 ( .A1(n333), .A2(n551), .ZN(n509) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_19 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n368, n370, n372, n374, n376, n378, n380,
         n382, n384, n386, n388, n390, n392, n394, n396, n398, n400, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n412, n414, n416,
         n418, n420, n422, n424, n426, n428, n430, n432, n434, n436, n438,
         n440, n442, n444, n446, n448, n450, n452, n454, n456, n458, n460,
         n462, n464, n466, n468, n470, n472, n474, n476, n478, n480, n482,
         n484, n486, n488, n490, n492, n494, n496, n498, n500, n502, n504,
         n506, n508, n510, n512, n514, n516, n518, n520, n522, n524, n525,
         n527, n528, n530, n531, n533, n534, n536, n537, n539, n540, n542,
         n543, n545, n547, n549, n551, n553, n555, n557, n559, n561, n562,
         n563, n564, n565;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n271), .SE(n522), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n410), .SE(n518), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n27) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n410), .SE(n516), .CK(clk), .Q(n562), 
        .QN(n30) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n410), .SE(n514), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n26) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n410), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n25) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n410), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n28) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n410), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n410), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n17) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n410), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n22) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n410), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n23) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n271), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n18) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n271), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n19) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n271), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n21) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n271), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n20) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n271), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n271), .SE(n488), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n271), .SE(n486), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n271), .SE(n484), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n271), .SE(n482), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n271), .SE(n480), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n271), .SE(n478), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n410), .SE(n476), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n410), .SE(n474), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n410), .SE(n472), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n410), .SE(n470), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n271), .SE(n468), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n410), .SE(n466), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n410), .SE(n464), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n271), .SE(n462), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n410), .SE(n460), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n410), .SE(n458), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n410), .SE(n456), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n410), .SE(n454), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n410), .SE(n450), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n271), .SE(n448), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n271), .SE(n446), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n410), .SE(n444), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n271), .SE(n442), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n410), .SE(n440), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n410), .SE(n438), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n410), .SE(n436), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n410), .SE(n434), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n410), .SE(n432), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n410), .SE(n430), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n410), .SE(n428), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n410), .SE(n426), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n410), .SE(n424), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n410), .SE(n422), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n410), .SE(n420), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n410), .SE(n418), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n410), .SE(n416), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n410), .SE(n414), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n410), .SE(n412), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n410), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n32) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n410), .SE(n520), .CK(clk), .Q(n563), 
        .QN(n29) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n565), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n365) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n565), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n364) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n565), .SE(n396), .CK(
        clk), .QN(n363) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n565), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n362), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n565), .SE(n392), .CK(
        clk), .Q(n408), .QN(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n565), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n360), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n565), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n359), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n565), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n565), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n357), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n565), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n565), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n355), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n565), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n354), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n565), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n353), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n565), .SE(n374), .CK(
        clk), .QN(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n565), .SE(n372), .CK(
        clk), .QN(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n565), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n350), .QN(n31) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n565), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n565), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n348) );
  SDFF_X2 clk_r_REG37_S2 ( .D(1'b0), .SI(n410), .SE(n452), .CK(clk), .Q(n543)
         );
  BUF_X1 U2 ( .A(n563), .Z(n11) );
  BUF_X1 U3 ( .A(\mult_x_1/n313 ), .Z(n128) );
  BUF_X1 U4 ( .A(n272), .Z(n268) );
  CLKBUF_X2 U5 ( .A(n272), .Z(n301) );
  CLKBUF_X2 U6 ( .A(n272), .Z(n303) );
  AND2_X1 U7 ( .A1(n115), .A2(n114), .ZN(n15) );
  NAND2_X1 U8 ( .A1(n71), .A2(n70), .ZN(n163) );
  INV_X1 U9 ( .A(n163), .ZN(n168) );
  OAI22_X1 U10 ( .A1(n211), .A2(n75), .B1(n209), .B2(n76), .ZN(n78) );
  NAND2_X1 U11 ( .A1(n63), .A2(n62), .ZN(n50) );
  NAND2_X1 U12 ( .A1(n126), .A2(n124), .ZN(n66) );
  CLKBUF_X1 U13 ( .A(n563), .Z(n346) );
  XNOR2_X1 U14 ( .A(n163), .B(n73), .ZN(n178) );
  NAND2_X1 U15 ( .A1(n138), .A2(n137), .ZN(n56) );
  NOR2_X1 U16 ( .A1(n138), .A2(n137), .ZN(n57) );
  INV_X1 U17 ( .A(n140), .ZN(n58) );
  NAND2_X1 U18 ( .A1(n84), .A2(n83), .ZN(n87) );
  NAND2_X1 U19 ( .A1(n92), .A2(n82), .ZN(n84) );
  XNOR2_X1 U20 ( .A(n92), .B(n91), .ZN(n118) );
  OAI21_X1 U21 ( .B1(n168), .B2(n167), .A(n166), .ZN(n236) );
  XNOR2_X1 U22 ( .A(n140), .B(n139), .ZN(n258) );
  XNOR2_X1 U23 ( .A(n138), .B(n137), .ZN(n139) );
  NAND2_X1 U24 ( .A1(n69), .A2(n68), .ZN(n370) );
  OR2_X1 U25 ( .A1(n268), .A2(n31), .ZN(n68) );
  BUF_X1 U26 ( .A(n37), .Z(n6) );
  NAND2_X2 U27 ( .A1(n7), .A2(n5), .ZN(n176) );
  NAND2_X1 U28 ( .A1(n36), .A2(n6), .ZN(n13) );
  INV_X1 U29 ( .A(n32), .ZN(n7) );
  INV_X1 U30 ( .A(n40), .ZN(n8) );
  OAI21_X1 U31 ( .B1(n292), .B2(n289), .A(n290), .ZN(n9) );
  OAI21_X1 U32 ( .B1(n292), .B2(n289), .A(n290), .ZN(n10) );
  XNOR2_X1 U33 ( .A(n25), .B(n17), .ZN(n55) );
  OAI21_X1 U34 ( .B1(n45), .B2(n213), .A(n42), .ZN(n12) );
  OAI21_X1 U35 ( .B1(n251), .B2(n250), .A(n268), .ZN(n69) );
  NAND2_X1 U36 ( .A1(n36), .A2(n6), .ZN(n189) );
  XNOR2_X1 U37 ( .A(n14), .B(n255), .ZN(n122) );
  NAND2_X1 U38 ( .A1(n253), .A2(n254), .ZN(n14) );
  XNOR2_X1 U39 ( .A(n90), .B(n89), .ZN(n91) );
  NAND2_X1 U40 ( .A1(n90), .A2(n89), .ZN(n83) );
  OR2_X1 U41 ( .A1(n90), .A2(n89), .ZN(n82) );
  NAND2_X1 U42 ( .A1(n165), .A2(n164), .ZN(n166) );
  NOR2_X1 U43 ( .A1(n165), .A2(n164), .ZN(n167) );
  AND2_X1 U44 ( .A1(n217), .A2(n216), .ZN(n227) );
  OAI21_X1 U45 ( .B1(n126), .B2(n124), .A(n123), .ZN(n67) );
  XOR2_X1 U46 ( .A(n115), .B(n114), .Z(n108) );
  AOI21_X1 U47 ( .B1(n296), .B2(n9), .A(n119), .ZN(n16) );
  NOR2_X2 U48 ( .A1(n110), .A2(n109), .ZN(n292) );
  AND2_X1 U49 ( .A1(n219), .A2(n218), .ZN(n24) );
  INV_X1 U50 ( .A(rst_n), .ZN(n565) );
  BUF_X2 U51 ( .A(n562), .Z(n345) );
  OR2_X1 U52 ( .A1(n63), .A2(n62), .ZN(n33) );
  XNOR2_X1 U53 ( .A(n562), .B(n26), .ZN(n34) );
  XNOR2_X1 U54 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n35) );
  NAND2_X2 U55 ( .A1(n34), .A2(n35), .ZN(n211) );
  XNOR2_X1 U56 ( .A(n345), .B(\mult_x_1/n281 ), .ZN(n48) );
  AND2_X1 U57 ( .A1(n564), .A2(\mult_x_1/n281 ), .ZN(n144) );
  XNOR2_X1 U58 ( .A(n144), .B(n345), .ZN(n147) );
  BUF_X2 U59 ( .A(n35), .Z(n209) );
  OAI22_X1 U60 ( .A1(n211), .A2(n48), .B1(n147), .B2(n209), .ZN(n152) );
  INV_X1 U61 ( .A(n152), .ZN(n151) );
  XNOR2_X1 U62 ( .A(n346), .B(n27), .ZN(n36) );
  XNOR2_X1 U63 ( .A(n562), .B(\mult_x_1/a[6] ), .ZN(n37) );
  XNOR2_X1 U64 ( .A(n11), .B(\mult_x_1/n283 ), .ZN(n39) );
  INV_X1 U65 ( .A(n37), .ZN(n72) );
  INV_X2 U66 ( .A(n72), .ZN(n190) );
  XNOR2_X1 U67 ( .A(n11), .B(\mult_x_1/n282 ), .ZN(n146) );
  OAI22_X1 U68 ( .A1(n13), .A2(n39), .B1(n190), .B2(n146), .ZN(n150) );
  AND2_X1 U69 ( .A1(n564), .A2(n563), .ZN(n38) );
  XNOR2_X1 U70 ( .A(n38), .B(n346), .ZN(n130) );
  BUF_X1 U71 ( .A(n130), .Z(n192) );
  NOR2_X1 U72 ( .A1(n18), .A2(n192), .ZN(n149) );
  XNOR2_X1 U73 ( .A(n11), .B(\mult_x_1/n284 ), .ZN(n47) );
  OAI22_X1 U74 ( .A1(n13), .A2(n47), .B1(n190), .B2(n39), .ZN(n61) );
  CLKBUF_X1 U75 ( .A(\mult_x_1/n312 ), .Z(n99) );
  XNOR2_X1 U76 ( .A(n144), .B(n99), .ZN(n45) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n44) );
  INV_X1 U78 ( .A(n44), .ZN(n40) );
  INV_X2 U79 ( .A(n40), .ZN(n213) );
  CLKBUF_X1 U80 ( .A(\mult_x_1/n312 ), .Z(n344) );
  INV_X1 U81 ( .A(n55), .ZN(n41) );
  XNOR2_X1 U82 ( .A(\mult_x_1/n312 ), .B(n28), .ZN(n43) );
  NAND3_X1 U83 ( .A1(n8), .A2(n41), .A3(n43), .ZN(n42) );
  OAI21_X1 U84 ( .B1(n45), .B2(n213), .A(n42), .ZN(n60) );
  NAND2_X1 U85 ( .A1(n44), .A2(n43), .ZN(n215) );
  AOI21_X1 U86 ( .B1(n213), .B2(n215), .A(n45), .ZN(n46) );
  INV_X1 U87 ( .A(n46), .ZN(n59) );
  XNOR2_X1 U88 ( .A(n11), .B(\mult_x_1/n285 ), .ZN(n53) );
  OAI22_X1 U89 ( .A1(n189), .A2(n53), .B1(n190), .B2(n47), .ZN(n136) );
  XNOR2_X1 U90 ( .A(n345), .B(\mult_x_1/n283 ), .ZN(n54) );
  XNOR2_X1 U91 ( .A(n345), .B(\mult_x_1/n282 ), .ZN(n49) );
  OAI22_X1 U92 ( .A1(n211), .A2(n54), .B1(n209), .B2(n49), .ZN(n135) );
  INV_X1 U93 ( .A(n60), .ZN(n134) );
  NOR2_X1 U94 ( .A1(n19), .A2(n192), .ZN(n63) );
  OAI22_X1 U95 ( .A1(n211), .A2(n49), .B1(n209), .B2(n48), .ZN(n62) );
  NAND2_X1 U96 ( .A1(n65), .A2(n33), .ZN(n51) );
  NAND2_X1 U97 ( .A1(n51), .A2(n50), .ZN(n159) );
  XNOR2_X1 U98 ( .A(n144), .B(n128), .ZN(n129) );
  AOI21_X1 U99 ( .B1(n176), .B2(n5), .A(n129), .ZN(n52) );
  INV_X1 U100 ( .A(n52), .ZN(n207) );
  XNOR2_X1 U101 ( .A(n11), .B(\mult_x_1/n286 ), .ZN(n127) );
  OAI22_X1 U102 ( .A1(n13), .A2(n127), .B1(n190), .B2(n53), .ZN(n206) );
  NOR2_X1 U103 ( .A1(n20), .A2(n192), .ZN(n205) );
  XNOR2_X1 U104 ( .A(n345), .B(\mult_x_1/n284 ), .ZN(n208) );
  OAI22_X1 U105 ( .A1(n211), .A2(n208), .B1(n209), .B2(n54), .ZN(n133) );
  XNOR2_X1 U106 ( .A(n344), .B(\mult_x_1/n282 ), .ZN(n212) );
  OAI22_X1 U107 ( .A1(n215), .A2(n212), .B1(n213), .B2(n55), .ZN(n132) );
  OR2_X1 U108 ( .A1(n133), .A2(n132), .ZN(n138) );
  NOR2_X1 U109 ( .A1(n21), .A2(n192), .ZN(n137) );
  OAI21_X1 U110 ( .B1(n58), .B2(n57), .A(n56), .ZN(n126) );
  FA_X1 U111 ( .A(n61), .B(n12), .CI(n59), .CO(n160), .S(n124) );
  XNOR2_X1 U112 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U113 ( .A(n65), .B(n64), .ZN(n123) );
  NAND2_X1 U114 ( .A1(n67), .A2(n66), .ZN(n250) );
  CLKBUF_X1 U115 ( .A(en), .Z(n272) );
  XNOR2_X1 U116 ( .A(n99), .B(\mult_x_1/n285 ), .ZN(n80) );
  OR2_X1 U117 ( .A1(n215), .A2(n80), .ZN(n71) );
  XNOR2_X1 U118 ( .A(n344), .B(\mult_x_1/n284 ), .ZN(n177) );
  OR2_X1 U119 ( .A1(n213), .A2(n177), .ZN(n70) );
  XNOR2_X1 U120 ( .A(n128), .B(\mult_x_1/n283 ), .ZN(n81) );
  XNOR2_X1 U121 ( .A(n128), .B(\mult_x_1/n282 ), .ZN(n175) );
  OAI22_X1 U122 ( .A1(n176), .A2(n81), .B1(n175), .B2(n5), .ZN(n165) );
  AND2_X1 U123 ( .A1(\mult_x_1/n288 ), .A2(n72), .ZN(n164) );
  XNOR2_X1 U124 ( .A(n165), .B(n164), .ZN(n73) );
  OR2_X1 U125 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n74) );
  OAI22_X1 U126 ( .A1(n211), .A2(n30), .B1(n74), .B2(n209), .ZN(n79) );
  XNOR2_X1 U127 ( .A(n345), .B(\mult_x_1/n288 ), .ZN(n75) );
  XNOR2_X1 U128 ( .A(n345), .B(\mult_x_1/n287 ), .ZN(n76) );
  XNOR2_X1 U129 ( .A(n345), .B(\mult_x_1/n286 ), .ZN(n172) );
  OAI22_X1 U130 ( .A1(n211), .A2(n76), .B1(n209), .B2(n172), .ZN(n179) );
  XNOR2_X1 U131 ( .A(n180), .B(n179), .ZN(n77) );
  XNOR2_X1 U132 ( .A(n178), .B(n77), .ZN(n88) );
  INV_X1 U133 ( .A(n88), .ZN(n86) );
  HA_X1 U134 ( .A(n79), .B(n78), .CO(n180), .S(n92) );
  XNOR2_X1 U135 ( .A(n99), .B(\mult_x_1/n286 ), .ZN(n95) );
  OAI22_X1 U136 ( .A1(n215), .A2(n95), .B1(n213), .B2(n80), .ZN(n90) );
  XNOR2_X1 U137 ( .A(n128), .B(\mult_x_1/n284 ), .ZN(n93) );
  OAI22_X1 U138 ( .A1(n176), .A2(n93), .B1(n81), .B2(n5), .ZN(n89) );
  INV_X1 U139 ( .A(n87), .ZN(n85) );
  NAND2_X1 U140 ( .A1(n86), .A2(n85), .ZN(n253) );
  NAND2_X1 U141 ( .A1(n88), .A2(n87), .ZN(n254) );
  XNOR2_X1 U142 ( .A(n128), .B(\mult_x_1/n285 ), .ZN(n98) );
  OAI22_X1 U143 ( .A1(n176), .A2(n98), .B1(n93), .B2(n5), .ZN(n113) );
  INV_X1 U144 ( .A(n209), .ZN(n94) );
  AND2_X1 U145 ( .A1(\mult_x_1/n288 ), .A2(n94), .ZN(n112) );
  XNOR2_X1 U146 ( .A(n99), .B(\mult_x_1/n287 ), .ZN(n96) );
  OAI22_X1 U147 ( .A1(n215), .A2(n96), .B1(n213), .B2(n95), .ZN(n111) );
  OR2_X1 U148 ( .A1(n118), .A2(n117), .ZN(n296) );
  XNOR2_X1 U149 ( .A(n344), .B(\mult_x_1/n288 ), .ZN(n97) );
  OAI22_X1 U150 ( .A1(n215), .A2(n97), .B1(n213), .B2(n96), .ZN(n115) );
  XNOR2_X1 U151 ( .A(n128), .B(\mult_x_1/n286 ), .ZN(n101) );
  OAI22_X1 U152 ( .A1(n176), .A2(n101), .B1(n98), .B2(n5), .ZN(n114) );
  OR2_X1 U153 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n100) );
  OAI22_X1 U154 ( .A1(n215), .A2(n25), .B1(n100), .B2(n213), .ZN(n107) );
  OR2_X1 U155 ( .A1(n108), .A2(n107), .ZN(n285) );
  XNOR2_X1 U156 ( .A(n128), .B(\mult_x_1/n287 ), .ZN(n103) );
  OAI22_X1 U157 ( .A1(n176), .A2(n103), .B1(n101), .B2(n5), .ZN(n106) );
  INV_X1 U158 ( .A(n213), .ZN(n102) );
  AND2_X1 U159 ( .A1(\mult_x_1/n288 ), .A2(n102), .ZN(n105) );
  NOR2_X1 U160 ( .A1(n106), .A2(n105), .ZN(n278) );
  OAI22_X1 U161 ( .A1(n176), .A2(\mult_x_1/n288 ), .B1(n103), .B2(n5), .ZN(
        n275) );
  OR2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n104) );
  NAND2_X1 U163 ( .A1(n104), .A2(n176), .ZN(n274) );
  NAND2_X1 U164 ( .A1(n275), .A2(n274), .ZN(n281) );
  NAND2_X1 U165 ( .A1(n106), .A2(n105), .ZN(n279) );
  OAI21_X1 U166 ( .B1(n278), .B2(n281), .A(n279), .ZN(n286) );
  AND2_X1 U167 ( .A1(n285), .A2(n286), .ZN(n110) );
  NAND2_X1 U168 ( .A1(n108), .A2(n107), .ZN(n284) );
  INV_X1 U169 ( .A(n284), .ZN(n109) );
  FA_X1 U170 ( .A(n113), .B(n112), .CI(n111), .CO(n117), .S(n116) );
  NOR2_X1 U171 ( .A1(n116), .A2(n15), .ZN(n289) );
  NAND2_X1 U172 ( .A1(n116), .A2(n15), .ZN(n290) );
  OAI21_X1 U173 ( .B1(n292), .B2(n289), .A(n290), .ZN(n297) );
  NAND2_X1 U174 ( .A1(n118), .A2(n117), .ZN(n295) );
  INV_X1 U175 ( .A(n295), .ZN(n119) );
  AOI21_X1 U176 ( .B1(n296), .B2(n10), .A(n119), .ZN(n255) );
  INV_X1 U177 ( .A(n303), .ZN(n121) );
  NAND2_X1 U178 ( .A1(n121), .A2(n543), .ZN(n120) );
  OAI21_X1 U179 ( .B1(n122), .B2(n121), .A(n120), .ZN(n452) );
  XNOR2_X1 U180 ( .A(n124), .B(n123), .ZN(n125) );
  XNOR2_X1 U181 ( .A(n126), .B(n125), .ZN(n248) );
  XNOR2_X1 U182 ( .A(n11), .B(\mult_x_1/n287 ), .ZN(n170) );
  OAI22_X1 U183 ( .A1(n13), .A2(n170), .B1(n190), .B2(n127), .ZN(n223) );
  XNOR2_X1 U184 ( .A(n128), .B(\mult_x_1/n281 ), .ZN(n174) );
  OAI22_X1 U185 ( .A1(n176), .A2(n174), .B1(n129), .B2(n5), .ZN(n222) );
  INV_X1 U186 ( .A(n130), .ZN(n131) );
  AND2_X1 U187 ( .A1(\mult_x_1/n288 ), .A2(n131), .ZN(n221) );
  XNOR2_X1 U188 ( .A(n133), .B(n132), .ZN(n218) );
  FA_X1 U189 ( .A(n136), .B(n135), .CI(n134), .CO(n65), .S(n259) );
  NAND2_X1 U190 ( .A1(n248), .A2(n247), .ZN(n141) );
  NAND2_X1 U191 ( .A1(n141), .A2(n268), .ZN(n143) );
  NAND2_X1 U192 ( .A1(n121), .A2(n354), .ZN(n142) );
  NAND2_X1 U193 ( .A1(n143), .A2(n142), .ZN(n378) );
  NOR2_X1 U212 ( .A1(n22), .A2(n192), .ZN(n187) );
  XNOR2_X1 U213 ( .A(n11), .B(\mult_x_1/n281 ), .ZN(n145) );
  XNOR2_X1 U214 ( .A(n144), .B(n11), .ZN(n188) );
  OAI22_X1 U215 ( .A1(n13), .A2(n145), .B1(n188), .B2(n190), .ZN(n196) );
  INV_X1 U216 ( .A(n196), .ZN(n186) );
  OAI22_X1 U217 ( .A1(n13), .A2(n146), .B1(n190), .B2(n145), .ZN(n154) );
  AOI21_X1 U218 ( .B1(n209), .B2(n211), .A(n147), .ZN(n148) );
  INV_X1 U219 ( .A(n148), .ZN(n153) );
  FA_X1 U220 ( .A(n151), .B(n150), .CI(n149), .CO(n158), .S(n161) );
  NOR2_X1 U221 ( .A1(n23), .A2(n192), .ZN(n157) );
  FA_X1 U222 ( .A(n154), .B(n153), .CI(n152), .CO(n185), .S(n156) );
  OR2_X1 U223 ( .A1(n203), .A2(n202), .ZN(n155) );
  MUX2_X1 U224 ( .A(n348), .B(n155), .S(n268), .Z(n366) );
  FA_X1 U225 ( .A(n158), .B(n157), .CI(n156), .CO(n202), .S(n245) );
  FA_X1 U226 ( .A(n161), .B(n160), .CI(n159), .CO(n244), .S(n251) );
  OR2_X1 U227 ( .A1(n245), .A2(n244), .ZN(n162) );
  MUX2_X1 U228 ( .A(n349), .B(n162), .S(n268), .Z(n368) );
  OR2_X1 U229 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n169) );
  OAI22_X1 U230 ( .A1(n189), .A2(n29), .B1(n169), .B2(n190), .ZN(n217) );
  XNOR2_X1 U231 ( .A(n11), .B(\mult_x_1/n288 ), .ZN(n171) );
  OAI22_X1 U232 ( .A1(n189), .A2(n171), .B1(n190), .B2(n170), .ZN(n216) );
  XOR2_X1 U233 ( .A(n217), .B(n216), .Z(n235) );
  XNOR2_X1 U234 ( .A(n345), .B(\mult_x_1/n285 ), .ZN(n210) );
  OAI22_X1 U235 ( .A1(n211), .A2(n172), .B1(n209), .B2(n210), .ZN(n226) );
  OAI22_X1 U236 ( .A1(n176), .A2(n175), .B1(n174), .B2(n5), .ZN(n225) );
  XNOR2_X1 U237 ( .A(n344), .B(\mult_x_1/n283 ), .ZN(n214) );
  OAI22_X1 U238 ( .A1(n215), .A2(n177), .B1(n213), .B2(n214), .ZN(n224) );
  NAND2_X1 U239 ( .A1(n178), .A2(n180), .ZN(n183) );
  NAND2_X1 U240 ( .A1(n178), .A2(n179), .ZN(n182) );
  NAND2_X1 U241 ( .A1(n180), .A2(n179), .ZN(n181) );
  NAND3_X1 U242 ( .A1(n183), .A2(n182), .A3(n181), .ZN(n241) );
  OR2_X1 U243 ( .A1(n242), .A2(n241), .ZN(n184) );
  MUX2_X1 U244 ( .A(n351), .B(n184), .S(n268), .Z(n372) );
  FA_X1 U245 ( .A(n187), .B(n186), .CI(n185), .CO(n198), .S(n203) );
  AOI21_X1 U246 ( .B1(n190), .B2(n13), .A(n188), .ZN(n191) );
  INV_X1 U247 ( .A(n191), .ZN(n194) );
  NOR2_X1 U248 ( .A1(n17), .A2(n192), .ZN(n193) );
  XOR2_X1 U249 ( .A(n194), .B(n193), .Z(n195) );
  XOR2_X1 U250 ( .A(n196), .B(n195), .Z(n197) );
  OR2_X1 U251 ( .A1(n198), .A2(n197), .ZN(n200) );
  NAND2_X1 U252 ( .A1(n198), .A2(n197), .ZN(n199) );
  NAND2_X1 U253 ( .A1(n200), .A2(n199), .ZN(n201) );
  MUX2_X1 U254 ( .A(n352), .B(n201), .S(n268), .Z(n374) );
  NAND2_X1 U255 ( .A1(n203), .A2(n202), .ZN(n204) );
  MUX2_X1 U256 ( .A(n353), .B(n204), .S(n268), .Z(n376) );
  FA_X1 U257 ( .A(n207), .B(n206), .CI(n205), .CO(n140), .S(n263) );
  OAI22_X1 U258 ( .A1(n211), .A2(n210), .B1(n209), .B2(n208), .ZN(n229) );
  OAI22_X1 U259 ( .A1(n215), .A2(n214), .B1(n213), .B2(n212), .ZN(n228) );
  INV_X1 U260 ( .A(n218), .ZN(n220) );
  XNOR2_X1 U261 ( .A(n220), .B(n219), .ZN(n261) );
  FA_X1 U262 ( .A(n223), .B(n222), .CI(n221), .CO(n219), .S(n233) );
  FA_X1 U263 ( .A(n226), .B(n225), .CI(n224), .CO(n232), .S(n234) );
  FA_X1 U264 ( .A(n229), .B(n228), .CI(n227), .CO(n262), .S(n231) );
  NOR2_X1 U265 ( .A1(n266), .A2(n265), .ZN(n230) );
  MUX2_X1 U266 ( .A(n355), .B(n230), .S(n268), .Z(n380) );
  FA_X1 U267 ( .A(n233), .B(n232), .CI(n231), .CO(n265), .S(n239) );
  FA_X1 U268 ( .A(n236), .B(n235), .CI(n234), .CO(n238), .S(n242) );
  NOR2_X1 U269 ( .A1(n239), .A2(n238), .ZN(n237) );
  MUX2_X1 U270 ( .A(n357), .B(n237), .S(n268), .Z(n384) );
  NAND2_X1 U271 ( .A1(n239), .A2(n238), .ZN(n240) );
  MUX2_X1 U272 ( .A(n358), .B(n240), .S(n268), .Z(n386) );
  NAND2_X1 U273 ( .A1(n242), .A2(n241), .ZN(n243) );
  MUX2_X1 U274 ( .A(n359), .B(n243), .S(n268), .Z(n388) );
  NAND2_X1 U275 ( .A1(n245), .A2(n244), .ZN(n246) );
  MUX2_X1 U276 ( .A(n360), .B(n246), .S(n301), .Z(n390) );
  NOR2_X1 U277 ( .A1(n248), .A2(n247), .ZN(n249) );
  MUX2_X1 U278 ( .A(n361), .B(n249), .S(n301), .Z(n392) );
  NAND2_X1 U279 ( .A1(n251), .A2(n250), .ZN(n252) );
  MUX2_X1 U280 ( .A(n362), .B(n252), .S(n301), .Z(n394) );
  INV_X1 U281 ( .A(n253), .ZN(n256) );
  OAI21_X1 U282 ( .B1(n256), .B2(n16), .A(n254), .ZN(n257) );
  MUX2_X1 U283 ( .A(n363), .B(n257), .S(n301), .Z(n396) );
  FA_X1 U284 ( .A(n24), .B(n259), .CI(n258), .CO(n247), .S(n260) );
  MUX2_X1 U285 ( .A(n364), .B(n260), .S(n268), .Z(n398) );
  FA_X1 U286 ( .A(n263), .B(n262), .CI(n261), .CO(n264), .S(n266) );
  MUX2_X1 U287 ( .A(n365), .B(n264), .S(n301), .Z(n400) );
  NAND2_X1 U288 ( .A1(n266), .A2(n265), .ZN(n267) );
  NAND2_X1 U289 ( .A1(n267), .A2(n268), .ZN(n270) );
  NAND2_X1 U290 ( .A1(n121), .A2(n356), .ZN(n269) );
  NAND2_X1 U291 ( .A1(n270), .A2(n269), .ZN(n382) );
  BUF_X2 U292 ( .A(rst_n), .Z(n410) );
  BUF_X1 U293 ( .A(rst_n), .Z(n271) );
  MUX2_X1 U294 ( .A(product[0]), .B(n524), .S(n301), .Z(n412) );
  MUX2_X1 U295 ( .A(n524), .B(n525), .S(n301), .Z(n414) );
  AND2_X1 U296 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n273) );
  MUX2_X1 U297 ( .A(n525), .B(n273), .S(n303), .Z(n416) );
  MUX2_X1 U298 ( .A(product[1]), .B(n527), .S(n301), .Z(n418) );
  MUX2_X1 U299 ( .A(n527), .B(n528), .S(n301), .Z(n420) );
  OR2_X1 U300 ( .A1(n275), .A2(n274), .ZN(n276) );
  AND2_X1 U301 ( .A1(n276), .A2(n281), .ZN(n277) );
  MUX2_X1 U302 ( .A(n528), .B(n277), .S(n303), .Z(n422) );
  MUX2_X1 U303 ( .A(product[2]), .B(n530), .S(n303), .Z(n424) );
  MUX2_X1 U304 ( .A(n530), .B(n531), .S(n301), .Z(n426) );
  INV_X1 U305 ( .A(n278), .ZN(n280) );
  NAND2_X1 U306 ( .A1(n280), .A2(n279), .ZN(n282) );
  XOR2_X1 U307 ( .A(n282), .B(n281), .Z(n283) );
  MUX2_X1 U308 ( .A(n531), .B(n283), .S(n303), .Z(n428) );
  MUX2_X1 U309 ( .A(product[3]), .B(n533), .S(n303), .Z(n430) );
  MUX2_X1 U310 ( .A(n533), .B(n534), .S(n301), .Z(n432) );
  NAND2_X1 U311 ( .A1(n285), .A2(n284), .ZN(n287) );
  XNOR2_X1 U312 ( .A(n287), .B(n286), .ZN(n288) );
  MUX2_X1 U313 ( .A(n534), .B(n288), .S(n303), .Z(n434) );
  MUX2_X1 U314 ( .A(product[4]), .B(n536), .S(n303), .Z(n436) );
  MUX2_X1 U315 ( .A(n536), .B(n537), .S(n301), .Z(n438) );
  INV_X1 U316 ( .A(n289), .ZN(n291) );
  NAND2_X1 U317 ( .A1(n291), .A2(n290), .ZN(n293) );
  XOR2_X1 U318 ( .A(n293), .B(n292), .Z(n294) );
  MUX2_X1 U319 ( .A(n537), .B(n294), .S(n303), .Z(n440) );
  MUX2_X1 U320 ( .A(product[5]), .B(n539), .S(n301), .Z(n442) );
  MUX2_X1 U321 ( .A(n539), .B(n540), .S(n303), .Z(n444) );
  NAND2_X1 U322 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U323 ( .A(n298), .B(n297), .ZN(n299) );
  MUX2_X1 U324 ( .A(n540), .B(n299), .S(n301), .Z(n446) );
  MUX2_X1 U325 ( .A(product[6]), .B(n542), .S(n303), .Z(n448) );
  MUX2_X1 U326 ( .A(n542), .B(n543), .S(n301), .Z(n450) );
  MUX2_X1 U327 ( .A(product[7]), .B(n545), .S(n301), .Z(n454) );
  NAND2_X1 U328 ( .A1(n351), .A2(n359), .ZN(n300) );
  XNOR2_X1 U329 ( .A(n363), .B(n300), .ZN(n302) );
  MUX2_X1 U330 ( .A(n545), .B(n302), .S(n301), .Z(n456) );
  MUX2_X1 U331 ( .A(product[8]), .B(n547), .S(n303), .Z(n458) );
  AOI21_X1 U332 ( .B1(n363), .B2(n351), .A(n405), .ZN(n306) );
  NAND2_X1 U333 ( .A1(n406), .A2(n358), .ZN(n304) );
  XOR2_X1 U334 ( .A(n306), .B(n304), .Z(n305) );
  BUF_X2 U335 ( .A(en), .Z(n347) );
  MUX2_X1 U336 ( .A(n547), .B(n305), .S(n347), .Z(n460) );
  MUX2_X1 U337 ( .A(product[9]), .B(n549), .S(n347), .Z(n462) );
  OAI21_X1 U338 ( .B1(n306), .B2(n357), .A(n358), .ZN(n317) );
  INV_X1 U339 ( .A(n317), .ZN(n309) );
  NAND2_X1 U340 ( .A1(n407), .A2(n356), .ZN(n307) );
  XOR2_X1 U341 ( .A(n309), .B(n307), .Z(n308) );
  MUX2_X1 U342 ( .A(n549), .B(n308), .S(n347), .Z(n464) );
  MUX2_X1 U343 ( .A(product[10]), .B(n551), .S(n347), .Z(n466) );
  OAI21_X1 U344 ( .B1(n309), .B2(n355), .A(n356), .ZN(n312) );
  NOR2_X1 U345 ( .A1(n364), .A2(n365), .ZN(n315) );
  INV_X1 U346 ( .A(n315), .ZN(n310) );
  NAND2_X1 U347 ( .A1(n364), .A2(n365), .ZN(n314) );
  NAND2_X1 U348 ( .A1(n310), .A2(n314), .ZN(n311) );
  XNOR2_X1 U349 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U350 ( .A(n551), .B(n313), .S(n347), .Z(n468) );
  MUX2_X1 U351 ( .A(product[11]), .B(n553), .S(n347), .Z(n470) );
  NOR2_X1 U352 ( .A1(n315), .A2(n355), .ZN(n318) );
  OAI21_X1 U353 ( .B1(n315), .B2(n356), .A(n314), .ZN(n316) );
  AOI21_X1 U354 ( .B1(n318), .B2(n317), .A(n316), .ZN(n341) );
  NAND2_X1 U355 ( .A1(n408), .A2(n354), .ZN(n319) );
  XOR2_X1 U356 ( .A(n341), .B(n319), .Z(n320) );
  MUX2_X1 U357 ( .A(n553), .B(n320), .S(n347), .Z(n472) );
  MUX2_X1 U358 ( .A(product[12]), .B(n555), .S(n347), .Z(n474) );
  OAI21_X1 U359 ( .B1(n341), .B2(n361), .A(n354), .ZN(n322) );
  NAND2_X1 U360 ( .A1(n350), .A2(n362), .ZN(n321) );
  XNOR2_X1 U361 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U362 ( .A(n555), .B(n323), .S(n347), .Z(n476) );
  MUX2_X1 U363 ( .A(product[13]), .B(n557), .S(n347), .Z(n478) );
  NAND2_X1 U364 ( .A1(n408), .A2(n350), .ZN(n325) );
  AOI21_X1 U365 ( .B1(n403), .B2(n350), .A(n409), .ZN(n324) );
  OAI21_X1 U366 ( .B1(n341), .B2(n325), .A(n324), .ZN(n327) );
  NAND2_X1 U367 ( .A1(n349), .A2(n360), .ZN(n326) );
  XNOR2_X1 U368 ( .A(n327), .B(n326), .ZN(n328) );
  MUX2_X1 U369 ( .A(n557), .B(n328), .S(n347), .Z(n480) );
  MUX2_X1 U370 ( .A(product[14]), .B(n559), .S(n347), .Z(n482) );
  NAND2_X1 U371 ( .A1(n350), .A2(n349), .ZN(n330) );
  INV_X1 U372 ( .A(n330), .ZN(n336) );
  NAND2_X1 U373 ( .A1(n408), .A2(n336), .ZN(n332) );
  AOI21_X1 U374 ( .B1(n409), .B2(n349), .A(n404), .ZN(n329) );
  OAI21_X1 U375 ( .B1(n330), .B2(n354), .A(n329), .ZN(n338) );
  INV_X1 U376 ( .A(n338), .ZN(n331) );
  OAI21_X1 U377 ( .B1(n341), .B2(n332), .A(n331), .ZN(n334) );
  NAND2_X1 U378 ( .A1(n348), .A2(n353), .ZN(n333) );
  XNOR2_X1 U379 ( .A(n334), .B(n333), .ZN(n335) );
  MUX2_X1 U380 ( .A(n559), .B(n335), .S(n347), .Z(n484) );
  MUX2_X1 U381 ( .A(product[15]), .B(n561), .S(n347), .Z(n486) );
  AND2_X1 U382 ( .A1(n408), .A2(n348), .ZN(n337) );
  NAND2_X1 U383 ( .A1(n337), .A2(n336), .ZN(n340) );
  AOI21_X1 U384 ( .B1(n338), .B2(n348), .A(n402), .ZN(n339) );
  OAI21_X1 U385 ( .B1(n341), .B2(n340), .A(n339), .ZN(n342) );
  XNOR2_X1 U386 ( .A(n342), .B(n352), .ZN(n343) );
  MUX2_X1 U387 ( .A(n561), .B(n343), .S(n347), .Z(n488) );
  MUX2_X1 U388 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n347), .Z(n490) );
  MUX2_X1 U389 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n347), .Z(n492) );
  MUX2_X1 U390 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n347), .Z(n494) );
  MUX2_X1 U391 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n347), .Z(n496) );
  MUX2_X1 U392 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n347), .Z(n498) );
  MUX2_X1 U393 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n347), .Z(n500) );
  MUX2_X1 U394 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n347), .Z(n502) );
  MUX2_X1 U395 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n347), .Z(n504) );
  MUX2_X1 U396 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n347), .Z(n506) );
  MUX2_X1 U397 ( .A(n7), .B(A_extended[1]), .S(n347), .Z(n508) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n347), .Z(n510) );
  MUX2_X1 U399 ( .A(n344), .B(A_extended[3]), .S(n347), .Z(n512) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n347), .Z(n514) );
  MUX2_X1 U401 ( .A(n345), .B(A_extended[5]), .S(n347), .Z(n516) );
  MUX2_X1 U402 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n347), .Z(n518) );
  MUX2_X1 U403 ( .A(n11), .B(A_extended[7]), .S(n347), .Z(n520) );
  OR2_X1 U404 ( .A1(n347), .A2(n564), .ZN(n522) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_20 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n347, n349,
         n351, n353, n355, n357, n359, n361, n363, n365, n367, n369, n371,
         n373, n375, n377, n379, n381, n383, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n396, n398, n400, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n420, n422, n424, n426, n428,
         n430, n432, n434, n436, n438, n440, n442, n444, n446, n448, n450,
         n452, n454, n456, n458, n460, n462, n464, n466, n468, n470, n472,
         n474, n476, n478, n480, n482, n484, n486, n488, n490, n492, n494,
         n496, n498, n500, n502, n504, n506, n507, n509, n510, n512, n513,
         n515, n516, n518, n519, n521, n522, n524, n526, n528, n530, n532,
         n534, n536, n538, n540, n542, n543, n544, n545;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n394), .SE(n504), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n394), .SE(n500), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n394), .SE(n496), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n25) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(n543), 
        .QN(n24) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n394), .SE(n492), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n8) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n394), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n22) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n394), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n23) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n394), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n394), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n19) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n394), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n21) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n394), .SE(n472), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n394), .SE(n470), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n394), .SE(n468), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(rst_n), .SE(n466), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n394), .SE(n464), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n394), .SE(n462), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n394), .SE(n460), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n394), .SE(n458), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n394), .SE(n456), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n394), .SE(n454), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n394), .SE(n450), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n394), .SE(n448), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n394), .SE(n444), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n394), .SE(n442), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n394), .SE(n440), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n438), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n434), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n430), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n428), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n426), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n420), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n418), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n394), .SE(n416), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n394), .SE(n414), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n394), .SE(n412), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n394), .SE(n410), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n394), .SE(n408), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n394), .SE(n406), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n394), .SE(n404), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n394), .SE(n402), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n394), .SE(n400), .CK(clk), .Q(n507)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n394), .SE(n398), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n394), .SE(n396), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n394), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n26) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n545), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n545), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n545), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n545), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n341), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n545), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n340), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n545), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n545), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n338), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n545), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n337), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n545), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n545), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n335), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n545), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n545), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n333), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n545), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n332), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n545), .SE(n357), .CK(
        clk), .Q(n392), .QN(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n545), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n330), .QN(n385) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n545), .SE(n353), .CK(
        clk), .QN(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n545), .SE(n351), .CK(
        clk), .QN(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n545), .SI(1'b1), .SE(n349), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n545), .SI(1'b1), .SE(n347), .CK(clk), 
        .Q(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n545), .SI(1'b1), .SE(n345), .CK(clk), 
        .Q(n325) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n324) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n394), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n323) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n394), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n20) );
  BUF_X1 U2 ( .A(\mult_x_1/n313 ), .Z(n215) );
  BUF_X2 U3 ( .A(en), .Z(n243) );
  INV_X1 U4 ( .A(n26), .ZN(n6) );
  CLKBUF_X1 U5 ( .A(n216), .Z(n12) );
  XNOR2_X1 U6 ( .A(n66), .B(n215), .ZN(n7) );
  XNOR2_X1 U7 ( .A(n8), .B(\mult_x_1/n313 ), .ZN(n37) );
  OR2_X1 U8 ( .A1(n88), .A2(n89), .ZN(n86) );
  OAI22_X1 U9 ( .A1(n139), .A2(n34), .B1(n199), .B2(n69), .ZN(n88) );
  NOR2_X1 U10 ( .A1(n124), .A2(n19), .ZN(n89) );
  OAI22_X1 U11 ( .A1(n122), .A2(n103), .B1(n121), .B2(n102), .ZN(n143) );
  NAND2_X1 U12 ( .A1(n233), .A2(n232), .ZN(n234) );
  INV_X1 U13 ( .A(n237), .ZN(n233) );
  INV_X1 U14 ( .A(n236), .ZN(n232) );
  XNOR2_X1 U15 ( .A(n149), .B(n148), .ZN(n235) );
  CLKBUF_X1 U16 ( .A(n44), .Z(n16) );
  AND2_X1 U17 ( .A1(n544), .A2(\mult_x_1/n310 ), .ZN(n27) );
  XNOR2_X1 U18 ( .A(n236), .B(n237), .ZN(n150) );
  NAND2_X1 U19 ( .A1(n162), .A2(n161), .ZN(n241) );
  NAND2_X1 U20 ( .A1(n165), .A2(n164), .ZN(n161) );
  NAND2_X1 U21 ( .A1(n166), .A2(n160), .ZN(n162) );
  OR2_X1 U22 ( .A1(n165), .A2(n164), .ZN(n160) );
  XNOR2_X1 U23 ( .A(n165), .B(n164), .ZN(n167) );
  NAND2_X1 U24 ( .A1(n89), .A2(n88), .ZN(n90) );
  NAND2_X1 U25 ( .A1(n239), .A2(n238), .ZN(n240) );
  NAND2_X1 U26 ( .A1(n237), .A2(n236), .ZN(n238) );
  NAND2_X1 U27 ( .A1(n235), .A2(n234), .ZN(n239) );
  BUF_X1 U28 ( .A(n73), .Z(n9) );
  AND2_X1 U29 ( .A1(n544), .A2(\mult_x_1/n281 ), .ZN(n66) );
  INV_X1 U30 ( .A(n26), .ZN(n10) );
  INV_X1 U31 ( .A(n20), .ZN(n11) );
  BUF_X2 U32 ( .A(n543), .Z(n13) );
  BUF_X1 U33 ( .A(n543), .Z(n319) );
  AOI21_X1 U34 ( .B1(n260), .B2(n261), .A(n222), .ZN(n14) );
  AOI21_X1 U35 ( .B1(n260), .B2(n261), .A(n222), .ZN(n267) );
  OAI21_X1 U36 ( .B1(n264), .B2(n14), .A(n265), .ZN(n15) );
  MUX2_X1 U37 ( .A(n116), .B(n328), .S(n245), .Z(n351) );
  NAND2_X1 U38 ( .A1(n28), .A2(n29), .ZN(n139) );
  INV_X1 U39 ( .A(n52), .ZN(n17) );
  AND2_X1 U40 ( .A1(n147), .A2(n148), .ZN(n18) );
  INV_X1 U41 ( .A(rst_n), .ZN(n545) );
  INV_X1 U42 ( .A(\mult_x_1/n310 ), .ZN(n102) );
  XNOR2_X1 U43 ( .A(n27), .B(n102), .ZN(n70) );
  INV_X1 U44 ( .A(n70), .ZN(n124) );
  XNOR2_X1 U45 ( .A(\mult_x_1/n311 ), .B(n25), .ZN(n28) );
  XNOR2_X1 U46 ( .A(n543), .B(\mult_x_1/a[4] ), .ZN(n29) );
  INV_X2 U47 ( .A(n323), .ZN(n320) );
  XNOR2_X1 U48 ( .A(n320), .B(\mult_x_1/n282 ), .ZN(n34) );
  INV_X1 U49 ( .A(n29), .ZN(n30) );
  INV_X2 U50 ( .A(n30), .ZN(n199) );
  XNOR2_X1 U51 ( .A(n320), .B(n11), .ZN(n69) );
  XNOR2_X1 U52 ( .A(n89), .B(n88), .ZN(n38) );
  XOR2_X1 U53 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n31) );
  XNOR2_X1 U54 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n32) );
  NAND2_X1 U55 ( .A1(n31), .A2(n32), .ZN(n121) );
  INV_X1 U56 ( .A(n324), .ZN(n321) );
  XNOR2_X1 U57 ( .A(n321), .B(\mult_x_1/n285 ), .ZN(n46) );
  INV_X1 U58 ( .A(n32), .ZN(n33) );
  INV_X2 U59 ( .A(n33), .ZN(n122) );
  XNOR2_X1 U60 ( .A(n321), .B(\mult_x_1/n284 ), .ZN(n39) );
  OAI22_X1 U61 ( .A1(n121), .A2(n46), .B1(n122), .B2(n39), .ZN(n54) );
  XNOR2_X1 U62 ( .A(n320), .B(\mult_x_1/n283 ), .ZN(n42) );
  OAI22_X1 U63 ( .A1(n139), .A2(n42), .B1(n199), .B2(n34), .ZN(n53) );
  XOR2_X1 U64 ( .A(\mult_x_1/a[2] ), .B(n319), .Z(n36) );
  INV_X1 U65 ( .A(n37), .ZN(n35) );
  NAND2_X1 U66 ( .A1(n36), .A2(n35), .ZN(n44) );
  XNOR2_X1 U67 ( .A(n13), .B(n11), .ZN(n43) );
  XNOR2_X1 U68 ( .A(n66), .B(n13), .ZN(n40) );
  INV_X2 U69 ( .A(n37), .ZN(n212) );
  OAI22_X1 U70 ( .A1(n44), .A2(n43), .B1(n40), .B2(n212), .ZN(n81) );
  INV_X1 U71 ( .A(n81), .ZN(n52) );
  XNOR2_X1 U72 ( .A(n38), .B(n87), .ZN(n96) );
  XNOR2_X1 U73 ( .A(n321), .B(\mult_x_1/n283 ), .ZN(n72) );
  OAI22_X1 U74 ( .A1(n121), .A2(n39), .B1(n122), .B2(n72), .ZN(n82) );
  CLKBUF_X2 U75 ( .A(n44), .Z(n210) );
  AOI21_X1 U76 ( .B1(n212), .B2(n210), .A(n40), .ZN(n41) );
  INV_X1 U77 ( .A(n41), .ZN(n80) );
  XNOR2_X1 U78 ( .A(n96), .B(n97), .ZN(n47) );
  XNOR2_X1 U79 ( .A(n320), .B(\mult_x_1/n284 ), .ZN(n137) );
  OAI22_X1 U80 ( .A1(n139), .A2(n137), .B1(n199), .B2(n42), .ZN(n49) );
  XNOR2_X1 U81 ( .A(n13), .B(\mult_x_1/n282 ), .ZN(n140) );
  OAI22_X1 U82 ( .A1(n16), .A2(n140), .B1(n212), .B2(n43), .ZN(n48) );
  OR2_X1 U83 ( .A1(n49), .A2(n48), .ZN(n57) );
  NOR2_X1 U84 ( .A1(n21), .A2(n124), .ZN(n56) );
  NAND2_X1 U85 ( .A1(n215), .A2(n5), .ZN(n216) );
  XNOR2_X1 U86 ( .A(n66), .B(n6), .ZN(n50) );
  AOI21_X1 U87 ( .B1(n216), .B2(n5), .A(n7), .ZN(n45) );
  INV_X1 U88 ( .A(n45), .ZN(n146) );
  AND2_X1 U89 ( .A1(n70), .A2(\mult_x_1/n287 ), .ZN(n145) );
  XNOR2_X1 U90 ( .A(n321), .B(\mult_x_1/n286 ), .ZN(n51) );
  OAI22_X1 U91 ( .A1(n121), .A2(n51), .B1(n122), .B2(n46), .ZN(n144) );
  XNOR2_X1 U92 ( .A(n47), .B(n98), .ZN(n63) );
  INV_X1 U93 ( .A(n243), .ZN(n245) );
  NAND2_X1 U94 ( .A1(n245), .A2(n332), .ZN(n59) );
  XNOR2_X1 U95 ( .A(n49), .B(n48), .ZN(n147) );
  AND2_X1 U96 ( .A1(\mult_x_1/n288 ), .A2(n70), .ZN(n156) );
  XNOR2_X1 U97 ( .A(n215), .B(n11), .ZN(n106) );
  OAI22_X1 U98 ( .A1(n216), .A2(n106), .B1(n50), .B2(n5), .ZN(n155) );
  XNOR2_X1 U99 ( .A(n321), .B(\mult_x_1/n287 ), .ZN(n104) );
  OAI22_X1 U100 ( .A1(n121), .A2(n104), .B1(n122), .B2(n51), .ZN(n154) );
  FA_X1 U101 ( .A(n54), .B(n53), .CI(n52), .CO(n87), .S(n230) );
  FA_X1 U102 ( .A(n57), .B(n56), .CI(n55), .CO(n98), .S(n229) );
  NAND2_X1 U103 ( .A1(n61), .A2(n243), .ZN(n58) );
  OAI211_X1 U104 ( .C1(n63), .C2(n245), .A(n59), .B(n58), .ZN(n359) );
  INV_X1 U105 ( .A(n60), .ZN(n61) );
  NAND2_X1 U106 ( .A1(n61), .A2(n243), .ZN(n64) );
  NAND2_X1 U107 ( .A1(n245), .A2(n331), .ZN(n62) );
  OAI21_X1 U108 ( .B1(n64), .B2(n63), .A(n62), .ZN(n357) );
  NOR2_X1 U129 ( .A1(n22), .A2(n124), .ZN(n119) );
  XNOR2_X1 U130 ( .A(n321), .B(n11), .ZN(n65) );
  XNOR2_X1 U131 ( .A(n66), .B(n321), .ZN(n120) );
  OAI22_X1 U132 ( .A1(n121), .A2(n65), .B1(n120), .B2(n122), .ZN(n128) );
  INV_X1 U133 ( .A(n128), .ZN(n118) );
  XNOR2_X1 U134 ( .A(n321), .B(\mult_x_1/n282 ), .ZN(n71) );
  OAI22_X1 U135 ( .A1(n121), .A2(n71), .B1(n122), .B2(n65), .ZN(n75) );
  XNOR2_X1 U136 ( .A(n66), .B(\mult_x_1/n311 ), .ZN(n68) );
  AOI21_X1 U137 ( .B1(n199), .B2(n139), .A(n68), .ZN(n67) );
  INV_X1 U138 ( .A(n67), .ZN(n74) );
  OAI22_X1 U139 ( .A1(n139), .A2(n69), .B1(n68), .B2(n199), .ZN(n73) );
  AND2_X1 U140 ( .A1(n70), .A2(\mult_x_1/n284 ), .ZN(n85) );
  OAI22_X1 U141 ( .A1(n121), .A2(n72), .B1(n122), .B2(n71), .ZN(n84) );
  INV_X1 U142 ( .A(n73), .ZN(n83) );
  NOR2_X1 U143 ( .A1(n23), .A2(n124), .ZN(n78) );
  FA_X1 U144 ( .A(n75), .B(n74), .CI(n9), .CO(n117), .S(n77) );
  OR2_X1 U145 ( .A1(n135), .A2(n134), .ZN(n76) );
  MUX2_X1 U146 ( .A(n325), .B(n76), .S(n243), .Z(n345) );
  FA_X1 U147 ( .A(n79), .B(n78), .CI(n77), .CO(n134), .S(n190) );
  FA_X1 U148 ( .A(n82), .B(n17), .CI(n80), .CO(n95), .S(n97) );
  FA_X1 U149 ( .A(n85), .B(n84), .CI(n83), .CO(n79), .S(n94) );
  NAND2_X1 U150 ( .A1(n87), .A2(n86), .ZN(n91) );
  NAND2_X1 U151 ( .A1(n91), .A2(n90), .ZN(n93) );
  OR2_X1 U152 ( .A1(n190), .A2(n189), .ZN(n92) );
  MUX2_X1 U153 ( .A(n326), .B(n92), .S(n243), .Z(n347) );
  FA_X1 U154 ( .A(n94), .B(n95), .CI(n93), .CO(n189), .S(n193) );
  OAI21_X1 U155 ( .B1(n98), .B2(n97), .A(n96), .ZN(n100) );
  NAND2_X1 U156 ( .A1(n98), .A2(n97), .ZN(n99) );
  NAND2_X1 U157 ( .A1(n100), .A2(n99), .ZN(n192) );
  OR2_X1 U158 ( .A1(n193), .A2(n192), .ZN(n101) );
  MUX2_X1 U159 ( .A(n327), .B(n101), .S(n243), .Z(n349) );
  XNOR2_X1 U160 ( .A(n6), .B(\mult_x_1/n283 ), .ZN(n182) );
  XNOR2_X1 U161 ( .A(n215), .B(\mult_x_1/n282 ), .ZN(n107) );
  OAI22_X1 U162 ( .A1(n216), .A2(n182), .B1(n107), .B2(n5), .ZN(n115) );
  AND2_X1 U163 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n114) );
  XNOR2_X1 U164 ( .A(n13), .B(\mult_x_1/n285 ), .ZN(n181) );
  XNOR2_X1 U165 ( .A(n13), .B(\mult_x_1/n284 ), .ZN(n108) );
  OAI22_X1 U166 ( .A1(n210), .A2(n181), .B1(n212), .B2(n108), .ZN(n113) );
  OR2_X1 U167 ( .A1(\mult_x_1/n288 ), .A2(n102), .ZN(n103) );
  XNOR2_X1 U168 ( .A(n321), .B(\mult_x_1/n288 ), .ZN(n105) );
  OAI22_X1 U169 ( .A1(n121), .A2(n105), .B1(n122), .B2(n104), .ZN(n142) );
  XNOR2_X1 U170 ( .A(n320), .B(\mult_x_1/n286 ), .ZN(n111) );
  XNOR2_X1 U171 ( .A(n320), .B(\mult_x_1/n285 ), .ZN(n138) );
  OAI22_X1 U172 ( .A1(n139), .A2(n111), .B1(n199), .B2(n138), .ZN(n159) );
  OAI22_X1 U173 ( .A1(n216), .A2(n107), .B1(n106), .B2(n5), .ZN(n158) );
  XNOR2_X1 U174 ( .A(n13), .B(\mult_x_1/n283 ), .ZN(n141) );
  OAI22_X1 U175 ( .A1(n44), .A2(n108), .B1(n212), .B2(n141), .ZN(n157) );
  OR2_X1 U176 ( .A1(\mult_x_1/n288 ), .A2(n323), .ZN(n109) );
  OAI22_X1 U177 ( .A1(n139), .A2(n323), .B1(n109), .B2(n199), .ZN(n184) );
  XNOR2_X1 U178 ( .A(n320), .B(\mult_x_1/n288 ), .ZN(n110) );
  XNOR2_X1 U179 ( .A(n320), .B(\mult_x_1/n287 ), .ZN(n112) );
  OAI22_X1 U180 ( .A1(n139), .A2(n110), .B1(n199), .B2(n112), .ZN(n183) );
  OAI22_X1 U181 ( .A1(n139), .A2(n112), .B1(n199), .B2(n111), .ZN(n179) );
  FA_X1 U182 ( .A(n115), .B(n114), .CI(n113), .CO(n170), .S(n178) );
  OR2_X1 U183 ( .A1(n176), .A2(n175), .ZN(n116) );
  FA_X1 U184 ( .A(n119), .B(n118), .CI(n117), .CO(n130), .S(n135) );
  AOI21_X1 U185 ( .B1(n122), .B2(n121), .A(n120), .ZN(n123) );
  INV_X1 U186 ( .A(n123), .ZN(n126) );
  NOR2_X1 U187 ( .A1(n20), .A2(n124), .ZN(n125) );
  XOR2_X1 U188 ( .A(n126), .B(n125), .Z(n127) );
  XOR2_X1 U189 ( .A(n128), .B(n127), .Z(n129) );
  OR2_X1 U190 ( .A1(n130), .A2(n129), .ZN(n132) );
  NAND2_X1 U191 ( .A1(n130), .A2(n129), .ZN(n131) );
  NAND2_X1 U192 ( .A1(n132), .A2(n131), .ZN(n133) );
  MUX2_X1 U193 ( .A(n329), .B(n133), .S(n243), .Z(n353) );
  NAND2_X1 U194 ( .A1(n135), .A2(n134), .ZN(n136) );
  MUX2_X1 U195 ( .A(n330), .B(n136), .S(n243), .Z(n355) );
  OAI22_X1 U196 ( .A1(n139), .A2(n138), .B1(n199), .B2(n137), .ZN(n153) );
  OAI22_X1 U197 ( .A1(n210), .A2(n141), .B1(n212), .B2(n140), .ZN(n152) );
  HA_X1 U198 ( .A(n143), .B(n142), .CO(n151), .S(n169) );
  FA_X1 U199 ( .A(n146), .B(n145), .CI(n144), .CO(n55), .S(n237) );
  INV_X1 U200 ( .A(n147), .ZN(n149) );
  XNOR2_X1 U201 ( .A(n150), .B(n235), .ZN(n242) );
  FA_X1 U202 ( .A(n153), .B(n152), .CI(n151), .CO(n236), .S(n166) );
  FA_X1 U203 ( .A(n156), .B(n155), .CI(n154), .CO(n148), .S(n165) );
  FA_X1 U204 ( .A(n159), .B(n158), .CI(n157), .CO(n164), .S(n168) );
  NOR2_X1 U205 ( .A1(n242), .A2(n241), .ZN(n163) );
  MUX2_X1 U206 ( .A(n333), .B(n163), .S(n243), .Z(n361) );
  XNOR2_X1 U207 ( .A(n167), .B(n166), .ZN(n173) );
  FA_X1 U208 ( .A(n170), .B(n169), .CI(n168), .CO(n172), .S(n176) );
  NOR2_X1 U209 ( .A1(n173), .A2(n172), .ZN(n171) );
  MUX2_X1 U210 ( .A(n335), .B(n171), .S(n243), .Z(n365) );
  NAND2_X1 U211 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2_X1 U212 ( .A(n336), .B(n174), .S(n243), .Z(n367) );
  NAND2_X1 U213 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U214 ( .A(n337), .B(n177), .S(n243), .Z(n369) );
  FA_X1 U215 ( .A(n180), .B(n179), .CI(n178), .CO(n175), .S(n187) );
  XNOR2_X1 U216 ( .A(n13), .B(\mult_x_1/n286 ), .ZN(n200) );
  OAI22_X1 U217 ( .A1(n210), .A2(n200), .B1(n212), .B2(n181), .ZN(n197) );
  XNOR2_X1 U218 ( .A(n215), .B(\mult_x_1/n284 ), .ZN(n198) );
  OAI22_X1 U219 ( .A1(n12), .A2(n198), .B1(n182), .B2(n5), .ZN(n196) );
  HA_X1 U220 ( .A(n184), .B(n183), .CO(n180), .S(n195) );
  NOR2_X1 U221 ( .A1(n187), .A2(n186), .ZN(n185) );
  MUX2_X1 U222 ( .A(n338), .B(n185), .S(n243), .Z(n371) );
  NAND2_X1 U223 ( .A1(n187), .A2(n186), .ZN(n188) );
  MUX2_X1 U224 ( .A(n339), .B(n188), .S(n243), .Z(n373) );
  NAND2_X1 U225 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U226 ( .A(n340), .B(n191), .S(n243), .Z(n375) );
  NAND2_X1 U227 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U228 ( .A(n341), .B(n194), .S(n243), .Z(n377) );
  FA_X1 U229 ( .A(n197), .B(n196), .CI(n195), .CO(n186), .S(n226) );
  XNOR2_X1 U230 ( .A(n10), .B(\mult_x_1/n285 ), .ZN(n206) );
  OAI22_X1 U231 ( .A1(n216), .A2(n206), .B1(n198), .B2(n5), .ZN(n203) );
  AND2_X1 U232 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n202) );
  XNOR2_X1 U233 ( .A(n13), .B(\mult_x_1/n287 ), .ZN(n204) );
  OAI22_X1 U234 ( .A1(n210), .A2(n204), .B1(n212), .B2(n200), .ZN(n201) );
  OR2_X1 U235 ( .A1(n226), .A2(n225), .ZN(n271) );
  FA_X1 U236 ( .A(n203), .B(n202), .CI(n201), .CO(n225), .S(n224) );
  XNOR2_X1 U237 ( .A(n13), .B(\mult_x_1/n288 ), .ZN(n205) );
  OAI22_X1 U238 ( .A1(n210), .A2(n205), .B1(n212), .B2(n204), .ZN(n208) );
  XNOR2_X1 U239 ( .A(n10), .B(\mult_x_1/n286 ), .ZN(n211) );
  OAI22_X1 U240 ( .A1(n12), .A2(n211), .B1(n206), .B2(n5), .ZN(n207) );
  NOR2_X1 U241 ( .A1(n224), .A2(n223), .ZN(n264) );
  HA_X1 U242 ( .A(n208), .B(n207), .CO(n223), .S(n221) );
  OR2_X1 U243 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n209) );
  OAI22_X1 U244 ( .A1(n210), .A2(n24), .B1(n209), .B2(n212), .ZN(n220) );
  OR2_X1 U245 ( .A1(n221), .A2(n220), .ZN(n260) );
  XNOR2_X1 U246 ( .A(n10), .B(\mult_x_1/n287 ), .ZN(n214) );
  OAI22_X1 U247 ( .A1(n12), .A2(n214), .B1(n211), .B2(n5), .ZN(n219) );
  INV_X1 U248 ( .A(n212), .ZN(n213) );
  AND2_X1 U249 ( .A1(\mult_x_1/n288 ), .A2(n213), .ZN(n218) );
  NOR2_X1 U250 ( .A1(n219), .A2(n218), .ZN(n253) );
  OAI22_X1 U251 ( .A1(n12), .A2(\mult_x_1/n288 ), .B1(n214), .B2(n5), .ZN(n250) );
  OR2_X1 U252 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n217) );
  NAND2_X1 U253 ( .A1(n217), .A2(n12), .ZN(n249) );
  NAND2_X1 U254 ( .A1(n250), .A2(n249), .ZN(n256) );
  NAND2_X1 U255 ( .A1(n219), .A2(n218), .ZN(n254) );
  OAI21_X1 U256 ( .B1(n253), .B2(n256), .A(n254), .ZN(n261) );
  NAND2_X1 U257 ( .A1(n221), .A2(n220), .ZN(n259) );
  INV_X1 U258 ( .A(n259), .ZN(n222) );
  NAND2_X1 U259 ( .A1(n224), .A2(n223), .ZN(n265) );
  OAI21_X1 U260 ( .B1(n264), .B2(n267), .A(n265), .ZN(n272) );
  NAND2_X1 U261 ( .A1(n226), .A2(n225), .ZN(n270) );
  INV_X1 U262 ( .A(n270), .ZN(n227) );
  AOI21_X1 U263 ( .B1(n271), .B2(n15), .A(n227), .ZN(n228) );
  MUX2_X1 U264 ( .A(n342), .B(n228), .S(n243), .Z(n379) );
  FA_X1 U265 ( .A(n18), .B(n230), .CI(n229), .CO(n60), .S(n231) );
  MUX2_X1 U266 ( .A(n343), .B(n231), .S(n243), .Z(n381) );
  MUX2_X1 U267 ( .A(n344), .B(n240), .S(n243), .Z(n383) );
  NAND2_X1 U268 ( .A1(n242), .A2(n241), .ZN(n244) );
  NAND2_X1 U269 ( .A1(n244), .A2(n243), .ZN(n247) );
  NAND2_X1 U270 ( .A1(n245), .A2(n334), .ZN(n246) );
  NAND2_X1 U271 ( .A1(n247), .A2(n246), .ZN(n363) );
  BUF_X2 U272 ( .A(rst_n), .Z(n394) );
  BUF_X4 U273 ( .A(en), .Z(n322) );
  MUX2_X1 U274 ( .A(product[0]), .B(n506), .S(n322), .Z(n396) );
  MUX2_X1 U275 ( .A(n506), .B(n507), .S(n322), .Z(n398) );
  AND2_X1 U276 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n248) );
  MUX2_X1 U277 ( .A(n507), .B(n248), .S(n322), .Z(n400) );
  MUX2_X1 U278 ( .A(product[1]), .B(n509), .S(n322), .Z(n402) );
  MUX2_X1 U279 ( .A(n509), .B(n510), .S(n322), .Z(n404) );
  OR2_X1 U280 ( .A1(n250), .A2(n249), .ZN(n251) );
  AND2_X1 U281 ( .A1(n251), .A2(n256), .ZN(n252) );
  MUX2_X1 U282 ( .A(n510), .B(n252), .S(n322), .Z(n406) );
  MUX2_X1 U283 ( .A(product[2]), .B(n512), .S(n322), .Z(n408) );
  MUX2_X1 U284 ( .A(n512), .B(n513), .S(n322), .Z(n410) );
  INV_X1 U285 ( .A(n253), .ZN(n255) );
  NAND2_X1 U286 ( .A1(n255), .A2(n254), .ZN(n257) );
  XOR2_X1 U287 ( .A(n257), .B(n256), .Z(n258) );
  MUX2_X1 U288 ( .A(n513), .B(n258), .S(n322), .Z(n412) );
  MUX2_X1 U289 ( .A(product[3]), .B(n515), .S(n322), .Z(n414) );
  MUX2_X1 U290 ( .A(n515), .B(n516), .S(n322), .Z(n416) );
  NAND2_X1 U291 ( .A1(n260), .A2(n259), .ZN(n262) );
  XNOR2_X1 U292 ( .A(n262), .B(n261), .ZN(n263) );
  MUX2_X1 U293 ( .A(n516), .B(n263), .S(n322), .Z(n418) );
  MUX2_X1 U294 ( .A(product[4]), .B(n518), .S(n322), .Z(n420) );
  MUX2_X1 U295 ( .A(n518), .B(n519), .S(n322), .Z(n422) );
  INV_X1 U296 ( .A(n264), .ZN(n266) );
  NAND2_X1 U297 ( .A1(n266), .A2(n265), .ZN(n268) );
  XOR2_X1 U298 ( .A(n268), .B(n14), .Z(n269) );
  MUX2_X1 U299 ( .A(n519), .B(n269), .S(n322), .Z(n424) );
  MUX2_X1 U300 ( .A(product[5]), .B(n521), .S(n322), .Z(n426) );
  MUX2_X1 U301 ( .A(n521), .B(n522), .S(n322), .Z(n428) );
  NAND2_X1 U302 ( .A1(n271), .A2(n270), .ZN(n273) );
  XNOR2_X1 U303 ( .A(n272), .B(n273), .ZN(n274) );
  MUX2_X1 U304 ( .A(n522), .B(n274), .S(n322), .Z(n430) );
  MUX2_X1 U305 ( .A(product[6]), .B(n524), .S(n322), .Z(n432) );
  NAND2_X1 U306 ( .A1(n388), .A2(n339), .ZN(n275) );
  XOR2_X1 U307 ( .A(n275), .B(n342), .Z(n276) );
  MUX2_X1 U308 ( .A(n524), .B(n276), .S(n322), .Z(n434) );
  MUX2_X1 U309 ( .A(product[7]), .B(n526), .S(n322), .Z(n436) );
  OAI21_X1 U310 ( .B1(n338), .B2(n342), .A(n339), .ZN(n279) );
  NAND2_X1 U311 ( .A1(n328), .A2(n337), .ZN(n277) );
  XNOR2_X1 U312 ( .A(n279), .B(n277), .ZN(n278) );
  MUX2_X1 U313 ( .A(n526), .B(n278), .S(n322), .Z(n438) );
  MUX2_X1 U314 ( .A(product[8]), .B(n528), .S(n322), .Z(n440) );
  AOI21_X1 U315 ( .B1(n279), .B2(n328), .A(n389), .ZN(n282) );
  NAND2_X1 U316 ( .A1(n390), .A2(n336), .ZN(n280) );
  XOR2_X1 U317 ( .A(n282), .B(n280), .Z(n281) );
  MUX2_X1 U318 ( .A(n528), .B(n281), .S(n322), .Z(n442) );
  MUX2_X1 U319 ( .A(product[9]), .B(n530), .S(n322), .Z(n444) );
  OAI21_X1 U320 ( .B1(n282), .B2(n335), .A(n336), .ZN(n293) );
  INV_X1 U321 ( .A(n293), .ZN(n285) );
  NAND2_X1 U322 ( .A1(n391), .A2(n334), .ZN(n283) );
  XOR2_X1 U323 ( .A(n285), .B(n283), .Z(n284) );
  MUX2_X1 U324 ( .A(n530), .B(n284), .S(n322), .Z(n446) );
  MUX2_X1 U325 ( .A(product[10]), .B(n532), .S(n322), .Z(n448) );
  OAI21_X1 U326 ( .B1(n285), .B2(n333), .A(n334), .ZN(n288) );
  NOR2_X1 U327 ( .A1(n343), .A2(n344), .ZN(n291) );
  INV_X1 U328 ( .A(n291), .ZN(n286) );
  NAND2_X1 U329 ( .A1(n343), .A2(n344), .ZN(n290) );
  NAND2_X1 U330 ( .A1(n286), .A2(n290), .ZN(n287) );
  XNOR2_X1 U331 ( .A(n288), .B(n287), .ZN(n289) );
  MUX2_X1 U332 ( .A(n532), .B(n289), .S(n322), .Z(n450) );
  MUX2_X1 U333 ( .A(product[11]), .B(n534), .S(n322), .Z(n452) );
  NOR2_X1 U334 ( .A1(n291), .A2(n333), .ZN(n294) );
  OAI21_X1 U335 ( .B1(n291), .B2(n334), .A(n290), .ZN(n292) );
  AOI21_X1 U336 ( .B1(n294), .B2(n293), .A(n292), .ZN(n316) );
  NAND2_X1 U337 ( .A1(n392), .A2(n332), .ZN(n295) );
  XOR2_X1 U338 ( .A(n316), .B(n295), .Z(n296) );
  MUX2_X1 U339 ( .A(n534), .B(n296), .S(n322), .Z(n454) );
  MUX2_X1 U340 ( .A(product[12]), .B(n536), .S(n322), .Z(n456) );
  OAI21_X1 U341 ( .B1(n316), .B2(n331), .A(n332), .ZN(n298) );
  NAND2_X1 U342 ( .A1(n327), .A2(n341), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  MUX2_X1 U344 ( .A(n536), .B(n299), .S(n322), .Z(n458) );
  MUX2_X1 U345 ( .A(product[13]), .B(n538), .S(n322), .Z(n460) );
  NAND2_X1 U346 ( .A1(n392), .A2(n327), .ZN(n301) );
  AOI21_X1 U347 ( .B1(n387), .B2(n327), .A(n393), .ZN(n300) );
  OAI21_X1 U348 ( .B1(n316), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U349 ( .A1(n326), .A2(n340), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U351 ( .A(n538), .B(n304), .S(n322), .Z(n462) );
  MUX2_X1 U352 ( .A(product[14]), .B(n540), .S(n322), .Z(n464) );
  NAND2_X1 U353 ( .A1(n327), .A2(n326), .ZN(n306) );
  NOR2_X1 U354 ( .A1(n331), .A2(n306), .ZN(n312) );
  INV_X1 U355 ( .A(n312), .ZN(n308) );
  AOI21_X1 U356 ( .B1(n393), .B2(n326), .A(n386), .ZN(n305) );
  OAI21_X1 U357 ( .B1(n306), .B2(n332), .A(n305), .ZN(n313) );
  INV_X1 U358 ( .A(n313), .ZN(n307) );
  OAI21_X1 U359 ( .B1(n316), .B2(n308), .A(n307), .ZN(n310) );
  NAND2_X1 U360 ( .A1(n325), .A2(n330), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  MUX2_X1 U362 ( .A(n540), .B(n311), .S(n322), .Z(n466) );
  MUX2_X1 U363 ( .A(product[15]), .B(n542), .S(n322), .Z(n468) );
  NAND2_X1 U364 ( .A1(n312), .A2(n325), .ZN(n315) );
  AOI21_X1 U365 ( .B1(n313), .B2(n325), .A(n385), .ZN(n314) );
  OAI21_X1 U366 ( .B1(n316), .B2(n315), .A(n314), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n317), .B(n329), .ZN(n318) );
  MUX2_X1 U368 ( .A(n542), .B(n318), .S(n322), .Z(n470) );
  MUX2_X1 U369 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n322), .Z(n472) );
  MUX2_X1 U370 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n322), .Z(n474) );
  MUX2_X1 U371 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n322), .Z(n476) );
  MUX2_X1 U372 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n322), .Z(n478) );
  MUX2_X1 U373 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n322), .Z(n480) );
  MUX2_X1 U374 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n322), .Z(n482) );
  MUX2_X1 U375 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n322), .Z(n484) );
  MUX2_X1 U376 ( .A(n11), .B(B_extended[7]), .S(n322), .Z(n486) );
  MUX2_X1 U377 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n322), .Z(n488) );
  MUX2_X1 U378 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n322), .Z(n490) );
  MUX2_X1 U379 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n322), .Z(n492) );
  MUX2_X1 U380 ( .A(n13), .B(A_extended[3]), .S(n322), .Z(n494) );
  MUX2_X1 U381 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n322), .Z(n496) );
  MUX2_X1 U382 ( .A(n320), .B(A_extended[5]), .S(n322), .Z(n498) );
  MUX2_X1 U383 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n322), .Z(n500) );
  MUX2_X1 U384 ( .A(n321), .B(A_extended[7]), .S(n322), .Z(n502) );
  OR2_X1 U385 ( .A1(n322), .A2(n544), .ZN(n504) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_21 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n361, n363, n365, n367, n369, n371, n373, n375, n377, n379,
         n381, n383, n385, n387, n389, n391, n393, n395, n397, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n411, n413,
         n415, n417, n419, n421, n423, n425, n427, n429, n431, n433, n435,
         n437, n439, n441, n443, n445, n447, n449, n451, n453, n455, n457,
         n459, n461, n463, n465, n467, n469, n471, n473, n475, n477, n479,
         n481, n483, n485, n487, n489, n491, n493, n495, n497, n499, n501,
         n503, n505, n507, n509, n511, n513, n515, n517, n519, n521, n522,
         n524, n525, n527, n528, n530, n531, n533, n534, n536, n537, n539,
         n541, n543, n545, n547, n549, n551, n553, n555, n557, n558, n559,
         n560;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n408), .SE(n519), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n337) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n409), .SE(n511), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n33) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n408), .SE(n509), .CK(clk), .Q(n558), 
        .QN(n25) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n409), .SE(n507), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n7) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n408), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n24) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n408), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n28) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n408), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n30) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n409), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n29) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n409), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n27) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n408), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n26) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n408), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n31) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n409), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n23) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n408), .SE(n485), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n409), .SE(n483), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n409), .SE(n481), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n408), .SE(n479), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n408), .SE(n477), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n409), .SE(n475), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n408), .SE(n473), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n409), .SE(n471), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n408), .SE(n469), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n409), .SE(n467), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG23_S3 ( .D(1'b0), .SI(n408), .SE(n465), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG24_S4 ( .D(1'b0), .SI(rst_n), .SE(n463), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG21_S3 ( .D(1'b0), .SI(rst_n), .SE(n461), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG22_S4 ( .D(1'b0), .SI(rst_n), .SE(n459), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n457), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(rst_n), .SE(n455), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n409), .SE(n453), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n409), .SE(n451), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n409), .SE(n449), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n409), .SE(n447), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n409), .SE(n445), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n409), .SE(n443), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n409), .SE(n441), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n409), .SE(n439), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n409), .SE(n437), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n409), .SE(n435), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n409), .SE(n433), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n408), .SE(n431), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n408), .SE(n429), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n408), .SE(n427), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n408), .SE(n425), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n408), .SE(n423), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n408), .SE(n421), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n408), .SE(n419), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n408), .SE(n417), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n408), .SE(n415), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n408), .SE(n413), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n408), .SE(n411), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n409), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n35) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n560), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n560), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n357), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n560), .SE(n393), .CK(
        clk), .QN(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n560), .SE(n391), .CK(
        clk), .Q(n406), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n560), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n560), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n353), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n560), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n352), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n560), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n560), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n350), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n560), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n560), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n348), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n560), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n347), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n560), .SE(n373), .CK(
        clk), .Q(n338), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n560), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n345), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n560), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n344), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n560), .SE(n367), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n560), .SE(n365), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n560), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n560), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n560), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n339) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n336) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n409), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n22) );
  BUF_X1 U2 ( .A(n269), .Z(n257) );
  NAND2_X1 U3 ( .A1(n90), .A2(n89), .ZN(n180) );
  XNOR2_X1 U4 ( .A(n80), .B(n79), .ZN(n181) );
  NAND2_X1 U5 ( .A1(n63), .A2(n62), .ZN(n50) );
  CLKBUF_X1 U6 ( .A(n68), .Z(n14) );
  XNOR2_X1 U7 ( .A(n78), .B(n77), .ZN(n79) );
  INV_X1 U8 ( .A(n188), .ZN(n86) );
  INV_X1 U9 ( .A(n189), .ZN(n87) );
  NAND2_X1 U10 ( .A1(n189), .A2(n188), .ZN(n89) );
  NAND2_X1 U11 ( .A1(n100), .A2(n355), .ZN(n95) );
  NAND2_X1 U12 ( .A1(n94), .A2(n295), .ZN(n96) );
  INV_X1 U13 ( .A(n260), .ZN(n94) );
  CLKBUF_X2 U14 ( .A(n43), .Z(n6) );
  XNOR2_X1 U15 ( .A(n7), .B(n558), .ZN(n44) );
  BUF_X1 U16 ( .A(n122), .Z(n8) );
  BUF_X1 U17 ( .A(n111), .Z(n9) );
  INV_X1 U18 ( .A(n53), .ZN(n10) );
  INV_X1 U19 ( .A(n10), .ZN(n11) );
  INV_X1 U20 ( .A(n10), .ZN(n12) );
  INV_X1 U21 ( .A(n22), .ZN(n13) );
  OAI22_X1 U22 ( .A1(n161), .A2(n81), .B1(n160), .B2(n22), .ZN(n141) );
  AND2_X1 U23 ( .A1(\mult_x_1/n310 ), .A2(n559), .ZN(n59) );
  XNOR2_X1 U24 ( .A(n15), .B(n14), .ZN(n75) );
  XNOR2_X1 U25 ( .A(n66), .B(n67), .ZN(n15) );
  NAND2_X1 U26 ( .A1(n42), .A2(n43), .ZN(n16) );
  CLKBUF_X2 U27 ( .A(\mult_x_1/n311 ), .Z(n17) );
  BUF_X1 U28 ( .A(n69), .Z(n18) );
  NAND2_X1 U29 ( .A1(n42), .A2(n43), .ZN(n151) );
  OR2_X1 U30 ( .A1(n70), .A2(n69), .ZN(n63) );
  NAND2_X1 U31 ( .A1(n66), .A2(n68), .ZN(n19) );
  NAND2_X1 U32 ( .A1(n68), .A2(n67), .ZN(n20) );
  NAND2_X1 U33 ( .A1(n66), .A2(n67), .ZN(n21) );
  NAND3_X1 U34 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n127) );
  BUF_X2 U35 ( .A(n269), .Z(n295) );
  BUF_X1 U36 ( .A(rst_n), .Z(n409) );
  BUF_X1 U37 ( .A(rst_n), .Z(n408) );
  INV_X1 U38 ( .A(rst_n), .ZN(n560) );
  AND2_X1 U39 ( .A1(n91), .A2(n93), .ZN(n32) );
  XNOR2_X1 U40 ( .A(n268), .B(n267), .ZN(n34) );
  XNOR2_X1 U41 ( .A(n337), .B(\mult_x_1/n310 ), .ZN(n36) );
  XNOR2_X1 U42 ( .A(n336), .B(n337), .ZN(n37) );
  NAND2_X2 U43 ( .A1(n36), .A2(n37), .ZN(n160) );
  XNOR2_X1 U44 ( .A(n13), .B(\mult_x_1/n286 ), .ZN(n71) );
  INV_X1 U45 ( .A(n37), .ZN(n38) );
  INV_X2 U46 ( .A(n38), .ZN(n161) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n57) );
  OAI22_X1 U48 ( .A1(n160), .A2(n71), .B1(n161), .B2(n57), .ZN(n80) );
  BUF_X2 U49 ( .A(\mult_x_1/n313 ), .Z(n239) );
  NAND2_X1 U50 ( .A1(n239), .A2(n5), .ZN(n240) );
  AND2_X1 U51 ( .A1(n559), .A2(\mult_x_1/n281 ), .ZN(n104) );
  XNOR2_X1 U52 ( .A(n104), .B(n239), .ZN(n72) );
  AOI21_X1 U53 ( .B1(n240), .B2(n5), .A(n72), .ZN(n39) );
  INV_X1 U54 ( .A(n39), .ZN(n77) );
  XNOR2_X1 U55 ( .A(n59), .B(\mult_x_1/n310 ), .ZN(n108) );
  NOR2_X1 U56 ( .A1(n108), .A2(n31), .ZN(n78) );
  OAI21_X1 U57 ( .B1(n80), .B2(n77), .A(n78), .ZN(n41) );
  NAND2_X1 U58 ( .A1(n80), .A2(n77), .ZN(n40) );
  NAND2_X1 U59 ( .A1(n41), .A2(n40), .ZN(n65) );
  XNOR2_X1 U60 ( .A(\mult_x_1/n311 ), .B(n33), .ZN(n42) );
  XNOR2_X1 U61 ( .A(n558), .B(\mult_x_1/a[4] ), .ZN(n43) );
  XNOR2_X1 U62 ( .A(n17), .B(\mult_x_1/n284 ), .ZN(n85) );
  XNOR2_X1 U63 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n58) );
  OAI22_X1 U64 ( .A1(n151), .A2(n85), .B1(n6), .B2(n58), .ZN(n69) );
  XNOR2_X1 U65 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n45) );
  NAND2_X1 U66 ( .A1(n44), .A2(n45), .ZN(n53) );
  CLKBUF_X2 U67 ( .A(n558), .Z(n334) );
  XNOR2_X1 U68 ( .A(n334), .B(\mult_x_1/n282 ), .ZN(n84) );
  INV_X1 U69 ( .A(n45), .ZN(n46) );
  INV_X2 U70 ( .A(n46), .ZN(n236) );
  XNOR2_X1 U71 ( .A(n334), .B(\mult_x_1/n281 ), .ZN(n52) );
  OAI22_X1 U72 ( .A1(n53), .A2(n84), .B1(n236), .B2(n52), .ZN(n70) );
  INV_X1 U73 ( .A(n63), .ZN(n48) );
  NOR2_X1 U74 ( .A1(n26), .A2(n108), .ZN(n62) );
  INV_X1 U75 ( .A(n62), .ZN(n47) );
  NAND2_X1 U76 ( .A1(n48), .A2(n47), .ZN(n49) );
  NAND2_X1 U77 ( .A1(n65), .A2(n49), .ZN(n51) );
  NAND2_X1 U78 ( .A1(n51), .A2(n50), .ZN(n138) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n56) );
  XNOR2_X1 U80 ( .A(n13), .B(\mult_x_1/n283 ), .ZN(n110) );
  OAI22_X1 U81 ( .A1(n160), .A2(n56), .B1(n161), .B2(n110), .ZN(n123) );
  XNOR2_X1 U82 ( .A(n104), .B(n334), .ZN(n54) );
  OAI22_X1 U83 ( .A1(n53), .A2(n52), .B1(n54), .B2(n236), .ZN(n122) );
  AOI21_X1 U84 ( .B1(n236), .B2(n11), .A(n54), .ZN(n55) );
  INV_X1 U85 ( .A(n55), .ZN(n121) );
  OAI22_X1 U86 ( .A1(n160), .A2(n57), .B1(n161), .B2(n56), .ZN(n68) );
  XNOR2_X1 U87 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n60) );
  OAI22_X1 U88 ( .A1(n16), .A2(n58), .B1(n6), .B2(n60), .ZN(n67) );
  INV_X1 U89 ( .A(n122), .ZN(n66) );
  XNOR2_X1 U90 ( .A(n59), .B(\mult_x_1/n310 ), .ZN(n163) );
  NOR2_X1 U91 ( .A1(n27), .A2(n163), .ZN(n129) );
  XNOR2_X1 U92 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n107) );
  OAI22_X1 U93 ( .A1(n16), .A2(n60), .B1(n6), .B2(n107), .ZN(n128) );
  XNOR2_X1 U94 ( .A(n129), .B(n128), .ZN(n61) );
  XNOR2_X1 U95 ( .A(n127), .B(n61), .ZN(n136) );
  XNOR2_X1 U96 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U97 ( .A(n65), .B(n64), .ZN(n76) );
  XNOR2_X1 U98 ( .A(n70), .B(n18), .ZN(n91) );
  XNOR2_X1 U99 ( .A(n13), .B(\mult_x_1/n287 ), .ZN(n82) );
  OAI22_X1 U100 ( .A1(n160), .A2(n82), .B1(n161), .B2(n71), .ZN(n184) );
  XNOR2_X1 U101 ( .A(n239), .B(\mult_x_1/n281 ), .ZN(n143) );
  OAI22_X1 U102 ( .A1(n240), .A2(n143), .B1(n72), .B2(n5), .ZN(n183) );
  NOR2_X1 U103 ( .A1(n163), .A2(n23), .ZN(n182) );
  INV_X1 U104 ( .A(n97), .ZN(n73) );
  CLKBUF_X1 U105 ( .A(en), .Z(n269) );
  NAND2_X1 U106 ( .A1(n73), .A2(n257), .ZN(n74) );
  OAI22_X1 U107 ( .A1(n98), .A2(n74), .B1(n257), .B2(n338), .ZN(n373) );
  FA_X1 U108 ( .A(n32), .B(n75), .CI(n76), .CO(n97), .S(n261) );
  OR2_X1 U109 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n81) );
  XNOR2_X1 U110 ( .A(n13), .B(\mult_x_1/n288 ), .ZN(n83) );
  OAI22_X1 U111 ( .A1(n160), .A2(n83), .B1(n161), .B2(n82), .ZN(n140) );
  XNOR2_X1 U112 ( .A(n334), .B(\mult_x_1/n283 ), .ZN(n145) );
  OAI22_X1 U113 ( .A1(n11), .A2(n145), .B1(n236), .B2(n84), .ZN(n189) );
  XNOR2_X1 U114 ( .A(n17), .B(\mult_x_1/n285 ), .ZN(n142) );
  OAI22_X1 U115 ( .A1(n16), .A2(n142), .B1(n6), .B2(n85), .ZN(n188) );
  NAND2_X1 U116 ( .A1(n87), .A2(n86), .ZN(n88) );
  NAND2_X1 U117 ( .A1(n191), .A2(n88), .ZN(n90) );
  INV_X1 U118 ( .A(n91), .ZN(n92) );
  XNOR2_X1 U119 ( .A(n93), .B(n92), .ZN(n179) );
  OAI21_X1 U120 ( .B1(n261), .B2(n96), .A(n95), .ZN(n391) );
  NAND2_X1 U121 ( .A1(n98), .A2(n97), .ZN(n99) );
  NAND2_X1 U122 ( .A1(n99), .A2(n257), .ZN(n102) );
  INV_X1 U123 ( .A(n257), .ZN(n100) );
  NAND2_X1 U124 ( .A1(n100), .A2(n347), .ZN(n101) );
  NAND2_X1 U125 ( .A1(n102), .A2(n101), .ZN(n375) );
  NOR2_X1 U146 ( .A1(n28), .A2(n163), .ZN(n158) );
  XNOR2_X1 U147 ( .A(n13), .B(\mult_x_1/n281 ), .ZN(n103) );
  XNOR2_X1 U148 ( .A(n104), .B(n13), .ZN(n159) );
  OAI22_X1 U149 ( .A1(n160), .A2(n103), .B1(n159), .B2(n161), .ZN(n167) );
  INV_X1 U150 ( .A(n167), .ZN(n157) );
  XNOR2_X1 U151 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n109) );
  OAI22_X1 U152 ( .A1(n160), .A2(n109), .B1(n161), .B2(n103), .ZN(n113) );
  XNOR2_X1 U153 ( .A(n104), .B(\mult_x_1/n311 ), .ZN(n106) );
  AOI21_X1 U154 ( .B1(n6), .B2(n151), .A(n106), .ZN(n105) );
  INV_X1 U155 ( .A(n105), .ZN(n112) );
  OAI22_X1 U156 ( .A1(n151), .A2(n107), .B1(n106), .B2(n6), .ZN(n111) );
  NOR2_X1 U157 ( .A1(n29), .A2(n108), .ZN(n120) );
  OAI22_X1 U158 ( .A1(n160), .A2(n110), .B1(n161), .B2(n109), .ZN(n119) );
  INV_X1 U159 ( .A(n111), .ZN(n118) );
  NOR2_X1 U160 ( .A1(n30), .A2(n163), .ZN(n116) );
  FA_X1 U161 ( .A(n113), .B(n112), .CI(n9), .CO(n156), .S(n115) );
  OR2_X1 U162 ( .A1(n174), .A2(n173), .ZN(n114) );
  MUX2_X1 U163 ( .A(n339), .B(n114), .S(n257), .Z(n359) );
  FA_X1 U164 ( .A(n117), .B(n116), .CI(n115), .CO(n173), .S(n218) );
  FA_X1 U165 ( .A(n119), .B(n120), .CI(n118), .CO(n117), .S(n135) );
  FA_X1 U166 ( .A(n123), .B(n8), .CI(n121), .CO(n134), .S(n137) );
  INV_X1 U167 ( .A(n129), .ZN(n125) );
  INV_X1 U168 ( .A(n128), .ZN(n124) );
  NAND2_X1 U169 ( .A1(n125), .A2(n124), .ZN(n126) );
  NAND2_X1 U170 ( .A1(n127), .A2(n126), .ZN(n131) );
  NAND2_X1 U171 ( .A1(n129), .A2(n128), .ZN(n130) );
  NAND2_X1 U172 ( .A1(n131), .A2(n130), .ZN(n133) );
  OR2_X1 U173 ( .A1(n218), .A2(n217), .ZN(n132) );
  MUX2_X1 U174 ( .A(n340), .B(n132), .S(n257), .Z(n361) );
  FA_X1 U175 ( .A(n135), .B(n134), .CI(n133), .CO(n217), .S(n177) );
  FA_X1 U176 ( .A(n138), .B(n137), .CI(n136), .CO(n176), .S(n98) );
  OR2_X1 U177 ( .A1(n177), .A2(n176), .ZN(n139) );
  MUX2_X1 U178 ( .A(n341), .B(n139), .S(n257), .Z(n363) );
  XNOR2_X1 U179 ( .A(n239), .B(\mult_x_1/n283 ), .ZN(n210) );
  XNOR2_X1 U180 ( .A(n239), .B(\mult_x_1/n282 ), .ZN(n144) );
  OAI22_X1 U181 ( .A1(n240), .A2(n210), .B1(n144), .B2(n5), .ZN(n154) );
  AND2_X1 U182 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n153) );
  XNOR2_X1 U183 ( .A(n334), .B(\mult_x_1/n285 ), .ZN(n209) );
  XNOR2_X1 U184 ( .A(n334), .B(\mult_x_1/n284 ), .ZN(n146) );
  OAI22_X1 U185 ( .A1(n11), .A2(n209), .B1(n236), .B2(n146), .ZN(n152) );
  HA_X1 U186 ( .A(n141), .B(n140), .CO(n191), .S(n197) );
  XNOR2_X1 U187 ( .A(n17), .B(\mult_x_1/n286 ), .ZN(n149) );
  OAI22_X1 U188 ( .A1(n16), .A2(n149), .B1(n6), .B2(n142), .ZN(n187) );
  OAI22_X1 U189 ( .A1(n240), .A2(n144), .B1(n143), .B2(n5), .ZN(n186) );
  OAI22_X1 U190 ( .A1(n12), .A2(n146), .B1(n236), .B2(n145), .ZN(n185) );
  OR2_X1 U191 ( .A1(\mult_x_1/n288 ), .A2(n336), .ZN(n147) );
  OAI22_X1 U192 ( .A1(n16), .A2(n336), .B1(n147), .B2(n6), .ZN(n212) );
  XNOR2_X1 U193 ( .A(n17), .B(\mult_x_1/n288 ), .ZN(n148) );
  XNOR2_X1 U194 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n150) );
  OAI22_X1 U195 ( .A1(n151), .A2(n148), .B1(n6), .B2(n150), .ZN(n211) );
  OAI22_X1 U196 ( .A1(n16), .A2(n150), .B1(n6), .B2(n149), .ZN(n207) );
  FA_X1 U197 ( .A(n154), .B(n153), .CI(n152), .CO(n198), .S(n206) );
  OR2_X1 U198 ( .A1(n204), .A2(n203), .ZN(n155) );
  MUX2_X1 U199 ( .A(n342), .B(n155), .S(n257), .Z(n365) );
  FA_X1 U200 ( .A(n158), .B(n157), .CI(n156), .CO(n169), .S(n174) );
  AOI21_X1 U201 ( .B1(n161), .B2(n160), .A(n159), .ZN(n162) );
  INV_X1 U202 ( .A(n162), .ZN(n165) );
  NOR2_X1 U203 ( .A1(n24), .A2(n163), .ZN(n164) );
  XOR2_X1 U204 ( .A(n165), .B(n164), .Z(n166) );
  XOR2_X1 U205 ( .A(n167), .B(n166), .Z(n168) );
  OR2_X1 U206 ( .A1(n169), .A2(n168), .ZN(n171) );
  NAND2_X1 U207 ( .A1(n169), .A2(n168), .ZN(n170) );
  NAND2_X1 U208 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U209 ( .A(n343), .B(n172), .S(n257), .Z(n367) );
  NAND2_X1 U210 ( .A1(n174), .A2(n173), .ZN(n175) );
  MUX2_X1 U211 ( .A(n344), .B(n175), .S(n257), .Z(n369) );
  NAND2_X1 U212 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2_X1 U213 ( .A(n345), .B(n178), .S(n257), .Z(n371) );
  FA_X1 U214 ( .A(n181), .B(n180), .CI(n179), .CO(n260), .S(n255) );
  FA_X1 U215 ( .A(n182), .B(n183), .CI(n184), .CO(n93), .S(n195) );
  FA_X1 U216 ( .A(n187), .B(n186), .CI(n185), .CO(n194), .S(n196) );
  XNOR2_X1 U217 ( .A(n189), .B(n188), .ZN(n190) );
  XNOR2_X1 U218 ( .A(n191), .B(n190), .ZN(n193) );
  NOR2_X1 U219 ( .A1(n255), .A2(n254), .ZN(n192) );
  MUX2_X1 U220 ( .A(n348), .B(n192), .S(n257), .Z(n377) );
  FA_X1 U221 ( .A(n195), .B(n194), .CI(n193), .CO(n254), .S(n201) );
  FA_X1 U222 ( .A(n198), .B(n197), .CI(n196), .CO(n200), .S(n204) );
  NOR2_X1 U223 ( .A1(n201), .A2(n200), .ZN(n199) );
  MUX2_X1 U224 ( .A(n350), .B(n199), .S(n257), .Z(n381) );
  NAND2_X1 U225 ( .A1(n201), .A2(n200), .ZN(n202) );
  MUX2_X1 U226 ( .A(n351), .B(n202), .S(n335), .Z(n383) );
  NAND2_X1 U227 ( .A1(n204), .A2(n203), .ZN(n205) );
  MUX2_X1 U228 ( .A(n352), .B(n205), .S(n335), .Z(n385) );
  FA_X1 U229 ( .A(n208), .B(n207), .CI(n206), .CO(n203), .S(n215) );
  XNOR2_X1 U230 ( .A(n334), .B(\mult_x_1/n286 ), .ZN(n225) );
  OAI22_X1 U231 ( .A1(n11), .A2(n225), .B1(n236), .B2(n209), .ZN(n222) );
  XNOR2_X1 U232 ( .A(n239), .B(\mult_x_1/n284 ), .ZN(n223) );
  OAI22_X1 U233 ( .A1(n240), .A2(n223), .B1(n210), .B2(n5), .ZN(n221) );
  HA_X1 U234 ( .A(n212), .B(n211), .CO(n208), .S(n220) );
  NOR2_X1 U235 ( .A1(n215), .A2(n214), .ZN(n213) );
  MUX2_X1 U236 ( .A(n353), .B(n213), .S(n295), .Z(n387) );
  NAND2_X1 U237 ( .A1(n215), .A2(n214), .ZN(n216) );
  MUX2_X1 U238 ( .A(n354), .B(n216), .S(n335), .Z(n389) );
  NAND2_X1 U239 ( .A1(n218), .A2(n217), .ZN(n219) );
  MUX2_X1 U240 ( .A(n357), .B(n219), .S(n295), .Z(n395) );
  FA_X1 U241 ( .A(n222), .B(n221), .CI(n220), .CO(n214), .S(n251) );
  XNOR2_X1 U242 ( .A(n239), .B(\mult_x_1/n285 ), .ZN(n231) );
  OAI22_X1 U243 ( .A1(n240), .A2(n231), .B1(n223), .B2(n5), .ZN(n228) );
  INV_X1 U244 ( .A(n6), .ZN(n224) );
  AND2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n224), .ZN(n227) );
  XNOR2_X1 U246 ( .A(n334), .B(\mult_x_1/n287 ), .ZN(n229) );
  OAI22_X1 U247 ( .A1(n12), .A2(n229), .B1(n236), .B2(n225), .ZN(n226) );
  OR2_X1 U248 ( .A1(n251), .A2(n250), .ZN(n288) );
  FA_X1 U249 ( .A(n228), .B(n227), .CI(n226), .CO(n250), .S(n248) );
  XNOR2_X1 U250 ( .A(n334), .B(\mult_x_1/n288 ), .ZN(n230) );
  OAI22_X1 U251 ( .A1(n12), .A2(n230), .B1(n236), .B2(n229), .ZN(n233) );
  XNOR2_X1 U252 ( .A(n239), .B(\mult_x_1/n286 ), .ZN(n235) );
  OAI22_X1 U253 ( .A1(n240), .A2(n235), .B1(n231), .B2(n5), .ZN(n232) );
  OR2_X1 U254 ( .A1(n248), .A2(n247), .ZN(n266) );
  INV_X1 U255 ( .A(n266), .ZN(n249) );
  HA_X1 U256 ( .A(n233), .B(n232), .CO(n247), .S(n245) );
  OR2_X1 U257 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n234) );
  OAI22_X1 U258 ( .A1(n12), .A2(n25), .B1(n234), .B2(n236), .ZN(n244) );
  OR2_X1 U259 ( .A1(n245), .A2(n244), .ZN(n283) );
  XNOR2_X1 U260 ( .A(n239), .B(\mult_x_1/n287 ), .ZN(n238) );
  OAI22_X1 U261 ( .A1(n240), .A2(n238), .B1(n235), .B2(n5), .ZN(n243) );
  INV_X1 U262 ( .A(n236), .ZN(n237) );
  AND2_X1 U263 ( .A1(\mult_x_1/n288 ), .A2(n237), .ZN(n242) );
  NOR2_X1 U264 ( .A1(n243), .A2(n242), .ZN(n276) );
  OAI22_X1 U265 ( .A1(n240), .A2(\mult_x_1/n288 ), .B1(n238), .B2(n5), .ZN(
        n273) );
  OR2_X1 U266 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n241) );
  NAND2_X1 U267 ( .A1(n241), .A2(n240), .ZN(n272) );
  NAND2_X1 U268 ( .A1(n273), .A2(n272), .ZN(n279) );
  NAND2_X1 U269 ( .A1(n243), .A2(n242), .ZN(n277) );
  OAI21_X1 U270 ( .B1(n276), .B2(n279), .A(n277), .ZN(n284) );
  NAND2_X1 U271 ( .A1(n245), .A2(n244), .ZN(n282) );
  INV_X1 U272 ( .A(n282), .ZN(n246) );
  AOI21_X1 U273 ( .B1(n283), .B2(n284), .A(n246), .ZN(n267) );
  NAND2_X1 U274 ( .A1(n248), .A2(n247), .ZN(n265) );
  OAI21_X1 U275 ( .B1(n249), .B2(n267), .A(n265), .ZN(n289) );
  NAND2_X1 U276 ( .A1(n251), .A2(n250), .ZN(n287) );
  INV_X1 U277 ( .A(n287), .ZN(n252) );
  AOI21_X1 U278 ( .B1(n288), .B2(n289), .A(n252), .ZN(n253) );
  MUX2_X1 U279 ( .A(n358), .B(n253), .S(n295), .Z(n397) );
  NAND2_X1 U280 ( .A1(n255), .A2(n254), .ZN(n256) );
  NAND2_X1 U281 ( .A1(n256), .A2(n257), .ZN(n259) );
  NAND2_X1 U282 ( .A1(n100), .A2(n349), .ZN(n258) );
  NAND2_X1 U283 ( .A1(n259), .A2(n258), .ZN(n379) );
  NAND2_X1 U284 ( .A1(n261), .A2(n260), .ZN(n262) );
  NAND2_X1 U285 ( .A1(n262), .A2(n335), .ZN(n264) );
  NAND2_X1 U286 ( .A1(n100), .A2(n356), .ZN(n263) );
  NAND2_X1 U287 ( .A1(n264), .A2(n263), .ZN(n393) );
  NAND2_X1 U288 ( .A1(n266), .A2(n265), .ZN(n268) );
  NAND2_X1 U289 ( .A1(n100), .A2(n534), .ZN(n270) );
  OAI21_X1 U290 ( .B1(n34), .B2(n100), .A(n270), .ZN(n439) );
  MUX2_X1 U291 ( .A(product[0]), .B(n521), .S(n295), .Z(n411) );
  MUX2_X1 U292 ( .A(n521), .B(n522), .S(n295), .Z(n413) );
  AND2_X1 U293 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n271) );
  MUX2_X1 U294 ( .A(n522), .B(n271), .S(n295), .Z(n415) );
  MUX2_X1 U295 ( .A(product[1]), .B(n524), .S(n295), .Z(n417) );
  MUX2_X1 U296 ( .A(n524), .B(n525), .S(n295), .Z(n419) );
  OR2_X1 U297 ( .A1(n273), .A2(n272), .ZN(n274) );
  AND2_X1 U298 ( .A1(n274), .A2(n279), .ZN(n275) );
  MUX2_X1 U299 ( .A(n525), .B(n275), .S(n295), .Z(n421) );
  MUX2_X1 U300 ( .A(product[2]), .B(n527), .S(n295), .Z(n423) );
  MUX2_X1 U301 ( .A(n527), .B(n528), .S(n295), .Z(n425) );
  INV_X1 U302 ( .A(n276), .ZN(n278) );
  NAND2_X1 U303 ( .A1(n278), .A2(n277), .ZN(n280) );
  XOR2_X1 U304 ( .A(n280), .B(n279), .Z(n281) );
  MUX2_X1 U305 ( .A(n528), .B(n281), .S(n295), .Z(n427) );
  MUX2_X1 U306 ( .A(product[3]), .B(n530), .S(n295), .Z(n429) );
  MUX2_X1 U307 ( .A(n530), .B(n531), .S(n295), .Z(n431) );
  NAND2_X1 U308 ( .A1(n283), .A2(n282), .ZN(n285) );
  XNOR2_X1 U309 ( .A(n285), .B(n284), .ZN(n286) );
  MUX2_X1 U310 ( .A(n531), .B(n286), .S(n295), .Z(n433) );
  MUX2_X1 U311 ( .A(product[4]), .B(n533), .S(n295), .Z(n435) );
  MUX2_X1 U312 ( .A(n533), .B(n534), .S(n295), .Z(n437) );
  MUX2_X1 U313 ( .A(product[5]), .B(n536), .S(n295), .Z(n441) );
  MUX2_X1 U314 ( .A(n536), .B(n537), .S(n295), .Z(n443) );
  NAND2_X1 U315 ( .A1(n288), .A2(n287), .ZN(n290) );
  XNOR2_X1 U316 ( .A(n290), .B(n289), .ZN(n291) );
  MUX2_X1 U317 ( .A(n537), .B(n291), .S(n295), .Z(n445) );
  MUX2_X1 U318 ( .A(product[6]), .B(n539), .S(n295), .Z(n447) );
  NAND2_X1 U319 ( .A1(n402), .A2(n354), .ZN(n292) );
  XOR2_X1 U320 ( .A(n292), .B(n358), .Z(n293) );
  MUX2_X1 U321 ( .A(n539), .B(n293), .S(n295), .Z(n449) );
  MUX2_X1 U322 ( .A(product[7]), .B(n541), .S(n295), .Z(n451) );
  OAI21_X1 U323 ( .B1(n353), .B2(n358), .A(n354), .ZN(n297) );
  NAND2_X1 U324 ( .A1(n342), .A2(n352), .ZN(n294) );
  XNOR2_X1 U325 ( .A(n297), .B(n294), .ZN(n296) );
  MUX2_X1 U326 ( .A(n541), .B(n296), .S(n295), .Z(n453) );
  BUF_X2 U327 ( .A(en), .Z(n335) );
  MUX2_X1 U328 ( .A(product[8]), .B(n543), .S(n335), .Z(n455) );
  AOI21_X1 U329 ( .B1(n297), .B2(n342), .A(n403), .ZN(n300) );
  NAND2_X1 U330 ( .A1(n404), .A2(n351), .ZN(n298) );
  XOR2_X1 U331 ( .A(n300), .B(n298), .Z(n299) );
  MUX2_X1 U332 ( .A(n543), .B(n299), .S(n335), .Z(n457) );
  MUX2_X1 U333 ( .A(product[9]), .B(n545), .S(n335), .Z(n459) );
  OAI21_X1 U334 ( .B1(n300), .B2(n350), .A(n351), .ZN(n308) );
  INV_X1 U335 ( .A(n308), .ZN(n303) );
  NAND2_X1 U336 ( .A1(n405), .A2(n349), .ZN(n301) );
  XOR2_X1 U337 ( .A(n303), .B(n301), .Z(n302) );
  MUX2_X1 U338 ( .A(n545), .B(n302), .S(n335), .Z(n461) );
  MUX2_X1 U339 ( .A(product[10]), .B(n547), .S(n335), .Z(n463) );
  OAI21_X1 U340 ( .B1(n303), .B2(n348), .A(n349), .ZN(n305) );
  NAND2_X1 U341 ( .A1(n406), .A2(n356), .ZN(n304) );
  XNOR2_X1 U342 ( .A(n305), .B(n304), .ZN(n306) );
  MUX2_X1 U343 ( .A(n547), .B(n306), .S(n335), .Z(n465) );
  MUX2_X1 U344 ( .A(product[11]), .B(n549), .S(n335), .Z(n467) );
  NOR2_X1 U345 ( .A1(n355), .A2(n348), .ZN(n309) );
  OAI21_X1 U346 ( .B1(n355), .B2(n349), .A(n356), .ZN(n307) );
  AOI21_X1 U347 ( .B1(n309), .B2(n308), .A(n307), .ZN(n331) );
  NAND2_X1 U348 ( .A1(n338), .A2(n347), .ZN(n310) );
  XOR2_X1 U349 ( .A(n331), .B(n310), .Z(n311) );
  MUX2_X1 U350 ( .A(n549), .B(n311), .S(n335), .Z(n469) );
  MUX2_X1 U351 ( .A(product[12]), .B(n551), .S(n335), .Z(n471) );
  OAI21_X1 U352 ( .B1(n331), .B2(n346), .A(n347), .ZN(n313) );
  NAND2_X1 U353 ( .A1(n341), .A2(n345), .ZN(n312) );
  XNOR2_X1 U354 ( .A(n313), .B(n312), .ZN(n314) );
  MUX2_X1 U355 ( .A(n551), .B(n314), .S(n335), .Z(n473) );
  MUX2_X1 U356 ( .A(product[13]), .B(n553), .S(n335), .Z(n475) );
  NAND2_X1 U357 ( .A1(n338), .A2(n341), .ZN(n316) );
  AOI21_X1 U358 ( .B1(n401), .B2(n341), .A(n407), .ZN(n315) );
  OAI21_X1 U359 ( .B1(n331), .B2(n316), .A(n315), .ZN(n318) );
  NAND2_X1 U360 ( .A1(n340), .A2(n357), .ZN(n317) );
  XNOR2_X1 U361 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U362 ( .A(n553), .B(n319), .S(n335), .Z(n477) );
  MUX2_X1 U363 ( .A(product[14]), .B(n555), .S(n335), .Z(n479) );
  NAND2_X1 U364 ( .A1(n341), .A2(n340), .ZN(n321) );
  NOR2_X1 U365 ( .A1(n346), .A2(n321), .ZN(n327) );
  INV_X1 U366 ( .A(n327), .ZN(n323) );
  AOI21_X1 U367 ( .B1(n407), .B2(n340), .A(n400), .ZN(n320) );
  OAI21_X1 U368 ( .B1(n321), .B2(n347), .A(n320), .ZN(n328) );
  INV_X1 U369 ( .A(n328), .ZN(n322) );
  OAI21_X1 U370 ( .B1(n331), .B2(n323), .A(n322), .ZN(n325) );
  NAND2_X1 U371 ( .A1(n339), .A2(n344), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U373 ( .A(n555), .B(n326), .S(n335), .Z(n481) );
  MUX2_X1 U374 ( .A(product[15]), .B(n557), .S(n335), .Z(n483) );
  NAND2_X1 U375 ( .A1(n327), .A2(n339), .ZN(n330) );
  AOI21_X1 U376 ( .B1(n328), .B2(n339), .A(n399), .ZN(n329) );
  OAI21_X1 U377 ( .B1(n331), .B2(n330), .A(n329), .ZN(n332) );
  XNOR2_X1 U378 ( .A(n332), .B(n343), .ZN(n333) );
  MUX2_X1 U379 ( .A(n557), .B(n333), .S(n335), .Z(n485) );
  MUX2_X1 U380 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n335), .Z(n487) );
  MUX2_X1 U381 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n335), .Z(n489) );
  MUX2_X1 U382 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n335), .Z(n491) );
  MUX2_X1 U383 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n335), .Z(n493) );
  MUX2_X1 U384 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n335), .Z(n495) );
  MUX2_X1 U385 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n335), .Z(n497) );
  MUX2_X1 U386 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n335), .Z(n499) );
  MUX2_X1 U387 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n335), .Z(n501) );
  MUX2_X1 U388 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n335), .Z(n503) );
  MUX2_X1 U389 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n335), .Z(n505) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n335), .Z(n507) );
  MUX2_X1 U391 ( .A(n334), .B(A_extended[3]), .S(n335), .Z(n509) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n335), .Z(n511) );
  MUX2_X1 U393 ( .A(n17), .B(A_extended[5]), .S(n335), .Z(n513) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n335), .Z(n515) );
  MUX2_X1 U395 ( .A(n13), .B(A_extended[7]), .S(n335), .Z(n517) );
  OR2_X1 U396 ( .A1(n335), .A2(n559), .ZN(n519) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_22 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n352, n354, n356, n358, n360, n362, n364, n366,
         n368, n370, n372, n374, n376, n378, n380, n382, n384, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n396, n398, n400, n402,
         n404, n406, n408, n410, n412, n414, n416, n418, n420, n422, n424,
         n426, n428, n430, n432, n434, n436, n438, n440, n442, n444, n446,
         n448, n450, n452, n454, n456, n458, n460, n462, n464, n466, n468,
         n470, n472, n474, n476, n478, n480, n482, n484, n486, n488, n490,
         n492, n494, n496, n498, n500, n502, n504, n506, n508, n509, n511,
         n512, n514, n515, n517, n518, n520, n521, n523, n524, n526, n527,
         n529, n531, n533, n535, n537, n539, n541, n543, n545, n546, n547,
         n548;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n252), .SE(n506), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n394), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n23) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n394), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n22) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n394), .SE(n498), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n11) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n394), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n21) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n394), .SE(n494), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n12) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n394), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n394), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n252), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n252), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n252), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n252), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n252), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n252), .SE(n472), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n252), .SE(n470), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n252), .SE(n468), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n252), .SE(n466), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n252), .SE(n464), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n252), .SE(n462), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n394), .SE(n460), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n394), .SE(n458), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n394), .SE(n456), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n394), .SE(n454), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n394), .SE(n452), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n252), .SE(n450), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n394), .SE(n448), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n394), .SE(n446), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n394), .SE(n444), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n252), .SE(n442), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n394), .SE(n440), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n394), .SE(n438), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n394), .SE(n436), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n394), .SE(n434), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n394), .SE(n432), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n394), .SE(n430), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n394), .SE(n428), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n394), .SE(n426), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n394), .SE(n424), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n394), .SE(n422), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n394), .SE(n420), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n394), .SE(n418), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n394), .SE(n416), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n394), .SE(n414), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n394), .SE(n412), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n394), .SE(n410), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n252), .SE(n408), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n394), .SE(n406), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n252), .SE(n404), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n394), .SE(n402), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n394), .SE(n400), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n252), .SE(n398), .CK(clk), .Q(n508)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n394), .SE(n396), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n394), .SE(n492), .CK(clk), .Q(n546), 
        .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n548), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n548), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n548), .SE(n380), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n548), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n346), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n548), .SE(n376), .CK(
        clk), .Q(n392), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n548), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n548), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n343), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n548), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n342), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n548), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n341), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n548), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n548), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n339), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n548), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n548), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n337), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n548), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n336), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n548), .SE(n356), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n548), .SE(n354), .CK(
        clk), .QN(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n548), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n548), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n332) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n394), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n331) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n394), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n394), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n20) );
  BUF_X1 U2 ( .A(en), .Z(n183) );
  INV_X1 U3 ( .A(n51), .ZN(n116) );
  BUF_X2 U4 ( .A(n32), .Z(n19) );
  CLKBUF_X1 U5 ( .A(n226), .Z(n5) );
  XNOR2_X1 U6 ( .A(n63), .B(n328), .ZN(n6) );
  CLKBUF_X1 U7 ( .A(n223), .Z(n7) );
  BUF_X1 U8 ( .A(n113), .Z(n8) );
  INV_X1 U9 ( .A(\mult_x_1/n180 ), .ZN(n9) );
  XNOR2_X1 U10 ( .A(n205), .B(n204), .ZN(n211) );
  XNOR2_X1 U11 ( .A(n203), .B(n202), .ZN(n205) );
  OR2_X1 U12 ( .A1(n248), .A2(n247), .ZN(n245) );
  NAND2_X1 U13 ( .A1(n142), .A2(n141), .ZN(n247) );
  NAND2_X1 U14 ( .A1(n154), .A2(n153), .ZN(n141) );
  NAND2_X1 U15 ( .A1(n156), .A2(n140), .ZN(n142) );
  OR2_X1 U16 ( .A1(n153), .A2(n154), .ZN(n140) );
  AND2_X1 U17 ( .A1(\mult_x_1/n310 ), .A2(n547), .ZN(n32) );
  CLKBUF_X1 U18 ( .A(n82), .Z(n18) );
  OAI21_X1 U19 ( .B1(n204), .B2(n200), .A(n199), .ZN(n236) );
  XNOR2_X1 U20 ( .A(n156), .B(n155), .ZN(n161) );
  XNOR2_X1 U21 ( .A(n154), .B(n153), .ZN(n155) );
  NAND2_X1 U22 ( .A1(n107), .A2(n106), .ZN(n171) );
  NAND2_X1 U23 ( .A1(n248), .A2(n247), .ZN(n249) );
  NAND2_X1 U24 ( .A1(n246), .A2(n245), .ZN(n250) );
  CLKBUF_X1 U25 ( .A(n272), .Z(n17) );
  CLKBUF_X1 U26 ( .A(n277), .Z(n13) );
  BUF_X1 U27 ( .A(n226), .Z(n10) );
  NAND2_X1 U28 ( .A1(n9), .A2(n327), .ZN(n226) );
  XNOR2_X1 U29 ( .A(n11), .B(\mult_x_1/n312 ), .ZN(n29) );
  XNOR2_X1 U30 ( .A(n194), .B(n193), .ZN(n237) );
  NAND2_X1 U31 ( .A1(n194), .A2(n105), .ZN(n107) );
  XNOR2_X1 U32 ( .A(n546), .B(n12), .ZN(n31) );
  NAND2_X1 U33 ( .A1(n27), .A2(n26), .ZN(n113) );
  BUF_X4 U34 ( .A(n546), .Z(n327) );
  XNOR2_X1 U35 ( .A(n327), .B(n63), .ZN(n14) );
  BUF_X1 U36 ( .A(\mult_x_1/n281 ), .Z(n15) );
  OAI22_X1 U37 ( .A1(n139), .A2(n64), .B1(n65), .B2(n207), .ZN(n16) );
  AND2_X2 U38 ( .A1(n547), .A2(\mult_x_1/n281 ), .ZN(n63) );
  OR2_X1 U39 ( .A1(n192), .A2(n191), .ZN(n105) );
  NAND2_X1 U40 ( .A1(n192), .A2(n191), .ZN(n106) );
  XNOR2_X1 U41 ( .A(n192), .B(n191), .ZN(n193) );
  XNOR2_X1 U42 ( .A(n196), .B(n195), .ZN(n204) );
  INV_X1 U43 ( .A(rst_n), .ZN(n548) );
  BUF_X2 U44 ( .A(\mult_x_1/n310 ), .Z(n329) );
  NOR2_X1 U45 ( .A1(n86), .A2(n85), .ZN(n24) );
  XNOR2_X1 U46 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n27) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(n23), .ZN(n26) );
  XNOR2_X1 U48 ( .A(n329), .B(\mult_x_1/n285 ), .ZN(n43) );
  BUF_X2 U49 ( .A(n27), .Z(n114) );
  XNOR2_X1 U50 ( .A(n329), .B(\mult_x_1/n284 ), .ZN(n36) );
  OAI22_X1 U51 ( .A1(n113), .A2(n43), .B1(n114), .B2(n36), .ZN(n54) );
  XNOR2_X1 U52 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[4] ), .ZN(n28) );
  OR2_X2 U53 ( .A1(n28), .A2(n29), .ZN(n139) );
  BUF_X2 U54 ( .A(\mult_x_1/n311 ), .Z(n101) );
  XNOR2_X1 U55 ( .A(n101), .B(\mult_x_1/n283 ), .ZN(n39) );
  INV_X2 U56 ( .A(n29), .ZN(n207) );
  XNOR2_X1 U57 ( .A(n101), .B(\mult_x_1/n282 ), .ZN(n34) );
  OAI22_X1 U58 ( .A1(n139), .A2(n39), .B1(n207), .B2(n34), .ZN(n53) );
  XNOR2_X1 U59 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n30) );
  OR2_X2 U60 ( .A1(n31), .A2(n30), .ZN(n221) );
  BUF_X2 U61 ( .A(\mult_x_1/n312 ), .Z(n328) );
  XNOR2_X1 U62 ( .A(n328), .B(n15), .ZN(n40) );
  XNOR2_X1 U63 ( .A(n63), .B(n328), .ZN(n37) );
  INV_X1 U64 ( .A(n31), .ZN(n223) );
  OAI22_X1 U65 ( .A1(n221), .A2(n40), .B1(n223), .B2(n37), .ZN(n82) );
  INV_X1 U66 ( .A(n82), .ZN(n52) );
  XNOR2_X1 U67 ( .A(n19), .B(\mult_x_1/n285 ), .ZN(n33) );
  XNOR2_X1 U68 ( .A(n32), .B(n331), .ZN(n51) );
  NOR2_X1 U69 ( .A1(n33), .A2(n116), .ZN(n86) );
  XNOR2_X1 U70 ( .A(n101), .B(n15), .ZN(n64) );
  OAI22_X1 U71 ( .A1(n139), .A2(n34), .B1(n207), .B2(n64), .ZN(n85) );
  XNOR2_X1 U72 ( .A(n86), .B(n85), .ZN(n35) );
  XNOR2_X1 U73 ( .A(n84), .B(n35), .ZN(n182) );
  XNOR2_X1 U74 ( .A(n329), .B(\mult_x_1/n283 ), .ZN(n68) );
  OAI22_X1 U75 ( .A1(n113), .A2(n36), .B1(n114), .B2(n68), .ZN(n83) );
  AOI21_X1 U76 ( .B1(n7), .B2(n221), .A(n6), .ZN(n38) );
  INV_X1 U77 ( .A(n38), .ZN(n81) );
  XNOR2_X1 U78 ( .A(n101), .B(\mult_x_1/n284 ), .ZN(n137) );
  OAI22_X1 U79 ( .A1(n139), .A2(n137), .B1(n207), .B2(n39), .ZN(n46) );
  XNOR2_X1 U80 ( .A(n328), .B(\mult_x_1/n282 ), .ZN(n135) );
  OAI22_X1 U81 ( .A1(n221), .A2(n135), .B1(n223), .B2(n40), .ZN(n45) );
  OR2_X1 U82 ( .A1(n46), .A2(n45), .ZN(n57) );
  XNOR2_X1 U83 ( .A(n19), .B(\mult_x_1/n286 ), .ZN(n41) );
  NOR2_X1 U84 ( .A1(n41), .A2(n116), .ZN(n56) );
  XNOR2_X1 U85 ( .A(n63), .B(n327), .ZN(n50) );
  AOI21_X1 U86 ( .B1(n226), .B2(n20), .A(n14), .ZN(n42) );
  INV_X1 U87 ( .A(n42), .ZN(n145) );
  XNOR2_X1 U88 ( .A(n329), .B(\mult_x_1/n286 ), .ZN(n49) );
  OAI22_X1 U89 ( .A1(n113), .A2(n49), .B1(n114), .B2(n43), .ZN(n144) );
  XNOR2_X1 U90 ( .A(n19), .B(\mult_x_1/n287 ), .ZN(n44) );
  NOR2_X1 U91 ( .A1(n44), .A2(n116), .ZN(n143) );
  XNOR2_X1 U92 ( .A(n46), .B(n45), .ZN(n132) );
  INV_X1 U93 ( .A(n19), .ZN(n47) );
  OR2_X1 U94 ( .A1(\mult_x_1/n288 ), .A2(n47), .ZN(n48) );
  NOR2_X1 U95 ( .A1(n48), .A2(n116), .ZN(n131) );
  XNOR2_X1 U96 ( .A(n329), .B(\mult_x_1/n287 ), .ZN(n92) );
  OAI22_X1 U97 ( .A1(n113), .A2(n92), .B1(n114), .B2(n49), .ZN(n149) );
  XNOR2_X1 U98 ( .A(n327), .B(n15), .ZN(n94) );
  OAI22_X1 U99 ( .A1(n5), .A2(n94), .B1(n50), .B2(n20), .ZN(n148) );
  AND2_X1 U100 ( .A1(n51), .A2(\mult_x_1/n288 ), .ZN(n147) );
  FA_X1 U101 ( .A(n54), .B(n53), .CI(n52), .CO(n84), .S(n242) );
  FA_X1 U102 ( .A(n57), .B(n56), .CI(n55), .CO(n180), .S(n241) );
  NAND2_X1 U103 ( .A1(n189), .A2(n188), .ZN(n58) );
  NAND2_X1 U104 ( .A1(n58), .A2(n330), .ZN(n60) );
  OR2_X1 U105 ( .A1(n183), .A2(n387), .ZN(n59) );
  NAND2_X1 U106 ( .A1(n60), .A2(n59), .ZN(n378) );
  XNOR2_X1 U125 ( .A(n19), .B(\mult_x_1/n282 ), .ZN(n61) );
  NOR2_X1 U126 ( .A1(n61), .A2(n116), .ZN(n111) );
  XNOR2_X1 U127 ( .A(n329), .B(n15), .ZN(n62) );
  XNOR2_X1 U128 ( .A(n63), .B(n329), .ZN(n112) );
  OAI22_X1 U129 ( .A1(n8), .A2(n62), .B1(n112), .B2(n114), .ZN(n121) );
  INV_X1 U130 ( .A(n121), .ZN(n110) );
  XNOR2_X1 U131 ( .A(n329), .B(\mult_x_1/n282 ), .ZN(n67) );
  OAI22_X1 U132 ( .A1(n8), .A2(n67), .B1(n114), .B2(n62), .ZN(n73) );
  XNOR2_X1 U133 ( .A(n63), .B(n101), .ZN(n65) );
  OAI22_X1 U134 ( .A1(n139), .A2(n64), .B1(n65), .B2(n207), .ZN(n72) );
  AOI21_X1 U135 ( .B1(n207), .B2(n139), .A(n65), .ZN(n66) );
  INV_X1 U136 ( .A(n66), .ZN(n71) );
  INV_X1 U137 ( .A(n72), .ZN(n80) );
  OAI22_X1 U138 ( .A1(n113), .A2(n68), .B1(n114), .B2(n67), .ZN(n79) );
  XNOR2_X1 U139 ( .A(n19), .B(\mult_x_1/n284 ), .ZN(n69) );
  NOR2_X1 U140 ( .A1(n69), .A2(n116), .ZN(n78) );
  XNOR2_X1 U141 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n70) );
  NOR2_X1 U142 ( .A1(n70), .A2(n116), .ZN(n76) );
  FA_X1 U143 ( .A(n73), .B(n16), .CI(n71), .CO(n109), .S(n75) );
  OR2_X1 U144 ( .A1(n128), .A2(n127), .ZN(n74) );
  MUX2_X1 U145 ( .A(n332), .B(n74), .S(n183), .Z(n350) );
  FA_X1 U146 ( .A(n77), .B(n76), .CI(n75), .CO(n127), .S(n175) );
  FA_X1 U147 ( .A(n80), .B(n79), .CI(n78), .CO(n77), .S(n179) );
  FA_X1 U148 ( .A(n83), .B(n18), .CI(n81), .CO(n178), .S(n181) );
  INV_X1 U149 ( .A(n84), .ZN(n88) );
  NAND2_X1 U150 ( .A1(n86), .A2(n85), .ZN(n87) );
  OAI21_X1 U151 ( .B1(n88), .B2(n24), .A(n87), .ZN(n177) );
  OR2_X1 U152 ( .A1(n175), .A2(n174), .ZN(n89) );
  MUX2_X1 U153 ( .A(n333), .B(n89), .S(n183), .Z(n352) );
  XNOR2_X1 U154 ( .A(n327), .B(\mult_x_1/n283 ), .ZN(n198) );
  XNOR2_X1 U155 ( .A(n327), .B(\mult_x_1/n282 ), .ZN(n95) );
  OAI22_X1 U156 ( .A1(n226), .A2(n198), .B1(n95), .B2(n20), .ZN(n99) );
  INV_X1 U157 ( .A(n114), .ZN(n90) );
  AND2_X1 U158 ( .A1(\mult_x_1/n288 ), .A2(n90), .ZN(n98) );
  XNOR2_X1 U159 ( .A(n328), .B(\mult_x_1/n285 ), .ZN(n197) );
  XNOR2_X1 U160 ( .A(n328), .B(\mult_x_1/n284 ), .ZN(n96) );
  OAI22_X1 U161 ( .A1(n221), .A2(n197), .B1(n223), .B2(n96), .ZN(n97) );
  OR2_X1 U162 ( .A1(\mult_x_1/n288 ), .A2(n331), .ZN(n91) );
  OAI22_X1 U163 ( .A1(n8), .A2(n331), .B1(n91), .B2(n114), .ZN(n134) );
  XNOR2_X1 U164 ( .A(n329), .B(\mult_x_1/n288 ), .ZN(n93) );
  OAI22_X1 U165 ( .A1(n8), .A2(n93), .B1(n114), .B2(n92), .ZN(n133) );
  XNOR2_X1 U166 ( .A(n101), .B(\mult_x_1/n286 ), .ZN(n103) );
  XNOR2_X1 U167 ( .A(n101), .B(\mult_x_1/n285 ), .ZN(n138) );
  OAI22_X1 U168 ( .A1(n139), .A2(n103), .B1(n207), .B2(n138), .ZN(n152) );
  OAI22_X1 U169 ( .A1(n10), .A2(n95), .B1(n94), .B2(n20), .ZN(n151) );
  XNOR2_X1 U170 ( .A(n328), .B(\mult_x_1/n283 ), .ZN(n136) );
  OAI22_X1 U171 ( .A1(n221), .A2(n96), .B1(n7), .B2(n136), .ZN(n150) );
  FA_X1 U172 ( .A(n99), .B(n98), .CI(n97), .CO(n166), .S(n194) );
  OR2_X1 U173 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n100) );
  OAI22_X1 U174 ( .A1(n139), .A2(n22), .B1(n100), .B2(n207), .ZN(n196) );
  XNOR2_X1 U175 ( .A(n101), .B(\mult_x_1/n288 ), .ZN(n102) );
  XNOR2_X1 U176 ( .A(n101), .B(\mult_x_1/n287 ), .ZN(n104) );
  OAI22_X1 U177 ( .A1(n139), .A2(n102), .B1(n207), .B2(n104), .ZN(n195) );
  AND2_X1 U178 ( .A1(n196), .A2(n195), .ZN(n192) );
  OAI22_X1 U179 ( .A1(n139), .A2(n104), .B1(n207), .B2(n103), .ZN(n191) );
  OR2_X1 U180 ( .A1(n172), .A2(n171), .ZN(n108) );
  MUX2_X1 U181 ( .A(n334), .B(n108), .S(n183), .Z(n354) );
  FA_X1 U182 ( .A(n111), .B(n110), .CI(n109), .CO(n123), .S(n128) );
  AOI21_X1 U183 ( .B1(n114), .B2(n8), .A(n112), .ZN(n115) );
  INV_X1 U184 ( .A(n115), .ZN(n119) );
  XNOR2_X1 U185 ( .A(n19), .B(n15), .ZN(n117) );
  NOR2_X1 U186 ( .A1(n117), .A2(n116), .ZN(n118) );
  XOR2_X1 U187 ( .A(n119), .B(n118), .Z(n120) );
  XOR2_X1 U188 ( .A(n121), .B(n120), .Z(n122) );
  OR2_X1 U189 ( .A1(n123), .A2(n122), .ZN(n125) );
  NAND2_X1 U190 ( .A1(n123), .A2(n122), .ZN(n124) );
  NAND2_X1 U191 ( .A1(n125), .A2(n124), .ZN(n126) );
  MUX2_X1 U192 ( .A(n335), .B(n126), .S(n183), .Z(n356) );
  NAND2_X1 U193 ( .A1(n128), .A2(n127), .ZN(n129) );
  MUX2_X1 U194 ( .A(n336), .B(n129), .S(n183), .Z(n358) );
  FA_X1 U195 ( .A(n132), .B(n131), .CI(n130), .CO(n243), .S(n246) );
  HA_X1 U196 ( .A(n134), .B(n133), .CO(n156), .S(n165) );
  OAI22_X1 U197 ( .A1(n221), .A2(n136), .B1(n223), .B2(n135), .ZN(n153) );
  OAI22_X1 U198 ( .A1(n139), .A2(n138), .B1(n207), .B2(n137), .ZN(n154) );
  FA_X1 U199 ( .A(n145), .B(n144), .CI(n143), .CO(n55), .S(n248) );
  XNOR2_X1 U200 ( .A(n247), .B(n248), .ZN(n146) );
  XNOR2_X1 U201 ( .A(n246), .B(n146), .ZN(n159) );
  FA_X1 U202 ( .A(n149), .B(n148), .CI(n147), .CO(n130), .S(n163) );
  FA_X1 U203 ( .A(n152), .B(n151), .CI(n150), .CO(n162), .S(n164) );
  NOR2_X1 U204 ( .A1(n159), .A2(n158), .ZN(n157) );
  MUX2_X1 U205 ( .A(n337), .B(n157), .S(n183), .Z(n360) );
  NAND2_X1 U206 ( .A1(n159), .A2(n158), .ZN(n160) );
  MUX2_X1 U207 ( .A(n338), .B(n160), .S(n183), .Z(n362) );
  FA_X1 U208 ( .A(n163), .B(n162), .CI(n161), .CO(n158), .S(n169) );
  FA_X1 U209 ( .A(n166), .B(n165), .CI(n164), .CO(n168), .S(n172) );
  NOR2_X1 U210 ( .A1(n169), .A2(n168), .ZN(n167) );
  MUX2_X1 U211 ( .A(n339), .B(n167), .S(n183), .Z(n364) );
  NAND2_X1 U212 ( .A1(n169), .A2(n168), .ZN(n170) );
  MUX2_X1 U213 ( .A(n340), .B(n170), .S(n183), .Z(n366) );
  NAND2_X1 U214 ( .A1(n172), .A2(n171), .ZN(n173) );
  MUX2_X1 U215 ( .A(n341), .B(n173), .S(n183), .Z(n368) );
  NAND2_X1 U216 ( .A1(n175), .A2(n174), .ZN(n176) );
  MUX2_X1 U217 ( .A(n342), .B(n176), .S(n183), .Z(n370) );
  FA_X1 U218 ( .A(n179), .B(n178), .CI(n177), .CO(n174), .S(n186) );
  FA_X1 U219 ( .A(n182), .B(n181), .CI(n180), .CO(n185), .S(n189) );
  NAND2_X1 U220 ( .A1(n186), .A2(n185), .ZN(n184) );
  MUX2_X1 U221 ( .A(n343), .B(n184), .S(n183), .Z(n372) );
  OR2_X1 U222 ( .A1(n186), .A2(n185), .ZN(n187) );
  MUX2_X1 U223 ( .A(n344), .B(n187), .S(n330), .Z(n374) );
  NOR2_X1 U224 ( .A1(n189), .A2(n188), .ZN(n190) );
  MUX2_X1 U225 ( .A(n345), .B(n190), .S(n183), .Z(n376) );
  XNOR2_X1 U226 ( .A(n328), .B(\mult_x_1/n286 ), .ZN(n209) );
  OAI22_X1 U227 ( .A1(n221), .A2(n209), .B1(n223), .B2(n197), .ZN(n203) );
  XNOR2_X1 U228 ( .A(n327), .B(\mult_x_1/n284 ), .ZN(n206) );
  OAI22_X1 U229 ( .A1(n226), .A2(n206), .B1(n198), .B2(n20), .ZN(n201) );
  NOR2_X1 U230 ( .A1(n203), .A2(n201), .ZN(n200) );
  NAND2_X1 U231 ( .A1(n203), .A2(n201), .ZN(n199) );
  OR2_X1 U232 ( .A1(n237), .A2(n236), .ZN(n281) );
  INV_X1 U233 ( .A(n281), .ZN(n239) );
  INV_X1 U234 ( .A(n201), .ZN(n202) );
  XNOR2_X1 U235 ( .A(n327), .B(\mult_x_1/n285 ), .ZN(n217) );
  OAI22_X1 U236 ( .A1(n226), .A2(n217), .B1(n206), .B2(n20), .ZN(n214) );
  INV_X1 U237 ( .A(n207), .ZN(n208) );
  AND2_X1 U238 ( .A1(\mult_x_1/n288 ), .A2(n208), .ZN(n213) );
  XNOR2_X1 U239 ( .A(n328), .B(\mult_x_1/n287 ), .ZN(n215) );
  OAI22_X1 U240 ( .A1(n221), .A2(n215), .B1(n223), .B2(n209), .ZN(n212) );
  NAND2_X1 U241 ( .A1(n211), .A2(n210), .ZN(n275) );
  OR2_X1 U242 ( .A1(n211), .A2(n210), .ZN(n276) );
  FA_X1 U243 ( .A(n214), .B(n213), .CI(n212), .CO(n210), .S(n234) );
  XNOR2_X1 U244 ( .A(n328), .B(\mult_x_1/n288 ), .ZN(n216) );
  OAI22_X1 U245 ( .A1(n221), .A2(n216), .B1(n223), .B2(n215), .ZN(n219) );
  XNOR2_X1 U246 ( .A(n327), .B(\mult_x_1/n286 ), .ZN(n222) );
  OAI22_X1 U247 ( .A1(n226), .A2(n222), .B1(n217), .B2(n20), .ZN(n218) );
  NOR2_X1 U248 ( .A1(n234), .A2(n233), .ZN(n269) );
  HA_X1 U249 ( .A(n219), .B(n218), .CO(n233), .S(n231) );
  OR2_X1 U250 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n220) );
  OAI22_X1 U251 ( .A1(n221), .A2(n21), .B1(n220), .B2(n7), .ZN(n230) );
  OR2_X1 U252 ( .A1(n231), .A2(n230), .ZN(n265) );
  XNOR2_X1 U253 ( .A(n327), .B(\mult_x_1/n287 ), .ZN(n225) );
  OAI22_X1 U254 ( .A1(n10), .A2(n225), .B1(n222), .B2(n20), .ZN(n229) );
  INV_X1 U255 ( .A(n223), .ZN(n224) );
  AND2_X1 U256 ( .A1(\mult_x_1/n288 ), .A2(n224), .ZN(n228) );
  NOR2_X1 U257 ( .A1(n229), .A2(n228), .ZN(n258) );
  OAI22_X1 U258 ( .A1(n10), .A2(\mult_x_1/n288 ), .B1(n225), .B2(n20), .ZN(
        n255) );
  OR2_X1 U259 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n227) );
  NAND2_X1 U260 ( .A1(n227), .A2(n10), .ZN(n254) );
  NAND2_X1 U261 ( .A1(n255), .A2(n254), .ZN(n261) );
  NAND2_X1 U262 ( .A1(n229), .A2(n228), .ZN(n259) );
  OAI21_X1 U263 ( .B1(n258), .B2(n261), .A(n259), .ZN(n266) );
  NAND2_X1 U264 ( .A1(n231), .A2(n230), .ZN(n264) );
  INV_X1 U265 ( .A(n264), .ZN(n232) );
  AOI21_X1 U266 ( .B1(n265), .B2(n266), .A(n232), .ZN(n272) );
  NAND2_X1 U267 ( .A1(n234), .A2(n233), .ZN(n270) );
  OAI21_X1 U268 ( .B1(n269), .B2(n272), .A(n270), .ZN(n277) );
  NAND2_X1 U269 ( .A1(n276), .A2(n277), .ZN(n235) );
  NAND2_X1 U270 ( .A1(n275), .A2(n235), .ZN(n283) );
  INV_X1 U271 ( .A(n283), .ZN(n238) );
  NAND2_X1 U272 ( .A1(n237), .A2(n236), .ZN(n280) );
  OAI21_X1 U273 ( .B1(n239), .B2(n238), .A(n280), .ZN(n240) );
  MUX2_X1 U274 ( .A(n347), .B(n240), .S(n330), .Z(n380) );
  FA_X1 U275 ( .A(n243), .B(n242), .CI(n241), .CO(n188), .S(n244) );
  MUX2_X1 U276 ( .A(n348), .B(n244), .S(n330), .Z(n382) );
  NAND2_X1 U277 ( .A1(n250), .A2(n249), .ZN(n251) );
  MUX2_X1 U278 ( .A(n349), .B(n251), .S(n183), .Z(n384) );
  BUF_X2 U279 ( .A(rst_n), .Z(n394) );
  BUF_X1 U280 ( .A(rst_n), .Z(n252) );
  BUF_X4 U281 ( .A(en), .Z(n287) );
  MUX2_X1 U282 ( .A(product[0]), .B(n508), .S(n287), .Z(n396) );
  MUX2_X1 U283 ( .A(n508), .B(n509), .S(n287), .Z(n398) );
  AND2_X1 U284 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n253) );
  MUX2_X1 U285 ( .A(n509), .B(n253), .S(n287), .Z(n400) );
  MUX2_X1 U286 ( .A(product[1]), .B(n511), .S(n287), .Z(n402) );
  MUX2_X1 U287 ( .A(n511), .B(n512), .S(n287), .Z(n404) );
  OR2_X1 U288 ( .A1(n255), .A2(n254), .ZN(n256) );
  AND2_X1 U289 ( .A1(n256), .A2(n261), .ZN(n257) );
  MUX2_X1 U290 ( .A(n512), .B(n257), .S(n287), .Z(n406) );
  MUX2_X1 U291 ( .A(product[2]), .B(n514), .S(n287), .Z(n408) );
  MUX2_X1 U292 ( .A(n514), .B(n515), .S(n287), .Z(n410) );
  INV_X1 U293 ( .A(n258), .ZN(n260) );
  NAND2_X1 U294 ( .A1(n260), .A2(n259), .ZN(n262) );
  XOR2_X1 U295 ( .A(n262), .B(n261), .Z(n263) );
  MUX2_X1 U296 ( .A(n515), .B(n263), .S(n287), .Z(n412) );
  MUX2_X1 U297 ( .A(product[3]), .B(n517), .S(n287), .Z(n414) );
  MUX2_X1 U298 ( .A(n517), .B(n518), .S(n287), .Z(n416) );
  NAND2_X1 U299 ( .A1(n265), .A2(n264), .ZN(n267) );
  XNOR2_X1 U300 ( .A(n267), .B(n266), .ZN(n268) );
  MUX2_X1 U301 ( .A(n518), .B(n268), .S(n287), .Z(n418) );
  MUX2_X1 U302 ( .A(product[4]), .B(n520), .S(n287), .Z(n420) );
  MUX2_X1 U303 ( .A(n520), .B(n521), .S(n287), .Z(n422) );
  INV_X1 U304 ( .A(n269), .ZN(n271) );
  NAND2_X1 U305 ( .A1(n271), .A2(n270), .ZN(n273) );
  XOR2_X1 U306 ( .A(n273), .B(n17), .Z(n274) );
  MUX2_X1 U307 ( .A(n521), .B(n274), .S(n287), .Z(n424) );
  MUX2_X1 U308 ( .A(product[5]), .B(n523), .S(n287), .Z(n426) );
  MUX2_X1 U309 ( .A(n523), .B(n524), .S(n287), .Z(n428) );
  NAND2_X1 U310 ( .A1(n276), .A2(n275), .ZN(n278) );
  XNOR2_X1 U311 ( .A(n278), .B(n13), .ZN(n279) );
  MUX2_X1 U312 ( .A(n524), .B(n279), .S(n287), .Z(n430) );
  MUX2_X1 U313 ( .A(product[6]), .B(n526), .S(n287), .Z(n432) );
  MUX2_X1 U314 ( .A(n526), .B(n527), .S(n287), .Z(n434) );
  NAND2_X1 U315 ( .A1(n281), .A2(n280), .ZN(n282) );
  XNOR2_X1 U316 ( .A(n283), .B(n282), .ZN(n284) );
  MUX2_X1 U317 ( .A(n527), .B(n284), .S(n287), .Z(n436) );
  MUX2_X1 U318 ( .A(product[7]), .B(n529), .S(n287), .Z(n438) );
  NAND2_X1 U319 ( .A1(n334), .A2(n341), .ZN(n285) );
  XNOR2_X1 U320 ( .A(n347), .B(n285), .ZN(n286) );
  MUX2_X1 U321 ( .A(n529), .B(n286), .S(n287), .Z(n440) );
  MUX2_X1 U322 ( .A(product[8]), .B(n531), .S(n287), .Z(n442) );
  AOI21_X1 U323 ( .B1(n347), .B2(n334), .A(n389), .ZN(n290) );
  NAND2_X1 U324 ( .A1(n390), .A2(n340), .ZN(n288) );
  XOR2_X1 U325 ( .A(n290), .B(n288), .Z(n289) );
  BUF_X4 U326 ( .A(en), .Z(n330) );
  MUX2_X1 U327 ( .A(n531), .B(n289), .S(n330), .Z(n444) );
  MUX2_X1 U328 ( .A(product[9]), .B(n533), .S(n330), .Z(n446) );
  OAI21_X1 U329 ( .B1(n290), .B2(n339), .A(n340), .ZN(n301) );
  INV_X1 U330 ( .A(n301), .ZN(n293) );
  NAND2_X1 U331 ( .A1(n391), .A2(n338), .ZN(n291) );
  XOR2_X1 U332 ( .A(n293), .B(n291), .Z(n292) );
  MUX2_X1 U333 ( .A(n533), .B(n292), .S(n330), .Z(n448) );
  MUX2_X1 U334 ( .A(product[10]), .B(n535), .S(n330), .Z(n450) );
  OAI21_X1 U335 ( .B1(n293), .B2(n337), .A(n338), .ZN(n296) );
  NOR2_X1 U336 ( .A1(n348), .A2(n349), .ZN(n299) );
  INV_X1 U337 ( .A(n299), .ZN(n294) );
  NAND2_X1 U338 ( .A1(n348), .A2(n349), .ZN(n298) );
  NAND2_X1 U339 ( .A1(n294), .A2(n298), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U341 ( .A(n535), .B(n297), .S(n330), .Z(n452) );
  MUX2_X1 U342 ( .A(product[11]), .B(n537), .S(n330), .Z(n454) );
  NOR2_X1 U343 ( .A1(n299), .A2(n337), .ZN(n302) );
  OAI21_X1 U344 ( .B1(n299), .B2(n338), .A(n298), .ZN(n300) );
  AOI21_X1 U345 ( .B1(n302), .B2(n301), .A(n300), .ZN(n324) );
  NAND2_X1 U346 ( .A1(n392), .A2(n346), .ZN(n303) );
  XOR2_X1 U347 ( .A(n324), .B(n303), .Z(n304) );
  MUX2_X1 U348 ( .A(n537), .B(n304), .S(n330), .Z(n456) );
  MUX2_X1 U349 ( .A(product[12]), .B(n539), .S(n330), .Z(n458) );
  OAI21_X1 U350 ( .B1(n324), .B2(n345), .A(n346), .ZN(n306) );
  NAND2_X1 U351 ( .A1(n344), .A2(n343), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U353 ( .A(n539), .B(n307), .S(n330), .Z(n460) );
  MUX2_X1 U354 ( .A(product[13]), .B(n541), .S(n330), .Z(n462) );
  NAND2_X1 U355 ( .A1(n392), .A2(n344), .ZN(n309) );
  AOI21_X1 U356 ( .B1(n387), .B2(n344), .A(n393), .ZN(n308) );
  OAI21_X1 U357 ( .B1(n324), .B2(n309), .A(n308), .ZN(n311) );
  NAND2_X1 U358 ( .A1(n333), .A2(n342), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  MUX2_X1 U360 ( .A(n541), .B(n312), .S(n330), .Z(n464) );
  MUX2_X1 U361 ( .A(product[14]), .B(n543), .S(n330), .Z(n466) );
  NAND2_X1 U362 ( .A1(n344), .A2(n333), .ZN(n314) );
  NOR2_X1 U363 ( .A1(n345), .A2(n314), .ZN(n320) );
  INV_X1 U364 ( .A(n320), .ZN(n316) );
  AOI21_X1 U365 ( .B1(n393), .B2(n333), .A(n388), .ZN(n313) );
  OAI21_X1 U366 ( .B1(n314), .B2(n346), .A(n313), .ZN(n321) );
  INV_X1 U367 ( .A(n321), .ZN(n315) );
  OAI21_X1 U368 ( .B1(n324), .B2(n316), .A(n315), .ZN(n318) );
  NAND2_X1 U369 ( .A1(n332), .A2(n336), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U371 ( .A(n543), .B(n319), .S(n330), .Z(n468) );
  MUX2_X1 U372 ( .A(product[15]), .B(n545), .S(n330), .Z(n470) );
  NAND2_X1 U373 ( .A1(n320), .A2(n332), .ZN(n323) );
  AOI21_X1 U374 ( .B1(n321), .B2(n332), .A(n386), .ZN(n322) );
  OAI21_X1 U375 ( .B1(n324), .B2(n323), .A(n322), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n325), .B(n335), .ZN(n326) );
  MUX2_X1 U377 ( .A(n545), .B(n326), .S(n330), .Z(n472) );
  MUX2_X1 U378 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n330), .Z(n474) );
  MUX2_X1 U379 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n330), .Z(n476) );
  MUX2_X1 U380 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n330), .Z(n478) );
  MUX2_X1 U381 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n330), .Z(n480) );
  MUX2_X1 U382 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n330), .Z(n482) );
  MUX2_X1 U383 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n330), .Z(n484) );
  MUX2_X1 U384 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n330), .Z(n486) );
  MUX2_X1 U385 ( .A(n15), .B(B_extended[7]), .S(n330), .Z(n488) );
  MUX2_X1 U386 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n330), .Z(n490) );
  MUX2_X1 U387 ( .A(n327), .B(A_extended[1]), .S(n330), .Z(n492) );
  MUX2_X1 U388 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n330), .Z(n494) );
  MUX2_X1 U389 ( .A(n328), .B(A_extended[3]), .S(n330), .Z(n496) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n330), .Z(n498) );
  MUX2_X1 U391 ( .A(\mult_x_1/n311 ), .B(A_extended[5]), .S(n330), .Z(n500) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n330), .Z(n502) );
  MUX2_X1 U393 ( .A(n329), .B(A_extended[7]), .S(n330), .Z(n504) );
  OR2_X1 U394 ( .A1(n330), .A2(n547), .ZN(n506) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_23 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n346, n348, n350, n352, n354, n356, n358,
         n360, n362, n364, n366, n368, n370, n372, n374, n376, n378, n380,
         n382, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n396, n398, n400, n402, n404, n406, n408, n410, n412, n414,
         n416, n418, n420, n422, n424, n426, n428, n430, n432, n434, n436,
         n438, n440, n442, n444, n446, n448, n450, n452, n454, n456, n458,
         n460, n462, n464, n466, n468, n470, n472, n474, n476, n478, n480,
         n482, n484, n486, n488, n490, n492, n494, n496, n498, n500, n502,
         n504, n506, n507, n509, n510, n512, n513, n515, n516, n518, n519,
         n521, n522, n524, n526, n528, n530, n532, n534, n536, n538, n540,
         n542, n543, n544, n545, n546;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n504), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n393), .SE(n500), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n27) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n393), .SE(n498), .CK(clk), .Q(n544), 
        .QN(n25) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n394), .SE(n496), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n16) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n394), .SE(n494), .CK(clk), .Q(n543), 
        .QN(n322) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n393), .SE(n492), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n14) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n393), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n18) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n394), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n23) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n394), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n24) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n393), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n21) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n393), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n22) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n394), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n19) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n394), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n20) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n393), .SE(n472), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n321) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n394), .SE(n470), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n393), .SE(n468), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n393), .SE(n466), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n394), .SE(n464), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n394), .SE(n462), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n393), .SE(n460), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n394), .SE(n458), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n393), .SE(n456), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n394), .SE(n454), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n393), .SE(n452), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n394), .SE(n450), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n393), .SE(n448), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n442), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n440), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n394), .SE(n438), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n394), .SE(n436), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n394), .SE(n434), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n394), .SE(n432), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n394), .SE(n430), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n394), .SE(n428), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n394), .SE(n426), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n394), .SE(n424), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n394), .SE(n422), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n394), .SE(n420), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n394), .SE(n418), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n393), .SE(n416), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n393), .SE(n414), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n393), .SE(n412), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n393), .SE(n410), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n393), .SE(n408), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n393), .SE(n406), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n393), .SE(n404), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n393), .SE(n402), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n393), .SE(n400), .CK(clk), .Q(n507)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n393), .SE(n398), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n393), .SE(n396), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n394), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n29) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n546), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n546), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n342), .QN(n384) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n546), .SE(n378), .CK(
        clk), .Q(n31), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n546), .SE(n376), .CK(
        clk), .Q(n323), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n546), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n339), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n546), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n546), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n337), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n546), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n336), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n546), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n546), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n334), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n546), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n546), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n332), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n546), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n331), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n546), .SE(n356), .CK(
        clk), .Q(n391), .QN(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n546), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n329), .QN(n385) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n546), .SE(n352), .CK(
        clk), .QN(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n546), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n546), .SE(n348), .CK(
        clk), .QN(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n546), .SI(1'b1), .SE(n346), .CK(clk), 
        .Q(n325), .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n546), .SI(1'b1), .SE(n344), .CK(clk), 
        .Q(n324) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n393), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n17) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n394), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  BUF_X1 U2 ( .A(en), .Z(n192) );
  MUX2_X1 U3 ( .A(n331), .B(n104), .S(n192), .Z(n358) );
  BUF_X1 U4 ( .A(n45), .Z(n151) );
  BUF_X1 U5 ( .A(n6), .Z(n11) );
  INV_X2 U6 ( .A(n10), .ZN(n149) );
  XNOR2_X1 U7 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n6) );
  OR2_X1 U8 ( .A1(n29), .A2(\mult_x_1/n180 ), .ZN(n236) );
  NAND2_X1 U9 ( .A1(n32), .A2(n12), .ZN(n7) );
  NAND2_X1 U10 ( .A1(n32), .A2(n12), .ZN(n132) );
  AND2_X1 U11 ( .A1(\mult_x_1/n310 ), .A2(n545), .ZN(n35) );
  INV_X1 U12 ( .A(n168), .ZN(n58) );
  INV_X1 U13 ( .A(n167), .ZN(n59) );
  NAND2_X1 U14 ( .A1(n112), .A2(n111), .ZN(n113) );
  XNOR2_X1 U15 ( .A(n168), .B(n167), .ZN(n169) );
  NAND2_X1 U16 ( .A1(n62), .A2(n61), .ZN(n95) );
  NAND2_X1 U17 ( .A1(n167), .A2(n168), .ZN(n61) );
  NAND2_X1 U18 ( .A1(n114), .A2(n113), .ZN(n139) );
  OAI21_X1 U19 ( .B1(n112), .B2(n111), .A(n110), .ZN(n114) );
  NAND2_X1 U20 ( .A1(n94), .A2(n93), .ZN(n346) );
  OR2_X1 U21 ( .A1(n192), .A2(n28), .ZN(n93) );
  OAI21_X1 U22 ( .B1(n210), .B2(n209), .A(n192), .ZN(n94) );
  BUF_X1 U23 ( .A(n125), .Z(n201) );
  CLKBUF_X1 U24 ( .A(n125), .Z(n231) );
  INV_X1 U25 ( .A(n18), .ZN(n8) );
  BUF_X2 U26 ( .A(n33), .Z(n9) );
  XOR2_X1 U27 ( .A(n544), .B(\mult_x_1/a[6] ), .Z(n10) );
  XNOR2_X1 U28 ( .A(n16), .B(n322), .ZN(n12) );
  INV_X1 U29 ( .A(n72), .ZN(n13) );
  XOR2_X1 U30 ( .A(n14), .B(n322), .Z(n34) );
  INV_X2 U31 ( .A(n17), .ZN(n15) );
  XNOR2_X1 U32 ( .A(n16), .B(n322), .ZN(n33) );
  BUF_X1 U33 ( .A(en), .Z(n248) );
  BUF_X1 U34 ( .A(rst_n), .Z(n393) );
  BUF_X1 U35 ( .A(rst_n), .Z(n394) );
  INV_X1 U36 ( .A(rst_n), .ZN(n546) );
  BUF_X2 U37 ( .A(n544), .Z(n319) );
  XOR2_X1 U38 ( .A(n49), .B(n48), .Z(n26) );
  AND2_X1 U39 ( .A1(n49), .A2(n48), .ZN(n30) );
  XOR2_X1 U40 ( .A(\mult_x_1/a[4] ), .B(n544), .Z(n32) );
  XNOR2_X1 U41 ( .A(n319), .B(\mult_x_1/n284 ), .ZN(n53) );
  XNOR2_X1 U42 ( .A(n319), .B(\mult_x_1/n283 ), .ZN(n41) );
  OAI22_X1 U43 ( .A1(n7), .A2(n53), .B1(n9), .B2(n41), .ZN(n44) );
  NAND2_X1 U44 ( .A1(n34), .A2(n6), .ZN(n125) );
  XNOR2_X1 U45 ( .A(n543), .B(\mult_x_1/n282 ), .ZN(n54) );
  XNOR2_X1 U46 ( .A(n543), .B(\mult_x_1/n281 ), .ZN(n42) );
  OAI22_X1 U47 ( .A1(n125), .A2(n54), .B1(n11), .B2(n42), .ZN(n43) );
  OR2_X1 U48 ( .A1(n44), .A2(n43), .ZN(n82) );
  XNOR2_X1 U49 ( .A(n35), .B(n15), .ZN(n45) );
  NOR2_X1 U50 ( .A1(n19), .A2(n151), .ZN(n81) );
  XNOR2_X1 U51 ( .A(n82), .B(n81), .ZN(n38) );
  BUF_X2 U52 ( .A(\mult_x_1/n313 ), .Z(n235) );
  AND2_X1 U53 ( .A1(n545), .A2(\mult_x_1/n281 ), .ZN(n105) );
  XNOR2_X1 U54 ( .A(n105), .B(n235), .ZN(n46) );
  AOI21_X1 U55 ( .B1(n236), .B2(n5), .A(n46), .ZN(n36) );
  INV_X1 U56 ( .A(n36), .ZN(n52) );
  NOR2_X1 U57 ( .A1(n20), .A2(n45), .ZN(n51) );
  XNOR2_X1 U58 ( .A(\mult_x_1/n310 ), .B(n27), .ZN(n37) );
  XNOR2_X1 U59 ( .A(n544), .B(\mult_x_1/a[6] ), .ZN(n39) );
  NAND2_X2 U60 ( .A1(n37), .A2(n39), .ZN(n148) );
  XNOR2_X1 U61 ( .A(n15), .B(\mult_x_1/n286 ), .ZN(n47) );
  XNOR2_X1 U62 ( .A(n15), .B(\mult_x_1/n285 ), .ZN(n40) );
  OAI22_X1 U63 ( .A1(n148), .A2(n47), .B1(n149), .B2(n40), .ZN(n50) );
  XNOR2_X1 U64 ( .A(n38), .B(n80), .ZN(n103) );
  XNOR2_X1 U65 ( .A(n15), .B(\mult_x_1/n284 ), .ZN(n69) );
  OAI22_X1 U66 ( .A1(n148), .A2(n40), .B1(n149), .B2(n69), .ZN(n74) );
  XNOR2_X1 U67 ( .A(n319), .B(\mult_x_1/n282 ), .ZN(n76) );
  OAI22_X1 U68 ( .A1(n7), .A2(n41), .B1(n9), .B2(n76), .ZN(n73) );
  XNOR2_X1 U69 ( .A(n105), .B(n543), .ZN(n70) );
  OAI22_X1 U70 ( .A1(n125), .A2(n42), .B1(n70), .B2(n6), .ZN(n87) );
  INV_X1 U71 ( .A(n87), .ZN(n72) );
  XNOR2_X1 U72 ( .A(n44), .B(n43), .ZN(n49) );
  NOR2_X1 U73 ( .A1(n321), .A2(n45), .ZN(n172) );
  XNOR2_X1 U74 ( .A(n235), .B(n8), .ZN(n123) );
  OAI22_X1 U75 ( .A1(n236), .A2(n123), .B1(n46), .B2(n5), .ZN(n171) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n56) );
  OAI22_X1 U77 ( .A1(n148), .A2(n56), .B1(n149), .B2(n47), .ZN(n170) );
  INV_X1 U78 ( .A(n248), .ZN(n66) );
  FA_X1 U79 ( .A(n52), .B(n51), .CI(n50), .CO(n80), .S(n167) );
  XNOR2_X1 U80 ( .A(n319), .B(\mult_x_1/n285 ), .ZN(n122) );
  OAI22_X1 U81 ( .A1(n7), .A2(n122), .B1(n9), .B2(n53), .ZN(n178) );
  XNOR2_X1 U82 ( .A(n543), .B(\mult_x_1/n283 ), .ZN(n126) );
  OAI22_X1 U83 ( .A1(n201), .A2(n126), .B1(n11), .B2(n54), .ZN(n177) );
  OR2_X1 U84 ( .A1(\mult_x_1/n288 ), .A2(n17), .ZN(n55) );
  OAI22_X1 U85 ( .A1(n148), .A2(n17), .B1(n149), .B2(n55), .ZN(n121) );
  XNOR2_X1 U86 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n57) );
  OAI22_X1 U87 ( .A1(n148), .A2(n57), .B1(n149), .B2(n56), .ZN(n120) );
  NAND2_X1 U88 ( .A1(n59), .A2(n58), .ZN(n60) );
  NAND2_X1 U89 ( .A1(n26), .A2(n60), .ZN(n62) );
  OR2_X1 U90 ( .A1(n248), .A2(n31), .ZN(n63) );
  OAI21_X1 U91 ( .B1(n95), .B2(n66), .A(n63), .ZN(n64) );
  INV_X1 U92 ( .A(n64), .ZN(n65) );
  OAI21_X1 U93 ( .B1(n98), .B2(n66), .A(n65), .ZN(n378) );
  XNOR2_X1 U94 ( .A(n15), .B(\mult_x_1/n283 ), .ZN(n68) );
  XNOR2_X1 U95 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n107) );
  OAI22_X1 U96 ( .A1(n148), .A2(n68), .B1(n149), .B2(n107), .ZN(n111) );
  XNOR2_X1 U97 ( .A(n319), .B(\mult_x_1/n281 ), .ZN(n75) );
  XNOR2_X1 U98 ( .A(n105), .B(n319), .ZN(n108) );
  OAI22_X1 U99 ( .A1(n132), .A2(n75), .B1(n108), .B2(n9), .ZN(n115) );
  INV_X1 U100 ( .A(n115), .ZN(n110) );
  XNOR2_X1 U101 ( .A(n111), .B(n110), .ZN(n67) );
  NOR2_X1 U102 ( .A1(n21), .A2(n151), .ZN(n112) );
  XNOR2_X1 U103 ( .A(n67), .B(n112), .ZN(n142) );
  OAI22_X1 U104 ( .A1(n148), .A2(n69), .B1(n149), .B2(n68), .ZN(n88) );
  AOI21_X1 U105 ( .B1(n11), .B2(n201), .A(n70), .ZN(n71) );
  INV_X1 U106 ( .A(n71), .ZN(n86) );
  FA_X1 U107 ( .A(n73), .B(n74), .CI(n72), .CO(n92), .S(n102) );
  NOR2_X1 U108 ( .A1(n22), .A2(n151), .ZN(n90) );
  OAI22_X1 U109 ( .A1(n7), .A2(n76), .B1(n9), .B2(n75), .ZN(n89) );
  OR2_X1 U110 ( .A1(n90), .A2(n89), .ZN(n77) );
  NAND2_X1 U111 ( .A1(n92), .A2(n77), .ZN(n79) );
  NAND2_X1 U112 ( .A1(n90), .A2(n89), .ZN(n78) );
  NAND2_X1 U113 ( .A1(n79), .A2(n78), .ZN(n140) );
  INV_X1 U114 ( .A(n80), .ZN(n85) );
  NOR2_X1 U115 ( .A1(n82), .A2(n81), .ZN(n84) );
  NAND2_X1 U116 ( .A1(n82), .A2(n81), .ZN(n83) );
  OAI21_X1 U117 ( .B1(n85), .B2(n84), .A(n83), .ZN(n101) );
  FA_X1 U118 ( .A(n88), .B(n13), .CI(n86), .CO(n141), .S(n100) );
  XNOR2_X1 U119 ( .A(n90), .B(n89), .ZN(n91) );
  XNOR2_X1 U120 ( .A(n92), .B(n91), .ZN(n99) );
  INV_X1 U121 ( .A(n95), .ZN(n96) );
  NAND2_X1 U122 ( .A1(n96), .A2(n248), .ZN(n97) );
  OAI22_X1 U123 ( .A1(n98), .A2(n97), .B1(n248), .B2(n323), .ZN(n376) );
  FA_X1 U124 ( .A(n101), .B(n100), .CI(n99), .CO(n209), .S(n165) );
  FA_X1 U125 ( .A(n103), .B(n102), .CI(n30), .CO(n164), .S(n98) );
  NAND2_X1 U126 ( .A1(n165), .A2(n164), .ZN(n104) );
  NOR2_X1 U147 ( .A1(n23), .A2(n151), .ZN(n146) );
  XNOR2_X1 U148 ( .A(n15), .B(n8), .ZN(n106) );
  XNOR2_X1 U149 ( .A(n105), .B(n15), .ZN(n147) );
  OAI22_X1 U150 ( .A1(n148), .A2(n106), .B1(n147), .B2(n149), .ZN(n155) );
  INV_X1 U151 ( .A(n155), .ZN(n145) );
  OAI22_X1 U152 ( .A1(n148), .A2(n107), .B1(n149), .B2(n106), .ZN(n117) );
  AOI21_X1 U153 ( .B1(n9), .B2(n132), .A(n108), .ZN(n109) );
  INV_X1 U154 ( .A(n109), .ZN(n116) );
  NOR2_X1 U155 ( .A1(n24), .A2(n151), .ZN(n138) );
  FA_X1 U156 ( .A(n117), .B(n116), .CI(n115), .CO(n144), .S(n137) );
  OR2_X1 U157 ( .A1(n162), .A2(n161), .ZN(n118) );
  MUX2_X1 U158 ( .A(n324), .B(n118), .S(n192), .Z(n344) );
  XNOR2_X1 U159 ( .A(n235), .B(\mult_x_1/n283 ), .ZN(n202) );
  XNOR2_X1 U160 ( .A(n235), .B(\mult_x_1/n282 ), .ZN(n124) );
  OAI22_X1 U161 ( .A1(n236), .A2(n202), .B1(n124), .B2(n5), .ZN(n135) );
  INV_X1 U162 ( .A(n149), .ZN(n119) );
  AND2_X1 U163 ( .A1(\mult_x_1/n288 ), .A2(n119), .ZN(n134) );
  XNOR2_X1 U164 ( .A(n543), .B(\mult_x_1/n285 ), .ZN(n200) );
  XNOR2_X1 U165 ( .A(n543), .B(\mult_x_1/n284 ), .ZN(n127) );
  OAI22_X1 U166 ( .A1(n201), .A2(n200), .B1(n11), .B2(n127), .ZN(n133) );
  HA_X1 U167 ( .A(n121), .B(n120), .CO(n176), .S(n187) );
  XNOR2_X1 U168 ( .A(n319), .B(\mult_x_1/n286 ), .ZN(n130) );
  OAI22_X1 U169 ( .A1(n7), .A2(n130), .B1(n9), .B2(n122), .ZN(n175) );
  OAI22_X1 U170 ( .A1(n236), .A2(n124), .B1(n123), .B2(n5), .ZN(n174) );
  OAI22_X1 U171 ( .A1(n231), .A2(n127), .B1(n11), .B2(n126), .ZN(n173) );
  OR2_X1 U172 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n128) );
  OAI22_X1 U173 ( .A1(n132), .A2(n25), .B1(n128), .B2(n9), .ZN(n204) );
  XNOR2_X1 U174 ( .A(n319), .B(\mult_x_1/n288 ), .ZN(n129) );
  XNOR2_X1 U175 ( .A(n319), .B(\mult_x_1/n287 ), .ZN(n131) );
  OAI22_X1 U176 ( .A1(n132), .A2(n129), .B1(n9), .B2(n131), .ZN(n203) );
  OAI22_X1 U177 ( .A1(n7), .A2(n131), .B1(n9), .B2(n130), .ZN(n198) );
  FA_X1 U178 ( .A(n135), .B(n134), .CI(n133), .CO(n188), .S(n197) );
  OR2_X1 U179 ( .A1(n195), .A2(n194), .ZN(n136) );
  MUX2_X1 U180 ( .A(n326), .B(n136), .S(n192), .Z(n348) );
  FA_X1 U181 ( .A(n139), .B(n138), .CI(n137), .CO(n161), .S(n213) );
  FA_X1 U182 ( .A(n140), .B(n141), .CI(n142), .CO(n212), .S(n210) );
  OR2_X1 U183 ( .A1(n213), .A2(n212), .ZN(n143) );
  MUX2_X1 U184 ( .A(n327), .B(n143), .S(n192), .Z(n350) );
  FA_X1 U185 ( .A(n146), .B(n145), .CI(n144), .CO(n157), .S(n162) );
  AOI21_X1 U186 ( .B1(n148), .B2(n149), .A(n147), .ZN(n150) );
  INV_X1 U187 ( .A(n150), .ZN(n153) );
  NOR2_X1 U188 ( .A1(n18), .A2(n151), .ZN(n152) );
  XOR2_X1 U189 ( .A(n153), .B(n152), .Z(n154) );
  XOR2_X1 U190 ( .A(n155), .B(n154), .Z(n156) );
  OR2_X1 U191 ( .A1(n157), .A2(n156), .ZN(n159) );
  NAND2_X1 U192 ( .A1(n157), .A2(n156), .ZN(n158) );
  NAND2_X1 U193 ( .A1(n159), .A2(n158), .ZN(n160) );
  MUX2_X1 U194 ( .A(n328), .B(n160), .S(n192), .Z(n352) );
  NAND2_X1 U195 ( .A1(n162), .A2(n161), .ZN(n163) );
  MUX2_X1 U196 ( .A(n329), .B(n163), .S(n192), .Z(n354) );
  NOR2_X1 U197 ( .A1(n165), .A2(n164), .ZN(n166) );
  MUX2_X1 U198 ( .A(n330), .B(n166), .S(n192), .Z(n356) );
  XNOR2_X1 U199 ( .A(n26), .B(n169), .ZN(n181) );
  FA_X1 U200 ( .A(n172), .B(n171), .CI(n170), .CO(n48), .S(n185) );
  FA_X1 U201 ( .A(n175), .B(n174), .CI(n173), .CO(n184), .S(n186) );
  FA_X1 U202 ( .A(n178), .B(n177), .CI(n176), .CO(n168), .S(n183) );
  NOR2_X1 U203 ( .A1(n181), .A2(n180), .ZN(n179) );
  MUX2_X1 U204 ( .A(n332), .B(n179), .S(n192), .Z(n360) );
  NAND2_X1 U205 ( .A1(n181), .A2(n180), .ZN(n182) );
  MUX2_X1 U206 ( .A(n333), .B(n182), .S(n192), .Z(n362) );
  FA_X1 U207 ( .A(n185), .B(n184), .CI(n183), .CO(n180), .S(n191) );
  FA_X1 U208 ( .A(n188), .B(n187), .CI(n186), .CO(n190), .S(n195) );
  NOR2_X1 U209 ( .A1(n191), .A2(n190), .ZN(n189) );
  MUX2_X1 U210 ( .A(n334), .B(n189), .S(n192), .Z(n364) );
  NAND2_X1 U211 ( .A1(n191), .A2(n190), .ZN(n193) );
  MUX2_X1 U212 ( .A(n335), .B(n193), .S(n192), .Z(n366) );
  NAND2_X1 U213 ( .A1(n195), .A2(n194), .ZN(n196) );
  MUX2_X1 U214 ( .A(n336), .B(n196), .S(n248), .Z(n368) );
  FA_X1 U215 ( .A(n199), .B(n198), .CI(n197), .CO(n194), .S(n207) );
  XNOR2_X1 U216 ( .A(n543), .B(\mult_x_1/n286 ), .ZN(n220) );
  OAI22_X1 U217 ( .A1(n201), .A2(n220), .B1(n11), .B2(n200), .ZN(n217) );
  XNOR2_X1 U218 ( .A(n235), .B(\mult_x_1/n284 ), .ZN(n218) );
  OAI22_X1 U219 ( .A1(n236), .A2(n218), .B1(n202), .B2(n5), .ZN(n216) );
  HA_X1 U220 ( .A(n204), .B(n203), .CO(n199), .S(n215) );
  NOR2_X1 U221 ( .A1(n207), .A2(n206), .ZN(n205) );
  MUX2_X1 U222 ( .A(n337), .B(n205), .S(n248), .Z(n370) );
  NAND2_X1 U223 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U224 ( .A(n338), .B(n208), .S(n248), .Z(n372) );
  NAND2_X1 U225 ( .A1(n210), .A2(n209), .ZN(n211) );
  MUX2_X1 U226 ( .A(n339), .B(n211), .S(n248), .Z(n374) );
  NAND2_X1 U227 ( .A1(n213), .A2(n212), .ZN(n214) );
  MUX2_X1 U228 ( .A(n342), .B(n214), .S(n248), .Z(n380) );
  FA_X1 U229 ( .A(n217), .B(n216), .CI(n215), .CO(n206), .S(n246) );
  XNOR2_X1 U230 ( .A(n235), .B(\mult_x_1/n285 ), .ZN(n226) );
  OAI22_X1 U231 ( .A1(n236), .A2(n226), .B1(n218), .B2(n5), .ZN(n223) );
  INV_X1 U232 ( .A(n9), .ZN(n219) );
  AND2_X1 U233 ( .A1(\mult_x_1/n288 ), .A2(n219), .ZN(n222) );
  XNOR2_X1 U234 ( .A(n543), .B(\mult_x_1/n287 ), .ZN(n224) );
  OAI22_X1 U235 ( .A1(n231), .A2(n224), .B1(n11), .B2(n220), .ZN(n221) );
  OR2_X1 U236 ( .A1(n246), .A2(n245), .ZN(n273) );
  FA_X1 U237 ( .A(n223), .B(n222), .CI(n221), .CO(n245), .S(n244) );
  XNOR2_X1 U238 ( .A(n543), .B(\mult_x_1/n288 ), .ZN(n225) );
  OAI22_X1 U239 ( .A1(n231), .A2(n225), .B1(n11), .B2(n224), .ZN(n228) );
  XNOR2_X1 U240 ( .A(n235), .B(\mult_x_1/n286 ), .ZN(n232) );
  OAI22_X1 U241 ( .A1(n236), .A2(n232), .B1(n226), .B2(n5), .ZN(n227) );
  NOR2_X1 U242 ( .A1(n244), .A2(n243), .ZN(n266) );
  HA_X1 U243 ( .A(n228), .B(n227), .CO(n243), .S(n241) );
  INV_X1 U244 ( .A(n543), .ZN(n230) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n230), .ZN(n229) );
  OAI22_X1 U246 ( .A1(n231), .A2(n230), .B1(n229), .B2(n11), .ZN(n240) );
  OR2_X1 U247 ( .A1(n241), .A2(n240), .ZN(n262) );
  XNOR2_X1 U248 ( .A(n235), .B(\mult_x_1/n287 ), .ZN(n234) );
  OAI22_X1 U249 ( .A1(n236), .A2(n234), .B1(n232), .B2(n5), .ZN(n239) );
  INV_X1 U250 ( .A(n11), .ZN(n233) );
  AND2_X1 U251 ( .A1(\mult_x_1/n288 ), .A2(n233), .ZN(n238) );
  NOR2_X1 U252 ( .A1(n239), .A2(n238), .ZN(n255) );
  OAI22_X1 U253 ( .A1(n236), .A2(\mult_x_1/n288 ), .B1(n234), .B2(n5), .ZN(
        n252) );
  OR2_X1 U254 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n237) );
  NAND2_X1 U255 ( .A1(n237), .A2(n236), .ZN(n251) );
  NAND2_X1 U256 ( .A1(n252), .A2(n251), .ZN(n258) );
  NAND2_X1 U257 ( .A1(n239), .A2(n238), .ZN(n256) );
  OAI21_X1 U258 ( .B1(n255), .B2(n258), .A(n256), .ZN(n263) );
  NAND2_X1 U259 ( .A1(n241), .A2(n240), .ZN(n261) );
  INV_X1 U260 ( .A(n261), .ZN(n242) );
  AOI21_X1 U261 ( .B1(n262), .B2(n263), .A(n242), .ZN(n269) );
  NAND2_X1 U262 ( .A1(n244), .A2(n243), .ZN(n267) );
  OAI21_X1 U263 ( .B1(n266), .B2(n269), .A(n267), .ZN(n274) );
  NAND2_X1 U264 ( .A1(n246), .A2(n245), .ZN(n272) );
  INV_X1 U265 ( .A(n272), .ZN(n247) );
  AOI21_X1 U266 ( .B1(n273), .B2(n274), .A(n247), .ZN(n249) );
  MUX2_X1 U267 ( .A(n343), .B(n249), .S(n248), .Z(n382) );
  MUX2_X1 U268 ( .A(product[0]), .B(n506), .S(n320), .Z(n396) );
  MUX2_X1 U269 ( .A(n506), .B(n507), .S(n320), .Z(n398) );
  AND2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n250) );
  MUX2_X1 U271 ( .A(n507), .B(n250), .S(n320), .Z(n400) );
  MUX2_X1 U272 ( .A(product[1]), .B(n509), .S(n320), .Z(n402) );
  MUX2_X1 U273 ( .A(n509), .B(n510), .S(n320), .Z(n404) );
  OR2_X1 U274 ( .A1(n252), .A2(n251), .ZN(n253) );
  AND2_X1 U275 ( .A1(n253), .A2(n258), .ZN(n254) );
  MUX2_X1 U276 ( .A(n510), .B(n254), .S(n320), .Z(n406) );
  MUX2_X1 U277 ( .A(product[2]), .B(n512), .S(n320), .Z(n408) );
  MUX2_X1 U278 ( .A(n512), .B(n513), .S(n320), .Z(n410) );
  INV_X1 U279 ( .A(n255), .ZN(n257) );
  NAND2_X1 U280 ( .A1(n257), .A2(n256), .ZN(n259) );
  XOR2_X1 U281 ( .A(n259), .B(n258), .Z(n260) );
  MUX2_X1 U282 ( .A(n513), .B(n260), .S(n320), .Z(n412) );
  MUX2_X1 U283 ( .A(product[3]), .B(n515), .S(n320), .Z(n414) );
  MUX2_X1 U284 ( .A(n515), .B(n516), .S(n192), .Z(n416) );
  NAND2_X1 U285 ( .A1(n262), .A2(n261), .ZN(n264) );
  XNOR2_X1 U286 ( .A(n264), .B(n263), .ZN(n265) );
  MUX2_X1 U287 ( .A(n516), .B(n265), .S(n320), .Z(n418) );
  MUX2_X1 U288 ( .A(product[4]), .B(n518), .S(n320), .Z(n420) );
  MUX2_X1 U289 ( .A(n518), .B(n519), .S(n192), .Z(n422) );
  INV_X1 U290 ( .A(n266), .ZN(n268) );
  NAND2_X1 U291 ( .A1(n268), .A2(n267), .ZN(n270) );
  XOR2_X1 U292 ( .A(n270), .B(n269), .Z(n271) );
  MUX2_X1 U293 ( .A(n519), .B(n271), .S(n320), .Z(n424) );
  MUX2_X1 U294 ( .A(product[5]), .B(n521), .S(n320), .Z(n426) );
  MUX2_X1 U295 ( .A(n521), .B(n522), .S(n320), .Z(n428) );
  NAND2_X1 U296 ( .A1(n273), .A2(n272), .ZN(n275) );
  XNOR2_X1 U297 ( .A(n275), .B(n274), .ZN(n276) );
  MUX2_X1 U298 ( .A(n522), .B(n276), .S(n192), .Z(n430) );
  MUX2_X1 U299 ( .A(product[6]), .B(n524), .S(n320), .Z(n432) );
  NAND2_X1 U300 ( .A1(n387), .A2(n338), .ZN(n277) );
  XOR2_X1 U301 ( .A(n277), .B(n343), .Z(n278) );
  MUX2_X1 U302 ( .A(n524), .B(n278), .S(n248), .Z(n434) );
  MUX2_X1 U303 ( .A(product[7]), .B(n526), .S(n320), .Z(n436) );
  OAI21_X1 U304 ( .B1(n337), .B2(n343), .A(n338), .ZN(n281) );
  NAND2_X1 U305 ( .A1(n326), .A2(n336), .ZN(n279) );
  XNOR2_X1 U306 ( .A(n281), .B(n279), .ZN(n280) );
  MUX2_X1 U307 ( .A(n526), .B(n280), .S(en), .Z(n438) );
  BUF_X4 U308 ( .A(en), .Z(n320) );
  MUX2_X1 U309 ( .A(product[8]), .B(n528), .S(n320), .Z(n440) );
  AOI21_X1 U310 ( .B1(n281), .B2(n326), .A(n388), .ZN(n284) );
  NAND2_X1 U311 ( .A1(n389), .A2(n335), .ZN(n282) );
  XOR2_X1 U312 ( .A(n284), .B(n282), .Z(n283) );
  MUX2_X1 U313 ( .A(n528), .B(n283), .S(n320), .Z(n442) );
  MUX2_X1 U314 ( .A(product[9]), .B(n530), .S(n320), .Z(n444) );
  OAI21_X1 U315 ( .B1(n284), .B2(n334), .A(n335), .ZN(n292) );
  INV_X1 U316 ( .A(n292), .ZN(n287) );
  NAND2_X1 U317 ( .A1(n390), .A2(n333), .ZN(n285) );
  XOR2_X1 U318 ( .A(n287), .B(n285), .Z(n286) );
  MUX2_X1 U319 ( .A(n530), .B(n286), .S(n320), .Z(n446) );
  MUX2_X1 U320 ( .A(product[10]), .B(n532), .S(n320), .Z(n448) );
  OAI21_X1 U321 ( .B1(n287), .B2(n332), .A(n333), .ZN(n289) );
  NAND2_X1 U322 ( .A1(n323), .A2(n341), .ZN(n288) );
  XNOR2_X1 U323 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U324 ( .A(n532), .B(n290), .S(n320), .Z(n450) );
  MUX2_X1 U325 ( .A(product[11]), .B(n534), .S(n320), .Z(n452) );
  NOR2_X1 U326 ( .A1(n340), .A2(n332), .ZN(n293) );
  OAI21_X1 U327 ( .B1(n340), .B2(n333), .A(n341), .ZN(n291) );
  AOI21_X1 U328 ( .B1(n293), .B2(n292), .A(n291), .ZN(n315) );
  NAND2_X1 U329 ( .A1(n391), .A2(n331), .ZN(n294) );
  XOR2_X1 U330 ( .A(n315), .B(n294), .Z(n295) );
  MUX2_X1 U331 ( .A(n534), .B(n295), .S(n320), .Z(n454) );
  MUX2_X1 U332 ( .A(product[12]), .B(n536), .S(n320), .Z(n456) );
  OAI21_X1 U333 ( .B1(n315), .B2(n330), .A(n331), .ZN(n297) );
  NAND2_X1 U334 ( .A1(n325), .A2(n339), .ZN(n296) );
  XNOR2_X1 U335 ( .A(n297), .B(n296), .ZN(n298) );
  MUX2_X1 U336 ( .A(n536), .B(n298), .S(n320), .Z(n458) );
  MUX2_X1 U337 ( .A(product[13]), .B(n538), .S(n320), .Z(n460) );
  NAND2_X1 U338 ( .A1(n391), .A2(n325), .ZN(n300) );
  AOI21_X1 U339 ( .B1(n386), .B2(n325), .A(n392), .ZN(n299) );
  OAI21_X1 U340 ( .B1(n315), .B2(n300), .A(n299), .ZN(n302) );
  NAND2_X1 U341 ( .A1(n327), .A2(n342), .ZN(n301) );
  XNOR2_X1 U342 ( .A(n302), .B(n301), .ZN(n303) );
  MUX2_X1 U343 ( .A(n538), .B(n303), .S(n320), .Z(n462) );
  MUX2_X1 U344 ( .A(product[14]), .B(n540), .S(n320), .Z(n464) );
  NAND2_X1 U345 ( .A1(n325), .A2(n327), .ZN(n305) );
  NOR2_X1 U346 ( .A1(n330), .A2(n305), .ZN(n311) );
  INV_X1 U347 ( .A(n311), .ZN(n307) );
  AOI21_X1 U348 ( .B1(n392), .B2(n327), .A(n384), .ZN(n304) );
  OAI21_X1 U349 ( .B1(n305), .B2(n331), .A(n304), .ZN(n312) );
  INV_X1 U350 ( .A(n312), .ZN(n306) );
  OAI21_X1 U351 ( .B1(n315), .B2(n307), .A(n306), .ZN(n309) );
  NAND2_X1 U352 ( .A1(n324), .A2(n329), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U354 ( .A(n540), .B(n310), .S(n320), .Z(n466) );
  MUX2_X1 U355 ( .A(product[15]), .B(n542), .S(n320), .Z(n468) );
  NAND2_X1 U356 ( .A1(n311), .A2(n324), .ZN(n314) );
  AOI21_X1 U357 ( .B1(n312), .B2(n324), .A(n385), .ZN(n313) );
  OAI21_X1 U358 ( .B1(n315), .B2(n314), .A(n313), .ZN(n316) );
  XNOR2_X1 U359 ( .A(n316), .B(n328), .ZN(n317) );
  MUX2_X1 U360 ( .A(n542), .B(n317), .S(n320), .Z(n470) );
  MUX2_X1 U361 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n320), .Z(n472) );
  MUX2_X1 U362 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n320), .Z(n474) );
  MUX2_X1 U363 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n320), .Z(n476) );
  MUX2_X1 U364 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n320), .Z(n478) );
  MUX2_X1 U365 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n320), .Z(n480) );
  MUX2_X1 U366 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n320), .Z(n482) );
  MUX2_X1 U367 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n320), .Z(n484) );
  MUX2_X1 U368 ( .A(n8), .B(B_extended[7]), .S(n320), .Z(n486) );
  MUX2_X1 U369 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n320), .Z(n488) );
  MUX2_X1 U370 ( .A(n235), .B(A_extended[1]), .S(n320), .Z(n490) );
  MUX2_X1 U371 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n320), .Z(n492) );
  MUX2_X1 U372 ( .A(n543), .B(A_extended[3]), .S(n320), .Z(n494) );
  MUX2_X1 U373 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n320), .Z(n496) );
  MUX2_X1 U374 ( .A(n319), .B(A_extended[5]), .S(n320), .Z(n498) );
  MUX2_X1 U375 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n320), .Z(n500) );
  MUX2_X1 U376 ( .A(\mult_x_1/n310 ), .B(A_extended[7]), .S(n320), .Z(n502) );
  OR2_X1 U377 ( .A1(n320), .A2(n545), .ZN(n504) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_24 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n311 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n351, n353,
         n355, n357, n359, n361, n363, n365, n367, n369, n371, n373, n375,
         n377, n379, n381, n383, n385, n387, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n420, n422, n424, n426, n428,
         n430, n432, n434, n436, n438, n440, n442, n444, n446, n448, n450,
         n452, n454, n456, n458, n460, n462, n464, n466, n468, n470, n472,
         n474, n476, n478, n480, n482, n484, n486, n488, n490, n492, n494,
         n496, n498, n500, n502, n504, n506, n508, n510, n512, n514, n515,
         n517, n518, n520, n521, n523, n524, n526, n527, n529, n530, n532,
         n534, n536, n538, n540, n542, n544, n546, n548, n550, n551, n552,
         n553, n554;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n402), .SE(n512), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n402), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n402), .SE(n504), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n28) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n402), .SE(n500), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n17) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n402), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n22) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n402), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n401), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n27) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n401), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n401), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n24) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n401), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n23) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n401), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n30) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n401), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n19) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n401), .SE(n478), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n401), .SE(n476), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n401), .SE(n474), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n401), .SE(n472), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n401), .SE(n470), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n400), .SE(n468), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n400), .SE(n466), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n400), .SE(n464), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n400), .SE(n462), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n400), .SE(n460), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n400), .SE(n458), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n400), .SE(n456), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n400), .SE(n454), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n400), .SE(n452), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n400), .SE(n450), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n400), .SE(n448), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n399), .SE(n446), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n399), .SE(n444), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n399), .SE(n442), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n399), .SE(n440), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n399), .SE(n438), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n399), .SE(n436), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n399), .SE(n434), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n399), .SE(n432), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n399), .SE(n430), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n399), .SE(n428), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n399), .SE(n426), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n398), .SE(n424), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n398), .SE(n422), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n398), .SE(n420), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n398), .SE(n418), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n398), .SE(n416), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n398), .SE(n414), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n398), .SE(n412), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n398), .SE(n410), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n398), .SE(n408), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n398), .SE(n406), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n398), .SE(n404), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n402), .SE(n502), .CK(clk), .Q(n551), 
        .QN(n29) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n402), .SE(n510), .CK(clk), .Q(n552), 
        .QN(n21) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n402), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n31) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n554), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n554), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n554), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n554), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n345), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n554), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n344), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n554), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n554), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n342), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n554), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n341), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n554), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n554), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n339), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n554), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n554), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n337), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n554), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n336), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n554), .SE(n361), .CK(
        clk), .Q(n395), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n554), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n334), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n554), .SE(n357), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n554), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n554), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n554), .SE(n351), .CK(
        clk), .QN(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n554), .SI(1'b1), .SE(n349), .CK(clk), 
        .Q(n329) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n402), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n328) );
  SDFF_X2 clk_r_REG62_S1 ( .D(1'b0), .SI(n402), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n18) );
  AND2_X1 U2 ( .A1(n553), .A2(\mult_x_1/n281 ), .ZN(n70) );
  NOR2_X1 U3 ( .A1(n141), .A2(n142), .ZN(n43) );
  NAND2_X1 U4 ( .A1(n6), .A2(n5), .ZN(n142) );
  NAND2_X1 U5 ( .A1(n227), .A2(n18), .ZN(n5) );
  INV_X1 U6 ( .A(n12), .ZN(n6) );
  CLKBUF_X2 U7 ( .A(n45), .Z(n222) );
  CLKBUF_X1 U8 ( .A(n250), .Z(n398) );
  CLKBUF_X1 U9 ( .A(n250), .Z(n402) );
  CLKBUF_X1 U10 ( .A(n250), .Z(n401) );
  CLKBUF_X1 U11 ( .A(n250), .Z(n400) );
  CLKBUF_X1 U12 ( .A(n250), .Z(n399) );
  OR2_X1 U13 ( .A1(n59), .A2(n58), .ZN(n65) );
  INV_X1 U14 ( .A(rst_n), .ZN(n554) );
  INV_X1 U15 ( .A(n33), .ZN(n211) );
  INV_X1 U16 ( .A(n31), .ZN(n7) );
  AND2_X1 U17 ( .A1(n552), .A2(n553), .ZN(n37) );
  CLKBUF_X1 U18 ( .A(n104), .Z(n16) );
  CLKBUF_X1 U19 ( .A(en), .Z(n251) );
  XNOR2_X1 U20 ( .A(n171), .B(n170), .ZN(n176) );
  XNOR2_X1 U21 ( .A(n169), .B(n168), .ZN(n170) );
  NAND2_X1 U22 ( .A1(n109), .A2(n108), .ZN(n110) );
  INV_X1 U23 ( .A(n554), .ZN(n250) );
  XOR2_X1 U24 ( .A(n37), .B(n21), .Z(n57) );
  XOR2_X1 U25 ( .A(n61), .B(n60), .Z(n8) );
  XOR2_X1 U26 ( .A(n62), .B(n8), .Z(n241) );
  NAND2_X1 U27 ( .A1(n62), .A2(n61), .ZN(n9) );
  NAND2_X1 U28 ( .A1(n62), .A2(n60), .ZN(n10) );
  NAND2_X1 U29 ( .A1(n61), .A2(n60), .ZN(n11) );
  NAND3_X1 U30 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n106) );
  XNOR2_X1 U31 ( .A(n70), .B(\mult_x_1/n313 ), .ZN(n12) );
  INV_X1 U32 ( .A(n22), .ZN(n13) );
  NAND2_X2 U33 ( .A1(n18), .A2(n7), .ZN(n227) );
  INV_X1 U34 ( .A(\mult_x_1/n313 ), .ZN(n14) );
  INV_X1 U35 ( .A(n36), .ZN(n15) );
  INV_X1 U36 ( .A(n36), .ZN(n224) );
  XNOR2_X1 U37 ( .A(n31), .B(n17), .ZN(n35) );
  AND2_X1 U38 ( .A1(n160), .A2(n158), .ZN(n20) );
  BUF_X2 U39 ( .A(n551), .Z(n324) );
  XNOR2_X1 U40 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .ZN(n32) );
  XNOR2_X1 U41 ( .A(n551), .B(n28), .ZN(n33) );
  OR2_X2 U42 ( .A1(n32), .A2(n33), .ZN(n152) );
  INV_X2 U43 ( .A(n328), .ZN(n325) );
  XNOR2_X1 U44 ( .A(n325), .B(\mult_x_1/n284 ), .ZN(n150) );
  XNOR2_X1 U45 ( .A(n325), .B(\mult_x_1/n283 ), .ZN(n49) );
  OAI22_X1 U46 ( .A1(n152), .A2(n150), .B1(n211), .B2(n49), .ZN(n59) );
  XOR2_X1 U47 ( .A(\mult_x_1/a[2] ), .B(n551), .Z(n34) );
  NAND2_X1 U48 ( .A1(n34), .A2(n35), .ZN(n45) );
  XNOR2_X1 U49 ( .A(n324), .B(\mult_x_1/n282 ), .ZN(n148) );
  INV_X1 U50 ( .A(n35), .ZN(n36) );
  XNOR2_X1 U51 ( .A(n324), .B(\mult_x_1/n281 ), .ZN(n44) );
  OAI22_X1 U52 ( .A1(n45), .A2(n148), .B1(n224), .B2(n44), .ZN(n58) );
  CLKBUF_X2 U53 ( .A(n552), .Z(n326) );
  NOR2_X1 U54 ( .A1(n23), .A2(n57), .ZN(n64) );
  XOR2_X1 U55 ( .A(\mult_x_1/a[6] ), .B(n552), .Z(n38) );
  XNOR2_X1 U56 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n39) );
  NAND2_X1 U57 ( .A1(n38), .A2(n39), .ZN(n85) );
  XNOR2_X1 U58 ( .A(n326), .B(\mult_x_1/n286 ), .ZN(n53) );
  INV_X1 U59 ( .A(n39), .ZN(n40) );
  INV_X2 U60 ( .A(n40), .ZN(n124) );
  XNOR2_X1 U61 ( .A(n326), .B(\mult_x_1/n285 ), .ZN(n51) );
  OAI22_X1 U62 ( .A1(n85), .A2(n53), .B1(n124), .B2(n51), .ZN(n141) );
  XNOR2_X1 U63 ( .A(n70), .B(\mult_x_1/n313 ), .ZN(n56) );
  OR2_X1 U64 ( .A1(n57), .A2(n30), .ZN(n143) );
  NAND2_X1 U65 ( .A1(n141), .A2(n142), .ZN(n42) );
  OAI21_X1 U66 ( .B1(n43), .B2(n143), .A(n42), .ZN(n63) );
  XNOR2_X1 U67 ( .A(n326), .B(\mult_x_1/n284 ), .ZN(n50) );
  XNOR2_X1 U68 ( .A(n326), .B(\mult_x_1/n283 ), .ZN(n73) );
  OAI22_X1 U69 ( .A1(n85), .A2(n50), .B1(n124), .B2(n73), .ZN(n105) );
  XNOR2_X1 U70 ( .A(n70), .B(n324), .ZN(n46) );
  OAI22_X1 U71 ( .A1(n46), .A2(n224), .B1(n45), .B2(n44), .ZN(n104) );
  AOI21_X1 U72 ( .B1(n15), .B2(n222), .A(n46), .ZN(n47) );
  INV_X1 U73 ( .A(n47), .ZN(n103) );
  NOR2_X1 U74 ( .A1(n24), .A2(n57), .ZN(n109) );
  XNOR2_X1 U75 ( .A(n325), .B(\mult_x_1/n282 ), .ZN(n48) );
  XNOR2_X1 U76 ( .A(n325), .B(\mult_x_1/n281 ), .ZN(n75) );
  OAI22_X1 U77 ( .A1(n152), .A2(n48), .B1(n211), .B2(n75), .ZN(n108) );
  XNOR2_X1 U78 ( .A(n109), .B(n108), .ZN(n52) );
  INV_X1 U79 ( .A(n104), .ZN(n62) );
  OAI22_X1 U80 ( .A1(n152), .A2(n49), .B1(n211), .B2(n48), .ZN(n61) );
  OAI22_X1 U81 ( .A1(n85), .A2(n51), .B1(n124), .B2(n50), .ZN(n60) );
  XNOR2_X1 U82 ( .A(n52), .B(n106), .ZN(n116) );
  XNOR2_X1 U83 ( .A(n326), .B(\mult_x_1/n287 ), .ZN(n83) );
  OR2_X1 U84 ( .A1(n85), .A2(n83), .ZN(n55) );
  OR2_X1 U85 ( .A1(n124), .A2(n53), .ZN(n54) );
  NAND2_X1 U86 ( .A1(n55), .A2(n54), .ZN(n164) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n313 ), .B(n13), .ZN(n86) );
  OAI22_X1 U88 ( .A1(n227), .A2(n86), .B1(n56), .B2(n18), .ZN(n163) );
  NOR2_X1 U89 ( .A1(n57), .A2(n19), .ZN(n162) );
  XNOR2_X1 U90 ( .A(n59), .B(n58), .ZN(n158) );
  FA_X1 U91 ( .A(n65), .B(n64), .CI(n63), .CO(n118), .S(n240) );
  NAND2_X1 U92 ( .A1(n139), .A2(n138), .ZN(n66) );
  BUF_X2 U93 ( .A(n251), .Z(n185) );
  NAND2_X1 U94 ( .A1(n66), .A2(n185), .ZN(n68) );
  OR2_X1 U95 ( .A1(n185), .A2(n391), .ZN(n67) );
  NAND2_X1 U96 ( .A1(n68), .A2(n67), .ZN(n363) );
  NOR2_X1 U117 ( .A1(n25), .A2(n57), .ZN(n122) );
  XNOR2_X1 U118 ( .A(n326), .B(\mult_x_1/n281 ), .ZN(n69) );
  XNOR2_X1 U119 ( .A(n70), .B(n326), .ZN(n123) );
  OAI22_X1 U120 ( .A1(n85), .A2(n69), .B1(n123), .B2(n124), .ZN(n129) );
  INV_X1 U121 ( .A(n129), .ZN(n121) );
  XNOR2_X1 U122 ( .A(n326), .B(\mult_x_1/n282 ), .ZN(n72) );
  OAI22_X1 U123 ( .A1(n85), .A2(n72), .B1(n124), .B2(n69), .ZN(n79) );
  XNOR2_X1 U124 ( .A(n70), .B(\mult_x_1/n311 ), .ZN(n74) );
  AOI21_X1 U125 ( .B1(n211), .B2(n152), .A(n74), .ZN(n71) );
  INV_X1 U126 ( .A(n71), .ZN(n78) );
  OAI22_X1 U127 ( .A1(n152), .A2(n75), .B1(n74), .B2(n211), .ZN(n77) );
  NOR2_X1 U128 ( .A1(n26), .A2(n57), .ZN(n102) );
  OAI22_X1 U129 ( .A1(n85), .A2(n73), .B1(n124), .B2(n72), .ZN(n101) );
  OAI22_X1 U130 ( .A1(n152), .A2(n75), .B1(n74), .B2(n211), .ZN(n76) );
  INV_X1 U131 ( .A(n76), .ZN(n100) );
  NOR2_X1 U132 ( .A1(n27), .A2(n57), .ZN(n98) );
  FA_X1 U133 ( .A(n79), .B(n78), .CI(n77), .CO(n120), .S(n97) );
  OR2_X1 U134 ( .A1(n136), .A2(n135), .ZN(n80) );
  MUX2_X1 U135 ( .A(n329), .B(n80), .S(n185), .Z(n349) );
  XNOR2_X1 U136 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n194) );
  XNOR2_X1 U137 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n87) );
  OAI22_X1 U138 ( .A1(n227), .A2(n194), .B1(n87), .B2(n18), .ZN(n95) );
  INV_X1 U139 ( .A(n124), .ZN(n81) );
  AND2_X1 U140 ( .A1(\mult_x_1/n288 ), .A2(n81), .ZN(n94) );
  XNOR2_X1 U141 ( .A(n324), .B(\mult_x_1/n285 ), .ZN(n193) );
  XNOR2_X1 U142 ( .A(n324), .B(\mult_x_1/n284 ), .ZN(n88) );
  OAI22_X1 U143 ( .A1(n222), .A2(n193), .B1(n15), .B2(n88), .ZN(n93) );
  OR2_X1 U144 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n82) );
  OAI22_X1 U145 ( .A1(n85), .A2(n21), .B1(n82), .B2(n124), .ZN(n147) );
  XNOR2_X1 U146 ( .A(n326), .B(\mult_x_1/n288 ), .ZN(n84) );
  OAI22_X1 U147 ( .A1(n85), .A2(n84), .B1(n124), .B2(n83), .ZN(n146) );
  XNOR2_X1 U148 ( .A(n325), .B(\mult_x_1/n286 ), .ZN(n91) );
  XNOR2_X1 U149 ( .A(n325), .B(\mult_x_1/n285 ), .ZN(n151) );
  OAI22_X1 U150 ( .A1(n152), .A2(n91), .B1(n211), .B2(n151), .ZN(n167) );
  OAI22_X1 U151 ( .A1(n227), .A2(n87), .B1(n86), .B2(n18), .ZN(n166) );
  XNOR2_X1 U152 ( .A(n324), .B(\mult_x_1/n283 ), .ZN(n149) );
  OAI22_X1 U153 ( .A1(n222), .A2(n88), .B1(n15), .B2(n149), .ZN(n165) );
  OR2_X1 U154 ( .A1(\mult_x_1/n288 ), .A2(n328), .ZN(n89) );
  OAI22_X1 U155 ( .A1(n152), .A2(n328), .B1(n89), .B2(n211), .ZN(n196) );
  XNOR2_X1 U156 ( .A(n325), .B(\mult_x_1/n288 ), .ZN(n90) );
  XNOR2_X1 U157 ( .A(n325), .B(\mult_x_1/n287 ), .ZN(n92) );
  OAI22_X1 U158 ( .A1(n152), .A2(n90), .B1(n211), .B2(n92), .ZN(n195) );
  OAI22_X1 U159 ( .A1(n152), .A2(n92), .B1(n211), .B2(n91), .ZN(n191) );
  FA_X1 U160 ( .A(n95), .B(n94), .CI(n93), .CO(n181), .S(n190) );
  OR2_X1 U161 ( .A1(n188), .A2(n187), .ZN(n96) );
  MUX2_X1 U162 ( .A(n330), .B(n96), .S(n185), .Z(n351) );
  FA_X1 U163 ( .A(n99), .B(n98), .CI(n97), .CO(n135), .S(n202) );
  FA_X1 U164 ( .A(n102), .B(n101), .CI(n100), .CO(n99), .S(n115) );
  FA_X1 U165 ( .A(n105), .B(n16), .CI(n103), .CO(n114), .S(n117) );
  OR2_X1 U166 ( .A1(n108), .A2(n109), .ZN(n107) );
  NAND2_X1 U167 ( .A1(n107), .A2(n106), .ZN(n111) );
  NAND2_X1 U168 ( .A1(n111), .A2(n110), .ZN(n113) );
  OR2_X1 U169 ( .A1(n202), .A2(n201), .ZN(n112) );
  MUX2_X1 U170 ( .A(n331), .B(n112), .S(n185), .Z(n353) );
  FA_X1 U171 ( .A(n115), .B(n114), .CI(n113), .CO(n201), .S(n205) );
  FA_X1 U172 ( .A(n118), .B(n117), .CI(n116), .CO(n204), .S(n139) );
  OR2_X1 U173 ( .A1(n205), .A2(n204), .ZN(n119) );
  MUX2_X1 U174 ( .A(n332), .B(n119), .S(n185), .Z(n355) );
  FA_X1 U175 ( .A(n122), .B(n121), .CI(n120), .CO(n131), .S(n136) );
  AOI21_X1 U176 ( .B1(n124), .B2(n85), .A(n123), .ZN(n125) );
  INV_X1 U177 ( .A(n125), .ZN(n127) );
  NOR2_X1 U178 ( .A1(n22), .A2(n57), .ZN(n126) );
  XOR2_X1 U179 ( .A(n127), .B(n126), .Z(n128) );
  XOR2_X1 U180 ( .A(n129), .B(n128), .Z(n130) );
  OR2_X1 U181 ( .A1(n131), .A2(n130), .ZN(n133) );
  NAND2_X1 U182 ( .A1(n131), .A2(n130), .ZN(n132) );
  NAND2_X1 U183 ( .A1(n133), .A2(n132), .ZN(n134) );
  MUX2_X1 U184 ( .A(n333), .B(n134), .S(n185), .Z(n357) );
  NAND2_X1 U185 ( .A1(n136), .A2(n135), .ZN(n137) );
  MUX2_X1 U186 ( .A(n334), .B(n137), .S(n185), .Z(n359) );
  NOR2_X1 U187 ( .A1(n139), .A2(n138), .ZN(n140) );
  MUX2_X1 U188 ( .A(n335), .B(n140), .S(n185), .Z(n361) );
  INV_X1 U189 ( .A(n141), .ZN(n145) );
  XNOR2_X1 U190 ( .A(n143), .B(n142), .ZN(n144) );
  XNOR2_X1 U191 ( .A(n145), .B(n144), .ZN(n245) );
  HA_X1 U192 ( .A(n147), .B(n146), .CO(n171), .S(n180) );
  OAI22_X1 U193 ( .A1(n222), .A2(n149), .B1(n15), .B2(n148), .ZN(n169) );
  INV_X1 U194 ( .A(n169), .ZN(n154) );
  OAI22_X1 U195 ( .A1(n152), .A2(n151), .B1(n211), .B2(n150), .ZN(n168) );
  INV_X1 U196 ( .A(n168), .ZN(n153) );
  NAND2_X1 U197 ( .A1(n154), .A2(n153), .ZN(n155) );
  NAND2_X1 U198 ( .A1(n171), .A2(n155), .ZN(n157) );
  NAND2_X1 U199 ( .A1(n169), .A2(n168), .ZN(n156) );
  NAND2_X1 U200 ( .A1(n157), .A2(n156), .ZN(n244) );
  XNOR2_X1 U201 ( .A(n245), .B(n244), .ZN(n161) );
  INV_X1 U202 ( .A(n158), .ZN(n159) );
  XNOR2_X1 U203 ( .A(n160), .B(n159), .ZN(n243) );
  XNOR2_X1 U204 ( .A(n161), .B(n243), .ZN(n174) );
  FA_X1 U205 ( .A(n164), .B(n163), .CI(n162), .CO(n160), .S(n178) );
  FA_X1 U206 ( .A(n167), .B(n166), .CI(n165), .CO(n177), .S(n179) );
  NOR2_X1 U207 ( .A1(n174), .A2(n173), .ZN(n172) );
  MUX2_X1 U208 ( .A(n337), .B(n172), .S(n185), .Z(n365) );
  NAND2_X1 U209 ( .A1(n174), .A2(n173), .ZN(n175) );
  MUX2_X1 U210 ( .A(n338), .B(n175), .S(n185), .Z(n367) );
  FA_X1 U211 ( .A(n178), .B(n177), .CI(n176), .CO(n173), .S(n184) );
  FA_X1 U212 ( .A(n181), .B(n180), .CI(n179), .CO(n183), .S(n188) );
  NOR2_X1 U213 ( .A1(n184), .A2(n183), .ZN(n182) );
  MUX2_X1 U214 ( .A(n339), .B(n182), .S(n185), .Z(n369) );
  NAND2_X1 U215 ( .A1(n184), .A2(n183), .ZN(n186) );
  MUX2_X1 U216 ( .A(n340), .B(n186), .S(n185), .Z(n371) );
  NAND2_X1 U217 ( .A1(n188), .A2(n187), .ZN(n189) );
  MUX2_X1 U218 ( .A(n341), .B(n189), .S(n185), .Z(n373) );
  FA_X1 U219 ( .A(n192), .B(n191), .CI(n190), .CO(n187), .S(n199) );
  XNOR2_X1 U220 ( .A(n324), .B(\mult_x_1/n286 ), .ZN(n212) );
  OAI22_X1 U221 ( .A1(n222), .A2(n212), .B1(n224), .B2(n193), .ZN(n209) );
  XNOR2_X1 U222 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n210) );
  OAI22_X1 U223 ( .A1(n227), .A2(n210), .B1(n194), .B2(n18), .ZN(n208) );
  HA_X1 U224 ( .A(n196), .B(n195), .CO(n192), .S(n207) );
  NOR2_X1 U225 ( .A1(n199), .A2(n198), .ZN(n197) );
  MUX2_X1 U226 ( .A(n342), .B(n197), .S(n185), .Z(n375) );
  NAND2_X1 U227 ( .A1(n199), .A2(n198), .ZN(n200) );
  MUX2_X1 U228 ( .A(n343), .B(n200), .S(n185), .Z(n377) );
  NAND2_X1 U229 ( .A1(n202), .A2(n201), .ZN(n203) );
  MUX2_X1 U230 ( .A(n344), .B(n203), .S(n185), .Z(n379) );
  NAND2_X1 U231 ( .A1(n205), .A2(n204), .ZN(n206) );
  MUX2_X1 U232 ( .A(n345), .B(n206), .S(n282), .Z(n381) );
  FA_X1 U233 ( .A(n209), .B(n208), .CI(n207), .CO(n198), .S(n237) );
  XNOR2_X1 U234 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n218) );
  OAI22_X1 U235 ( .A1(n227), .A2(n218), .B1(n210), .B2(n18), .ZN(n215) );
  AND2_X1 U236 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n214) );
  XNOR2_X1 U237 ( .A(n324), .B(\mult_x_1/n287 ), .ZN(n216) );
  OAI22_X1 U238 ( .A1(n222), .A2(n216), .B1(n15), .B2(n212), .ZN(n213) );
  OR2_X1 U239 ( .A1(n237), .A2(n236), .ZN(n275) );
  FA_X1 U240 ( .A(n215), .B(n214), .CI(n213), .CO(n236), .S(n235) );
  XNOR2_X1 U241 ( .A(n324), .B(\mult_x_1/n288 ), .ZN(n217) );
  OAI22_X1 U242 ( .A1(n222), .A2(n217), .B1(n15), .B2(n216), .ZN(n220) );
  XNOR2_X1 U243 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n223) );
  OAI22_X1 U244 ( .A1(n227), .A2(n223), .B1(n218), .B2(n18), .ZN(n219) );
  NOR2_X1 U245 ( .A1(n235), .A2(n234), .ZN(n268) );
  HA_X1 U246 ( .A(n220), .B(n219), .CO(n234), .S(n232) );
  OR2_X1 U247 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n221) );
  OAI22_X1 U248 ( .A1(n222), .A2(n29), .B1(n221), .B2(n15), .ZN(n231) );
  OR2_X1 U249 ( .A1(n232), .A2(n231), .ZN(n264) );
  XNOR2_X1 U250 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n226) );
  OAI22_X1 U251 ( .A1(n227), .A2(n226), .B1(n223), .B2(n18), .ZN(n230) );
  INV_X1 U252 ( .A(n15), .ZN(n225) );
  AND2_X1 U253 ( .A1(\mult_x_1/n288 ), .A2(n225), .ZN(n229) );
  NOR2_X1 U254 ( .A1(n230), .A2(n229), .ZN(n257) );
  OAI22_X1 U255 ( .A1(n227), .A2(\mult_x_1/n288 ), .B1(n226), .B2(n18), .ZN(
        n254) );
  OR2_X1 U256 ( .A1(\mult_x_1/n288 ), .A2(n14), .ZN(n228) );
  NAND2_X1 U257 ( .A1(n228), .A2(n227), .ZN(n253) );
  NAND2_X1 U258 ( .A1(n254), .A2(n253), .ZN(n260) );
  NAND2_X1 U259 ( .A1(n230), .A2(n229), .ZN(n258) );
  OAI21_X1 U260 ( .B1(n257), .B2(n260), .A(n258), .ZN(n265) );
  NAND2_X1 U261 ( .A1(n232), .A2(n231), .ZN(n263) );
  INV_X1 U262 ( .A(n263), .ZN(n233) );
  AOI21_X1 U263 ( .B1(n264), .B2(n265), .A(n233), .ZN(n271) );
  NAND2_X1 U264 ( .A1(n235), .A2(n234), .ZN(n269) );
  OAI21_X1 U265 ( .B1(n268), .B2(n271), .A(n269), .ZN(n276) );
  NAND2_X1 U266 ( .A1(n237), .A2(n236), .ZN(n274) );
  INV_X1 U267 ( .A(n274), .ZN(n238) );
  AOI21_X1 U268 ( .B1(n275), .B2(n276), .A(n238), .ZN(n239) );
  MUX2_X1 U269 ( .A(n346), .B(n239), .S(n282), .Z(n383) );
  FA_X1 U270 ( .A(n20), .B(n241), .CI(n240), .CO(n138), .S(n242) );
  MUX2_X1 U271 ( .A(n347), .B(n242), .S(n185), .Z(n385) );
  NAND2_X1 U272 ( .A1(n243), .A2(n245), .ZN(n248) );
  NAND2_X1 U273 ( .A1(n243), .A2(n244), .ZN(n247) );
  NAND2_X1 U274 ( .A1(n245), .A2(n244), .ZN(n246) );
  NAND3_X1 U275 ( .A1(n248), .A2(n247), .A3(n246), .ZN(n249) );
  MUX2_X1 U276 ( .A(n348), .B(n249), .S(n282), .Z(n387) );
  BUF_X4 U277 ( .A(n251), .Z(n282) );
  MUX2_X1 U278 ( .A(product[0]), .B(n514), .S(n282), .Z(n404) );
  MUX2_X1 U279 ( .A(n514), .B(n515), .S(n282), .Z(n406) );
  AND2_X1 U280 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n252) );
  MUX2_X1 U281 ( .A(n515), .B(n252), .S(n282), .Z(n408) );
  MUX2_X1 U282 ( .A(product[1]), .B(n517), .S(n282), .Z(n410) );
  MUX2_X1 U283 ( .A(n517), .B(n518), .S(n282), .Z(n412) );
  OR2_X1 U284 ( .A1(n254), .A2(n253), .ZN(n255) );
  AND2_X1 U285 ( .A1(n255), .A2(n260), .ZN(n256) );
  MUX2_X1 U286 ( .A(n518), .B(n256), .S(n282), .Z(n414) );
  MUX2_X1 U287 ( .A(product[2]), .B(n520), .S(n282), .Z(n416) );
  MUX2_X1 U288 ( .A(n520), .B(n521), .S(n282), .Z(n418) );
  INV_X1 U289 ( .A(n257), .ZN(n259) );
  NAND2_X1 U290 ( .A1(n259), .A2(n258), .ZN(n261) );
  XOR2_X1 U291 ( .A(n261), .B(n260), .Z(n262) );
  MUX2_X1 U292 ( .A(n521), .B(n262), .S(n282), .Z(n420) );
  MUX2_X1 U293 ( .A(product[3]), .B(n523), .S(n282), .Z(n422) );
  MUX2_X1 U294 ( .A(n523), .B(n524), .S(n282), .Z(n424) );
  NAND2_X1 U295 ( .A1(n264), .A2(n263), .ZN(n266) );
  XNOR2_X1 U296 ( .A(n266), .B(n265), .ZN(n267) );
  MUX2_X1 U297 ( .A(n524), .B(n267), .S(n282), .Z(n426) );
  MUX2_X1 U298 ( .A(product[4]), .B(n526), .S(n282), .Z(n428) );
  MUX2_X1 U299 ( .A(n526), .B(n527), .S(n282), .Z(n430) );
  INV_X1 U300 ( .A(n268), .ZN(n270) );
  NAND2_X1 U301 ( .A1(n270), .A2(n269), .ZN(n272) );
  XOR2_X1 U302 ( .A(n272), .B(n271), .Z(n273) );
  MUX2_X1 U303 ( .A(n527), .B(n273), .S(n282), .Z(n432) );
  MUX2_X1 U304 ( .A(product[5]), .B(n529), .S(n282), .Z(n434) );
  MUX2_X1 U305 ( .A(n529), .B(n530), .S(n282), .Z(n436) );
  NAND2_X1 U306 ( .A1(n275), .A2(n274), .ZN(n277) );
  XNOR2_X1 U307 ( .A(n277), .B(n276), .ZN(n278) );
  MUX2_X1 U308 ( .A(n530), .B(n278), .S(n282), .Z(n438) );
  MUX2_X1 U309 ( .A(product[6]), .B(n532), .S(n282), .Z(n440) );
  NAND2_X1 U310 ( .A1(n392), .A2(n343), .ZN(n279) );
  XOR2_X1 U311 ( .A(n279), .B(n346), .Z(n280) );
  MUX2_X1 U312 ( .A(n532), .B(n280), .S(n282), .Z(n442) );
  MUX2_X1 U313 ( .A(product[7]), .B(n534), .S(n282), .Z(n444) );
  OAI21_X1 U314 ( .B1(n342), .B2(n346), .A(n343), .ZN(n284) );
  NAND2_X1 U315 ( .A1(n330), .A2(n341), .ZN(n281) );
  XNOR2_X1 U316 ( .A(n284), .B(n281), .ZN(n283) );
  MUX2_X1 U317 ( .A(n534), .B(n283), .S(n282), .Z(n446) );
  BUF_X2 U318 ( .A(en), .Z(n327) );
  MUX2_X1 U319 ( .A(product[8]), .B(n536), .S(n327), .Z(n448) );
  AOI21_X1 U320 ( .B1(n284), .B2(n330), .A(n393), .ZN(n287) );
  NAND2_X1 U321 ( .A1(n394), .A2(n340), .ZN(n285) );
  XOR2_X1 U322 ( .A(n287), .B(n285), .Z(n286) );
  MUX2_X1 U323 ( .A(n536), .B(n286), .S(n327), .Z(n450) );
  MUX2_X1 U324 ( .A(product[9]), .B(n538), .S(n327), .Z(n452) );
  OAI21_X1 U325 ( .B1(n287), .B2(n339), .A(n340), .ZN(n298) );
  INV_X1 U326 ( .A(n298), .ZN(n290) );
  NAND2_X1 U327 ( .A1(n396), .A2(n338), .ZN(n288) );
  XOR2_X1 U328 ( .A(n290), .B(n288), .Z(n289) );
  MUX2_X1 U329 ( .A(n538), .B(n289), .S(n327), .Z(n454) );
  MUX2_X1 U330 ( .A(product[10]), .B(n540), .S(n327), .Z(n456) );
  OAI21_X1 U331 ( .B1(n290), .B2(n337), .A(n338), .ZN(n293) );
  NOR2_X1 U332 ( .A1(n347), .A2(n348), .ZN(n296) );
  INV_X1 U333 ( .A(n296), .ZN(n291) );
  NAND2_X1 U334 ( .A1(n347), .A2(n348), .ZN(n295) );
  NAND2_X1 U335 ( .A1(n291), .A2(n295), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  MUX2_X1 U337 ( .A(n540), .B(n294), .S(n327), .Z(n458) );
  MUX2_X1 U338 ( .A(product[11]), .B(n542), .S(n327), .Z(n460) );
  NOR2_X1 U339 ( .A1(n296), .A2(n337), .ZN(n299) );
  OAI21_X1 U340 ( .B1(n296), .B2(n338), .A(n295), .ZN(n297) );
  AOI21_X1 U341 ( .B1(n299), .B2(n298), .A(n297), .ZN(n321) );
  NAND2_X1 U342 ( .A1(n395), .A2(n336), .ZN(n300) );
  XOR2_X1 U343 ( .A(n321), .B(n300), .Z(n301) );
  MUX2_X1 U344 ( .A(n542), .B(n301), .S(n327), .Z(n462) );
  MUX2_X1 U345 ( .A(product[12]), .B(n544), .S(n327), .Z(n464) );
  OAI21_X1 U346 ( .B1(n321), .B2(n335), .A(n336), .ZN(n303) );
  NAND2_X1 U347 ( .A1(n332), .A2(n345), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U349 ( .A(n544), .B(n304), .S(n327), .Z(n466) );
  MUX2_X1 U350 ( .A(product[13]), .B(n546), .S(n327), .Z(n468) );
  NAND2_X1 U351 ( .A1(n395), .A2(n332), .ZN(n306) );
  AOI21_X1 U352 ( .B1(n391), .B2(n332), .A(n397), .ZN(n305) );
  OAI21_X1 U353 ( .B1(n321), .B2(n306), .A(n305), .ZN(n308) );
  NAND2_X1 U354 ( .A1(n331), .A2(n344), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U356 ( .A(n546), .B(n309), .S(n327), .Z(n470) );
  MUX2_X1 U357 ( .A(product[14]), .B(n548), .S(n327), .Z(n472) );
  NAND2_X1 U358 ( .A1(n332), .A2(n331), .ZN(n311) );
  NOR2_X1 U359 ( .A1(n335), .A2(n311), .ZN(n317) );
  INV_X1 U360 ( .A(n317), .ZN(n313) );
  AOI21_X1 U361 ( .B1(n397), .B2(n331), .A(n389), .ZN(n310) );
  OAI21_X1 U362 ( .B1(n311), .B2(n336), .A(n310), .ZN(n318) );
  INV_X1 U363 ( .A(n318), .ZN(n312) );
  OAI21_X1 U364 ( .B1(n321), .B2(n313), .A(n312), .ZN(n315) );
  NAND2_X1 U365 ( .A1(n329), .A2(n334), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U367 ( .A(n548), .B(n316), .S(n327), .Z(n474) );
  MUX2_X1 U368 ( .A(product[15]), .B(n550), .S(n327), .Z(n476) );
  NAND2_X1 U369 ( .A1(n317), .A2(n329), .ZN(n320) );
  AOI21_X1 U370 ( .B1(n318), .B2(n329), .A(n390), .ZN(n319) );
  OAI21_X1 U371 ( .B1(n321), .B2(n320), .A(n319), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n322), .B(n333), .ZN(n323) );
  MUX2_X1 U373 ( .A(n550), .B(n323), .S(n327), .Z(n478) );
  MUX2_X1 U374 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n327), .Z(n480) );
  MUX2_X1 U375 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n327), .Z(n482) );
  MUX2_X1 U376 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n327), .Z(n484) );
  MUX2_X1 U377 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n327), .Z(n486) );
  MUX2_X1 U378 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n327), .Z(n488) );
  MUX2_X1 U379 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n327), .Z(n490) );
  MUX2_X1 U380 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n327), .Z(n492) );
  MUX2_X1 U381 ( .A(n13), .B(B_extended[7]), .S(n327), .Z(n494) );
  MUX2_X1 U382 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n327), .Z(n496) );
  MUX2_X1 U383 ( .A(n7), .B(A_extended[1]), .S(n327), .Z(n498) );
  MUX2_X1 U384 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n327), .Z(n500) );
  MUX2_X1 U385 ( .A(n324), .B(A_extended[3]), .S(n327), .Z(n502) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n327), .Z(n504) );
  MUX2_X1 U387 ( .A(n325), .B(A_extended[5]), .S(n327), .Z(n506) );
  MUX2_X1 U388 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n327), .Z(n508) );
  MUX2_X1 U389 ( .A(n326), .B(A_extended[7]), .S(n327), .Z(n510) );
  OR2_X1 U390 ( .A1(n327), .A2(n553), .ZN(n512) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_25 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n397, n399, n401, n403, n405, n407, n409, n411, n413, n415, n417,
         n419, n421, n423, n425, n427, n429, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n448, n450, n452, n454, n456, n458, n460, n462, n464, n466, n468,
         n470, n472, n474, n476, n478, n480, n482, n484, n486, n488, n490,
         n492, n494, n496, n498, n500, n502, n504, n506, n508, n510, n512,
         n514, n516, n518, n520, n522, n524, n526, n528, n530, n532, n534,
         n536, n538, n540, n542, n544, n546, n548, n550, n552, n554, n556,
         n558, n560, n561, n563, n564, n566, n567, n569, n570, n572, n573,
         n575, n576, n578, n579, n581, n583, n585, n587, n589, n591, n593,
         n595, n597, n598, n599, n600, n601;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n445), .SE(n558), .CK(clk), .Q(n600), 
        .QN(n440) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n446), .SE(n554), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n446), .SE(n552), .CK(clk), .Q(n598), 
        .QN(n41) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n446), .SE(n550), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n22) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n446), .SE(n546), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n40) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n446), .SE(n542), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n31) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n446), .SE(n540), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n32) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n446), .SE(n538), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n35) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n446), .SE(n536), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n37) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n445), .SE(n534), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n36) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n445), .SE(n532), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n38) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n445), .SE(n530), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n33) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n445), .SE(n528), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n34) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n445), .SE(n526), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n445), .SE(n524), .CK(clk), .Q(n597)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n445), .SE(n522), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n445), .SE(n520), .CK(clk), .Q(n595)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n445), .SE(n518), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n445), .SE(n516), .CK(clk), .Q(n593)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n445), .SE(n514), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n444), .SE(n512), .CK(clk), .Q(n591)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n444), .SE(n510), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n444), .SE(n508), .CK(clk), .Q(n589)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n444), .SE(n506), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n444), .SE(n504), .CK(clk), .Q(n587)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n444), .SE(n502), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n444), .SE(n500), .CK(clk), .Q(n585)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n444), .SE(n498), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n444), .SE(n496), .CK(clk), .Q(n583)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n444), .SE(n494), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n444), .SE(n492), .CK(clk), .Q(n581)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n443), .SE(n490), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n443), .SE(n486), .CK(clk), .Q(n578)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n443), .SE(n484), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n443), .SE(n482), .CK(clk), .Q(n576)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n443), .SE(n480), .CK(clk), .Q(n575)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n443), .SE(n478), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n443), .SE(n476), .CK(clk), .Q(n573)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n443), .SE(n474), .CK(clk), .Q(n572)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n443), .SE(n472), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n443), .SE(n470), .CK(clk), .Q(n570)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n442), .SE(n468), .CK(clk), .Q(n569)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n442), .SE(n466), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n442), .SE(n464), .CK(clk), .Q(n567)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n442), .SE(n462), .CK(clk), .Q(n566)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n442), .SE(n460), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n442), .SE(n458), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n442), .SE(n456), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n442), .SE(n454), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n442), .SE(n452), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n442), .SE(n450), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n442), .SE(n448), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n446), .SE(n556), .CK(clk), .Q(n599), 
        .QN(n441) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n446), .SE(n544), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n43) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n446), .SE(n548), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n39) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n601), .SE(n429), .CK(
        clk), .Q(n44), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n601), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n393), .QN(n439) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n601), .SI(1'b1), .SE(n425), .CK(clk), 
        .Q(n392), .QN(n432) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n601), .SE(n423), .CK(
        clk), .Q(n45), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n601), .SE(n421), .CK(
        clk), .Q(n438), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n601), .SI(1'b1), .SE(n419), .CK(clk), 
        .Q(n389), .QN(n434) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n601), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n601), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n387), .QN(n437) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n601), .SI(1'b1), .SE(n411), .CK(clk), 
        .Q(n385), .QN(n435) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n601), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n384), .QN(n433) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n601), .SE(n407), .CK(
        clk), .Q(n436), .QN(n383) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n601), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n382), .QN(n431) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n601), .SE(n403), .CK(
        clk), .QN(n381) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n601), .SE(n401), .CK(
        clk), .QN(n380) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n601), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n379) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n601), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n378) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n601), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n377) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n601), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n386), .QN(n42) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n443), .SE(n488), .CK(clk), .Q(n579), 
        .QN(n376) );
  CLKBUF_X1 U2 ( .A(n12), .Z(n445) );
  CLKBUF_X1 U3 ( .A(n305), .Z(n12) );
  NAND2_X1 U4 ( .A1(n6), .A2(n5), .ZN(n286) );
  NAND2_X1 U5 ( .A1(n145), .A2(n146), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n144), .A2(n7), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n9), .A2(n8), .ZN(n7) );
  INV_X1 U8 ( .A(n146), .ZN(n8) );
  INV_X1 U9 ( .A(n145), .ZN(n9) );
  AND2_X1 U10 ( .A1(n600), .A2(\mult_x_1/n281 ), .ZN(n166) );
  NAND2_X1 U11 ( .A1(n273), .A2(n274), .ZN(n160) );
  XNOR2_X1 U12 ( .A(n144), .B(n10), .ZN(n274) );
  XNOR2_X1 U13 ( .A(n145), .B(n146), .ZN(n10) );
  OR2_X1 U14 ( .A1(n15), .A2(n23), .ZN(n11) );
  INV_X1 U15 ( .A(rst_n), .ZN(n601) );
  BUF_X1 U16 ( .A(n104), .Z(n165) );
  NAND2_X1 U17 ( .A1(n104), .A2(n103), .ZN(n244) );
  BUF_X1 U18 ( .A(n599), .Z(n374) );
  XNOR2_X2 U19 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n14) );
  NOR2_X1 U20 ( .A1(n80), .A2(n79), .ZN(n139) );
  OR2_X1 U21 ( .A1(n46), .A2(n47), .ZN(n30) );
  INV_X1 U22 ( .A(n269), .ZN(n265) );
  NAND2_X1 U23 ( .A1(n221), .A2(n220), .ZN(n222) );
  INV_X1 U24 ( .A(n225), .ZN(n221) );
  INV_X1 U25 ( .A(n224), .ZN(n220) );
  AND2_X1 U26 ( .A1(n81), .A2(\mult_x_1/n288 ), .ZN(n225) );
  NAND2_X1 U27 ( .A1(n113), .A2(n112), .ZN(n269) );
  XNOR2_X1 U28 ( .A(n27), .B(n36), .ZN(n169) );
  XNOR2_X1 U29 ( .A(n26), .B(n38), .ZN(n185) );
  XNOR2_X1 U30 ( .A(n27), .B(n33), .ZN(n116) );
  XNOR2_X1 U31 ( .A(n246), .B(n34), .ZN(n119) );
  OAI22_X1 U32 ( .A1(n244), .A2(n120), .B1(n165), .B2(n198), .ZN(n181) );
  INV_X1 U33 ( .A(n94), .ZN(n90) );
  INV_X1 U34 ( .A(n93), .ZN(n89) );
  XNOR2_X1 U35 ( .A(n50), .B(n85), .ZN(n92) );
  XNOR2_X1 U36 ( .A(n26), .B(n32), .ZN(n248) );
  XNOR2_X1 U37 ( .A(n84), .B(n223), .ZN(n234) );
  XNOR2_X1 U38 ( .A(n234), .B(n88), .ZN(n98) );
  XNOR2_X1 U39 ( .A(n236), .B(n235), .ZN(n88) );
  NAND2_X1 U40 ( .A1(n96), .A2(n95), .ZN(n97) );
  NAND2_X1 U41 ( .A1(n94), .A2(n93), .ZN(n95) );
  NAND2_X1 U42 ( .A1(n92), .A2(n91), .ZN(n96) );
  NAND2_X1 U43 ( .A1(n90), .A2(n89), .ZN(n91) );
  XNOR2_X1 U44 ( .A(n92), .B(n53), .ZN(n78) );
  XNOR2_X1 U45 ( .A(n94), .B(n93), .ZN(n53) );
  XNOR2_X1 U46 ( .A(n27), .B(n35), .ZN(n163) );
  NAND2_X1 U47 ( .A1(n271), .A2(n270), .ZN(n295) );
  NAND2_X1 U48 ( .A1(n227), .A2(n226), .ZN(n281) );
  NAND2_X1 U49 ( .A1(n225), .A2(n224), .ZN(n226) );
  NAND2_X1 U50 ( .A1(n223), .A2(n222), .ZN(n227) );
  NAND2_X1 U51 ( .A1(n238), .A2(n237), .ZN(n283) );
  NAND2_X1 U52 ( .A1(n236), .A2(n235), .ZN(n237) );
  NAND2_X1 U53 ( .A1(n234), .A2(n233), .ZN(n238) );
  OR2_X1 U54 ( .A1(n236), .A2(n235), .ZN(n233) );
  XNOR2_X1 U55 ( .A(n26), .B(n37), .ZN(n171) );
  OAI21_X1 U56 ( .B1(n193), .B2(n203), .A(n202), .ZN(n289) );
  NAND2_X1 U57 ( .A1(n25), .A2(n205), .ZN(n202) );
  NOR2_X1 U58 ( .A1(n25), .A2(n205), .ZN(n203) );
  NAND2_X1 U59 ( .A1(n98), .A2(n97), .ZN(n137) );
  BUF_X1 U60 ( .A(n12), .Z(n442) );
  CLKBUF_X1 U61 ( .A(n325), .Z(n21) );
  BUF_X1 U62 ( .A(n12), .Z(n443) );
  BUF_X1 U63 ( .A(n12), .Z(n444) );
  BUF_X1 U64 ( .A(n12), .Z(n446) );
  AND2_X1 U65 ( .A1(n154), .A2(n31), .ZN(n15) );
  INV_X1 U66 ( .A(n43), .ZN(n16) );
  OAI22_X1 U67 ( .A1(n200), .A2(n109), .B1(n199), .B2(n14), .ZN(n214) );
  XOR2_X1 U68 ( .A(n278), .B(n277), .Z(n17) );
  XOR2_X1 U69 ( .A(n276), .B(n17), .Z(n304) );
  NAND2_X1 U70 ( .A1(n276), .A2(n278), .ZN(n18) );
  NAND2_X1 U71 ( .A1(n276), .A2(n277), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n278), .A2(n277), .ZN(n20) );
  NAND3_X1 U73 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n273) );
  NAND2_X1 U74 ( .A1(n183), .A2(n182), .ZN(n212) );
  XNOR2_X1 U75 ( .A(n22), .B(\mult_x_1/n312 ), .ZN(n47) );
  XNOR2_X1 U76 ( .A(n166), .B(n106), .ZN(n23) );
  INV_X1 U77 ( .A(n32), .ZN(n24) );
  FA_X1 U78 ( .A(n196), .B(n195), .CI(n194), .S(n25) );
  OR2_X1 U79 ( .A1(n440), .A2(n441), .ZN(n26) );
  OR2_X1 U80 ( .A1(n440), .A2(n441), .ZN(n27) );
  OR2_X1 U81 ( .A1(n440), .A2(n441), .ZN(n246) );
  OR2_X2 U82 ( .A1(\mult_x_1/n180 ), .A2(n43), .ZN(n154) );
  INV_X1 U83 ( .A(n599), .ZN(n28) );
  INV_X1 U84 ( .A(n28), .ZN(n29) );
  OR2_X1 U85 ( .A1(n46), .A2(n47), .ZN(n189) );
  BUF_X2 U86 ( .A(n598), .Z(n373) );
  BUF_X4 U87 ( .A(en), .Z(n335) );
  XNOR2_X1 U88 ( .A(n598), .B(\mult_x_1/a[4] ), .ZN(n46) );
  OR2_X1 U89 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n48) );
  INV_X2 U90 ( .A(n47), .ZN(n187) );
  OAI22_X1 U91 ( .A1(n30), .A2(n41), .B1(n48), .B2(n187), .ZN(n86) );
  INV_X1 U92 ( .A(n86), .ZN(n50) );
  XNOR2_X1 U93 ( .A(n373), .B(\mult_x_1/n288 ), .ZN(n49) );
  XNOR2_X1 U94 ( .A(n373), .B(\mult_x_1/n287 ), .ZN(n87) );
  OAI22_X1 U95 ( .A1(n30), .A2(n49), .B1(n187), .B2(n87), .ZN(n85) );
  XNOR2_X1 U96 ( .A(\mult_x_1/n312 ), .B(n40), .ZN(n51) );
  XNOR2_X1 U97 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n52) );
  NAND2_X2 U98 ( .A1(n51), .A2(n52), .ZN(n200) );
  BUF_X2 U99 ( .A(\mult_x_1/n312 ), .Z(n372) );
  XNOR2_X1 U100 ( .A(n372), .B(\mult_x_1/n286 ), .ZN(n56) );
  XNOR2_X1 U101 ( .A(n372), .B(\mult_x_1/n285 ), .ZN(n83) );
  OAI22_X1 U102 ( .A1(n200), .A2(n56), .B1(n14), .B2(n83), .ZN(n94) );
  BUF_X2 U103 ( .A(\mult_x_1/n313 ), .Z(n106) );
  XNOR2_X1 U104 ( .A(n106), .B(\mult_x_1/n284 ), .ZN(n54) );
  XNOR2_X1 U105 ( .A(n106), .B(\mult_x_1/n283 ), .ZN(n82) );
  OAI22_X1 U106 ( .A1(n154), .A2(n54), .B1(n82), .B2(n31), .ZN(n93) );
  XNOR2_X1 U107 ( .A(n106), .B(\mult_x_1/n285 ), .ZN(n62) );
  OAI22_X1 U108 ( .A1(n154), .A2(n62), .B1(n54), .B2(n31), .ZN(n59) );
  INV_X1 U109 ( .A(n187), .ZN(n55) );
  AND2_X1 U110 ( .A1(\mult_x_1/n288 ), .A2(n55), .ZN(n58) );
  XNOR2_X1 U111 ( .A(n372), .B(\mult_x_1/n287 ), .ZN(n60) );
  OAI22_X1 U112 ( .A1(n200), .A2(n60), .B1(n14), .B2(n56), .ZN(n57) );
  OR2_X1 U113 ( .A1(n78), .A2(n77), .ZN(n329) );
  FA_X1 U114 ( .A(n59), .B(n58), .CI(n57), .CO(n77), .S(n76) );
  XNOR2_X1 U115 ( .A(n372), .B(\mult_x_1/n288 ), .ZN(n61) );
  OAI22_X1 U116 ( .A1(n200), .A2(n61), .B1(n14), .B2(n60), .ZN(n64) );
  XNOR2_X1 U117 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n66) );
  OAI22_X1 U118 ( .A1(n154), .A2(n66), .B1(n62), .B2(n31), .ZN(n63) );
  NOR2_X1 U119 ( .A1(n76), .A2(n75), .ZN(n322) );
  HA_X1 U120 ( .A(n64), .B(n63), .CO(n75), .S(n73) );
  OR2_X1 U121 ( .A1(\mult_x_1/n288 ), .A2(n39), .ZN(n65) );
  OAI22_X1 U122 ( .A1(n200), .A2(n39), .B1(n65), .B2(n14), .ZN(n72) );
  OR2_X1 U123 ( .A1(n73), .A2(n72), .ZN(n318) );
  XNOR2_X1 U124 ( .A(n16), .B(\mult_x_1/n287 ), .ZN(n68) );
  OAI22_X1 U125 ( .A1(n154), .A2(n68), .B1(n66), .B2(n31), .ZN(n71) );
  INV_X1 U126 ( .A(n14), .ZN(n67) );
  AND2_X1 U127 ( .A1(\mult_x_1/n288 ), .A2(n67), .ZN(n70) );
  NOR2_X1 U128 ( .A1(n71), .A2(n70), .ZN(n311) );
  OAI22_X1 U129 ( .A1(n154), .A2(\mult_x_1/n288 ), .B1(n68), .B2(n31), .ZN(
        n308) );
  OR2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n43), .ZN(n69) );
  NAND2_X1 U131 ( .A1(n69), .A2(n154), .ZN(n307) );
  NAND2_X1 U132 ( .A1(n308), .A2(n307), .ZN(n314) );
  NAND2_X1 U133 ( .A1(n71), .A2(n70), .ZN(n312) );
  OAI21_X1 U134 ( .B1(n311), .B2(n314), .A(n312), .ZN(n319) );
  NAND2_X1 U135 ( .A1(n73), .A2(n72), .ZN(n317) );
  INV_X1 U136 ( .A(n317), .ZN(n74) );
  AOI21_X1 U137 ( .B1(n318), .B2(n319), .A(n74), .ZN(n325) );
  NAND2_X1 U138 ( .A1(n76), .A2(n75), .ZN(n323) );
  OAI21_X1 U139 ( .B1(n322), .B2(n325), .A(n323), .ZN(n330) );
  AND2_X1 U140 ( .A1(n329), .A2(n330), .ZN(n80) );
  NAND2_X1 U141 ( .A1(n78), .A2(n77), .ZN(n328) );
  INV_X1 U142 ( .A(n328), .ZN(n79) );
  XNOR2_X1 U143 ( .A(n598), .B(\mult_x_1/a[6] ), .ZN(n104) );
  INV_X1 U144 ( .A(n165), .ZN(n81) );
  XNOR2_X1 U145 ( .A(n106), .B(\mult_x_1/n282 ), .ZN(n153) );
  OAI22_X1 U146 ( .A1(n154), .A2(n82), .B1(n153), .B2(n31), .ZN(n224) );
  XNOR2_X1 U147 ( .A(n225), .B(n224), .ZN(n84) );
  XNOR2_X1 U148 ( .A(n372), .B(\mult_x_1/n284 ), .ZN(n156) );
  OAI22_X1 U149 ( .A1(n200), .A2(n83), .B1(n14), .B2(n156), .ZN(n223) );
  AND2_X1 U150 ( .A1(n86), .A2(n85), .ZN(n236) );
  XNOR2_X1 U151 ( .A(n373), .B(\mult_x_1/n286 ), .ZN(n151) );
  OAI22_X1 U152 ( .A1(n30), .A2(n87), .B1(n187), .B2(n151), .ZN(n235) );
  OR2_X1 U153 ( .A1(n98), .A2(n97), .ZN(n138) );
  INV_X1 U154 ( .A(n138), .ZN(n99) );
  OAI21_X1 U155 ( .B1(n139), .B2(n99), .A(n137), .ZN(n100) );
  NAND2_X1 U156 ( .A1(n100), .A2(n375), .ZN(n102) );
  OR2_X1 U157 ( .A1(n375), .A2(n44), .ZN(n101) );
  NAND2_X1 U158 ( .A1(n102), .A2(n101), .ZN(n429) );
  XOR2_X1 U159 ( .A(\mult_x_1/a[6] ), .B(n599), .Z(n103) );
  XNOR2_X1 U160 ( .A(n374), .B(\mult_x_1/n285 ), .ZN(n120) );
  XNOR2_X1 U161 ( .A(n374), .B(\mult_x_1/n284 ), .ZN(n198) );
  XNOR2_X1 U162 ( .A(n373), .B(\mult_x_1/n283 ), .ZN(n108) );
  XNOR2_X1 U163 ( .A(n373), .B(\mult_x_1/n282 ), .ZN(n188) );
  OAI22_X1 U164 ( .A1(n30), .A2(n108), .B1(n187), .B2(n188), .ZN(n180) );
  XNOR2_X1 U165 ( .A(n181), .B(n180), .ZN(n105) );
  XNOR2_X1 U166 ( .A(n372), .B(\mult_x_1/n281 ), .ZN(n109) );
  XNOR2_X1 U167 ( .A(n166), .B(n372), .ZN(n199) );
  INV_X1 U168 ( .A(n214), .ZN(n179) );
  XNOR2_X1 U169 ( .A(n105), .B(n179), .ZN(n268) );
  XNOR2_X1 U170 ( .A(n374), .B(\mult_x_1/n287 ), .ZN(n128) );
  XNOR2_X1 U171 ( .A(n29), .B(\mult_x_1/n286 ), .ZN(n121) );
  OAI22_X1 U172 ( .A1(n244), .A2(n128), .B1(n165), .B2(n121), .ZN(n149) );
  XNOR2_X1 U173 ( .A(n16), .B(\mult_x_1/n281 ), .ZN(n152) );
  XNOR2_X1 U174 ( .A(n166), .B(n16), .ZN(n117) );
  OAI22_X1 U175 ( .A1(n154), .A2(n152), .B1(n117), .B2(n31), .ZN(n148) );
  XNOR2_X1 U176 ( .A(n246), .B(n441), .ZN(n118) );
  INV_X1 U177 ( .A(n118), .ZN(n107) );
  AND2_X1 U178 ( .A1(\mult_x_1/n288 ), .A2(n107), .ZN(n147) );
  XNOR2_X1 U179 ( .A(n373), .B(\mult_x_1/n284 ), .ZN(n125) );
  OAI22_X1 U180 ( .A1(n189), .A2(n125), .B1(n187), .B2(n108), .ZN(n115) );
  XNOR2_X1 U181 ( .A(n372), .B(\mult_x_1/n282 ), .ZN(n126) );
  OAI22_X1 U182 ( .A1(n200), .A2(n126), .B1(n14), .B2(n109), .ZN(n114) );
  XNOR2_X1 U183 ( .A(n115), .B(n114), .ZN(n131) );
  OR2_X1 U184 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n110) );
  XNOR2_X1 U185 ( .A(n246), .B(n441), .ZN(n247) );
  NOR2_X1 U186 ( .A1(n110), .A2(n247), .ZN(n130) );
  OR2_X1 U187 ( .A1(n130), .A2(n131), .ZN(n111) );
  NAND2_X1 U188 ( .A1(n132), .A2(n111), .ZN(n113) );
  NAND2_X1 U189 ( .A1(n131), .A2(n130), .ZN(n112) );
  XNOR2_X1 U190 ( .A(n268), .B(n269), .ZN(n122) );
  OR2_X1 U191 ( .A1(n115), .A2(n114), .ZN(n218) );
  XNOR2_X1 U192 ( .A(n26), .B(n28), .ZN(n184) );
  NOR2_X1 U193 ( .A1(n116), .A2(n184), .ZN(n217) );
  NOR2_X1 U194 ( .A1(n119), .A2(n118), .ZN(n124) );
  OAI22_X1 U195 ( .A1(n244), .A2(n121), .B1(n165), .B2(n120), .ZN(n123) );
  XNOR2_X1 U196 ( .A(n122), .B(n267), .ZN(n287) );
  FA_X1 U197 ( .A(n11), .B(n124), .CI(n123), .CO(n216), .S(n146) );
  XNOR2_X1 U198 ( .A(n373), .B(\mult_x_1/n285 ), .ZN(n150) );
  OAI22_X1 U199 ( .A1(n30), .A2(n150), .B1(n187), .B2(n125), .ZN(n159) );
  XNOR2_X1 U200 ( .A(n372), .B(\mult_x_1/n283 ), .ZN(n155) );
  OAI22_X1 U201 ( .A1(n200), .A2(n155), .B1(n14), .B2(n126), .ZN(n158) );
  OR2_X1 U202 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n127) );
  OAI22_X1 U203 ( .A1(n244), .A2(n28), .B1(n127), .B2(n165), .ZN(n229) );
  XNOR2_X1 U204 ( .A(n374), .B(\mult_x_1/n288 ), .ZN(n129) );
  OAI22_X1 U205 ( .A1(n244), .A2(n129), .B1(n165), .B2(n128), .ZN(n228) );
  XNOR2_X1 U206 ( .A(n131), .B(n130), .ZN(n133) );
  XNOR2_X1 U207 ( .A(n133), .B(n132), .ZN(n144) );
  NAND2_X1 U208 ( .A1(n287), .A2(n286), .ZN(n134) );
  NAND2_X1 U209 ( .A1(n134), .A2(n375), .ZN(n136) );
  OR2_X1 U210 ( .A1(n375), .A2(n45), .ZN(n135) );
  NAND2_X1 U211 ( .A1(n136), .A2(n135), .ZN(n423) );
  NAND2_X1 U212 ( .A1(n138), .A2(n137), .ZN(n140) );
  XNOR2_X1 U213 ( .A(n140), .B(n139), .ZN(n143) );
  INV_X1 U214 ( .A(n335), .ZN(n142) );
  OR2_X1 U215 ( .A1(n335), .A2(n376), .ZN(n141) );
  OAI21_X1 U216 ( .B1(n143), .B2(n142), .A(n141), .ZN(n488) );
  FA_X1 U217 ( .A(n149), .B(n148), .CI(n147), .CO(n132), .S(n278) );
  OAI22_X1 U218 ( .A1(n30), .A2(n151), .B1(n187), .B2(n150), .ZN(n232) );
  OAI22_X1 U219 ( .A1(n154), .A2(n153), .B1(n152), .B2(n31), .ZN(n231) );
  OAI22_X1 U220 ( .A1(n200), .A2(n156), .B1(n14), .B2(n155), .ZN(n230) );
  FA_X1 U221 ( .A(n159), .B(n158), .CI(n157), .CO(n145), .S(n276) );
  NAND2_X1 U222 ( .A1(n160), .A2(n335), .ZN(n162) );
  OR2_X1 U223 ( .A1(n335), .A2(n42), .ZN(n161) );
  NAND2_X1 U224 ( .A1(n162), .A2(n161), .ZN(n413) );
  NOR2_X1 U243 ( .A1(n163), .A2(n247), .ZN(n242) );
  XNOR2_X1 U244 ( .A(n374), .B(n24), .ZN(n164) );
  XNOR2_X1 U245 ( .A(n166), .B(n29), .ZN(n243) );
  OAI22_X1 U246 ( .A1(n244), .A2(n164), .B1(n243), .B2(n165), .ZN(n252) );
  INV_X1 U247 ( .A(n252), .ZN(n241) );
  XNOR2_X1 U248 ( .A(n374), .B(\mult_x_1/n282 ), .ZN(n170) );
  OAI22_X1 U249 ( .A1(n244), .A2(n170), .B1(n165), .B2(n164), .ZN(n174) );
  XNOR2_X1 U250 ( .A(n373), .B(n166), .ZN(n168) );
  AOI21_X1 U251 ( .B1(n187), .B2(n189), .A(n168), .ZN(n167) );
  INV_X1 U252 ( .A(n167), .ZN(n173) );
  XNOR2_X1 U253 ( .A(n373), .B(\mult_x_1/n281 ), .ZN(n186) );
  OAI22_X1 U254 ( .A1(n189), .A2(n186), .B1(n168), .B2(n187), .ZN(n172) );
  NOR2_X1 U255 ( .A1(n169), .A2(n247), .ZN(n196) );
  XNOR2_X1 U256 ( .A(n29), .B(\mult_x_1/n283 ), .ZN(n197) );
  OAI22_X1 U257 ( .A1(n244), .A2(n197), .B1(n165), .B2(n170), .ZN(n195) );
  INV_X1 U258 ( .A(n172), .ZN(n194) );
  NOR2_X1 U259 ( .A1(n171), .A2(n184), .ZN(n177) );
  FA_X1 U260 ( .A(n174), .B(n173), .CI(n172), .CO(n240), .S(n176) );
  OR2_X1 U261 ( .A1(n259), .A2(n258), .ZN(n175) );
  MUX2_X1 U262 ( .A(n377), .B(n175), .S(n335), .Z(n395) );
  FA_X1 U263 ( .A(n178), .B(n177), .CI(n176), .CO(n258), .S(n290) );
  OAI21_X1 U264 ( .B1(n181), .B2(n180), .A(n179), .ZN(n183) );
  NAND2_X1 U265 ( .A1(n181), .A2(n180), .ZN(n182) );
  NOR2_X1 U266 ( .A1(n185), .A2(n184), .ZN(n210) );
  INV_X1 U267 ( .A(n210), .ZN(n191) );
  OAI22_X1 U268 ( .A1(n30), .A2(n188), .B1(n187), .B2(n186), .ZN(n209) );
  INV_X1 U269 ( .A(n209), .ZN(n190) );
  NAND2_X1 U270 ( .A1(n191), .A2(n190), .ZN(n192) );
  AOI22_X1 U271 ( .A1(n212), .A2(n192), .B1(n209), .B2(n210), .ZN(n193) );
  INV_X1 U272 ( .A(n193), .ZN(n208) );
  FA_X1 U273 ( .A(n196), .B(n195), .CI(n194), .CO(n178), .S(n206) );
  OAI22_X1 U274 ( .A1(n244), .A2(n198), .B1(n165), .B2(n197), .ZN(n215) );
  AOI21_X1 U275 ( .B1(n14), .B2(n200), .A(n199), .ZN(n201) );
  INV_X1 U276 ( .A(n201), .ZN(n213) );
  OR2_X1 U277 ( .A1(n290), .A2(n289), .ZN(n204) );
  MUX2_X1 U278 ( .A(n378), .B(n204), .S(n335), .Z(n397) );
  XNOR2_X1 U279 ( .A(n206), .B(n205), .ZN(n207) );
  XNOR2_X1 U280 ( .A(n208), .B(n207), .ZN(n293) );
  XNOR2_X1 U281 ( .A(n210), .B(n209), .ZN(n211) );
  XNOR2_X1 U282 ( .A(n212), .B(n211), .ZN(n263) );
  FA_X1 U283 ( .A(n215), .B(n214), .CI(n213), .CO(n205), .S(n262) );
  FA_X1 U284 ( .A(n218), .B(n217), .CI(n216), .CO(n261), .S(n267) );
  OR2_X1 U285 ( .A1(n293), .A2(n292), .ZN(n219) );
  MUX2_X1 U286 ( .A(n379), .B(n219), .S(n335), .Z(n399) );
  HA_X1 U287 ( .A(n229), .B(n228), .CO(n157), .S(n280) );
  FA_X1 U288 ( .A(n232), .B(n231), .CI(n230), .CO(n277), .S(n279) );
  OR2_X1 U289 ( .A1(n284), .A2(n283), .ZN(n239) );
  MUX2_X1 U290 ( .A(n380), .B(n239), .S(n335), .Z(n401) );
  FA_X1 U291 ( .A(n242), .B(n241), .CI(n240), .CO(n254), .S(n259) );
  AOI21_X1 U292 ( .B1(n165), .B2(n244), .A(n243), .ZN(n245) );
  INV_X1 U293 ( .A(n245), .ZN(n250) );
  NOR2_X1 U294 ( .A1(n248), .A2(n247), .ZN(n249) );
  XOR2_X1 U295 ( .A(n250), .B(n249), .Z(n251) );
  XOR2_X1 U296 ( .A(n252), .B(n251), .Z(n253) );
  OR2_X1 U297 ( .A1(n254), .A2(n253), .ZN(n256) );
  NAND2_X1 U298 ( .A1(n254), .A2(n253), .ZN(n255) );
  NAND2_X1 U299 ( .A1(n256), .A2(n255), .ZN(n257) );
  MUX2_X1 U300 ( .A(n381), .B(n257), .S(n335), .Z(n403) );
  NAND2_X1 U301 ( .A1(n259), .A2(n258), .ZN(n260) );
  MUX2_X1 U302 ( .A(n382), .B(n260), .S(n335), .Z(n405) );
  FA_X1 U303 ( .A(n263), .B(n262), .CI(n261), .CO(n292), .S(n296) );
  INV_X1 U304 ( .A(n268), .ZN(n264) );
  NAND2_X1 U305 ( .A1(n265), .A2(n264), .ZN(n266) );
  NAND2_X1 U306 ( .A1(n267), .A2(n266), .ZN(n271) );
  NAND2_X1 U307 ( .A1(n269), .A2(n268), .ZN(n270) );
  NOR2_X1 U308 ( .A1(n296), .A2(n295), .ZN(n272) );
  MUX2_X1 U309 ( .A(n383), .B(n272), .S(n335), .Z(n407) );
  NOR2_X1 U310 ( .A1(n274), .A2(n273), .ZN(n275) );
  MUX2_X1 U311 ( .A(n385), .B(n275), .S(n335), .Z(n411) );
  FA_X1 U312 ( .A(n281), .B(n280), .CI(n279), .CO(n300), .S(n284) );
  NAND2_X1 U313 ( .A1(n304), .A2(n300), .ZN(n282) );
  MUX2_X1 U314 ( .A(n388), .B(n282), .S(n335), .Z(n417) );
  NAND2_X1 U315 ( .A1(n284), .A2(n283), .ZN(n285) );
  MUX2_X1 U316 ( .A(n389), .B(n285), .S(n375), .Z(n419) );
  NOR2_X1 U317 ( .A1(n287), .A2(n286), .ZN(n288) );
  MUX2_X1 U318 ( .A(n390), .B(n288), .S(n375), .Z(n421) );
  NAND2_X1 U319 ( .A1(n290), .A2(n289), .ZN(n291) );
  MUX2_X1 U320 ( .A(n392), .B(n291), .S(n375), .Z(n425) );
  NAND2_X1 U321 ( .A1(n293), .A2(n292), .ZN(n294) );
  MUX2_X1 U322 ( .A(n393), .B(n294), .S(n375), .Z(n427) );
  NAND2_X1 U323 ( .A1(n296), .A2(n295), .ZN(n297) );
  NAND2_X1 U324 ( .A1(n297), .A2(n335), .ZN(n299) );
  NAND2_X1 U325 ( .A1(n142), .A2(n384), .ZN(n298) );
  NAND2_X1 U326 ( .A1(n299), .A2(n298), .ZN(n409) );
  INV_X1 U327 ( .A(n300), .ZN(n301) );
  NAND2_X1 U328 ( .A1(n301), .A2(n335), .ZN(n303) );
  NAND2_X1 U329 ( .A1(n142), .A2(n387), .ZN(n302) );
  OAI21_X1 U330 ( .B1(n304), .B2(n303), .A(n302), .ZN(n415) );
  INV_X1 U331 ( .A(n601), .ZN(n305) );
  MUX2_X1 U332 ( .A(product[0]), .B(n560), .S(n335), .Z(n448) );
  MUX2_X1 U333 ( .A(n560), .B(n561), .S(n335), .Z(n450) );
  AND2_X1 U334 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n306) );
  MUX2_X1 U335 ( .A(n561), .B(n306), .S(n335), .Z(n452) );
  MUX2_X1 U336 ( .A(product[1]), .B(n563), .S(n335), .Z(n454) );
  MUX2_X1 U337 ( .A(n563), .B(n564), .S(n335), .Z(n456) );
  OR2_X1 U338 ( .A1(n308), .A2(n307), .ZN(n309) );
  AND2_X1 U339 ( .A1(n309), .A2(n314), .ZN(n310) );
  MUX2_X1 U340 ( .A(n564), .B(n310), .S(n335), .Z(n458) );
  MUX2_X1 U341 ( .A(product[2]), .B(n566), .S(n335), .Z(n460) );
  MUX2_X1 U342 ( .A(n566), .B(n567), .S(n335), .Z(n462) );
  INV_X1 U343 ( .A(n311), .ZN(n313) );
  NAND2_X1 U344 ( .A1(n313), .A2(n312), .ZN(n315) );
  XOR2_X1 U345 ( .A(n315), .B(n314), .Z(n316) );
  MUX2_X1 U346 ( .A(n567), .B(n316), .S(n335), .Z(n464) );
  MUX2_X1 U347 ( .A(product[3]), .B(n569), .S(n335), .Z(n466) );
  MUX2_X1 U348 ( .A(n569), .B(n570), .S(n335), .Z(n468) );
  NAND2_X1 U349 ( .A1(n318), .A2(n317), .ZN(n320) );
  XNOR2_X1 U350 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U351 ( .A(n570), .B(n321), .S(n335), .Z(n470) );
  MUX2_X1 U352 ( .A(product[4]), .B(n572), .S(n335), .Z(n472) );
  MUX2_X1 U353 ( .A(n572), .B(n573), .S(n335), .Z(n474) );
  INV_X1 U354 ( .A(n322), .ZN(n324) );
  NAND2_X1 U355 ( .A1(n324), .A2(n323), .ZN(n326) );
  XOR2_X1 U356 ( .A(n326), .B(n21), .Z(n327) );
  MUX2_X1 U357 ( .A(n573), .B(n327), .S(n335), .Z(n476) );
  MUX2_X1 U358 ( .A(product[5]), .B(n575), .S(n335), .Z(n478) );
  MUX2_X1 U359 ( .A(n575), .B(n576), .S(n335), .Z(n480) );
  NAND2_X1 U360 ( .A1(n329), .A2(n328), .ZN(n331) );
  XNOR2_X1 U361 ( .A(n331), .B(n330), .ZN(n332) );
  MUX2_X1 U362 ( .A(n576), .B(n332), .S(n335), .Z(n482) );
  MUX2_X1 U363 ( .A(product[6]), .B(n578), .S(n335), .Z(n484) );
  MUX2_X1 U364 ( .A(n578), .B(n579), .S(n335), .Z(n486) );
  MUX2_X1 U365 ( .A(product[7]), .B(n581), .S(n335), .Z(n490) );
  NAND2_X1 U366 ( .A1(n380), .A2(n389), .ZN(n333) );
  XNOR2_X1 U367 ( .A(n394), .B(n333), .ZN(n334) );
  MUX2_X1 U368 ( .A(n581), .B(n334), .S(n335), .Z(n492) );
  MUX2_X1 U369 ( .A(product[8]), .B(n583), .S(n335), .Z(n494) );
  AOI21_X1 U370 ( .B1(n394), .B2(n380), .A(n434), .ZN(n338) );
  NAND2_X1 U371 ( .A1(n437), .A2(n388), .ZN(n336) );
  XOR2_X1 U372 ( .A(n338), .B(n336), .Z(n337) );
  BUF_X4 U373 ( .A(en), .Z(n375) );
  MUX2_X1 U374 ( .A(n583), .B(n337), .S(n375), .Z(n496) );
  MUX2_X1 U375 ( .A(product[9]), .B(n585), .S(n375), .Z(n498) );
  OAI21_X1 U376 ( .B1(n338), .B2(n387), .A(n388), .ZN(n346) );
  INV_X1 U377 ( .A(n346), .ZN(n341) );
  NAND2_X1 U378 ( .A1(n435), .A2(n386), .ZN(n339) );
  XOR2_X1 U379 ( .A(n341), .B(n339), .Z(n340) );
  MUX2_X1 U380 ( .A(n585), .B(n340), .S(n375), .Z(n500) );
  MUX2_X1 U381 ( .A(product[10]), .B(n587), .S(n375), .Z(n502) );
  OAI21_X1 U382 ( .B1(n341), .B2(n385), .A(n386), .ZN(n343) );
  NAND2_X1 U383 ( .A1(n438), .A2(n391), .ZN(n342) );
  XNOR2_X1 U384 ( .A(n343), .B(n342), .ZN(n344) );
  MUX2_X1 U385 ( .A(n587), .B(n344), .S(n375), .Z(n504) );
  MUX2_X1 U386 ( .A(product[11]), .B(n589), .S(n375), .Z(n506) );
  NOR2_X1 U387 ( .A1(n390), .A2(n385), .ZN(n347) );
  OAI21_X1 U388 ( .B1(n390), .B2(n386), .A(n391), .ZN(n345) );
  AOI21_X1 U389 ( .B1(n347), .B2(n346), .A(n345), .ZN(n369) );
  NAND2_X1 U390 ( .A1(n436), .A2(n384), .ZN(n348) );
  XOR2_X1 U391 ( .A(n369), .B(n348), .Z(n349) );
  MUX2_X1 U392 ( .A(n589), .B(n349), .S(n375), .Z(n508) );
  MUX2_X1 U393 ( .A(product[12]), .B(n591), .S(n375), .Z(n510) );
  OAI21_X1 U394 ( .B1(n369), .B2(n383), .A(n384), .ZN(n351) );
  NAND2_X1 U395 ( .A1(n379), .A2(n393), .ZN(n350) );
  XNOR2_X1 U396 ( .A(n351), .B(n350), .ZN(n352) );
  MUX2_X1 U397 ( .A(n591), .B(n352), .S(n375), .Z(n512) );
  MUX2_X1 U398 ( .A(product[13]), .B(n593), .S(n375), .Z(n514) );
  NAND2_X1 U399 ( .A1(n436), .A2(n379), .ZN(n354) );
  AOI21_X1 U400 ( .B1(n433), .B2(n379), .A(n439), .ZN(n353) );
  OAI21_X1 U401 ( .B1(n369), .B2(n354), .A(n353), .ZN(n356) );
  NAND2_X1 U402 ( .A1(n378), .A2(n392), .ZN(n355) );
  XNOR2_X1 U403 ( .A(n356), .B(n355), .ZN(n357) );
  MUX2_X1 U404 ( .A(n593), .B(n357), .S(n375), .Z(n516) );
  MUX2_X1 U405 ( .A(product[14]), .B(n595), .S(n375), .Z(n518) );
  NAND2_X1 U406 ( .A1(n379), .A2(n378), .ZN(n359) );
  NOR2_X1 U407 ( .A1(n383), .A2(n359), .ZN(n365) );
  INV_X1 U408 ( .A(n365), .ZN(n361) );
  AOI21_X1 U409 ( .B1(n439), .B2(n378), .A(n432), .ZN(n358) );
  OAI21_X1 U410 ( .B1(n359), .B2(n384), .A(n358), .ZN(n366) );
  INV_X1 U411 ( .A(n366), .ZN(n360) );
  OAI21_X1 U412 ( .B1(n369), .B2(n361), .A(n360), .ZN(n363) );
  NAND2_X1 U413 ( .A1(n377), .A2(n382), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n364) );
  MUX2_X1 U415 ( .A(n595), .B(n364), .S(n375), .Z(n520) );
  MUX2_X1 U416 ( .A(product[15]), .B(n597), .S(n375), .Z(n522) );
  NAND2_X1 U417 ( .A1(n365), .A2(n377), .ZN(n368) );
  AOI21_X1 U418 ( .B1(n366), .B2(n377), .A(n431), .ZN(n367) );
  OAI21_X1 U419 ( .B1(n369), .B2(n368), .A(n367), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n370), .B(n381), .ZN(n371) );
  MUX2_X1 U421 ( .A(n597), .B(n371), .S(n375), .Z(n524) );
  MUX2_X1 U422 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n375), .Z(n526) );
  MUX2_X1 U423 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n375), .Z(n528) );
  MUX2_X1 U424 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n375), .Z(n530) );
  MUX2_X1 U425 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n375), .Z(n532) );
  MUX2_X1 U426 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n375), .Z(n534) );
  MUX2_X1 U427 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n375), .Z(n536) );
  MUX2_X1 U428 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n375), .Z(n538) );
  MUX2_X1 U429 ( .A(n24), .B(B_extended[7]), .S(n375), .Z(n540) );
  MUX2_X1 U430 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n375), .Z(n542) );
  MUX2_X1 U431 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n375), .Z(n544) );
  MUX2_X1 U432 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n375), .Z(n546) );
  MUX2_X1 U433 ( .A(n372), .B(A_extended[3]), .S(n375), .Z(n548) );
  MUX2_X1 U434 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n375), .Z(n550) );
  MUX2_X1 U435 ( .A(n373), .B(A_extended[5]), .S(n375), .Z(n552) );
  MUX2_X1 U436 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n375), .Z(n554) );
  MUX2_X1 U437 ( .A(n374), .B(A_extended[7]), .S(n375), .Z(n556) );
  OR2_X1 U438 ( .A1(n375), .A2(n600), .ZN(n558) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_26 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n403, n405, n407,
         n409, n411, n413, n415, n417, n419, n421, n423, n425, n427, n429,
         n431, n433, n435, n437, n439, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n522, n524, n526,
         n528, n530, n532, n534, n536, n538, n540, n542, n544, n546, n548,
         n550, n552, n554, n556, n558, n560, n562, n564, n566, n568, n570,
         n572, n574, n576, n578, n580, n582, n584, n586, n588, n590, n592,
         n594, n596, n598, n600, n602, n604, n606, n608, n610, n612, n614,
         n616, n618, n620, n622, n624, n626, n628, n630, n647, n648, n649;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n465), .SE(n630), .CK(clk), .Q(n648), 
        .QN(n466) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n465), .SE(n626), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n468) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n465), .SE(n624), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n469) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n465), .SE(n622), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n470) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n465), .SE(n620), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n471) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n465), .SE(n618), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n472) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n465), .SE(n616), .CK(clk), .Q(n647), 
        .QN(n473) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n465), .SE(n614), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n474) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n465), .SE(n612), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n475) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n465), .SE(n610), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n476) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n464), .SE(n608), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n477) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n464), .SE(n606), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n478) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n464), .SE(n604), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n479) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n464), .SE(n602), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n480) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n464), .SE(n600), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n481) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n464), .SE(n598), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n482) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n464), .SE(n596), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n464), .SE(n594), .CK(clk), .Q(
        product[15]), .QN(n484) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n464), .SE(n592), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n464), .SE(n590), .CK(clk), .Q(
        product[14]), .QN(n486) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n464), .SE(n588), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n463), .SE(n586), .CK(clk), .Q(
        product[13]), .QN(n488) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n463), .SE(n584), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n463), .SE(n582), .CK(clk), .Q(
        product[12]), .QN(n490) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n463), .SE(n580), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n463), .SE(n578), .CK(clk), .Q(
        product[11]), .QN(n492) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n463), .SE(n576), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n463), .SE(n574), .CK(clk), .Q(
        product[10]), .QN(n494) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n463), .SE(n572), .CK(clk), .QN(n495)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n463), .SE(n570), .CK(clk), .Q(
        product[9]), .QN(n496) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n463), .SE(n568), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n463), .SE(n566), .CK(clk), .Q(
        product[8]), .QN(n498) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n462), .SE(n564), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n462), .SE(n562), .CK(clk), .Q(
        product[7]), .QN(n500) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n462), .SE(n560), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n462), .SE(n558), .CK(clk), .Q(
        product[6]), .QN(n502) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n462), .SE(n554), .CK(clk), .QN(n504)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n462), .SE(n552), .CK(clk), .Q(
        product[5]), .QN(n505) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n462), .SE(n550), .CK(clk), .QN(n506)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n462), .SE(n548), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n462), .SE(n546), .CK(clk), .Q(
        product[4]), .QN(n508) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n462), .SE(n544), .CK(clk), .QN(n509)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n461), .SE(n542), .CK(clk), .QN(n510)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n461), .SE(n540), .CK(clk), .Q(
        product[3]), .QN(n511) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n461), .SE(n538), .CK(clk), .QN(n512)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n461), .SE(n536), .CK(clk), .QN(n513)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n461), .SE(n534), .CK(clk), .Q(
        product[2]), .QN(n514) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n461), .SE(n532), .CK(clk), .QN(n515)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n461), .SE(n530), .CK(clk), .QN(n516)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n461), .SE(n528), .CK(clk), .Q(
        product[1]), .QN(n517) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n461), .SE(n526), .CK(clk), .QN(n518)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n461), .SE(n524), .CK(clk), .QN(n519)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n461), .SE(n522), .CK(clk), .Q(
        product[0]), .QN(n520) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n649), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n381), .QN(n460) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n649), .SI(1'b1), .SE(n439), .CK(clk), 
        .Q(n400), .QN(n441) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n649), .SI(1'b1), .SE(n437), .CK(clk), 
        .Q(n399), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n649), .SI(1'b1), .SE(n433), .CK(clk), 
        .Q(n397), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n649), .SI(1'b1), .SE(n431), .CK(clk), 
        .Q(n396), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n649), .SI(1'b1), .SE(n429), .CK(clk), 
        .Q(n395), .QN(n446) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n649), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n394), .QN(n447) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n649), .SE(n425), .CK(
        clk), .Q(n448), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n649), .SE(n423), .CK(
        clk), .Q(n449), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n649), .SI(1'b1), .SE(n421), .CK(clk), 
        .Q(n391), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n649), .SI(1'b1), .SE(n419), .CK(clk), 
        .Q(n390), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n649), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n389), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n649), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n388), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n649), .SI(1'b1), .SE(n411), .CK(clk), 
        .Q(n386), .QN(n455) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n649), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n385), .QN(n456) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n649), .SE(n407), .CK(
        clk), .Q(n457), .QN(n384) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n649), .SE(n405), .CK(
        clk), .Q(n458), .QN(n383) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n649), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n382), .QN(n459) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n465), .SE(n628), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n467) );
  SDFF_X2 clk_r_REG42_S2 ( .D(1'b0), .SI(n462), .SE(n556), .CK(clk), .QN(n503)
         );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n649), .SE(n435), .CK(
        clk), .Q(n443), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n649), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n387), .QN(n454) );
  BUF_X1 U2 ( .A(n273), .Z(n380) );
  BUF_X1 U3 ( .A(n273), .Z(n288) );
  INV_X1 U4 ( .A(n146), .ZN(n5) );
  AND2_X1 U5 ( .A1(n145), .A2(n146), .ZN(n48) );
  XNOR2_X1 U6 ( .A(n5), .B(n145), .ZN(n189) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(n413) );
  OR2_X1 U8 ( .A1(n267), .A2(n454), .ZN(n6) );
  NAND2_X1 U9 ( .A1(n191), .A2(n377), .ZN(n7) );
  BUF_X2 U10 ( .A(\mult_x_1/n310 ), .Z(n18) );
  CLKBUF_X2 U11 ( .A(n351), .Z(n213) );
  CLKBUF_X1 U12 ( .A(n272), .Z(n461) );
  CLKBUF_X1 U13 ( .A(n272), .Z(n462) );
  CLKBUF_X1 U14 ( .A(n272), .Z(n463) );
  CLKBUF_X1 U15 ( .A(n272), .Z(n464) );
  CLKBUF_X1 U16 ( .A(n272), .Z(n465) );
  INV_X1 U17 ( .A(rst_n), .ZN(n649) );
  CLKBUF_X1 U18 ( .A(n155), .Z(n8) );
  BUF_X1 U19 ( .A(n31), .Z(n168) );
  XNOR2_X1 U20 ( .A(\mult_x_1/a[2] ), .B(n471), .ZN(n24) );
  BUF_X1 U21 ( .A(n155), .Z(n9) );
  XNOR2_X1 U22 ( .A(n120), .B(n647), .ZN(n10) );
  INV_X1 U23 ( .A(n66), .ZN(n11) );
  INV_X1 U24 ( .A(n475), .ZN(n12) );
  OR2_X1 U25 ( .A1(n373), .A2(n446), .ZN(n13) );
  NAND2_X1 U26 ( .A1(n13), .A2(n222), .ZN(n429) );
  CLKBUF_X1 U27 ( .A(n95), .Z(n14) );
  OR2_X1 U28 ( .A1(n98), .A2(n97), .ZN(n88) );
  INV_X2 U29 ( .A(n288), .ZN(n371) );
  NAND2_X1 U30 ( .A1(n98), .A2(n97), .ZN(n89) );
  NAND2_X1 U31 ( .A1(n102), .A2(n101), .ZN(n219) );
  NAND2_X1 U32 ( .A1(n112), .A2(n110), .ZN(n101) );
  INV_X1 U33 ( .A(n649), .ZN(n272) );
  OR2_X1 U34 ( .A1(n373), .A2(n453), .ZN(n17) );
  NAND2_X1 U35 ( .A1(n66), .A2(n65), .ZN(n68) );
  OAI22_X1 U36 ( .A1(n165), .A2(n38), .B1(n57), .B2(n166), .ZN(n65) );
  XNOR2_X1 U37 ( .A(n473), .B(n472), .ZN(n15) );
  NAND2_X1 U38 ( .A1(n25), .A2(n26), .ZN(n165) );
  INV_X1 U39 ( .A(n23), .ZN(n16) );
  INV_X1 U40 ( .A(n23), .ZN(n227) );
  NAND2_X1 U41 ( .A1(n17), .A2(n196), .ZN(n415) );
  AND2_X2 U42 ( .A1(n648), .A2(\mult_x_1/n281 ), .ZN(n120) );
  OAI21_X1 U43 ( .B1(n112), .B2(n110), .A(n109), .ZN(n102) );
  BUF_X2 U44 ( .A(n60), .Z(n241) );
  INV_X2 U45 ( .A(n288), .ZN(n379) );
  INV_X2 U46 ( .A(n273), .ZN(n351) );
  XOR2_X1 U47 ( .A(n71), .B(n69), .Z(n19) );
  AND3_X1 U48 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n20) );
  BUF_X1 U49 ( .A(n351), .Z(n267) );
  XOR2_X1 U50 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[4] ), .Z(n21) );
  XNOR2_X1 U51 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n22) );
  NAND2_X1 U52 ( .A1(n21), .A2(n22), .ZN(n155) );
  BUF_X2 U53 ( .A(\mult_x_1/n311 ), .Z(n151) );
  XNOR2_X1 U54 ( .A(n151), .B(\mult_x_1/n285 ), .ZN(n45) );
  INV_X1 U55 ( .A(n22), .ZN(n23) );
  XNOR2_X1 U56 ( .A(n151), .B(\mult_x_1/n284 ), .ZN(n34) );
  OAI22_X1 U57 ( .A1(n9), .A2(n45), .B1(n16), .B2(n34), .ZN(n50) );
  NAND2_X1 U58 ( .A1(n24), .A2(n15), .ZN(n60) );
  CLKBUF_X2 U59 ( .A(\mult_x_1/n312 ), .Z(n239) );
  XNOR2_X1 U60 ( .A(n239), .B(\mult_x_1/n283 ), .ZN(n47) );
  BUF_X1 U61 ( .A(n15), .Z(n243) );
  XNOR2_X1 U62 ( .A(n239), .B(\mult_x_1/n282 ), .ZN(n35) );
  OAI22_X1 U63 ( .A1(n241), .A2(n47), .B1(n243), .B2(n35), .ZN(n49) );
  XNOR2_X1 U64 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n26) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n310 ), .B(n468), .ZN(n25) );
  OR2_X1 U66 ( .A1(\mult_x_1/n288 ), .A2(n467), .ZN(n28) );
  INV_X1 U67 ( .A(n26), .ZN(n27) );
  INV_X2 U68 ( .A(n27), .ZN(n166) );
  OAI22_X1 U69 ( .A1(n165), .A2(n467), .B1(n28), .B2(n166), .ZN(n146) );
  XNOR2_X1 U70 ( .A(n18), .B(\mult_x_1/n288 ), .ZN(n29) );
  XNOR2_X1 U71 ( .A(n18), .B(\mult_x_1/n287 ), .ZN(n39) );
  OAI22_X1 U72 ( .A1(n165), .A2(n29), .B1(n166), .B2(n39), .ZN(n145) );
  XNOR2_X1 U73 ( .A(n18), .B(\mult_x_1/n286 ), .ZN(n38) );
  XNOR2_X1 U74 ( .A(n18), .B(\mult_x_1/n285 ), .ZN(n57) );
  NAND2_X1 U75 ( .A1(n647), .A2(n474), .ZN(n247) );
  XNOR2_X1 U76 ( .A(n120), .B(n647), .ZN(n40) );
  AOI21_X1 U77 ( .B1(n247), .B2(n474), .A(n10), .ZN(n30) );
  INV_X1 U78 ( .A(n30), .ZN(n66) );
  XNOR2_X1 U79 ( .A(n65), .B(n11), .ZN(n33) );
  AND2_X1 U80 ( .A1(n648), .A2(\mult_x_1/n310 ), .ZN(n31) );
  XNOR2_X1 U81 ( .A(n168), .B(\mult_x_1/n287 ), .ZN(n32) );
  XNOR2_X1 U82 ( .A(n31), .B(n467), .ZN(n41) );
  INV_X1 U83 ( .A(n41), .ZN(n169) );
  NOR2_X1 U84 ( .A1(n32), .A2(n169), .ZN(n64) );
  XNOR2_X1 U85 ( .A(n33), .B(n64), .ZN(n69) );
  XNOR2_X1 U86 ( .A(n151), .B(\mult_x_1/n283 ), .ZN(n58) );
  OAI22_X1 U87 ( .A1(n9), .A2(n34), .B1(n16), .B2(n58), .ZN(n62) );
  CLKBUF_X1 U88 ( .A(n60), .Z(n235) );
  XNOR2_X1 U89 ( .A(n239), .B(\mult_x_1/n281 ), .ZN(n59) );
  OAI22_X1 U90 ( .A1(n235), .A2(n35), .B1(n243), .B2(n59), .ZN(n61) );
  XNOR2_X1 U91 ( .A(n62), .B(n61), .ZN(n56) );
  INV_X1 U92 ( .A(n168), .ZN(n36) );
  OR2_X1 U93 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n37) );
  NOR2_X1 U94 ( .A1(n37), .A2(n169), .ZN(n55) );
  OAI22_X1 U95 ( .A1(n165), .A2(n39), .B1(n166), .B2(n38), .ZN(n44) );
  XNOR2_X1 U96 ( .A(n647), .B(\mult_x_1/n281 ), .ZN(n46) );
  OAI22_X1 U97 ( .A1(n247), .A2(n46), .B1(n40), .B2(n474), .ZN(n43) );
  AND2_X1 U98 ( .A1(n41), .A2(\mult_x_1/n288 ), .ZN(n42) );
  XNOR2_X1 U99 ( .A(n19), .B(n70), .ZN(n262) );
  FA_X1 U100 ( .A(n44), .B(n43), .CI(n42), .CO(n54), .S(n187) );
  XNOR2_X1 U101 ( .A(n151), .B(\mult_x_1/n286 ), .ZN(n153) );
  OAI22_X1 U102 ( .A1(n9), .A2(n153), .B1(n16), .B2(n45), .ZN(n149) );
  XNOR2_X1 U103 ( .A(n647), .B(\mult_x_1/n282 ), .ZN(n142) );
  OAI22_X1 U104 ( .A1(n247), .A2(n142), .B1(n46), .B2(n474), .ZN(n148) );
  XNOR2_X1 U105 ( .A(n239), .B(\mult_x_1/n284 ), .ZN(n144) );
  OAI22_X1 U106 ( .A1(n241), .A2(n144), .B1(n243), .B2(n47), .ZN(n147) );
  FA_X1 U107 ( .A(n50), .B(n49), .CI(n48), .CO(n71), .S(n185) );
  NAND2_X1 U108 ( .A1(n262), .A2(n261), .ZN(n51) );
  INV_X1 U109 ( .A(en), .ZN(n273) );
  NAND2_X1 U110 ( .A1(n51), .A2(n371), .ZN(n53) );
  OR2_X1 U111 ( .A1(n373), .A2(n455), .ZN(n52) );
  NAND2_X1 U112 ( .A1(n53), .A2(n52), .ZN(n411) );
  FA_X1 U113 ( .A(n56), .B(n55), .CI(n54), .CO(n115), .S(n70) );
  XNOR2_X1 U114 ( .A(n18), .B(\mult_x_1/n284 ), .ZN(n79) );
  OAI22_X1 U115 ( .A1(n165), .A2(n57), .B1(n166), .B2(n79), .ZN(n84) );
  XNOR2_X1 U116 ( .A(n151), .B(\mult_x_1/n282 ), .ZN(n87) );
  OAI22_X1 U117 ( .A1(n9), .A2(n58), .B1(n227), .B2(n87), .ZN(n83) );
  XNOR2_X1 U118 ( .A(n120), .B(n239), .ZN(n80) );
  OAI22_X1 U119 ( .A1(n60), .A2(n59), .B1(n80), .B2(n15), .ZN(n95) );
  INV_X1 U120 ( .A(n95), .ZN(n82) );
  OR2_X1 U121 ( .A1(n61), .A2(n62), .ZN(n93) );
  XNOR2_X1 U122 ( .A(n168), .B(\mult_x_1/n286 ), .ZN(n63) );
  NOR2_X1 U123 ( .A1(n63), .A2(n169), .ZN(n92) );
  OAI21_X1 U124 ( .B1(n66), .B2(n65), .A(n64), .ZN(n67) );
  NAND2_X1 U125 ( .A1(n68), .A2(n67), .ZN(n91) );
  INV_X1 U126 ( .A(n69), .ZN(n72) );
  NAND2_X1 U127 ( .A1(n70), .A2(n72), .ZN(n75) );
  NAND2_X1 U128 ( .A1(n70), .A2(n71), .ZN(n74) );
  NAND2_X1 U129 ( .A1(n72), .A2(n71), .ZN(n73) );
  NAND2_X1 U130 ( .A1(n20), .A2(n213), .ZN(n76) );
  OAI22_X1 U131 ( .A1(n108), .A2(n76), .B1(n373), .B2(n449), .ZN(n423) );
  XNOR2_X1 U132 ( .A(n151), .B(\mult_x_1/n281 ), .ZN(n86) );
  XNOR2_X1 U133 ( .A(n120), .B(n151), .ZN(n123) );
  OAI22_X1 U134 ( .A1(n8), .A2(n86), .B1(n123), .B2(n227), .ZN(n130) );
  INV_X1 U135 ( .A(n130), .ZN(n127) );
  XNOR2_X1 U136 ( .A(n18), .B(\mult_x_1/n283 ), .ZN(n78) );
  XNOR2_X1 U137 ( .A(n18), .B(\mult_x_1/n282 ), .ZN(n122) );
  OAI22_X1 U138 ( .A1(n165), .A2(n78), .B1(n166), .B2(n122), .ZN(n126) );
  XNOR2_X1 U139 ( .A(n168), .B(\mult_x_1/n284 ), .ZN(n77) );
  NOR2_X1 U140 ( .A1(n77), .A2(n169), .ZN(n125) );
  OAI22_X1 U141 ( .A1(n165), .A2(n79), .B1(n166), .B2(n78), .ZN(n96) );
  AOI21_X1 U142 ( .B1(n243), .B2(n241), .A(n80), .ZN(n81) );
  INV_X1 U143 ( .A(n81), .ZN(n94) );
  FA_X1 U144 ( .A(n84), .B(n83), .CI(n82), .CO(n100), .S(n114) );
  XNOR2_X1 U145 ( .A(n168), .B(\mult_x_1/n285 ), .ZN(n85) );
  NOR2_X1 U146 ( .A1(n85), .A2(n169), .ZN(n98) );
  OAI22_X1 U147 ( .A1(n9), .A2(n87), .B1(n227), .B2(n86), .ZN(n97) );
  NAND2_X1 U148 ( .A1(n100), .A2(n88), .ZN(n90) );
  NAND2_X1 U149 ( .A1(n90), .A2(n89), .ZN(n137) );
  FA_X1 U150 ( .A(n93), .B(n92), .CI(n91), .CO(n112), .S(n113) );
  FA_X1 U151 ( .A(n96), .B(n14), .CI(n94), .CO(n138), .S(n110) );
  XNOR2_X1 U152 ( .A(n98), .B(n97), .ZN(n99) );
  XNOR2_X1 U153 ( .A(n100), .B(n99), .ZN(n109) );
  OR2_X1 U154 ( .A1(n220), .A2(n219), .ZN(n103) );
  NAND2_X1 U155 ( .A1(n103), .A2(n267), .ZN(n105) );
  OR2_X1 U156 ( .A1(n213), .A2(n444), .ZN(n104) );
  NAND2_X1 U157 ( .A1(n105), .A2(n104), .ZN(n433) );
  OR2_X1 U158 ( .A1(n213), .A2(n448), .ZN(n107) );
  NAND2_X1 U159 ( .A1(n20), .A2(n213), .ZN(n106) );
  OAI211_X1 U160 ( .C1(n108), .C2(n380), .A(n107), .B(n106), .ZN(n425) );
  XNOR2_X1 U161 ( .A(n110), .B(n109), .ZN(n111) );
  XNOR2_X1 U162 ( .A(n112), .B(n111), .ZN(n271) );
  FA_X1 U163 ( .A(n115), .B(n114), .CI(n113), .CO(n266), .S(n108) );
  NAND2_X1 U164 ( .A1(n271), .A2(n266), .ZN(n116) );
  NAND2_X1 U165 ( .A1(n116), .A2(n267), .ZN(n118) );
  OR2_X1 U166 ( .A1(n213), .A2(n442), .ZN(n117) );
  NAND2_X1 U167 ( .A1(n118), .A2(n117), .ZN(n437) );
  XNOR2_X1 U188 ( .A(n168), .B(\mult_x_1/n282 ), .ZN(n119) );
  NOR2_X1 U189 ( .A1(n119), .A2(n169), .ZN(n163) );
  XNOR2_X1 U190 ( .A(n18), .B(\mult_x_1/n281 ), .ZN(n121) );
  XNOR2_X1 U191 ( .A(n120), .B(n18), .ZN(n164) );
  OAI22_X1 U192 ( .A1(n165), .A2(n121), .B1(n164), .B2(n166), .ZN(n174) );
  INV_X1 U193 ( .A(n174), .ZN(n162) );
  OAI22_X1 U194 ( .A1(n165), .A2(n122), .B1(n166), .B2(n121), .ZN(n131) );
  AOI21_X1 U195 ( .B1(n9), .B2(n227), .A(n123), .ZN(n124) );
  INV_X1 U196 ( .A(n124), .ZN(n129) );
  FA_X1 U197 ( .A(n127), .B(n126), .CI(n125), .CO(n136), .S(n139) );
  XNOR2_X1 U198 ( .A(n168), .B(\mult_x_1/n283 ), .ZN(n128) );
  NOR2_X1 U199 ( .A1(n128), .A2(n169), .ZN(n135) );
  FA_X1 U200 ( .A(n131), .B(n130), .CI(n129), .CO(n161), .S(n134) );
  OR2_X1 U201 ( .A1(n182), .A2(n181), .ZN(n132) );
  NAND2_X1 U202 ( .A1(n267), .A2(n132), .ZN(n133) );
  OAI21_X1 U203 ( .B1(n267), .B2(n460), .A(n133), .ZN(n401) );
  FA_X1 U204 ( .A(n136), .B(n135), .CI(n134), .CO(n181), .S(n216) );
  FA_X1 U205 ( .A(n139), .B(n138), .CI(n137), .CO(n215), .S(n220) );
  OR2_X1 U206 ( .A1(n216), .A2(n215), .ZN(n140) );
  NAND2_X1 U207 ( .A1(n267), .A2(n140), .ZN(n141) );
  OAI21_X1 U208 ( .B1(n373), .B2(n459), .A(n141), .ZN(n403) );
  XNOR2_X1 U209 ( .A(n647), .B(\mult_x_1/n283 ), .ZN(n205) );
  OAI22_X1 U210 ( .A1(n247), .A2(n205), .B1(n142), .B2(n474), .ZN(n158) );
  INV_X1 U211 ( .A(n166), .ZN(n143) );
  AND2_X1 U212 ( .A1(\mult_x_1/n288 ), .A2(n143), .ZN(n157) );
  XNOR2_X1 U213 ( .A(n239), .B(\mult_x_1/n285 ), .ZN(n204) );
  OAI22_X1 U214 ( .A1(n241), .A2(n204), .B1(n243), .B2(n144), .ZN(n156) );
  FA_X1 U215 ( .A(n149), .B(n148), .CI(n147), .CO(n186), .S(n188) );
  OR2_X1 U216 ( .A1(\mult_x_1/n288 ), .A2(n469), .ZN(n150) );
  OAI22_X1 U217 ( .A1(n8), .A2(n469), .B1(n150), .B2(n227), .ZN(n207) );
  XNOR2_X1 U218 ( .A(n151), .B(\mult_x_1/n288 ), .ZN(n152) );
  XNOR2_X1 U219 ( .A(n151), .B(\mult_x_1/n287 ), .ZN(n154) );
  OAI22_X1 U220 ( .A1(n8), .A2(n152), .B1(n227), .B2(n154), .ZN(n206) );
  OAI22_X1 U221 ( .A1(n9), .A2(n154), .B1(n16), .B2(n153), .ZN(n202) );
  FA_X1 U222 ( .A(n158), .B(n157), .CI(n156), .CO(n190), .S(n201) );
  OR2_X1 U223 ( .A1(n198), .A2(n197), .ZN(n159) );
  NAND2_X1 U224 ( .A1(n267), .A2(n159), .ZN(n160) );
  OAI21_X1 U225 ( .B1(n373), .B2(n458), .A(n160), .ZN(n405) );
  FA_X1 U226 ( .A(n163), .B(n162), .CI(n161), .CO(n176), .S(n182) );
  AOI21_X1 U227 ( .B1(n166), .B2(n165), .A(n164), .ZN(n167) );
  INV_X1 U228 ( .A(n167), .ZN(n172) );
  XNOR2_X1 U229 ( .A(n168), .B(n12), .ZN(n170) );
  NOR2_X1 U230 ( .A1(n170), .A2(n169), .ZN(n171) );
  XOR2_X1 U231 ( .A(n172), .B(n171), .Z(n173) );
  XOR2_X1 U232 ( .A(n174), .B(n173), .Z(n175) );
  OR2_X1 U233 ( .A1(n176), .A2(n175), .ZN(n178) );
  NAND2_X1 U234 ( .A1(n176), .A2(n175), .ZN(n177) );
  NAND2_X1 U235 ( .A1(n178), .A2(n177), .ZN(n179) );
  NAND2_X1 U236 ( .A1(n213), .A2(n179), .ZN(n180) );
  OAI21_X1 U237 ( .B1(n267), .B2(n457), .A(n180), .ZN(n407) );
  NAND2_X1 U238 ( .A1(n182), .A2(n181), .ZN(n183) );
  NAND2_X1 U239 ( .A1(n213), .A2(n183), .ZN(n184) );
  OAI21_X1 U240 ( .B1(n377), .B2(n456), .A(n184), .ZN(n409) );
  FA_X1 U241 ( .A(n187), .B(n186), .CI(n185), .CO(n261), .S(n194) );
  FA_X1 U242 ( .A(n190), .B(n189), .CI(n188), .CO(n193), .S(n198) );
  NOR2_X1 U243 ( .A1(n194), .A2(n193), .ZN(n191) );
  NAND2_X1 U244 ( .A1(n194), .A2(n193), .ZN(n195) );
  NAND2_X1 U245 ( .A1(n371), .A2(n195), .ZN(n196) );
  NAND2_X1 U246 ( .A1(n198), .A2(n197), .ZN(n199) );
  NAND2_X1 U247 ( .A1(n379), .A2(n199), .ZN(n200) );
  OAI21_X1 U248 ( .B1(n267), .B2(n452), .A(n200), .ZN(n417) );
  FA_X1 U249 ( .A(n203), .B(n202), .CI(n201), .CO(n197), .S(n211) );
  XNOR2_X1 U250 ( .A(n239), .B(\mult_x_1/n286 ), .ZN(n229) );
  OAI22_X1 U251 ( .A1(n241), .A2(n229), .B1(n243), .B2(n204), .ZN(n225) );
  XNOR2_X1 U252 ( .A(n647), .B(\mult_x_1/n284 ), .ZN(n226) );
  OAI22_X1 U253 ( .A1(n247), .A2(n226), .B1(n205), .B2(n474), .ZN(n224) );
  HA_X1 U254 ( .A(n206), .B(n207), .CO(n203), .S(n223) );
  NOR2_X1 U255 ( .A1(n211), .A2(n210), .ZN(n208) );
  NAND2_X1 U256 ( .A1(n213), .A2(n208), .ZN(n209) );
  OAI21_X1 U257 ( .B1(n267), .B2(n451), .A(n209), .ZN(n419) );
  NAND2_X1 U258 ( .A1(n211), .A2(n210), .ZN(n212) );
  NAND2_X1 U259 ( .A1(n267), .A2(n212), .ZN(n214) );
  OAI21_X1 U260 ( .B1(n373), .B2(n450), .A(n214), .ZN(n421) );
  NAND2_X1 U261 ( .A1(n216), .A2(n215), .ZN(n217) );
  NAND2_X1 U262 ( .A1(n213), .A2(n217), .ZN(n218) );
  OAI21_X1 U263 ( .B1(n377), .B2(n447), .A(n218), .ZN(n427) );
  NAND2_X1 U264 ( .A1(n220), .A2(n219), .ZN(n221) );
  NAND2_X1 U265 ( .A1(n213), .A2(n221), .ZN(n222) );
  FA_X1 U266 ( .A(n225), .B(n224), .CI(n223), .CO(n210), .S(n257) );
  XNOR2_X1 U267 ( .A(n647), .B(\mult_x_1/n285 ), .ZN(n236) );
  OAI22_X1 U268 ( .A1(n247), .A2(n236), .B1(n226), .B2(n474), .ZN(n232) );
  INV_X1 U269 ( .A(n16), .ZN(n228) );
  AND2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(n228), .ZN(n231) );
  XNOR2_X1 U271 ( .A(n239), .B(\mult_x_1/n287 ), .ZN(n233) );
  OAI22_X1 U272 ( .A1(n235), .A2(n233), .B1(n243), .B2(n229), .ZN(n230) );
  OR2_X1 U273 ( .A1(n257), .A2(n256), .ZN(n303) );
  FA_X1 U274 ( .A(n232), .B(n231), .CI(n230), .CO(n256), .S(n255) );
  XNOR2_X1 U275 ( .A(n239), .B(\mult_x_1/n288 ), .ZN(n234) );
  OAI22_X1 U276 ( .A1(n235), .A2(n234), .B1(n243), .B2(n233), .ZN(n238) );
  XNOR2_X1 U277 ( .A(n647), .B(\mult_x_1/n286 ), .ZN(n242) );
  OAI22_X1 U278 ( .A1(n247), .A2(n242), .B1(n236), .B2(n474), .ZN(n237) );
  NOR2_X1 U279 ( .A1(n255), .A2(n254), .ZN(n295) );
  HA_X1 U280 ( .A(n238), .B(n237), .CO(n254), .S(n252) );
  OR2_X1 U281 ( .A1(\mult_x_1/n288 ), .A2(n471), .ZN(n240) );
  OAI22_X1 U282 ( .A1(n241), .A2(n471), .B1(n240), .B2(n243), .ZN(n251) );
  OR2_X1 U283 ( .A1(n252), .A2(n251), .ZN(n290) );
  XNOR2_X1 U284 ( .A(n647), .B(\mult_x_1/n287 ), .ZN(n246) );
  OAI22_X1 U285 ( .A1(n247), .A2(n246), .B1(n242), .B2(n474), .ZN(n250) );
  INV_X1 U286 ( .A(n243), .ZN(n244) );
  AND2_X1 U287 ( .A1(\mult_x_1/n288 ), .A2(n244), .ZN(n249) );
  NOR2_X1 U288 ( .A1(n250), .A2(n249), .ZN(n281) );
  OAI22_X1 U289 ( .A1(n247), .A2(\mult_x_1/n288 ), .B1(n246), .B2(n474), .ZN(
        n277) );
  OR2_X1 U290 ( .A1(\mult_x_1/n288 ), .A2(n473), .ZN(n248) );
  NAND2_X1 U291 ( .A1(n248), .A2(n247), .ZN(n276) );
  NAND2_X1 U292 ( .A1(n277), .A2(n276), .ZN(n284) );
  NAND2_X1 U293 ( .A1(n250), .A2(n249), .ZN(n282) );
  OAI21_X1 U294 ( .B1(n281), .B2(n284), .A(n282), .ZN(n291) );
  NAND2_X1 U295 ( .A1(n252), .A2(n251), .ZN(n289) );
  INV_X1 U296 ( .A(n289), .ZN(n253) );
  AOI21_X1 U297 ( .B1(n290), .B2(n291), .A(n253), .ZN(n298) );
  NAND2_X1 U298 ( .A1(n255), .A2(n254), .ZN(n296) );
  OAI21_X1 U299 ( .B1(n295), .B2(n298), .A(n296), .ZN(n304) );
  NAND2_X1 U300 ( .A1(n257), .A2(n256), .ZN(n302) );
  INV_X1 U301 ( .A(n302), .ZN(n258) );
  AOI21_X1 U302 ( .B1(n303), .B2(n304), .A(n258), .ZN(n259) );
  NAND2_X1 U303 ( .A1(n379), .A2(n259), .ZN(n260) );
  OAI21_X1 U304 ( .B1(n373), .B2(n441), .A(n260), .ZN(n439) );
  OR2_X1 U305 ( .A1(n377), .A2(n445), .ZN(n265) );
  NOR2_X1 U306 ( .A1(n262), .A2(n261), .ZN(n263) );
  NAND2_X1 U307 ( .A1(n213), .A2(n263), .ZN(n264) );
  NAND2_X1 U308 ( .A1(n265), .A2(n264), .ZN(n431) );
  INV_X1 U309 ( .A(n266), .ZN(n268) );
  NAND2_X1 U310 ( .A1(n268), .A2(n213), .ZN(n270) );
  OR2_X1 U311 ( .A1(n377), .A2(n443), .ZN(n269) );
  OAI21_X1 U312 ( .B1(n271), .B2(n270), .A(n269), .ZN(n435) );
  AOI22_X1 U313 ( .A1(n351), .A2(n519), .B1(n520), .B2(n380), .ZN(n522) );
  AOI22_X1 U314 ( .A1(n351), .A2(n518), .B1(n519), .B2(n380), .ZN(n524) );
  AND2_X1 U315 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n274) );
  NAND2_X1 U316 ( .A1(n377), .A2(n274), .ZN(n275) );
  OAI21_X1 U317 ( .B1(n379), .B2(n518), .A(n275), .ZN(n526) );
  AOI22_X1 U318 ( .A1(n351), .A2(n516), .B1(n517), .B2(n380), .ZN(n528) );
  AOI22_X1 U319 ( .A1(n351), .A2(n515), .B1(n516), .B2(n380), .ZN(n530) );
  INV_X2 U320 ( .A(n288), .ZN(n377) );
  OR2_X1 U321 ( .A1(n277), .A2(n276), .ZN(n278) );
  AND2_X1 U322 ( .A1(n278), .A2(n284), .ZN(n279) );
  NAND2_X1 U323 ( .A1(n377), .A2(n279), .ZN(n280) );
  OAI21_X1 U324 ( .B1(n377), .B2(n515), .A(n280), .ZN(n532) );
  AOI22_X1 U325 ( .A1(n351), .A2(n513), .B1(n514), .B2(n380), .ZN(n534) );
  AOI22_X1 U326 ( .A1(n351), .A2(n512), .B1(n513), .B2(n380), .ZN(n536) );
  INV_X1 U327 ( .A(n281), .ZN(n283) );
  NAND2_X1 U328 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U329 ( .A(n285), .B(n284), .Z(n286) );
  NAND2_X1 U330 ( .A1(n371), .A2(n286), .ZN(n287) );
  OAI21_X1 U331 ( .B1(n377), .B2(n512), .A(n287), .ZN(n538) );
  AOI22_X1 U332 ( .A1(n351), .A2(n510), .B1(n511), .B2(n380), .ZN(n540) );
  AOI22_X1 U333 ( .A1(n351), .A2(n509), .B1(n510), .B2(n380), .ZN(n542) );
  INV_X2 U334 ( .A(n288), .ZN(n373) );
  NAND2_X1 U335 ( .A1(n290), .A2(n289), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n293) );
  NAND2_X1 U337 ( .A1(n371), .A2(n293), .ZN(n294) );
  OAI21_X1 U338 ( .B1(n373), .B2(n509), .A(n294), .ZN(n544) );
  AOI22_X1 U339 ( .A1(n351), .A2(n507), .B1(n508), .B2(n380), .ZN(n546) );
  AOI22_X1 U340 ( .A1(n351), .A2(n506), .B1(n507), .B2(n380), .ZN(n548) );
  INV_X1 U341 ( .A(n295), .ZN(n297) );
  NAND2_X1 U342 ( .A1(n297), .A2(n296), .ZN(n299) );
  XOR2_X1 U343 ( .A(n299), .B(n298), .Z(n300) );
  NAND2_X1 U344 ( .A1(n371), .A2(n300), .ZN(n301) );
  OAI21_X1 U345 ( .B1(n377), .B2(n506), .A(n301), .ZN(n550) );
  AOI22_X1 U346 ( .A1(n351), .A2(n504), .B1(n505), .B2(n380), .ZN(n552) );
  AOI22_X1 U347 ( .A1(n379), .A2(n503), .B1(n504), .B2(n380), .ZN(n554) );
  NAND2_X1 U348 ( .A1(n303), .A2(n302), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n306) );
  NAND2_X1 U350 ( .A1(n306), .A2(n371), .ZN(n307) );
  OAI21_X1 U351 ( .B1(n377), .B2(n503), .A(n307), .ZN(n556) );
  AOI22_X1 U352 ( .A1(n379), .A2(n501), .B1(n502), .B2(n380), .ZN(n558) );
  NAND2_X1 U353 ( .A1(n451), .A2(n391), .ZN(n308) );
  XOR2_X1 U354 ( .A(n308), .B(n400), .Z(n309) );
  NAND2_X1 U355 ( .A1(n371), .A2(n309), .ZN(n310) );
  OAI21_X1 U356 ( .B1(n373), .B2(n501), .A(n310), .ZN(n560) );
  AOI22_X1 U357 ( .A1(n379), .A2(n499), .B1(n500), .B2(n380), .ZN(n562) );
  OAI21_X1 U358 ( .B1(n390), .B2(n400), .A(n391), .ZN(n314) );
  NAND2_X1 U359 ( .A1(n383), .A2(n389), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n314), .B(n311), .ZN(n312) );
  NAND2_X1 U361 ( .A1(n371), .A2(n312), .ZN(n313) );
  OAI21_X1 U362 ( .B1(n377), .B2(n499), .A(n313), .ZN(n564) );
  AOI22_X1 U363 ( .A1(n379), .A2(n497), .B1(n498), .B2(n380), .ZN(n566) );
  AOI21_X1 U364 ( .B1(n314), .B2(n383), .A(n452), .ZN(n318) );
  NAND2_X1 U365 ( .A1(n454), .A2(n388), .ZN(n315) );
  XOR2_X1 U366 ( .A(n318), .B(n315), .Z(n316) );
  NAND2_X1 U367 ( .A1(n377), .A2(n316), .ZN(n317) );
  OAI21_X1 U368 ( .B1(n377), .B2(n497), .A(n317), .ZN(n568) );
  AOI22_X1 U369 ( .A1(n379), .A2(n495), .B1(n496), .B2(n380), .ZN(n570) );
  OAI21_X1 U370 ( .B1(n318), .B2(n387), .A(n388), .ZN(n328) );
  INV_X1 U371 ( .A(n328), .ZN(n322) );
  NAND2_X1 U372 ( .A1(n445), .A2(n386), .ZN(n319) );
  XOR2_X1 U373 ( .A(n322), .B(n319), .Z(n320) );
  NAND2_X1 U374 ( .A1(n377), .A2(n320), .ZN(n321) );
  OAI21_X1 U375 ( .B1(n377), .B2(n495), .A(n321), .ZN(n572) );
  AOI22_X1 U376 ( .A1(n379), .A2(n493), .B1(n494), .B2(n380), .ZN(n574) );
  OAI21_X1 U377 ( .B1(n322), .B2(n396), .A(n386), .ZN(n324) );
  NAND2_X1 U378 ( .A1(n449), .A2(n393), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  NAND2_X1 U380 ( .A1(n377), .A2(n325), .ZN(n326) );
  OAI21_X1 U381 ( .B1(n373), .B2(n493), .A(n326), .ZN(n576) );
  AOI22_X1 U382 ( .A1(n379), .A2(n491), .B1(n492), .B2(n380), .ZN(n578) );
  NOR2_X1 U383 ( .A1(n392), .A2(n396), .ZN(n329) );
  OAI21_X1 U384 ( .B1(n392), .B2(n386), .A(n393), .ZN(n327) );
  AOI21_X1 U385 ( .B1(n329), .B2(n328), .A(n327), .ZN(n356) );
  NAND2_X1 U386 ( .A1(n443), .A2(n399), .ZN(n330) );
  XOR2_X1 U387 ( .A(n356), .B(n330), .Z(n331) );
  NAND2_X1 U388 ( .A1(n377), .A2(n331), .ZN(n332) );
  OAI21_X1 U389 ( .B1(n373), .B2(n491), .A(n332), .ZN(n580) );
  AOI22_X1 U390 ( .A1(n351), .A2(n489), .B1(n490), .B2(n380), .ZN(n582) );
  OAI21_X1 U391 ( .B1(n356), .B2(n398), .A(n399), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n397), .A2(n395), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  NAND2_X1 U394 ( .A1(n377), .A2(n335), .ZN(n336) );
  OAI21_X1 U395 ( .B1(n373), .B2(n489), .A(n336), .ZN(n584) );
  AOI22_X1 U396 ( .A1(n379), .A2(n487), .B1(n488), .B2(n380), .ZN(n586) );
  NAND2_X1 U397 ( .A1(n443), .A2(n397), .ZN(n338) );
  AOI21_X1 U398 ( .B1(n442), .B2(n397), .A(n446), .ZN(n337) );
  OAI21_X1 U399 ( .B1(n356), .B2(n338), .A(n337), .ZN(n340) );
  NAND2_X1 U400 ( .A1(n382), .A2(n394), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  NAND2_X1 U402 ( .A1(n377), .A2(n341), .ZN(n342) );
  OAI21_X1 U403 ( .B1(n373), .B2(n487), .A(n342), .ZN(n588) );
  AOI22_X1 U404 ( .A1(n351), .A2(n485), .B1(n486), .B2(n380), .ZN(n590) );
  NAND2_X1 U405 ( .A1(n397), .A2(n382), .ZN(n344) );
  NOR2_X1 U406 ( .A1(n398), .A2(n344), .ZN(n352) );
  INV_X1 U407 ( .A(n352), .ZN(n346) );
  AOI21_X1 U408 ( .B1(n446), .B2(n382), .A(n447), .ZN(n343) );
  OAI21_X1 U409 ( .B1(n344), .B2(n399), .A(n343), .ZN(n353) );
  INV_X1 U410 ( .A(n353), .ZN(n345) );
  OAI21_X1 U411 ( .B1(n356), .B2(n346), .A(n345), .ZN(n348) );
  NAND2_X1 U412 ( .A1(n381), .A2(n385), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  NAND2_X1 U414 ( .A1(n377), .A2(n349), .ZN(n350) );
  OAI21_X1 U415 ( .B1(n373), .B2(n485), .A(n350), .ZN(n592) );
  AOI22_X1 U416 ( .A1(n351), .A2(n483), .B1(n484), .B2(n380), .ZN(n594) );
  NAND2_X1 U417 ( .A1(n352), .A2(n381), .ZN(n355) );
  AOI21_X1 U418 ( .B1(n353), .B2(n381), .A(n456), .ZN(n354) );
  OAI21_X1 U419 ( .B1(n356), .B2(n355), .A(n354), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n357), .B(n384), .ZN(n358) );
  NAND2_X1 U421 ( .A1(n377), .A2(n358), .ZN(n359) );
  OAI21_X1 U422 ( .B1(n373), .B2(n483), .A(n359), .ZN(n596) );
  NAND2_X1 U423 ( .A1(n371), .A2(B_extended[0]), .ZN(n360) );
  OAI21_X1 U424 ( .B1(n373), .B2(n482), .A(n360), .ZN(n598) );
  NAND2_X1 U425 ( .A1(n377), .A2(B_extended[1]), .ZN(n361) );
  OAI21_X1 U426 ( .B1(n373), .B2(n481), .A(n361), .ZN(n600) );
  NAND2_X1 U427 ( .A1(n371), .A2(B_extended[2]), .ZN(n362) );
  OAI21_X1 U428 ( .B1(n373), .B2(n480), .A(n362), .ZN(n602) );
  NAND2_X1 U429 ( .A1(n371), .A2(B_extended[3]), .ZN(n363) );
  OAI21_X1 U430 ( .B1(n373), .B2(n479), .A(n363), .ZN(n604) );
  NAND2_X1 U431 ( .A1(n371), .A2(B_extended[4]), .ZN(n364) );
  OAI21_X1 U432 ( .B1(n373), .B2(n478), .A(n364), .ZN(n606) );
  NAND2_X1 U433 ( .A1(n371), .A2(B_extended[5]), .ZN(n365) );
  OAI21_X1 U434 ( .B1(n373), .B2(n477), .A(n365), .ZN(n608) );
  NAND2_X1 U435 ( .A1(n371), .A2(B_extended[6]), .ZN(n366) );
  OAI21_X1 U436 ( .B1(n373), .B2(n476), .A(n366), .ZN(n610) );
  NAND2_X1 U437 ( .A1(n371), .A2(B_extended[7]), .ZN(n367) );
  OAI21_X1 U438 ( .B1(n379), .B2(n475), .A(n367), .ZN(n612) );
  NAND2_X1 U439 ( .A1(n371), .A2(A_extended[0]), .ZN(n368) );
  OAI21_X1 U440 ( .B1(n379), .B2(n474), .A(n368), .ZN(n614) );
  NAND2_X1 U441 ( .A1(n371), .A2(A_extended[1]), .ZN(n369) );
  OAI21_X1 U442 ( .B1(n379), .B2(n473), .A(n369), .ZN(n616) );
  NAND2_X1 U443 ( .A1(n371), .A2(A_extended[2]), .ZN(n370) );
  OAI21_X1 U444 ( .B1(n373), .B2(n472), .A(n370), .ZN(n618) );
  NAND2_X1 U445 ( .A1(n371), .A2(A_extended[3]), .ZN(n372) );
  OAI21_X1 U446 ( .B1(n373), .B2(n471), .A(n372), .ZN(n620) );
  NAND2_X1 U447 ( .A1(n377), .A2(A_extended[4]), .ZN(n374) );
  OAI21_X1 U448 ( .B1(n379), .B2(n470), .A(n374), .ZN(n622) );
  NAND2_X1 U449 ( .A1(n377), .A2(A_extended[5]), .ZN(n375) );
  OAI21_X1 U450 ( .B1(n379), .B2(n469), .A(n375), .ZN(n624) );
  NAND2_X1 U451 ( .A1(n373), .A2(A_extended[6]), .ZN(n376) );
  OAI21_X1 U452 ( .B1(n379), .B2(n468), .A(n376), .ZN(n626) );
  NAND2_X1 U453 ( .A1(n377), .A2(A_extended[7]), .ZN(n378) );
  OAI21_X1 U454 ( .B1(n379), .B2(n467), .A(n378), .ZN(n628) );
  NAND2_X1 U455 ( .A1(n466), .A2(n380), .ZN(n630) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_27 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n397, n399, n401, n403, n405, n407, n409, n411,
         n413, n415, n417, n419, n421, n423, n425, n427, n429, n431, n433,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n514, n516, n518, n520, n522, n524, n526, n528, n530, n532,
         n534, n536, n538, n540, n542, n544, n546, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n567, n569, n571, n573, n575,
         n577, n579, n581, n583, n585, n587, n589, n591, n593, n595, n597,
         n599, n601, n603, n605, n607, n609, n611, n613, n615, n617, n619,
         n621, n638, n639, n640;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n457), .SE(n621), .CK(clk), .Q(n639), 
        .QN(n458) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n457), .SE(n617), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n460) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n457), .SE(n615), .CK(clk), .Q(n638), 
        .QN(n461) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n457), .SE(n609), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n464) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n457), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n466) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n457), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n467) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n457), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n468) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n456), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n469) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n456), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n470) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n456), .SE(n595), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n471) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n456), .SE(n593), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n472) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n456), .SE(n591), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n473) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n456), .SE(n589), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n474) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n456), .SE(n587), .CK(clk), .QN(n475)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n456), .SE(n585), .CK(clk), .Q(
        product[15]), .QN(n476) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n456), .SE(n583), .CK(clk), .QN(n477)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n456), .SE(n581), .CK(clk), .Q(
        product[14]), .QN(n478) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n456), .SE(n579), .CK(clk), .QN(n479)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n455), .SE(n577), .CK(clk), .Q(
        product[13]), .QN(n480) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n455), .SE(n575), .CK(clk), .QN(n481)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n455), .SE(n573), .CK(clk), .Q(
        product[12]), .QN(n482) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n455), .SE(n571), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n455), .SE(n569), .CK(clk), .Q(
        product[11]), .QN(n484) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n455), .SE(n567), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n455), .SE(n565), .CK(clk), .Q(
        product[10]), .QN(n486) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n455), .SE(n563), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n455), .SE(n561), .CK(clk), .Q(
        product[9]), .QN(n488) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n455), .SE(n559), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n455), .SE(n557), .CK(clk), .Q(
        product[8]), .QN(n490) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n454), .SE(n555), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n454), .SE(n553), .CK(clk), .Q(
        product[7]), .QN(n492) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n454), .SE(n551), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n454), .SE(n549), .CK(clk), .Q(
        product[6]), .QN(n494) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n454), .SE(n546), .CK(clk), .QN(n496)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n454), .SE(n544), .CK(clk), .Q(
        product[5]), .QN(n497) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n454), .SE(n542), .CK(clk), .QN(n498)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n454), .SE(n540), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n454), .SE(n538), .CK(clk), .Q(
        product[4]), .QN(n500) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n454), .SE(n536), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n453), .SE(n534), .CK(clk), .QN(n502)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n453), .SE(n532), .CK(clk), .Q(
        product[3]), .QN(n503) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n453), .SE(n530), .CK(clk), .QN(n504)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n453), .SE(n528), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n453), .SE(n526), .CK(clk), .Q(
        product[2]), .QN(n506) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n453), .SE(n524), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n453), .SE(n522), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n453), .SE(n520), .CK(clk), .Q(
        product[1]), .QN(n509) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n453), .SE(n518), .CK(clk), .QN(n510)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n453), .SE(n516), .CK(clk), .QN(n511)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n453), .SE(n514), .CK(clk), .Q(
        product[0]), .QN(n512) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n457), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n465) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n640), .SI(1'b1), .SE(n433), .CK(clk), 
        .Q(n394), .QN(n435) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n640), .SI(1'b1), .SE(n431), .CK(clk), 
        .Q(n393), .QN(n436) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n640), .SI(1'b1), .SE(n429), .CK(clk), 
        .Q(n392), .QN(n437) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n640), .SE(n427), .CK(
        clk), .QN(n376) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n640), .SE(n425), .CK(
        clk), .Q(n438), .QN(n375) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n640), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n391), .QN(n439) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n640), .SI(1'b1), .SE(n421), .CK(clk), 
        .Q(n390), .QN(n440) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n640), .SI(1'b1), .SE(n419), .CK(clk), 
        .Q(n389), .QN(n441) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n640), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n388), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n640), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n387), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n640), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n377) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n640), .SI(1'b1), .SE(n411), .CK(clk), 
        .Q(n386), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n640), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n385), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n640), .SE(n407), .CK(
        clk), .Q(n446), .QN(n384) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n640), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n383), .QN(n447) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n640), .SE(n403), .CK(
        clk), .Q(n448), .QN(n382) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n640), .SE(n401), .CK(
        clk), .Q(n449), .QN(n381) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n640), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n380), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n640), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n379), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n640), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n378), .QN(n452) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n457), .SE(n619), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n459) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n457), .SE(n611), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n463) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n454), .SE(n547), .CK(clk), .Q(n23), 
        .QN(n495) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n457), .SE(n613), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n462) );
  BUF_X1 U2 ( .A(n638), .Z(n141) );
  OR2_X1 U3 ( .A1(\mult_x_1/n180 ), .A2(n465), .ZN(n181) );
  BUF_X1 U4 ( .A(\mult_x_1/n313 ), .Z(n143) );
  CLKBUF_X1 U5 ( .A(n276), .Z(n454) );
  CLKBUF_X1 U6 ( .A(n276), .Z(n455) );
  CLKBUF_X1 U7 ( .A(n276), .Z(n456) );
  CLKBUF_X1 U8 ( .A(n276), .Z(n457) );
  CLKBUF_X1 U9 ( .A(n276), .Z(n453) );
  INV_X1 U10 ( .A(rst_n), .ZN(n640) );
  BUF_X1 U11 ( .A(n96), .Z(n209) );
  OR2_X1 U12 ( .A1(n11), .A2(n95), .ZN(n84) );
  INV_X1 U13 ( .A(n459), .ZN(n5) );
  INV_X1 U14 ( .A(n459), .ZN(n155) );
  OR2_X1 U15 ( .A1(n269), .A2(n451), .ZN(n6) );
  NAND2_X1 U16 ( .A1(n6), .A2(n178), .ZN(n397) );
  OR2_X2 U17 ( .A1(n25), .A2(n26), .ZN(n7) );
  OR2_X1 U18 ( .A1(n25), .A2(n26), .ZN(n196) );
  CLKBUF_X1 U19 ( .A(\mult_x_1/n312 ), .Z(n16) );
  INV_X1 U20 ( .A(n207), .ZN(n8) );
  XOR2_X1 U21 ( .A(n156), .B(n461), .Z(n159) );
  CLKBUF_X1 U22 ( .A(n207), .Z(n9) );
  INV_X2 U23 ( .A(n17), .ZN(n14) );
  BUF_X1 U24 ( .A(\mult_x_1/n313 ), .Z(n10) );
  AND2_X1 U25 ( .A1(n181), .A2(n466), .ZN(n11) );
  BUF_X1 U26 ( .A(n83), .Z(n146) );
  NAND2_X1 U27 ( .A1(n77), .A2(n71), .ZN(n73) );
  OR2_X1 U28 ( .A1(n75), .A2(n74), .ZN(n71) );
  NAND2_X1 U29 ( .A1(n75), .A2(n74), .ZN(n72) );
  XNOR2_X1 U30 ( .A(n20), .B(n137), .ZN(n154) );
  XNOR2_X1 U31 ( .A(n136), .B(n135), .ZN(n137) );
  CLKBUF_X1 U32 ( .A(n207), .Z(n12) );
  INV_X1 U33 ( .A(n135), .ZN(n111) );
  INV_X1 U34 ( .A(n136), .ZN(n112) );
  XNOR2_X1 U35 ( .A(n243), .B(n31), .ZN(n35) );
  XNOR2_X1 U36 ( .A(n245), .B(n244), .ZN(n31) );
  NAND2_X1 U37 ( .A1(n19), .A2(n124), .ZN(n125) );
  NAND2_X1 U38 ( .A1(n247), .A2(n246), .ZN(n250) );
  NAND2_X1 U39 ( .A1(n245), .A2(n244), .ZN(n246) );
  NAND2_X1 U40 ( .A1(n243), .A2(n21), .ZN(n247) );
  NAND2_X1 U41 ( .A1(n115), .A2(n114), .ZN(n130) );
  NAND2_X1 U42 ( .A1(n136), .A2(n135), .ZN(n114) );
  NAND2_X1 U43 ( .A1(n20), .A2(n113), .ZN(n115) );
  NAND2_X1 U44 ( .A1(n112), .A2(n111), .ZN(n113) );
  NAND2_X1 U45 ( .A1(n73), .A2(n72), .ZN(n174) );
  INV_X1 U46 ( .A(n640), .ZN(n276) );
  OAI22_X1 U47 ( .A1(n154), .A2(n24), .B1(n271), .B2(n444), .ZN(n411) );
  OAI22_X1 U48 ( .A1(n83), .A2(n82), .B1(n66), .B2(n183), .ZN(n13) );
  XNOR2_X1 U49 ( .A(n161), .B(n15), .ZN(n176) );
  XNOR2_X1 U50 ( .A(n163), .B(n162), .ZN(n15) );
  INV_X1 U51 ( .A(n17), .ZN(n183) );
  AND2_X1 U52 ( .A1(n639), .A2(\mult_x_1/n281 ), .ZN(n156) );
  INV_X1 U53 ( .A(n64), .ZN(n207) );
  XOR2_X1 U54 ( .A(n10), .B(\mult_x_1/a[2] ), .Z(n17) );
  XNOR2_X1 U55 ( .A(n463), .B(\mult_x_1/a[4] ), .ZN(n18) );
  XNOR2_X1 U56 ( .A(n462), .B(n461), .ZN(n25) );
  INV_X1 U57 ( .A(en), .ZN(n311) );
  BUF_X2 U58 ( .A(en), .Z(n269) );
  INV_X1 U59 ( .A(n311), .ZN(n372) );
  INV_X2 U60 ( .A(en), .ZN(n307) );
  AND2_X1 U61 ( .A1(n103), .A2(n102), .ZN(n19) );
  XOR2_X1 U62 ( .A(n103), .B(n102), .Z(n20) );
  OR2_X1 U63 ( .A1(n245), .A2(n244), .ZN(n21) );
  OR2_X1 U64 ( .A1(n19), .A2(n124), .ZN(n22) );
  OR2_X1 U65 ( .A1(n153), .A2(n307), .ZN(n24) );
  XNOR2_X1 U67 ( .A(n463), .B(\mult_x_1/a[4] ), .ZN(n26) );
  OR2_X1 U68 ( .A1(\mult_x_1/n288 ), .A2(n461), .ZN(n27) );
  INV_X1 U69 ( .A(n18), .ZN(n194) );
  OAI22_X1 U70 ( .A1(n7), .A2(n461), .B1(n27), .B2(n194), .ZN(n192) );
  XNOR2_X1 U71 ( .A(n141), .B(\mult_x_1/n288 ), .ZN(n28) );
  XNOR2_X1 U72 ( .A(n141), .B(\mult_x_1/n287 ), .ZN(n195) );
  OAI22_X1 U73 ( .A1(n7), .A2(n28), .B1(n194), .B2(n195), .ZN(n191) );
  XOR2_X1 U74 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n29) );
  XNOR2_X1 U75 ( .A(n10), .B(\mult_x_1/a[2] ), .ZN(n30) );
  NAND2_X1 U76 ( .A1(n29), .A2(n30), .ZN(n83) );
  XNOR2_X1 U77 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n33) );
  XNOR2_X1 U78 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n184) );
  OAI22_X1 U79 ( .A1(n146), .A2(n33), .B1(n14), .B2(n184), .ZN(n245) );
  XNOR2_X1 U80 ( .A(n143), .B(\mult_x_1/n284 ), .ZN(n32) );
  XNOR2_X1 U81 ( .A(n143), .B(\mult_x_1/n283 ), .ZN(n180) );
  OAI22_X1 U82 ( .A1(n181), .A2(n32), .B1(n180), .B2(n466), .ZN(n244) );
  XNOR2_X1 U83 ( .A(n143), .B(\mult_x_1/n285 ), .ZN(n41) );
  OAI22_X1 U84 ( .A1(n181), .A2(n41), .B1(n32), .B2(n466), .ZN(n38) );
  AND2_X1 U85 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n37) );
  XNOR2_X1 U86 ( .A(n16), .B(\mult_x_1/n287 ), .ZN(n39) );
  OAI22_X1 U87 ( .A1(n146), .A2(n39), .B1(n14), .B2(n33), .ZN(n36) );
  OR2_X1 U88 ( .A1(n35), .A2(n34), .ZN(n266) );
  NAND2_X1 U89 ( .A1(n35), .A2(n34), .ZN(n263) );
  NAND2_X1 U90 ( .A1(n266), .A2(n263), .ZN(n56) );
  FA_X1 U91 ( .A(n38), .B(n37), .CI(n36), .CO(n34), .S(n55) );
  XNOR2_X1 U92 ( .A(n16), .B(\mult_x_1/n288 ), .ZN(n40) );
  OAI22_X1 U93 ( .A1(n146), .A2(n40), .B1(n14), .B2(n39), .ZN(n43) );
  XNOR2_X1 U94 ( .A(n143), .B(\mult_x_1/n286 ), .ZN(n45) );
  OAI22_X1 U95 ( .A1(n181), .A2(n45), .B1(n41), .B2(n466), .ZN(n42) );
  NOR2_X1 U96 ( .A1(n55), .A2(n54), .ZN(n297) );
  HA_X1 U97 ( .A(n43), .B(n42), .CO(n54), .S(n52) );
  OR2_X1 U98 ( .A1(\mult_x_1/n288 ), .A2(n463), .ZN(n44) );
  OAI22_X1 U99 ( .A1(n146), .A2(n463), .B1(n44), .B2(n14), .ZN(n51) );
  OR2_X1 U100 ( .A1(n52), .A2(n51), .ZN(n292) );
  XNOR2_X1 U101 ( .A(n143), .B(\mult_x_1/n287 ), .ZN(n47) );
  OAI22_X1 U102 ( .A1(n181), .A2(n47), .B1(n45), .B2(n466), .ZN(n50) );
  INV_X1 U103 ( .A(n14), .ZN(n46) );
  AND2_X1 U104 ( .A1(\mult_x_1/n288 ), .A2(n46), .ZN(n49) );
  NOR2_X1 U105 ( .A1(n50), .A2(n49), .ZN(n284) );
  OAI22_X1 U106 ( .A1(n181), .A2(\mult_x_1/n288 ), .B1(n47), .B2(n466), .ZN(
        n280) );
  OR2_X1 U107 ( .A1(\mult_x_1/n288 ), .A2(n465), .ZN(n48) );
  NAND2_X1 U108 ( .A1(n48), .A2(n181), .ZN(n279) );
  NAND2_X1 U109 ( .A1(n280), .A2(n279), .ZN(n287) );
  NAND2_X1 U110 ( .A1(n50), .A2(n49), .ZN(n285) );
  OAI21_X1 U111 ( .B1(n284), .B2(n287), .A(n285), .ZN(n293) );
  NAND2_X1 U112 ( .A1(n52), .A2(n51), .ZN(n291) );
  INV_X1 U113 ( .A(n291), .ZN(n53) );
  AOI21_X1 U114 ( .B1(n292), .B2(n293), .A(n53), .ZN(n300) );
  NAND2_X1 U115 ( .A1(n55), .A2(n54), .ZN(n298) );
  OAI21_X1 U116 ( .B1(n297), .B2(n300), .A(n298), .ZN(n265) );
  XNOR2_X1 U117 ( .A(n56), .B(n265), .ZN(n57) );
  NAND2_X1 U118 ( .A1(n57), .A2(n271), .ZN(n59) );
  NAND2_X1 U119 ( .A1(n307), .A2(n23), .ZN(n58) );
  NAND2_X1 U120 ( .A1(n59), .A2(n58), .ZN(n547) );
  XNOR2_X1 U121 ( .A(n141), .B(\mult_x_1/n281 ), .ZN(n69) );
  OR2_X1 U122 ( .A1(n196), .A2(n69), .ZN(n61) );
  OR2_X1 U123 ( .A1(n159), .A2(n194), .ZN(n60) );
  NAND2_X1 U124 ( .A1(n61), .A2(n60), .ZN(n167) );
  INV_X1 U125 ( .A(n167), .ZN(n161) );
  AND2_X1 U126 ( .A1(n639), .A2(\mult_x_1/n310 ), .ZN(n62) );
  XNOR2_X1 U127 ( .A(n62), .B(\mult_x_1/n310 ), .ZN(n96) );
  NOR2_X1 U128 ( .A1(n470), .A2(n209), .ZN(n163) );
  XNOR2_X1 U129 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/a[6] ), .ZN(n63) );
  XOR2_X1 U130 ( .A(\mult_x_1/a[6] ), .B(n638), .Z(n64) );
  OR2_X2 U131 ( .A1(n64), .A2(n63), .ZN(n206) );
  XNOR2_X1 U132 ( .A(n5), .B(\mult_x_1/n283 ), .ZN(n65) );
  XNOR2_X1 U133 ( .A(n155), .B(\mult_x_1/n282 ), .ZN(n158) );
  OAI22_X1 U134 ( .A1(n206), .A2(n65), .B1(n207), .B2(n158), .ZN(n162) );
  XNOR2_X1 U135 ( .A(n155), .B(\mult_x_1/n284 ), .ZN(n68) );
  OAI22_X1 U136 ( .A1(n206), .A2(n68), .B1(n12), .B2(n65), .ZN(n80) );
  XNOR2_X1 U137 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n82) );
  XNOR2_X1 U138 ( .A(n156), .B(\mult_x_1/n312 ), .ZN(n66) );
  OAI22_X1 U139 ( .A1(n83), .A2(n82), .B1(n66), .B2(n183), .ZN(n79) );
  CLKBUF_X1 U140 ( .A(n83), .Z(n185) );
  AOI21_X1 U141 ( .B1(n14), .B2(n185), .A(n66), .ZN(n67) );
  INV_X1 U142 ( .A(n67), .ZN(n78) );
  XNOR2_X1 U143 ( .A(n155), .B(\mult_x_1/n285 ), .ZN(n85) );
  OAI22_X1 U144 ( .A1(n206), .A2(n85), .B1(n207), .B2(n68), .ZN(n100) );
  XNOR2_X1 U145 ( .A(n141), .B(\mult_x_1/n283 ), .ZN(n81) );
  XNOR2_X1 U146 ( .A(n141), .B(\mult_x_1/n282 ), .ZN(n70) );
  OAI22_X1 U147 ( .A1(n7), .A2(n81), .B1(n194), .B2(n70), .ZN(n99) );
  INV_X1 U148 ( .A(n79), .ZN(n98) );
  NOR2_X1 U149 ( .A1(n471), .A2(n209), .ZN(n75) );
  OAI22_X1 U150 ( .A1(n7), .A2(n70), .B1(n194), .B2(n69), .ZN(n74) );
  XNOR2_X1 U151 ( .A(n75), .B(n74), .ZN(n76) );
  XNOR2_X1 U152 ( .A(n77), .B(n76), .ZN(n122) );
  FA_X1 U153 ( .A(n80), .B(n13), .CI(n78), .CO(n175), .S(n121) );
  XNOR2_X1 U154 ( .A(n141), .B(\mult_x_1/n284 ), .ZN(n106) );
  OAI22_X1 U155 ( .A1(n7), .A2(n106), .B1(n194), .B2(n81), .ZN(n93) );
  XNOR2_X1 U156 ( .A(n16), .B(\mult_x_1/n282 ), .ZN(n107) );
  OAI22_X1 U157 ( .A1(n83), .A2(n107), .B1(n14), .B2(n82), .ZN(n92) );
  OR2_X1 U158 ( .A1(n93), .A2(n92), .ZN(n91) );
  NOR2_X1 U159 ( .A1(n472), .A2(n209), .ZN(n90) );
  XNOR2_X1 U160 ( .A(n156), .B(n143), .ZN(n95) );
  XNOR2_X1 U161 ( .A(n155), .B(\mult_x_1/n286 ), .ZN(n94) );
  OAI22_X1 U162 ( .A1(n206), .A2(n94), .B1(n207), .B2(n85), .ZN(n105) );
  NOR2_X1 U163 ( .A1(n473), .A2(n96), .ZN(n104) );
  OR2_X1 U164 ( .A1(n255), .A2(n254), .ZN(n86) );
  BUF_X1 U165 ( .A(en), .Z(n271) );
  NAND2_X1 U166 ( .A1(n86), .A2(n271), .ZN(n88) );
  OR2_X1 U167 ( .A1(n271), .A2(n450), .ZN(n87) );
  NAND2_X1 U168 ( .A1(n88), .A2(n87), .ZN(n399) );
  FA_X1 U169 ( .A(n91), .B(n90), .CI(n89), .CO(n120), .S(n123) );
  XNOR2_X1 U170 ( .A(n93), .B(n92), .ZN(n103) );
  XNOR2_X1 U171 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n109) );
  OAI22_X1 U172 ( .A1(n206), .A2(n109), .B1(n9), .B2(n94), .ZN(n140) );
  XNOR2_X1 U173 ( .A(n143), .B(\mult_x_1/n281 ), .ZN(n144) );
  OAI22_X1 U174 ( .A1(n181), .A2(n144), .B1(n95), .B2(n466), .ZN(n139) );
  INV_X1 U175 ( .A(n96), .ZN(n97) );
  AND2_X1 U176 ( .A1(\mult_x_1/n288 ), .A2(n97), .ZN(n138) );
  FA_X1 U177 ( .A(n99), .B(n100), .CI(n98), .CO(n77), .S(n124) );
  XNOR2_X1 U178 ( .A(n19), .B(n124), .ZN(n101) );
  XNOR2_X1 U179 ( .A(n123), .B(n101), .ZN(n131) );
  INV_X1 U180 ( .A(n131), .ZN(n117) );
  FA_X1 U181 ( .A(n84), .B(n105), .CI(n104), .CO(n89), .S(n136) );
  XNOR2_X1 U182 ( .A(n141), .B(\mult_x_1/n285 ), .ZN(n142) );
  OAI22_X1 U183 ( .A1(n7), .A2(n142), .B1(n194), .B2(n106), .ZN(n149) );
  XNOR2_X1 U184 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n145) );
  OAI22_X1 U185 ( .A1(n185), .A2(n145), .B1(n14), .B2(n107), .ZN(n148) );
  OR2_X1 U186 ( .A1(\mult_x_1/n288 ), .A2(n459), .ZN(n108) );
  OAI22_X1 U187 ( .A1(n206), .A2(n459), .B1(n108), .B2(n207), .ZN(n187) );
  XNOR2_X1 U188 ( .A(n155), .B(\mult_x_1/n288 ), .ZN(n110) );
  OAI22_X1 U189 ( .A1(n206), .A2(n110), .B1(n207), .B2(n109), .ZN(n186) );
  BUF_X1 U190 ( .A(en), .Z(n261) );
  NOR2_X1 U191 ( .A1(n130), .A2(n307), .ZN(n116) );
  NAND2_X1 U192 ( .A1(n117), .A2(n116), .ZN(n119) );
  NAND2_X1 U193 ( .A1(n307), .A2(n375), .ZN(n118) );
  NAND2_X1 U194 ( .A1(n119), .A2(n118), .ZN(n425) );
  FA_X1 U195 ( .A(n122), .B(n121), .CI(n120), .CO(n254), .S(n275) );
  NAND2_X1 U196 ( .A1(n123), .A2(n22), .ZN(n126) );
  NAND2_X1 U197 ( .A1(n126), .A2(n125), .ZN(n270) );
  NAND2_X1 U198 ( .A1(n275), .A2(n270), .ZN(n127) );
  NAND2_X1 U199 ( .A1(n127), .A2(n269), .ZN(n129) );
  NAND2_X1 U200 ( .A1(n307), .A2(n385), .ZN(n128) );
  NAND2_X1 U201 ( .A1(n129), .A2(n128), .ZN(n409) );
  NAND2_X1 U202 ( .A1(n131), .A2(n130), .ZN(n132) );
  NAND2_X1 U203 ( .A1(n132), .A2(n261), .ZN(n134) );
  BUF_X1 U204 ( .A(en), .Z(n273) );
  NAND2_X1 U205 ( .A1(n307), .A2(n376), .ZN(n133) );
  NAND2_X1 U206 ( .A1(n134), .A2(n133), .ZN(n427) );
  FA_X1 U207 ( .A(n140), .B(n139), .CI(n138), .CO(n102), .S(n226) );
  XNOR2_X1 U208 ( .A(n141), .B(\mult_x_1/n286 ), .ZN(n193) );
  OAI22_X1 U209 ( .A1(n7), .A2(n193), .B1(n194), .B2(n142), .ZN(n190) );
  XNOR2_X1 U210 ( .A(n143), .B(\mult_x_1/n282 ), .ZN(n179) );
  OAI22_X1 U211 ( .A1(n181), .A2(n179), .B1(n144), .B2(n466), .ZN(n189) );
  XNOR2_X1 U212 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n182) );
  OAI22_X1 U213 ( .A1(n146), .A2(n182), .B1(n14), .B2(n145), .ZN(n188) );
  FA_X1 U214 ( .A(n149), .B(n148), .CI(n147), .CO(n135), .S(n224) );
  NAND2_X1 U215 ( .A1(n154), .A2(n153), .ZN(n150) );
  NAND2_X1 U216 ( .A1(n150), .A2(n261), .ZN(n152) );
  NAND2_X1 U217 ( .A1(n307), .A2(n377), .ZN(n151) );
  NAND2_X1 U218 ( .A1(n152), .A2(n151), .ZN(n413) );
  NOR2_X1 U239 ( .A1(n468), .A2(n209), .ZN(n204) );
  XNOR2_X1 U240 ( .A(n5), .B(\mult_x_1/n281 ), .ZN(n157) );
  XNOR2_X1 U241 ( .A(n156), .B(n5), .ZN(n205) );
  OAI22_X1 U242 ( .A1(n206), .A2(n157), .B1(n205), .B2(n12), .ZN(n213) );
  INV_X1 U243 ( .A(n213), .ZN(n203) );
  OAI22_X1 U244 ( .A1(n206), .A2(n158), .B1(n9), .B2(n157), .ZN(n169) );
  AOI21_X1 U245 ( .B1(n194), .B2(n196), .A(n159), .ZN(n160) );
  INV_X1 U246 ( .A(n160), .ZN(n168) );
  NAND2_X1 U247 ( .A1(n161), .A2(n163), .ZN(n166) );
  NAND2_X1 U248 ( .A1(n161), .A2(n162), .ZN(n165) );
  NAND2_X1 U249 ( .A1(n163), .A2(n162), .ZN(n164) );
  NAND3_X1 U250 ( .A1(n166), .A2(n165), .A3(n164), .ZN(n173) );
  NOR2_X1 U251 ( .A1(n469), .A2(n209), .ZN(n172) );
  FA_X1 U252 ( .A(n169), .B(n168), .CI(n167), .CO(n202), .S(n171) );
  OAI21_X1 U253 ( .B1(n221), .B2(n220), .A(n273), .ZN(n170) );
  OAI21_X1 U254 ( .B1(n273), .B2(n452), .A(n170), .ZN(n395) );
  FA_X1 U255 ( .A(n173), .B(n172), .CI(n171), .CO(n220), .S(n259) );
  FA_X1 U256 ( .A(n176), .B(n175), .CI(n174), .CO(n258), .S(n255) );
  OR2_X1 U257 ( .A1(n259), .A2(n258), .ZN(n177) );
  NAND2_X1 U258 ( .A1(n271), .A2(n177), .ZN(n178) );
  OAI22_X1 U259 ( .A1(n181), .A2(n180), .B1(n179), .B2(n466), .ZN(n199) );
  AND2_X1 U260 ( .A1(\mult_x_1/n288 ), .A2(n8), .ZN(n198) );
  OAI22_X1 U261 ( .A1(n185), .A2(n184), .B1(n14), .B2(n182), .ZN(n197) );
  HA_X1 U262 ( .A(n186), .B(n187), .CO(n147), .S(n228) );
  FA_X1 U263 ( .A(n190), .B(n189), .CI(n188), .CO(n225), .S(n227) );
  HA_X1 U264 ( .A(n192), .B(n191), .CO(n242), .S(n243) );
  OAI22_X1 U265 ( .A1(n7), .A2(n195), .B1(n194), .B2(n193), .ZN(n241) );
  FA_X1 U266 ( .A(n199), .B(n198), .CI(n197), .CO(n229), .S(n240) );
  OR2_X1 U267 ( .A1(n237), .A2(n236), .ZN(n200) );
  NAND2_X1 U268 ( .A1(n261), .A2(n200), .ZN(n201) );
  OAI21_X1 U269 ( .B1(n273), .B2(n449), .A(n201), .ZN(n401) );
  FA_X1 U270 ( .A(n204), .B(n203), .CI(n202), .CO(n215), .S(n221) );
  AOI21_X1 U271 ( .B1(n12), .B2(n206), .A(n205), .ZN(n208) );
  INV_X1 U272 ( .A(n208), .ZN(n211) );
  NOR2_X1 U273 ( .A1(n467), .A2(n209), .ZN(n210) );
  XOR2_X1 U274 ( .A(n211), .B(n210), .Z(n212) );
  XOR2_X1 U275 ( .A(n213), .B(n212), .Z(n214) );
  OR2_X1 U276 ( .A1(n215), .A2(n214), .ZN(n217) );
  NAND2_X1 U277 ( .A1(n215), .A2(n214), .ZN(n216) );
  NAND2_X1 U278 ( .A1(n217), .A2(n216), .ZN(n218) );
  NAND2_X1 U279 ( .A1(n261), .A2(n218), .ZN(n219) );
  OAI21_X1 U280 ( .B1(n269), .B2(n448), .A(n219), .ZN(n403) );
  NAND2_X1 U281 ( .A1(n221), .A2(n220), .ZN(n222) );
  NAND2_X1 U282 ( .A1(n269), .A2(n222), .ZN(n223) );
  OAI21_X1 U283 ( .B1(n271), .B2(n447), .A(n223), .ZN(n405) );
  FA_X1 U284 ( .A(n226), .B(n225), .CI(n224), .CO(n153), .S(n233) );
  FA_X1 U285 ( .A(n229), .B(n228), .CI(n227), .CO(n232), .S(n237) );
  NOR2_X1 U286 ( .A1(n233), .A2(n232), .ZN(n230) );
  NAND2_X1 U287 ( .A1(n273), .A2(n230), .ZN(n231) );
  OAI21_X1 U288 ( .B1(n269), .B2(n443), .A(n231), .ZN(n415) );
  NAND2_X1 U289 ( .A1(n233), .A2(n232), .ZN(n234) );
  NAND2_X1 U290 ( .A1(n234), .A2(n273), .ZN(n235) );
  OAI21_X1 U291 ( .B1(n271), .B2(n442), .A(n235), .ZN(n417) );
  NAND2_X1 U292 ( .A1(n237), .A2(n236), .ZN(n238) );
  NAND2_X1 U293 ( .A1(n261), .A2(n238), .ZN(n239) );
  OAI21_X1 U294 ( .B1(n273), .B2(n441), .A(n239), .ZN(n419) );
  FA_X1 U295 ( .A(n242), .B(n241), .CI(n240), .CO(n236), .S(n251) );
  NOR2_X1 U296 ( .A1(n251), .A2(n250), .ZN(n248) );
  NAND2_X1 U297 ( .A1(n261), .A2(n248), .ZN(n249) );
  OAI21_X1 U298 ( .B1(n269), .B2(n440), .A(n249), .ZN(n421) );
  NAND2_X1 U299 ( .A1(n251), .A2(n250), .ZN(n252) );
  NAND2_X1 U300 ( .A1(n261), .A2(n252), .ZN(n253) );
  OAI21_X1 U301 ( .B1(n269), .B2(n439), .A(n253), .ZN(n423) );
  NAND2_X1 U302 ( .A1(n255), .A2(n254), .ZN(n256) );
  NAND2_X1 U303 ( .A1(n261), .A2(n256), .ZN(n257) );
  OAI21_X1 U304 ( .B1(n271), .B2(n437), .A(n257), .ZN(n429) );
  NAND2_X1 U305 ( .A1(n259), .A2(n258), .ZN(n260) );
  NAND2_X1 U306 ( .A1(n261), .A2(n260), .ZN(n262) );
  OAI21_X1 U307 ( .B1(n273), .B2(n436), .A(n262), .ZN(n431) );
  INV_X1 U308 ( .A(n263), .ZN(n264) );
  AOI21_X1 U309 ( .B1(n266), .B2(n265), .A(n264), .ZN(n267) );
  NAND2_X1 U310 ( .A1(n269), .A2(n267), .ZN(n268) );
  OAI21_X1 U311 ( .B1(n269), .B2(n435), .A(n268), .ZN(n433) );
  INV_X1 U312 ( .A(n270), .ZN(n272) );
  NAND2_X1 U313 ( .A1(n272), .A2(n271), .ZN(n274) );
  OAI22_X1 U314 ( .A1(n275), .A2(n274), .B1(n273), .B2(n446), .ZN(n407) );
  AOI22_X1 U315 ( .A1(n269), .A2(n511), .B1(n512), .B2(n307), .ZN(n514) );
  AOI22_X1 U316 ( .A1(n372), .A2(n510), .B1(n511), .B2(n307), .ZN(n516) );
  AND2_X1 U317 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n277) );
  NAND2_X1 U318 ( .A1(n269), .A2(n277), .ZN(n278) );
  OAI21_X1 U319 ( .B1(n261), .B2(n510), .A(n278), .ZN(n518) );
  AOI22_X1 U320 ( .A1(n269), .A2(n508), .B1(n509), .B2(n307), .ZN(n520) );
  AOI22_X1 U321 ( .A1(n261), .A2(n507), .B1(n508), .B2(n307), .ZN(n522) );
  OR2_X1 U322 ( .A1(n280), .A2(n279), .ZN(n281) );
  AND2_X1 U323 ( .A1(n281), .A2(n287), .ZN(n282) );
  NAND2_X1 U324 ( .A1(n273), .A2(n282), .ZN(n283) );
  OAI21_X1 U325 ( .B1(n372), .B2(n507), .A(n283), .ZN(n524) );
  AOI22_X1 U326 ( .A1(n269), .A2(n505), .B1(n506), .B2(n307), .ZN(n526) );
  AOI22_X1 U327 ( .A1(n269), .A2(n504), .B1(n505), .B2(n307), .ZN(n528) );
  INV_X1 U328 ( .A(n284), .ZN(n286) );
  NAND2_X1 U329 ( .A1(n286), .A2(n285), .ZN(n288) );
  XOR2_X1 U330 ( .A(n288), .B(n287), .Z(n289) );
  NAND2_X1 U331 ( .A1(n269), .A2(n289), .ZN(n290) );
  OAI21_X1 U332 ( .B1(n372), .B2(n504), .A(n290), .ZN(n530) );
  AOI22_X1 U333 ( .A1(n372), .A2(n502), .B1(n503), .B2(n307), .ZN(n532) );
  AOI22_X1 U334 ( .A1(n269), .A2(n501), .B1(n502), .B2(n307), .ZN(n534) );
  NAND2_X1 U335 ( .A1(n292), .A2(n291), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  NAND2_X1 U337 ( .A1(n261), .A2(n295), .ZN(n296) );
  OAI21_X1 U338 ( .B1(n269), .B2(n501), .A(n296), .ZN(n536) );
  AOI22_X1 U339 ( .A1(n273), .A2(n499), .B1(n500), .B2(n307), .ZN(n538) );
  AOI22_X1 U340 ( .A1(n269), .A2(n498), .B1(n499), .B2(n307), .ZN(n540) );
  INV_X1 U341 ( .A(n297), .ZN(n299) );
  NAND2_X1 U342 ( .A1(n299), .A2(n298), .ZN(n301) );
  XOR2_X1 U343 ( .A(n301), .B(n300), .Z(n302) );
  NAND2_X1 U344 ( .A1(n271), .A2(n302), .ZN(n303) );
  OAI21_X1 U345 ( .B1(n372), .B2(n498), .A(n303), .ZN(n542) );
  AOI22_X1 U346 ( .A1(n261), .A2(n496), .B1(n497), .B2(n307), .ZN(n544) );
  AOI22_X1 U347 ( .A1(n269), .A2(n495), .B1(n496), .B2(n307), .ZN(n546) );
  AOI22_X1 U348 ( .A1(n273), .A2(n493), .B1(n494), .B2(n307), .ZN(n549) );
  NAND2_X1 U349 ( .A1(n440), .A2(n391), .ZN(n304) );
  XOR2_X1 U350 ( .A(n304), .B(n394), .Z(n305) );
  NAND2_X1 U351 ( .A1(n269), .A2(n305), .ZN(n306) );
  OAI21_X1 U352 ( .B1(n269), .B2(n493), .A(n306), .ZN(n551) );
  AOI22_X1 U353 ( .A1(n273), .A2(n491), .B1(n492), .B2(n307), .ZN(n553) );
  OAI21_X1 U354 ( .B1(n390), .B2(n394), .A(n391), .ZN(n312) );
  NAND2_X1 U355 ( .A1(n381), .A2(n389), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n312), .B(n308), .ZN(n309) );
  NAND2_X1 U357 ( .A1(n269), .A2(n309), .ZN(n310) );
  OAI21_X1 U358 ( .B1(n372), .B2(n491), .A(n310), .ZN(n555) );
  AOI22_X1 U359 ( .A1(n273), .A2(n489), .B1(n490), .B2(n307), .ZN(n557) );
  AOI21_X1 U360 ( .B1(n312), .B2(n381), .A(n441), .ZN(n316) );
  NAND2_X1 U361 ( .A1(n443), .A2(n388), .ZN(n313) );
  XOR2_X1 U362 ( .A(n316), .B(n313), .Z(n314) );
  NAND2_X1 U363 ( .A1(n372), .A2(n314), .ZN(n315) );
  OAI21_X1 U364 ( .B1(n372), .B2(n489), .A(n315), .ZN(n559) );
  AOI22_X1 U365 ( .A1(n261), .A2(n487), .B1(n488), .B2(n307), .ZN(n561) );
  OAI21_X1 U366 ( .B1(n316), .B2(n387), .A(n388), .ZN(n326) );
  INV_X1 U367 ( .A(n326), .ZN(n320) );
  NAND2_X1 U368 ( .A1(n444), .A2(n377), .ZN(n317) );
  XOR2_X1 U369 ( .A(n320), .B(n317), .Z(n318) );
  NAND2_X1 U370 ( .A1(n372), .A2(n318), .ZN(n319) );
  OAI21_X1 U371 ( .B1(n372), .B2(n487), .A(n319), .ZN(n563) );
  AOI22_X1 U372 ( .A1(n269), .A2(n485), .B1(n486), .B2(n307), .ZN(n565) );
  OAI21_X1 U373 ( .B1(n320), .B2(n386), .A(n377), .ZN(n322) );
  NAND2_X1 U374 ( .A1(n438), .A2(n376), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  NAND2_X1 U376 ( .A1(n372), .A2(n323), .ZN(n324) );
  OAI21_X1 U377 ( .B1(n269), .B2(n485), .A(n324), .ZN(n567) );
  AOI22_X1 U378 ( .A1(n271), .A2(n483), .B1(n484), .B2(n307), .ZN(n569) );
  NOR2_X1 U379 ( .A1(n375), .A2(n386), .ZN(n327) );
  OAI21_X1 U380 ( .B1(n375), .B2(n377), .A(n376), .ZN(n325) );
  AOI21_X1 U381 ( .B1(n327), .B2(n326), .A(n325), .ZN(n353) );
  NAND2_X1 U382 ( .A1(n446), .A2(n385), .ZN(n328) );
  XOR2_X1 U383 ( .A(n353), .B(n328), .Z(n329) );
  NAND2_X1 U384 ( .A1(n372), .A2(n329), .ZN(n330) );
  OAI21_X1 U385 ( .B1(n269), .B2(n483), .A(n330), .ZN(n571) );
  AOI22_X1 U386 ( .A1(n372), .A2(n481), .B1(n482), .B2(n307), .ZN(n573) );
  OAI21_X1 U387 ( .B1(n353), .B2(n384), .A(n385), .ZN(n332) );
  NAND2_X1 U388 ( .A1(n380), .A2(n392), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  NAND2_X1 U390 ( .A1(n372), .A2(n333), .ZN(n334) );
  OAI21_X1 U391 ( .B1(n261), .B2(n481), .A(n334), .ZN(n575) );
  AOI22_X1 U392 ( .A1(n271), .A2(n479), .B1(n480), .B2(n307), .ZN(n577) );
  NAND2_X1 U393 ( .A1(n446), .A2(n380), .ZN(n336) );
  AOI21_X1 U394 ( .B1(n445), .B2(n380), .A(n437), .ZN(n335) );
  OAI21_X1 U395 ( .B1(n353), .B2(n336), .A(n335), .ZN(n338) );
  NAND2_X1 U396 ( .A1(n379), .A2(n393), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  NAND2_X1 U398 ( .A1(n372), .A2(n339), .ZN(n340) );
  OAI21_X1 U399 ( .B1(n269), .B2(n479), .A(n340), .ZN(n579) );
  AOI22_X1 U400 ( .A1(n261), .A2(n477), .B1(n478), .B2(n307), .ZN(n581) );
  NAND2_X1 U401 ( .A1(n380), .A2(n379), .ZN(n342) );
  NOR2_X1 U402 ( .A1(n384), .A2(n342), .ZN(n349) );
  INV_X1 U403 ( .A(n349), .ZN(n344) );
  AOI21_X1 U404 ( .B1(n437), .B2(n379), .A(n436), .ZN(n341) );
  OAI21_X1 U405 ( .B1(n342), .B2(n385), .A(n341), .ZN(n350) );
  INV_X1 U406 ( .A(n350), .ZN(n343) );
  OAI21_X1 U407 ( .B1(n353), .B2(n344), .A(n343), .ZN(n346) );
  NAND2_X1 U408 ( .A1(n378), .A2(n383), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n347) );
  NAND2_X1 U410 ( .A1(n372), .A2(n347), .ZN(n348) );
  OAI21_X1 U411 ( .B1(n271), .B2(n477), .A(n348), .ZN(n583) );
  AOI22_X1 U412 ( .A1(n273), .A2(n475), .B1(n476), .B2(n307), .ZN(n585) );
  NAND2_X1 U413 ( .A1(n349), .A2(n378), .ZN(n352) );
  AOI21_X1 U414 ( .B1(n350), .B2(n378), .A(n447), .ZN(n351) );
  OAI21_X1 U415 ( .B1(n353), .B2(n352), .A(n351), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n354), .B(n382), .ZN(n355) );
  NAND2_X1 U417 ( .A1(n372), .A2(n355), .ZN(n356) );
  OAI21_X1 U418 ( .B1(n269), .B2(n475), .A(n356), .ZN(n587) );
  NAND2_X1 U419 ( .A1(n273), .A2(B_extended[0]), .ZN(n357) );
  OAI21_X1 U420 ( .B1(n273), .B2(n474), .A(n357), .ZN(n589) );
  NAND2_X1 U421 ( .A1(n372), .A2(B_extended[1]), .ZN(n358) );
  OAI21_X1 U422 ( .B1(n261), .B2(n473), .A(n358), .ZN(n591) );
  NAND2_X1 U423 ( .A1(n261), .A2(B_extended[2]), .ZN(n359) );
  OAI21_X1 U424 ( .B1(n269), .B2(n472), .A(n359), .ZN(n593) );
  NAND2_X1 U425 ( .A1(n271), .A2(B_extended[3]), .ZN(n360) );
  OAI21_X1 U426 ( .B1(n271), .B2(n471), .A(n360), .ZN(n595) );
  NAND2_X1 U427 ( .A1(n269), .A2(B_extended[4]), .ZN(n361) );
  OAI21_X1 U428 ( .B1(n269), .B2(n470), .A(n361), .ZN(n597) );
  NAND2_X1 U429 ( .A1(n269), .A2(B_extended[5]), .ZN(n362) );
  OAI21_X1 U430 ( .B1(n261), .B2(n469), .A(n362), .ZN(n599) );
  NAND2_X1 U431 ( .A1(n273), .A2(B_extended[6]), .ZN(n363) );
  OAI21_X1 U432 ( .B1(n273), .B2(n468), .A(n363), .ZN(n601) );
  NAND2_X1 U433 ( .A1(n271), .A2(B_extended[7]), .ZN(n364) );
  OAI21_X1 U434 ( .B1(n271), .B2(n467), .A(n364), .ZN(n603) );
  NAND2_X1 U435 ( .A1(n261), .A2(A_extended[0]), .ZN(n365) );
  OAI21_X1 U436 ( .B1(n273), .B2(n466), .A(n365), .ZN(n605) );
  NAND2_X1 U437 ( .A1(n269), .A2(A_extended[1]), .ZN(n366) );
  OAI21_X1 U438 ( .B1(n269), .B2(n465), .A(n366), .ZN(n607) );
  NAND2_X1 U439 ( .A1(n261), .A2(A_extended[2]), .ZN(n367) );
  OAI21_X1 U440 ( .B1(n269), .B2(n464), .A(n367), .ZN(n609) );
  NAND2_X1 U441 ( .A1(n269), .A2(A_extended[3]), .ZN(n368) );
  OAI21_X1 U442 ( .B1(n271), .B2(n463), .A(n368), .ZN(n611) );
  NAND2_X1 U443 ( .A1(n372), .A2(A_extended[4]), .ZN(n369) );
  OAI21_X1 U444 ( .B1(n273), .B2(n462), .A(n369), .ZN(n613) );
  NAND2_X1 U445 ( .A1(n273), .A2(A_extended[5]), .ZN(n370) );
  OAI21_X1 U446 ( .B1(n261), .B2(n461), .A(n370), .ZN(n615) );
  NAND2_X1 U447 ( .A1(n372), .A2(A_extended[6]), .ZN(n371) );
  OAI21_X1 U448 ( .B1(n269), .B2(n460), .A(n371), .ZN(n617) );
  NAND2_X1 U449 ( .A1(n372), .A2(A_extended[7]), .ZN(n373) );
  OAI21_X1 U450 ( .B1(n271), .B2(n459), .A(n373), .ZN(n619) );
  NAND2_X1 U451 ( .A1(n458), .A2(n307), .ZN(n621) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_28 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n397, n399, n401, n403, n405, n407, n409, n411,
         n413, n415, n417, n419, n421, n423, n425, n427, n429, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n511, n513, n515, n517, n519, n521, n523, n525, n527, n529, n531,
         n533, n535, n537, n539, n541, n543, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n567, n569, n571, n573, n575,
         n577, n579, n581, n583, n585, n587, n589, n591, n593, n595, n597,
         n599, n601, n603, n605, n607, n609, n611, n613, n615, n617, n619,
         n621, n638, n639, n640;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n452), .SE(n621), .CK(clk), .Q(n639), 
        .QN(n454) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n453), .SE(n617), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n456) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n453), .SE(n615), .CK(clk), .Q(n638), 
        .QN(n457) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n453), .SE(n613), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n458) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n453), .SE(n609), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n460) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n453), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n463) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n453), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n464) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n453), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n465) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n452), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n466) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n452), .SE(n595), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n467) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n452), .SE(n593), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n468) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n452), .SE(n591), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n469) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n452), .SE(n589), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n470) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n452), .SE(n587), .CK(clk), .QN(n471)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n452), .SE(n585), .CK(clk), .Q(
        product[15]), .QN(n472) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n452), .SE(n583), .CK(clk), .QN(n473)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n452), .SE(n581), .CK(clk), .Q(
        product[14]), .QN(n474) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n452), .SE(n579), .CK(clk), .QN(n475)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n452), .SE(n577), .CK(clk), .Q(
        product[13]), .QN(n476) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n451), .SE(n575), .CK(clk), .QN(n477)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n451), .SE(n573), .CK(clk), .Q(
        product[12]), .QN(n478) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n451), .SE(n571), .CK(clk), .QN(n479)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n451), .SE(n569), .CK(clk), .Q(
        product[11]), .QN(n480) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n451), .SE(n567), .CK(clk), .QN(n481)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n451), .SE(n565), .CK(clk), .Q(
        product[10]), .QN(n482) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n451), .SE(n563), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n451), .SE(n561), .CK(clk), .Q(
        product[9]), .QN(n484) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n451), .SE(n559), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n451), .SE(n557), .CK(clk), .Q(
        product[8]), .QN(n486) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n451), .SE(n555), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n450), .SE(n553), .CK(clk), .Q(
        product[7]), .QN(n488) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n450), .SE(n551), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n450), .SE(n549), .CK(clk), .QN(n490)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n450), .SE(n547), .CK(clk), .Q(
        product[6]), .QN(n491) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n450), .SE(n545), .CK(clk), .QN(n492)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n450), .SE(n543), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n450), .SE(n541), .CK(clk), .Q(
        product[5]), .QN(n494) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n450), .SE(n539), .CK(clk), .QN(n495)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n450), .SE(n537), .CK(clk), .QN(n496)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n450), .SE(n535), .CK(clk), .Q(
        product[4]), .QN(n497) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n450), .SE(n533), .CK(clk), .QN(n498)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n449), .SE(n531), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n449), .SE(n529), .CK(clk), .Q(
        product[3]), .QN(n500) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n449), .SE(n527), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n449), .SE(n525), .CK(clk), .QN(n502)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n449), .SE(n523), .CK(clk), .Q(
        product[2]), .QN(n503) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n449), .SE(n521), .CK(clk), .QN(n504)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n449), .SE(n519), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n449), .SE(n517), .CK(clk), .Q(
        product[1]), .QN(n506) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n449), .SE(n515), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n449), .SE(n513), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n449), .SE(n511), .CK(clk), .Q(
        product[0]), .QN(n509) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n453), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n461) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n453), .SE(n611), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n640), .SI(1'b1), .SE(n429), .CK(clk), 
        .Q(n394), .QN(n431) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n640), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n393), .QN(n432) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n640), .SE(n425), .CK(
        clk), .Q(n433), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n640), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n391), .QN(n434) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n640), .SI(1'b1), .SE(n421), .CK(clk), 
        .Q(n390), .QN(n435) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n640), .SE(n419), .CK(
        clk), .Q(n436), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n640), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n388), .QN(n437) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n640), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n387), .QN(n438) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n640), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n386), .QN(n439) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n640), .SI(1'b1), .SE(n411), .CK(clk), 
        .Q(n385), .QN(n440) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n640), .SI(1'b1), .SE(n409), .CK(clk), 
        .Q(n384), .QN(n441) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n640), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n383), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n640), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n382), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n640), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n381), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n640), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n380), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n640), .SE(n399), .CK(
        clk), .Q(n446), .QN(n379) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n640), .SE(n397), .CK(
        clk), .Q(n447), .QN(n378) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n640), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n377), .QN(n448) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n453), .SE(n619), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n455) );
  SDFF_X2 clk_r_REG61_S1 ( .D(1'b0), .SI(n453), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n462) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n452) );
  BUF_X2 U3 ( .A(n276), .Z(n376) );
  CLKBUF_X1 U4 ( .A(n266), .Z(n5) );
  CLKBUF_X2 U5 ( .A(\mult_x_1/n313 ), .Z(n215) );
  INV_X1 U6 ( .A(n14), .ZN(n15) );
  INV_X1 U7 ( .A(rst_n), .ZN(n640) );
  BUF_X2 U8 ( .A(n91), .Z(n6) );
  XNOR2_X1 U9 ( .A(\mult_x_1/a[6] ), .B(n638), .ZN(n7) );
  CLKBUF_X1 U10 ( .A(n234), .Z(n8) );
  OAI21_X1 U11 ( .B1(n232), .B2(n304), .A(n303), .ZN(n9) );
  OAI21_X1 U12 ( .B1(n298), .B2(n295), .A(n296), .ZN(n10) );
  NOR2_X1 U13 ( .A1(n72), .A2(n71), .ZN(n49) );
  NAND2_X1 U14 ( .A1(n72), .A2(n71), .ZN(n48) );
  CLKBUF_X1 U15 ( .A(n52), .Z(n11) );
  NAND2_X1 U16 ( .A1(n242), .A2(n241), .ZN(n243) );
  NAND2_X1 U17 ( .A1(n240), .A2(n239), .ZN(n241) );
  NAND2_X1 U18 ( .A1(n238), .A2(n237), .ZN(n242) );
  OR2_X1 U19 ( .A1(n240), .A2(n239), .ZN(n237) );
  XNOR2_X1 U20 ( .A(n238), .B(n199), .ZN(n231) );
  XNOR2_X1 U21 ( .A(n240), .B(n239), .ZN(n199) );
  INV_X1 U22 ( .A(n368), .ZN(n14) );
  OAI21_X1 U23 ( .B1(n50), .B2(n49), .A(n48), .ZN(n62) );
  NAND2_X1 U24 ( .A1(n184), .A2(n183), .ZN(n191) );
  NAND2_X1 U25 ( .A1(n182), .A2(n181), .ZN(n183) );
  OAI21_X1 U26 ( .B1(n182), .B2(n181), .A(n180), .ZN(n184) );
  XNOR2_X1 U27 ( .A(n72), .B(n71), .ZN(n73) );
  AND2_X1 U28 ( .A1(n268), .A2(n267), .ZN(n269) );
  BUF_X1 U29 ( .A(n5), .Z(n449) );
  BUF_X1 U30 ( .A(n5), .Z(n450) );
  BUF_X1 U31 ( .A(n5), .Z(n451) );
  BUF_X1 U32 ( .A(n5), .Z(n453) );
  NAND2_X1 U33 ( .A1(n462), .A2(\mult_x_1/n313 ), .ZN(n216) );
  XNOR2_X1 U34 ( .A(n461), .B(n467), .ZN(n206) );
  XOR2_X1 U35 ( .A(n227), .B(n226), .Z(n221) );
  AND2_X1 U36 ( .A1(n227), .A2(n226), .ZN(n228) );
  CLKBUF_X1 U37 ( .A(n210), .Z(n12) );
  INV_X1 U38 ( .A(n455), .ZN(n13) );
  NAND2_X1 U39 ( .A1(n454), .A2(n13), .ZN(n119) );
  INV_X1 U40 ( .A(n276), .ZN(n368) );
  INV_X4 U41 ( .A(n276), .ZN(n374) );
  INV_X2 U42 ( .A(n14), .ZN(n16) );
  INV_X2 U43 ( .A(n14), .ZN(n17) );
  AOI21_X1 U44 ( .B1(n290), .B2(n291), .A(n222), .ZN(n298) );
  BUF_X1 U45 ( .A(n91), .Z(n18) );
  BUF_X1 U46 ( .A(n91), .Z(n19) );
  INV_X1 U47 ( .A(n74), .ZN(n50) );
  XNOR2_X1 U48 ( .A(n74), .B(n73), .ZN(n248) );
  INV_X1 U49 ( .A(n212), .ZN(n20) );
  INV_X1 U50 ( .A(n212), .ZN(n208) );
  XOR2_X1 U51 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[2] ), .Z(n30) );
  XOR2_X1 U52 ( .A(n135), .B(n134), .Z(n21) );
  INV_X1 U53 ( .A(en), .ZN(n276) );
  XNOR2_X1 U54 ( .A(n254), .B(n253), .ZN(n22) );
  AND2_X1 U55 ( .A1(n135), .A2(n134), .ZN(n23) );
  OR2_X1 U56 ( .A1(n188), .A2(n187), .ZN(n24) );
  INV_X1 U57 ( .A(n276), .ZN(n91) );
  BUF_X2 U58 ( .A(n91), .Z(n252) );
  OR2_X1 U59 ( .A1(n259), .A2(n437), .ZN(n59) );
  XNOR2_X1 U60 ( .A(n638), .B(n458), .ZN(n25) );
  XNOR2_X1 U61 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n26) );
  NAND2_X1 U62 ( .A1(n25), .A2(n26), .ZN(n141) );
  BUF_X2 U63 ( .A(n638), .Z(n103) );
  XNOR2_X1 U64 ( .A(n103), .B(\mult_x_1/n281 ), .ZN(n32) );
  AND2_X1 U65 ( .A1(n639), .A2(\mult_x_1/n281 ), .ZN(n78) );
  XNOR2_X1 U66 ( .A(n78), .B(n103), .ZN(n81) );
  INV_X1 U67 ( .A(n26), .ZN(n27) );
  INV_X2 U68 ( .A(n27), .ZN(n201) );
  OAI22_X1 U69 ( .A1(n141), .A2(n32), .B1(n81), .B2(n201), .ZN(n86) );
  INV_X1 U70 ( .A(n86), .ZN(n85) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n310 ), .B(n456), .ZN(n28) );
  XNOR2_X1 U72 ( .A(\mult_x_1/a[6] ), .B(n638), .ZN(n29) );
  NAND2_X2 U73 ( .A1(n28), .A2(n7), .ZN(n116) );
  XNOR2_X1 U74 ( .A(n13), .B(\mult_x_1/n283 ), .ZN(n39) );
  BUF_X2 U75 ( .A(n29), .Z(n117) );
  XNOR2_X1 U76 ( .A(n13), .B(\mult_x_1/n282 ), .ZN(n80) );
  OAI22_X1 U77 ( .A1(n116), .A2(n39), .B1(n117), .B2(n80), .ZN(n84) );
  NOR2_X1 U78 ( .A1(n466), .A2(n119), .ZN(n83) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n45) );
  XNOR2_X1 U80 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n40) );
  OAI22_X1 U81 ( .A1(n116), .A2(n45), .B1(n117), .B2(n40), .ZN(n70) );
  XNOR2_X1 U82 ( .A(n103), .B(\mult_x_1/n283 ), .ZN(n46) );
  XNOR2_X1 U83 ( .A(n103), .B(\mult_x_1/n282 ), .ZN(n33) );
  OAI22_X1 U84 ( .A1(n141), .A2(n46), .B1(n201), .B2(n33), .ZN(n69) );
  BUF_X2 U85 ( .A(\mult_x_1/n312 ), .Z(n207) );
  XNOR2_X1 U86 ( .A(n207), .B(\mult_x_1/n281 ), .ZN(n47) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n31) );
  NAND2_X1 U88 ( .A1(n30), .A2(n31), .ZN(n210) );
  XNOR2_X1 U89 ( .A(n78), .B(n207), .ZN(n41) );
  INV_X1 U90 ( .A(n31), .ZN(n212) );
  OAI22_X1 U91 ( .A1(n47), .A2(n210), .B1(n41), .B2(n208), .ZN(n52) );
  INV_X1 U92 ( .A(n52), .ZN(n68) );
  NOR2_X1 U93 ( .A1(n467), .A2(n119), .ZN(n55) );
  INV_X1 U94 ( .A(n55), .ZN(n35) );
  OAI22_X1 U95 ( .A1(n141), .A2(n33), .B1(n201), .B2(n32), .ZN(n54) );
  INV_X1 U96 ( .A(n54), .ZN(n34) );
  NAND2_X1 U97 ( .A1(n35), .A2(n34), .ZN(n36) );
  NAND2_X1 U98 ( .A1(n57), .A2(n36), .ZN(n38) );
  NAND2_X1 U99 ( .A1(n55), .A2(n54), .ZN(n37) );
  NAND2_X1 U100 ( .A1(n38), .A2(n37), .ZN(n180) );
  OAI22_X1 U101 ( .A1(n116), .A2(n40), .B1(n117), .B2(n39), .ZN(n53) );
  AOI21_X1 U102 ( .B1(n20), .B2(n210), .A(n41), .ZN(n42) );
  INV_X1 U103 ( .A(n42), .ZN(n51) );
  XNOR2_X1 U104 ( .A(n180), .B(n181), .ZN(n43) );
  XNOR2_X1 U105 ( .A(n43), .B(n182), .ZN(n188) );
  XNOR2_X1 U106 ( .A(n78), .B(n215), .ZN(n66) );
  AOI21_X1 U107 ( .B1(n216), .B2(n462), .A(n66), .ZN(n44) );
  INV_X1 U108 ( .A(n44), .ZN(n138) );
  XNOR2_X1 U109 ( .A(n13), .B(\mult_x_1/n286 ), .ZN(n65) );
  OAI22_X1 U110 ( .A1(n116), .A2(n65), .B1(n117), .B2(n45), .ZN(n137) );
  NOR2_X1 U111 ( .A1(n469), .A2(n119), .ZN(n136) );
  XNOR2_X1 U112 ( .A(n103), .B(\mult_x_1/n284 ), .ZN(n139) );
  OAI22_X1 U113 ( .A1(n141), .A2(n139), .B1(n201), .B2(n46), .ZN(n64) );
  XNOR2_X1 U114 ( .A(n207), .B(\mult_x_1/n282 ), .ZN(n142) );
  OAI22_X1 U115 ( .A1(n210), .A2(n142), .B1(n208), .B2(n47), .ZN(n63) );
  OR2_X1 U116 ( .A1(n64), .A2(n63), .ZN(n72) );
  NOR2_X1 U117 ( .A1(n468), .A2(n119), .ZN(n71) );
  FA_X1 U118 ( .A(n53), .B(n11), .CI(n51), .CO(n181), .S(n61) );
  XNOR2_X1 U119 ( .A(n55), .B(n54), .ZN(n56) );
  XNOR2_X1 U120 ( .A(n57), .B(n56), .ZN(n60) );
  NAND2_X1 U121 ( .A1(n252), .A2(n24), .ZN(n58) );
  NAND2_X1 U122 ( .A1(n59), .A2(n58), .ZN(n417) );
  FA_X1 U123 ( .A(n62), .B(n61), .CI(n60), .CO(n187), .S(n262) );
  XNOR2_X1 U124 ( .A(n64), .B(n63), .ZN(n135) );
  XNOR2_X1 U125 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n94) );
  OAI22_X1 U126 ( .A1(n116), .A2(n94), .B1(n117), .B2(n65), .ZN(n148) );
  XNOR2_X1 U127 ( .A(n215), .B(\mult_x_1/n281 ), .ZN(n96) );
  OAI22_X1 U128 ( .A1(n216), .A2(n96), .B1(n66), .B2(n462), .ZN(n147) );
  INV_X1 U129 ( .A(n119), .ZN(n67) );
  AND2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n67), .ZN(n146) );
  FA_X1 U131 ( .A(n70), .B(n69), .CI(n68), .CO(n57), .S(n249) );
  NOR2_X1 U132 ( .A1(n262), .A2(n261), .ZN(n75) );
  NAND2_X1 U133 ( .A1(n75), .A2(n6), .ZN(n77) );
  OR2_X1 U134 ( .A1(n259), .A2(n436), .ZN(n76) );
  NAND2_X1 U135 ( .A1(n77), .A2(n76), .ZN(n419) );
  NOR2_X1 U154 ( .A1(n464), .A2(n119), .ZN(n114) );
  XNOR2_X1 U155 ( .A(n13), .B(\mult_x_1/n281 ), .ZN(n79) );
  XNOR2_X1 U156 ( .A(n78), .B(n13), .ZN(n115) );
  OAI22_X1 U157 ( .A1(n116), .A2(n79), .B1(n115), .B2(n117), .ZN(n123) );
  INV_X1 U158 ( .A(n123), .ZN(n113) );
  OAI22_X1 U159 ( .A1(n116), .A2(n80), .B1(n117), .B2(n79), .ZN(n88) );
  AOI21_X1 U160 ( .B1(n201), .B2(n141), .A(n81), .ZN(n82) );
  INV_X1 U161 ( .A(n82), .ZN(n87) );
  FA_X1 U162 ( .A(n85), .B(n84), .CI(n83), .CO(n179), .S(n182) );
  NOR2_X1 U163 ( .A1(n465), .A2(n119), .ZN(n178) );
  FA_X1 U164 ( .A(n88), .B(n87), .CI(n86), .CO(n112), .S(n177) );
  OR2_X1 U165 ( .A1(n131), .A2(n130), .ZN(n89) );
  NAND2_X1 U166 ( .A1(n252), .A2(n89), .ZN(n90) );
  OAI21_X1 U167 ( .B1(n19), .B2(n448), .A(n90), .ZN(n395) );
  BUF_X2 U168 ( .A(n91), .Z(n259) );
  XNOR2_X1 U169 ( .A(n215), .B(\mult_x_1/n283 ), .ZN(n198) );
  XNOR2_X1 U170 ( .A(n215), .B(\mult_x_1/n282 ), .ZN(n97) );
  OAI22_X1 U171 ( .A1(n216), .A2(n198), .B1(n97), .B2(n462), .ZN(n101) );
  XNOR2_X1 U172 ( .A(n207), .B(\mult_x_1/n285 ), .ZN(n197) );
  XNOR2_X1 U173 ( .A(n207), .B(\mult_x_1/n284 ), .ZN(n98) );
  OAI22_X1 U174 ( .A1(n210), .A2(n197), .B1(n208), .B2(n98), .ZN(n100) );
  INV_X1 U175 ( .A(n117), .ZN(n92) );
  AND2_X1 U176 ( .A1(\mult_x_1/n288 ), .A2(n92), .ZN(n99) );
  OR2_X1 U177 ( .A1(\mult_x_1/n288 ), .A2(n455), .ZN(n93) );
  OAI22_X1 U178 ( .A1(n116), .A2(n455), .B1(n93), .B2(n117), .ZN(n145) );
  XNOR2_X1 U179 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n95) );
  OAI22_X1 U180 ( .A1(n116), .A2(n95), .B1(n117), .B2(n94), .ZN(n144) );
  XNOR2_X1 U181 ( .A(n103), .B(\mult_x_1/n286 ), .ZN(n105) );
  XNOR2_X1 U182 ( .A(n103), .B(\mult_x_1/n285 ), .ZN(n140) );
  OAI22_X1 U183 ( .A1(n141), .A2(n105), .B1(n201), .B2(n140), .ZN(n151) );
  OAI22_X1 U184 ( .A1(n216), .A2(n97), .B1(n96), .B2(n462), .ZN(n150) );
  XNOR2_X1 U185 ( .A(n207), .B(\mult_x_1/n283 ), .ZN(n143) );
  OAI22_X1 U186 ( .A1(n12), .A2(n98), .B1(n20), .B2(n143), .ZN(n149) );
  FA_X1 U187 ( .A(n101), .B(n100), .CI(n99), .CO(n166), .S(n236) );
  OR2_X1 U188 ( .A1(\mult_x_1/n288 ), .A2(n457), .ZN(n102) );
  OAI22_X1 U189 ( .A1(n141), .A2(n457), .B1(n102), .B2(n201), .ZN(n196) );
  XNOR2_X1 U190 ( .A(n103), .B(\mult_x_1/n288 ), .ZN(n104) );
  XNOR2_X1 U191 ( .A(n103), .B(\mult_x_1/n287 ), .ZN(n106) );
  OAI22_X1 U192 ( .A1(n141), .A2(n104), .B1(n201), .B2(n106), .ZN(n195) );
  NAND2_X1 U193 ( .A1(n236), .A2(n8), .ZN(n109) );
  OAI22_X1 U194 ( .A1(n141), .A2(n106), .B1(n201), .B2(n105), .ZN(n233) );
  NAND2_X1 U195 ( .A1(n236), .A2(n233), .ZN(n108) );
  NAND2_X1 U196 ( .A1(n8), .A2(n233), .ZN(n107) );
  NAND3_X1 U197 ( .A1(n109), .A2(n108), .A3(n107), .ZN(n173) );
  OR2_X1 U198 ( .A1(n174), .A2(n173), .ZN(n110) );
  NAND2_X1 U199 ( .A1(n259), .A2(n110), .ZN(n111) );
  OAI21_X1 U200 ( .B1(n6), .B2(n447), .A(n111), .ZN(n397) );
  FA_X1 U201 ( .A(n114), .B(n113), .CI(n112), .CO(n125), .S(n131) );
  AOI21_X1 U202 ( .B1(n117), .B2(n116), .A(n115), .ZN(n118) );
  INV_X1 U203 ( .A(n118), .ZN(n121) );
  NOR2_X1 U204 ( .A1(n463), .A2(n119), .ZN(n120) );
  XOR2_X1 U205 ( .A(n121), .B(n120), .Z(n122) );
  XOR2_X1 U206 ( .A(n123), .B(n122), .Z(n124) );
  OR2_X1 U207 ( .A1(n125), .A2(n124), .ZN(n127) );
  NAND2_X1 U208 ( .A1(n125), .A2(n124), .ZN(n126) );
  NAND2_X1 U209 ( .A1(n127), .A2(n126), .ZN(n128) );
  NAND2_X1 U210 ( .A1(n18), .A2(n128), .ZN(n129) );
  OAI21_X1 U211 ( .B1(n252), .B2(n446), .A(n129), .ZN(n399) );
  NAND2_X1 U212 ( .A1(n131), .A2(n130), .ZN(n132) );
  NAND2_X1 U213 ( .A1(n252), .A2(n132), .ZN(n133) );
  OAI21_X1 U214 ( .B1(n17), .B2(n445), .A(n133), .ZN(n401) );
  FA_X1 U215 ( .A(n138), .B(n137), .CI(n136), .CO(n74), .S(n254) );
  OAI22_X1 U216 ( .A1(n141), .A2(n140), .B1(n201), .B2(n139), .ZN(n154) );
  OAI22_X1 U217 ( .A1(n12), .A2(n143), .B1(n20), .B2(n142), .ZN(n153) );
  HA_X1 U218 ( .A(n145), .B(n144), .CO(n152), .S(n165) );
  XNOR2_X1 U219 ( .A(n21), .B(n22), .ZN(n158) );
  FA_X1 U220 ( .A(n148), .B(n147), .CI(n146), .CO(n134), .S(n163) );
  FA_X1 U221 ( .A(n151), .B(n150), .CI(n149), .CO(n162), .S(n164) );
  FA_X1 U222 ( .A(n154), .B(n153), .CI(n152), .CO(n253), .S(n161) );
  NOR2_X1 U223 ( .A1(n158), .A2(n157), .ZN(n155) );
  NAND2_X1 U224 ( .A1(n6), .A2(n155), .ZN(n156) );
  OAI21_X1 U225 ( .B1(n252), .B2(n444), .A(n156), .ZN(n403) );
  NAND2_X1 U226 ( .A1(n158), .A2(n157), .ZN(n159) );
  NAND2_X1 U227 ( .A1(n159), .A2(n6), .ZN(n160) );
  OAI21_X1 U228 ( .B1(n19), .B2(n443), .A(n160), .ZN(n405) );
  FA_X1 U229 ( .A(n163), .B(n162), .CI(n161), .CO(n157), .S(n170) );
  FA_X1 U230 ( .A(n166), .B(n165), .CI(n164), .CO(n169), .S(n174) );
  NOR2_X1 U231 ( .A1(n170), .A2(n169), .ZN(n167) );
  NAND2_X1 U232 ( .A1(n259), .A2(n167), .ZN(n168) );
  OAI21_X1 U233 ( .B1(n259), .B2(n442), .A(n168), .ZN(n407) );
  NAND2_X1 U234 ( .A1(n170), .A2(n169), .ZN(n171) );
  NAND2_X1 U235 ( .A1(n171), .A2(n19), .ZN(n172) );
  OAI21_X1 U236 ( .B1(n6), .B2(n441), .A(n172), .ZN(n409) );
  NAND2_X1 U237 ( .A1(n174), .A2(n173), .ZN(n175) );
  NAND2_X1 U238 ( .A1(n6), .A2(n175), .ZN(n176) );
  OAI21_X1 U239 ( .B1(n6), .B2(n440), .A(n176), .ZN(n411) );
  FA_X1 U240 ( .A(n179), .B(n178), .CI(n177), .CO(n130), .S(n192) );
  NAND2_X1 U241 ( .A1(n192), .A2(n191), .ZN(n185) );
  NAND2_X1 U242 ( .A1(n259), .A2(n185), .ZN(n186) );
  OAI21_X1 U243 ( .B1(n18), .B2(n439), .A(n186), .ZN(n413) );
  NAND2_X1 U244 ( .A1(n188), .A2(n187), .ZN(n189) );
  NAND2_X1 U245 ( .A1(n259), .A2(n189), .ZN(n190) );
  OAI21_X1 U246 ( .B1(n252), .B2(n438), .A(n190), .ZN(n415) );
  OR2_X1 U247 ( .A1(n192), .A2(n191), .ZN(n193) );
  NAND2_X1 U248 ( .A1(n252), .A2(n193), .ZN(n194) );
  OAI21_X1 U249 ( .B1(n6), .B2(n434), .A(n194), .ZN(n423) );
  HA_X1 U250 ( .A(n196), .B(n195), .CO(n234), .S(n238) );
  XNOR2_X1 U251 ( .A(n207), .B(\mult_x_1/n286 ), .ZN(n203) );
  OAI22_X1 U252 ( .A1(n210), .A2(n203), .B1(n208), .B2(n197), .ZN(n240) );
  XNOR2_X1 U253 ( .A(n215), .B(\mult_x_1/n284 ), .ZN(n200) );
  OAI22_X1 U254 ( .A1(n216), .A2(n200), .B1(n198), .B2(n462), .ZN(n239) );
  OAI22_X1 U255 ( .A1(n216), .A2(n206), .B1(n200), .B2(n462), .ZN(n225) );
  INV_X1 U256 ( .A(n201), .ZN(n202) );
  AND2_X1 U257 ( .A1(\mult_x_1/n288 ), .A2(n202), .ZN(n224) );
  XNOR2_X1 U258 ( .A(n207), .B(\mult_x_1/n287 ), .ZN(n204) );
  OAI22_X1 U259 ( .A1(n210), .A2(n204), .B1(n20), .B2(n203), .ZN(n223) );
  NAND2_X1 U260 ( .A1(n231), .A2(n230), .ZN(n302) );
  INV_X1 U261 ( .A(n302), .ZN(n232) );
  XNOR2_X1 U262 ( .A(n207), .B(\mult_x_1/n288 ), .ZN(n205) );
  OAI22_X1 U263 ( .A1(n210), .A2(n205), .B1(n208), .B2(n204), .ZN(n227) );
  XNOR2_X1 U264 ( .A(n215), .B(\mult_x_1/n286 ), .ZN(n211) );
  OAI22_X1 U265 ( .A1(n216), .A2(n211), .B1(n206), .B2(n462), .ZN(n226) );
  OR2_X1 U266 ( .A1(\mult_x_1/n288 ), .A2(n459), .ZN(n209) );
  OAI22_X1 U267 ( .A1(n12), .A2(n459), .B1(n209), .B2(n20), .ZN(n220) );
  OR2_X1 U268 ( .A1(n221), .A2(n220), .ZN(n290) );
  XNOR2_X1 U269 ( .A(n215), .B(\mult_x_1/n287 ), .ZN(n214) );
  OAI22_X1 U270 ( .A1(n216), .A2(n214), .B1(n211), .B2(n462), .ZN(n219) );
  AND2_X1 U271 ( .A1(\mult_x_1/n288 ), .A2(n212), .ZN(n218) );
  NOR2_X1 U272 ( .A1(n219), .A2(n218), .ZN(n282) );
  OAI22_X1 U273 ( .A1(n216), .A2(\mult_x_1/n288 ), .B1(n214), .B2(n462), .ZN(
        n278) );
  OR2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(n461), .ZN(n217) );
  NAND2_X1 U275 ( .A1(n217), .A2(n216), .ZN(n277) );
  NAND2_X1 U276 ( .A1(n278), .A2(n277), .ZN(n285) );
  NAND2_X1 U277 ( .A1(n219), .A2(n218), .ZN(n283) );
  OAI21_X1 U278 ( .B1(n282), .B2(n285), .A(n283), .ZN(n291) );
  NAND2_X1 U279 ( .A1(n221), .A2(n220), .ZN(n289) );
  INV_X1 U280 ( .A(n289), .ZN(n222) );
  FA_X1 U281 ( .A(n225), .B(n224), .CI(n223), .CO(n230), .S(n229) );
  NOR2_X1 U282 ( .A1(n229), .A2(n228), .ZN(n295) );
  NAND2_X1 U283 ( .A1(n229), .A2(n228), .ZN(n296) );
  OAI21_X1 U284 ( .B1(n298), .B2(n295), .A(n296), .ZN(n304) );
  OR2_X1 U285 ( .A1(n231), .A2(n230), .ZN(n303) );
  OAI21_X1 U286 ( .B1(n232), .B2(n10), .A(n303), .ZN(n270) );
  XNOR2_X1 U287 ( .A(n234), .B(n233), .ZN(n235) );
  XNOR2_X1 U288 ( .A(n236), .B(n235), .ZN(n244) );
  OR2_X1 U289 ( .A1(n244), .A2(n243), .ZN(n268) );
  INV_X1 U290 ( .A(n268), .ZN(n245) );
  NAND2_X1 U291 ( .A1(n244), .A2(n243), .ZN(n267) );
  OAI21_X1 U292 ( .B1(n270), .B2(n245), .A(n267), .ZN(n246) );
  NAND2_X1 U293 ( .A1(n259), .A2(n246), .ZN(n247) );
  OAI21_X1 U294 ( .B1(n18), .B2(n433), .A(n247), .ZN(n425) );
  FA_X1 U295 ( .A(n23), .B(n249), .CI(n248), .CO(n261), .S(n250) );
  NAND2_X1 U296 ( .A1(n259), .A2(n250), .ZN(n251) );
  OAI21_X1 U297 ( .B1(n252), .B2(n432), .A(n251), .ZN(n427) );
  NAND2_X1 U298 ( .A1(n21), .A2(n254), .ZN(n257) );
  NAND2_X1 U299 ( .A1(n21), .A2(n253), .ZN(n256) );
  NAND2_X1 U300 ( .A1(n254), .A2(n253), .ZN(n255) );
  NAND3_X1 U301 ( .A1(n257), .A2(n256), .A3(n255), .ZN(n258) );
  NAND2_X1 U302 ( .A1(n6), .A2(n258), .ZN(n260) );
  OAI21_X1 U303 ( .B1(n18), .B2(n431), .A(n260), .ZN(n429) );
  OR2_X1 U304 ( .A1(n259), .A2(n435), .ZN(n265) );
  NAND2_X1 U305 ( .A1(n262), .A2(n261), .ZN(n263) );
  NAND2_X1 U306 ( .A1(n252), .A2(n263), .ZN(n264) );
  NAND2_X1 U307 ( .A1(n265), .A2(n264), .ZN(n421) );
  INV_X1 U308 ( .A(n640), .ZN(n266) );
  XNOR2_X1 U309 ( .A(n9), .B(n269), .ZN(n271) );
  NAND2_X1 U310 ( .A1(n271), .A2(n374), .ZN(n273) );
  OR2_X1 U311 ( .A1(n374), .A2(n489), .ZN(n272) );
  NAND2_X1 U312 ( .A1(n273), .A2(n272), .ZN(n551) );
  AOI22_X1 U313 ( .A1(n374), .A2(n508), .B1(n509), .B2(n376), .ZN(n511) );
  AOI22_X1 U314 ( .A1(n19), .A2(n507), .B1(n508), .B2(n376), .ZN(n513) );
  AND2_X1 U315 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n274) );
  NAND2_X1 U316 ( .A1(n374), .A2(n274), .ZN(n275) );
  OAI21_X1 U317 ( .B1(n19), .B2(n507), .A(n275), .ZN(n515) );
  AOI22_X1 U318 ( .A1(n19), .A2(n505), .B1(n506), .B2(n376), .ZN(n517) );
  AOI22_X1 U319 ( .A1(n6), .A2(n504), .B1(n505), .B2(n376), .ZN(n519) );
  OR2_X1 U320 ( .A1(n278), .A2(n277), .ZN(n279) );
  AND2_X1 U321 ( .A1(n279), .A2(n285), .ZN(n280) );
  NAND2_X1 U322 ( .A1(n374), .A2(n280), .ZN(n281) );
  OAI21_X1 U323 ( .B1(n17), .B2(n504), .A(n281), .ZN(n521) );
  AOI22_X1 U324 ( .A1(n374), .A2(n502), .B1(n503), .B2(n376), .ZN(n523) );
  AOI22_X1 U325 ( .A1(n17), .A2(n501), .B1(n502), .B2(n376), .ZN(n525) );
  INV_X1 U326 ( .A(n282), .ZN(n284) );
  NAND2_X1 U327 ( .A1(n284), .A2(n283), .ZN(n286) );
  XOR2_X1 U328 ( .A(n286), .B(n285), .Z(n287) );
  NAND2_X1 U329 ( .A1(n374), .A2(n287), .ZN(n288) );
  OAI21_X1 U330 ( .B1(n19), .B2(n501), .A(n288), .ZN(n527) );
  AOI22_X1 U331 ( .A1(n17), .A2(n499), .B1(n500), .B2(n376), .ZN(n529) );
  AOI22_X1 U332 ( .A1(n374), .A2(n498), .B1(n499), .B2(n376), .ZN(n531) );
  NAND2_X1 U333 ( .A1(n290), .A2(n289), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n293) );
  NAND2_X1 U335 ( .A1(n16), .A2(n293), .ZN(n294) );
  OAI21_X1 U336 ( .B1(n16), .B2(n498), .A(n294), .ZN(n533) );
  AOI22_X1 U337 ( .A1(n17), .A2(n496), .B1(n497), .B2(n376), .ZN(n535) );
  AOI22_X1 U338 ( .A1(n17), .A2(n495), .B1(n496), .B2(n376), .ZN(n537) );
  INV_X1 U339 ( .A(n295), .ZN(n297) );
  NAND2_X1 U340 ( .A1(n297), .A2(n296), .ZN(n299) );
  XOR2_X1 U341 ( .A(n299), .B(n298), .Z(n300) );
  NAND2_X1 U342 ( .A1(n15), .A2(n300), .ZN(n301) );
  OAI21_X1 U343 ( .B1(n17), .B2(n495), .A(n301), .ZN(n539) );
  AOI22_X1 U344 ( .A1(n374), .A2(n493), .B1(n494), .B2(n376), .ZN(n541) );
  AOI22_X1 U345 ( .A1(n18), .A2(n492), .B1(n493), .B2(n376), .ZN(n543) );
  NAND2_X1 U346 ( .A1(n303), .A2(n302), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n305), .B(n10), .ZN(n306) );
  NAND2_X1 U348 ( .A1(n15), .A2(n306), .ZN(n307) );
  OAI21_X1 U349 ( .B1(n374), .B2(n492), .A(n307), .ZN(n545) );
  AOI22_X1 U350 ( .A1(n252), .A2(n490), .B1(n491), .B2(n376), .ZN(n547) );
  AOI22_X1 U351 ( .A1(n17), .A2(n489), .B1(n490), .B2(n376), .ZN(n549) );
  AOI22_X1 U352 ( .A1(n259), .A2(n487), .B1(n488), .B2(n376), .ZN(n553) );
  NAND2_X1 U353 ( .A1(n378), .A2(n385), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n392), .B(n308), .ZN(n309) );
  NAND2_X1 U355 ( .A1(n252), .A2(n309), .ZN(n310) );
  OAI21_X1 U356 ( .B1(n16), .B2(n487), .A(n310), .ZN(n555) );
  AOI22_X1 U357 ( .A1(n17), .A2(n485), .B1(n486), .B2(n376), .ZN(n557) );
  AOI21_X1 U358 ( .B1(n392), .B2(n378), .A(n440), .ZN(n314) );
  NAND2_X1 U359 ( .A1(n442), .A2(n384), .ZN(n311) );
  XOR2_X1 U360 ( .A(n314), .B(n311), .Z(n312) );
  NAND2_X1 U361 ( .A1(n374), .A2(n312), .ZN(n313) );
  OAI21_X1 U362 ( .B1(n18), .B2(n485), .A(n313), .ZN(n559) );
  AOI22_X1 U363 ( .A1(n374), .A2(n483), .B1(n484), .B2(n376), .ZN(n561) );
  OAI21_X1 U364 ( .B1(n314), .B2(n383), .A(n384), .ZN(n327) );
  INV_X1 U365 ( .A(n327), .ZN(n318) );
  NAND2_X1 U366 ( .A1(n444), .A2(n382), .ZN(n315) );
  XOR2_X1 U367 ( .A(n318), .B(n315), .Z(n316) );
  NAND2_X1 U368 ( .A1(n16), .A2(n316), .ZN(n317) );
  OAI21_X1 U369 ( .B1(n252), .B2(n483), .A(n317), .ZN(n563) );
  AOI22_X1 U370 ( .A1(n374), .A2(n481), .B1(n482), .B2(n376), .ZN(n565) );
  OAI21_X1 U371 ( .B1(n318), .B2(n381), .A(n382), .ZN(n321) );
  NOR2_X1 U372 ( .A1(n393), .A2(n394), .ZN(n325) );
  INV_X1 U373 ( .A(n325), .ZN(n319) );
  NAND2_X1 U374 ( .A1(n393), .A2(n394), .ZN(n324) );
  NAND2_X1 U375 ( .A1(n319), .A2(n324), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  NAND2_X1 U377 ( .A1(n15), .A2(n322), .ZN(n323) );
  OAI21_X1 U378 ( .B1(n17), .B2(n481), .A(n323), .ZN(n567) );
  AOI22_X1 U379 ( .A1(n17), .A2(n479), .B1(n480), .B2(n376), .ZN(n569) );
  NOR2_X1 U380 ( .A1(n325), .A2(n381), .ZN(n328) );
  OAI21_X1 U381 ( .B1(n325), .B2(n382), .A(n324), .ZN(n326) );
  AOI21_X1 U382 ( .B1(n328), .B2(n327), .A(n326), .ZN(n354) );
  NAND2_X1 U383 ( .A1(n436), .A2(n390), .ZN(n329) );
  XOR2_X1 U384 ( .A(n354), .B(n329), .Z(n330) );
  NAND2_X1 U385 ( .A1(n374), .A2(n330), .ZN(n331) );
  OAI21_X1 U386 ( .B1(n374), .B2(n479), .A(n331), .ZN(n571) );
  AOI22_X1 U387 ( .A1(n16), .A2(n477), .B1(n478), .B2(n376), .ZN(n573) );
  OAI21_X1 U388 ( .B1(n354), .B2(n389), .A(n390), .ZN(n333) );
  NAND2_X1 U389 ( .A1(n388), .A2(n387), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  NAND2_X1 U391 ( .A1(n16), .A2(n334), .ZN(n335) );
  OAI21_X1 U392 ( .B1(n15), .B2(n477), .A(n335), .ZN(n575) );
  AOI22_X1 U393 ( .A1(n17), .A2(n475), .B1(n476), .B2(n376), .ZN(n577) );
  NAND2_X1 U394 ( .A1(n436), .A2(n388), .ZN(n337) );
  AOI21_X1 U395 ( .B1(n435), .B2(n388), .A(n438), .ZN(n336) );
  OAI21_X1 U396 ( .B1(n354), .B2(n337), .A(n336), .ZN(n339) );
  NAND2_X1 U397 ( .A1(n391), .A2(n386), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  NAND2_X1 U399 ( .A1(n15), .A2(n340), .ZN(n341) );
  OAI21_X1 U400 ( .B1(n6), .B2(n475), .A(n341), .ZN(n579) );
  AOI22_X1 U401 ( .A1(n17), .A2(n473), .B1(n474), .B2(n376), .ZN(n581) );
  NAND2_X1 U402 ( .A1(n388), .A2(n391), .ZN(n343) );
  NOR2_X1 U403 ( .A1(n389), .A2(n343), .ZN(n350) );
  INV_X1 U404 ( .A(n350), .ZN(n345) );
  AOI21_X1 U405 ( .B1(n438), .B2(n391), .A(n439), .ZN(n342) );
  OAI21_X1 U406 ( .B1(n343), .B2(n390), .A(n342), .ZN(n351) );
  INV_X1 U407 ( .A(n351), .ZN(n344) );
  OAI21_X1 U408 ( .B1(n354), .B2(n345), .A(n344), .ZN(n347) );
  NAND2_X1 U409 ( .A1(n377), .A2(n380), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  NAND2_X1 U411 ( .A1(n374), .A2(n348), .ZN(n349) );
  OAI21_X1 U412 ( .B1(n16), .B2(n473), .A(n349), .ZN(n583) );
  AOI22_X1 U413 ( .A1(n374), .A2(n471), .B1(n472), .B2(n376), .ZN(n585) );
  NAND2_X1 U414 ( .A1(n350), .A2(n377), .ZN(n353) );
  AOI21_X1 U415 ( .B1(n351), .B2(n377), .A(n445), .ZN(n352) );
  OAI21_X1 U416 ( .B1(n354), .B2(n353), .A(n352), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n355), .B(n379), .ZN(n356) );
  NAND2_X1 U418 ( .A1(n15), .A2(n356), .ZN(n357) );
  OAI21_X1 U419 ( .B1(n16), .B2(n471), .A(n357), .ZN(n587) );
  NAND2_X1 U420 ( .A1(n15), .A2(B_extended[0]), .ZN(n358) );
  OAI21_X1 U421 ( .B1(n374), .B2(n470), .A(n358), .ZN(n589) );
  NAND2_X1 U422 ( .A1(n6), .A2(B_extended[1]), .ZN(n359) );
  OAI21_X1 U423 ( .B1(n374), .B2(n469), .A(n359), .ZN(n591) );
  NAND2_X1 U424 ( .A1(n374), .A2(B_extended[2]), .ZN(n360) );
  OAI21_X1 U425 ( .B1(n16), .B2(n468), .A(n360), .ZN(n593) );
  NAND2_X1 U426 ( .A1(n374), .A2(B_extended[3]), .ZN(n361) );
  OAI21_X1 U427 ( .B1(n374), .B2(n467), .A(n361), .ZN(n595) );
  NAND2_X1 U428 ( .A1(n15), .A2(B_extended[4]), .ZN(n362) );
  OAI21_X1 U429 ( .B1(n17), .B2(n466), .A(n362), .ZN(n597) );
  NAND2_X1 U430 ( .A1(n374), .A2(B_extended[5]), .ZN(n363) );
  OAI21_X1 U431 ( .B1(n16), .B2(n465), .A(n363), .ZN(n599) );
  NAND2_X1 U432 ( .A1(n259), .A2(B_extended[6]), .ZN(n364) );
  OAI21_X1 U433 ( .B1(n18), .B2(n464), .A(n364), .ZN(n601) );
  NAND2_X1 U434 ( .A1(n374), .A2(B_extended[7]), .ZN(n365) );
  OAI21_X1 U435 ( .B1(n17), .B2(n463), .A(n365), .ZN(n603) );
  NAND2_X1 U436 ( .A1(n374), .A2(A_extended[0]), .ZN(n366) );
  OAI21_X1 U437 ( .B1(n16), .B2(n462), .A(n366), .ZN(n605) );
  NAND2_X1 U438 ( .A1(n259), .A2(A_extended[1]), .ZN(n367) );
  OAI21_X1 U439 ( .B1(n17), .B2(n461), .A(n367), .ZN(n607) );
  NAND2_X1 U440 ( .A1(n16), .A2(A_extended[2]), .ZN(n369) );
  OAI21_X1 U441 ( .B1(n91), .B2(n460), .A(n369), .ZN(n609) );
  NAND2_X1 U442 ( .A1(n374), .A2(A_extended[3]), .ZN(n370) );
  OAI21_X1 U443 ( .B1(n17), .B2(n459), .A(n370), .ZN(n611) );
  NAND2_X1 U444 ( .A1(n374), .A2(A_extended[4]), .ZN(n371) );
  OAI21_X1 U445 ( .B1(n374), .B2(n458), .A(n371), .ZN(n613) );
  NAND2_X1 U446 ( .A1(n374), .A2(A_extended[5]), .ZN(n372) );
  OAI21_X1 U447 ( .B1(n374), .B2(n457), .A(n372), .ZN(n615) );
  NAND2_X1 U448 ( .A1(n374), .A2(A_extended[6]), .ZN(n373) );
  OAI21_X1 U449 ( .B1(n374), .B2(n456), .A(n373), .ZN(n617) );
  NAND2_X1 U450 ( .A1(n374), .A2(A_extended[7]), .ZN(n375) );
  OAI21_X1 U451 ( .B1(n374), .B2(n455), .A(n375), .ZN(n619) );
  NAND2_X1 U452 ( .A1(n454), .A2(n376), .ZN(n621) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_29 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[2] , \mult_x_1/n312 , \mult_x_1/n311 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n405, n407, n409, n411,
         n413, n415, n417, n419, n421, n423, n425, n427, n429, n431, n433,
         n435, n437, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n515, n517, n519, n521, n523, n525, n527, n529, n531, n533, n535,
         n537, n539, n541, n543, n545, n547, n548, n550, n552, n554, n556,
         n558, n560, n562, n564, n566, n568, n570, n572, n574, n576, n578,
         n580, n582, n584, n586, n588, n590, n592, n594, n596, n598, n600,
         n602, n604, n606, n608, n610, n612, n614, n616, n618, n620, n622,
         n624, n641, n642, n643;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n624), .CK(clk), .Q(n642), 
        .QN(n458) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n620), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n460) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(rst_n), .SE(n616), .CK(clk), .QN(n462) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(rst_n), .SE(n612), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n464) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(rst_n), .SE(n610), .CK(clk), .Q(n641), 
        .QN(n465) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(rst_n), .SE(n606), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n467) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n604), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n468) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n602), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n469) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n457), .SE(n600), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n470) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n456), .SE(n598), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n471) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n596), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n472) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n457), .SE(n594), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n473) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n456), .SE(n592), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n474) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n590), .CK(clk), .QN(n475)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n588), .CK(clk), .Q(
        product[15]), .QN(n476) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n456), .SE(n586), .CK(clk), .QN(n477)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n457), .SE(n584), .CK(clk), .Q(
        product[14]), .QN(n478) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n457), .SE(n582), .CK(clk), .QN(n479)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n456), .SE(n580), .CK(clk), .Q(
        product[13]), .QN(n480) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n457), .SE(n578), .CK(clk), .QN(n481)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n457), .SE(n576), .CK(clk), .Q(
        product[12]), .QN(n482) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n457), .SE(n574), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n457), .SE(n572), .CK(clk), .Q(
        product[11]), .QN(n484) );
  SDFF_X1 clk_r_REG23_S3 ( .D(1'b0), .SI(n457), .SE(n570), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG24_S4 ( .D(1'b0), .SI(n457), .SE(n568), .CK(clk), .Q(
        product[10]), .QN(n486) );
  SDFF_X1 clk_r_REG21_S3 ( .D(1'b0), .SI(n457), .SE(n566), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG22_S4 ( .D(1'b0), .SI(n457), .SE(n564), .CK(clk), .Q(
        product[9]), .QN(n488) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n457), .SE(n562), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n457), .SE(n560), .CK(clk), .Q(
        product[8]), .QN(n490) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n457), .SE(n558), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n456), .SE(n556), .CK(clk), .Q(
        product[7]), .QN(n492) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n456), .SE(n552), .CK(clk), .QN(n494)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n456), .SE(n550), .CK(clk), .Q(
        product[6]), .QN(n495) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n456), .SE(n547), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n456), .SE(n545), .CK(clk), .Q(
        product[5]), .QN(n498) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n456), .SE(n543), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n456), .SE(n541), .CK(clk), .QN(n500)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n456), .SE(n539), .CK(clk), .Q(
        product[4]), .QN(n501) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n456), .SE(n537), .CK(clk), .QN(n502)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(rst_n), .SE(n535), .CK(clk), .QN(n503) );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(rst_n), .SE(n533), .CK(clk), .Q(
        product[3]), .QN(n504) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(rst_n), .SE(n531), .CK(clk), .QN(n505) );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(rst_n), .SE(n529), .CK(clk), .QN(n506) );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(rst_n), .SE(n527), .CK(clk), .Q(
        product[2]), .QN(n507) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(rst_n), .SE(n525), .CK(clk), .QN(n508) );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(rst_n), .SE(n523), .CK(clk), .QN(n509) );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(rst_n), .SE(n521), .CK(clk), .Q(
        product[1]), .QN(n510) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(rst_n), .SE(n519), .CK(clk), .QN(n511) );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(rst_n), .SE(n517), .CK(clk), .QN(n512) );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(rst_n), .SE(n515), .CK(clk), .Q(
        product[0]), .QN(n513) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n456), .SE(n554), .CK(clk), .Q(n455), 
        .QN(n493) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n643), .SE(n417), .CK(
        clk), .Q(n447), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n643), .SE(n437), .CK(
        clk), .Q(n439), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n643), .SI(1'b1), .SE(n435), .CK(clk), 
        .Q(n401), .QN(n440) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n643), .SE(n431), .CK(
        clk), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n643), .SI(1'b1), .SE(n429), .CK(clk), 
        .Q(n398), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n643), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n643), .SI(1'b1), .SE(n425), .CK(clk), 
        .Q(n396), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n643), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n395), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n643), .SI(1'b1), .SE(n421), .CK(clk), 
        .Q(n394), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n643), .SI(1'b1), .SE(n419), .CK(clk), 
        .Q(n393), .QN(n446) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n643), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n391), .QN(n448) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n643), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n390), .QN(n449) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n643), .SE(n411), .CK(
        clk), .Q(n450), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n643), .SE(n409), .CK(
        clk), .Q(n451), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n643), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n387), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n643), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n386), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n643), .SI(1'b1), .SE(n403), .CK(clk), 
        .Q(n385), .QN(n454) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n622), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n459) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n618), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n461) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n643), .SE(n433), .CK(
        clk), .Q(n441), .QN(n400) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n456), .SE(n548), .CK(clk), .QN(n496)
         );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(rst_n), .SE(n614), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n463) );
  SDFF_X2 clk_r_REG61_S1 ( .D(1'b0), .SI(rst_n), .SE(n608), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n466) );
  INV_X1 U2 ( .A(n356), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(rst_n), .Z(n456) );
  CLKBUF_X1 U4 ( .A(rst_n), .Z(n457) );
  INV_X1 U5 ( .A(n459), .ZN(n11) );
  INV_X2 U6 ( .A(n281), .ZN(n6) );
  INV_X2 U7 ( .A(en), .ZN(n281) );
  NAND2_X2 U8 ( .A1(n641), .A2(n466), .ZN(n162) );
  INV_X1 U9 ( .A(n463), .ZN(n7) );
  INV_X1 U10 ( .A(n141), .ZN(n15) );
  CLKBUF_X1 U11 ( .A(n141), .Z(n14) );
  INV_X1 U12 ( .A(n39), .ZN(n40) );
  NAND2_X1 U13 ( .A1(n126), .A2(n36), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n71), .B(n70), .ZN(n104) );
  AND2_X1 U15 ( .A1(n41), .A2(n39), .ZN(n110) );
  NAND2_X1 U16 ( .A1(n134), .A2(n133), .ZN(n174) );
  NAND2_X1 U17 ( .A1(n136), .A2(n135), .ZN(n133) );
  NAND2_X1 U18 ( .A1(n138), .A2(n132), .ZN(n134) );
  OR2_X1 U19 ( .A1(n136), .A2(n135), .ZN(n132) );
  INV_X1 U20 ( .A(n461), .ZN(n13) );
  AND2_X1 U21 ( .A1(\mult_x_1/n310 ), .A2(n642), .ZN(n21) );
  XNOR2_X1 U22 ( .A(n136), .B(n135), .ZN(n137) );
  NAND2_X1 U23 ( .A1(n144), .A2(n143), .ZN(n171) );
  INV_X1 U24 ( .A(n146), .ZN(n142) );
  CLKBUF_X1 U25 ( .A(n87), .Z(n17) );
  NAND2_X1 U26 ( .A1(n78), .A2(n77), .ZN(n256) );
  NAND2_X1 U27 ( .A1(n267), .A2(n266), .ZN(n268) );
  NAND2_X1 U28 ( .A1(n265), .A2(n264), .ZN(n269) );
  OR2_X1 U29 ( .A1(n267), .A2(n266), .ZN(n264) );
  XNOR2_X1 U30 ( .A(n32), .B(n265), .ZN(n221) );
  XNOR2_X1 U31 ( .A(n267), .B(n266), .ZN(n32) );
  NAND2_X1 U32 ( .A1(n38), .A2(n37), .ZN(n207) );
  NAND2_X1 U33 ( .A1(n213), .A2(n212), .ZN(n224) );
  NAND2_X1 U34 ( .A1(n211), .A2(n210), .ZN(n212) );
  OR2_X1 U35 ( .A1(n211), .A2(n210), .ZN(n208) );
  OAI22_X1 U36 ( .A1(n177), .A2(n5), .B1(n378), .B2(n439), .ZN(n437) );
  INV_X1 U37 ( .A(n274), .ZN(n176) );
  AOI21_X1 U38 ( .B1(n275), .B2(n277), .A(n176), .ZN(n177) );
  NAND2_X1 U39 ( .A1(n23), .A2(n22), .ZN(n8) );
  NAND2_X1 U40 ( .A1(n23), .A2(n22), .ZN(n9) );
  NAND2_X1 U41 ( .A1(n23), .A2(n22), .ZN(n186) );
  NAND2_X1 U42 ( .A1(n105), .A2(n104), .ZN(n77) );
  OAI21_X1 U43 ( .B1(n105), .B2(n104), .A(n18), .ZN(n78) );
  OR2_X1 U44 ( .A1(n75), .A2(n76), .ZN(n65) );
  NAND2_X1 U45 ( .A1(n209), .A2(n208), .ZN(n213) );
  OR2_X1 U46 ( .A1(n124), .A2(n123), .ZN(n36) );
  NAND2_X1 U47 ( .A1(n124), .A2(n123), .ZN(n37) );
  NAND2_X1 U48 ( .A1(n172), .A2(n171), .ZN(n310) );
  OR2_X1 U49 ( .A1(n172), .A2(n171), .ZN(n311) );
  NAND2_X1 U50 ( .A1(n25), .A2(n26), .ZN(n12) );
  INV_X1 U51 ( .A(n141), .ZN(n187) );
  OAI21_X1 U52 ( .B1(n302), .B2(n305), .A(n303), .ZN(n10) );
  INV_X4 U53 ( .A(n316), .ZN(n356) );
  NAND2_X1 U54 ( .A1(n147), .A2(n145), .ZN(n143) );
  OAI21_X1 U55 ( .B1(n147), .B2(n145), .A(n142), .ZN(n144) );
  NAND2_X1 U56 ( .A1(n25), .A2(n26), .ZN(n155) );
  XNOR2_X1 U57 ( .A(n463), .B(n462), .ZN(n16) );
  OAI22_X1 U58 ( .A1(n236), .A2(n31), .B1(n237), .B2(n30), .ZN(n39) );
  INV_X1 U59 ( .A(n35), .ZN(n237) );
  AND2_X1 U60 ( .A1(n114), .A2(n113), .ZN(n18) );
  AND2_X1 U61 ( .A1(n269), .A2(n268), .ZN(n19) );
  XNOR2_X1 U63 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n20) );
  XNOR2_X1 U64 ( .A(\mult_x_1/n311 ), .B(n460), .ZN(n35) );
  OR2_X2 U65 ( .A1(n20), .A2(n35), .ZN(n236) );
  XNOR2_X1 U66 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n30) );
  XNOR2_X1 U67 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n50) );
  OAI22_X1 U68 ( .A1(n236), .A2(n30), .B1(n237), .B2(n50), .ZN(n74) );
  BUF_X2 U69 ( .A(n641), .Z(n161) );
  XNOR2_X1 U70 ( .A(n161), .B(\mult_x_1/n281 ), .ZN(n24) );
  AND2_X1 U71 ( .A1(n642), .A2(\mult_x_1/n281 ), .ZN(n182) );
  XNOR2_X1 U72 ( .A(n182), .B(n161), .ZN(n48) );
  OAI22_X1 U73 ( .A1(n162), .A2(n24), .B1(n48), .B2(n466), .ZN(n73) );
  XNOR2_X1 U74 ( .A(n21), .B(n11), .ZN(n83) );
  NOR2_X1 U75 ( .A1(n83), .A2(n474), .ZN(n72) );
  XNOR2_X1 U76 ( .A(n463), .B(n462), .ZN(n23) );
  XNOR2_X1 U77 ( .A(n462), .B(\mult_x_1/n311 ), .ZN(n22) );
  XNOR2_X1 U78 ( .A(n13), .B(\mult_x_1/n286 ), .ZN(n121) );
  INV_X1 U79 ( .A(n16), .ZN(n141) );
  XNOR2_X1 U80 ( .A(n13), .B(\mult_x_1/n285 ), .ZN(n27) );
  OAI22_X1 U81 ( .A1(n9), .A2(n121), .B1(n15), .B2(n27), .ZN(n44) );
  XNOR2_X1 U82 ( .A(n161), .B(\mult_x_1/n282 ), .ZN(n34) );
  OAI22_X1 U83 ( .A1(n162), .A2(n34), .B1(n24), .B2(n466), .ZN(n43) );
  XNOR2_X1 U84 ( .A(\mult_x_1/n312 ), .B(n464), .ZN(n25) );
  XNOR2_X1 U85 ( .A(n641), .B(\mult_x_1/a[2] ), .ZN(n26) );
  XNOR2_X1 U86 ( .A(n7), .B(\mult_x_1/n284 ), .ZN(n33) );
  BUF_X2 U87 ( .A(n26), .Z(n157) );
  XNOR2_X1 U88 ( .A(n7), .B(\mult_x_1/n283 ), .ZN(n28) );
  OAI22_X1 U89 ( .A1(n12), .A2(n33), .B1(n157), .B2(n28), .ZN(n42) );
  XNOR2_X1 U90 ( .A(n13), .B(\mult_x_1/n284 ), .ZN(n52) );
  OAI22_X1 U91 ( .A1(n9), .A2(n27), .B1(n15), .B2(n52), .ZN(n112) );
  XNOR2_X1 U92 ( .A(n7), .B(\mult_x_1/n282 ), .ZN(n51) );
  OAI22_X1 U93 ( .A1(n12), .A2(n28), .B1(n157), .B2(n51), .ZN(n111) );
  OR2_X1 U94 ( .A1(\mult_x_1/n288 ), .A2(n459), .ZN(n29) );
  OAI22_X1 U95 ( .A1(n236), .A2(n459), .B1(n29), .B2(n237), .ZN(n41) );
  XNOR2_X1 U96 ( .A(n11), .B(\mult_x_1/n288 ), .ZN(n31) );
  XNOR2_X1 U97 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n130) );
  OAI22_X1 U98 ( .A1(n12), .A2(n130), .B1(n157), .B2(n33), .ZN(n126) );
  XNOR2_X1 U99 ( .A(n161), .B(\mult_x_1/n283 ), .ZN(n131) );
  OAI22_X1 U100 ( .A1(n162), .A2(n131), .B1(n34), .B2(n466), .ZN(n124) );
  AND2_X1 U101 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n123) );
  XNOR2_X1 U102 ( .A(n41), .B(n40), .ZN(n206) );
  FA_X1 U103 ( .A(n44), .B(n43), .CI(n42), .CO(n266), .S(n205) );
  NAND2_X1 U104 ( .A1(n221), .A2(n220), .ZN(n45) );
  INV_X1 U105 ( .A(en), .ZN(n316) );
  NAND2_X1 U106 ( .A1(n45), .A2(n356), .ZN(n47) );
  NAND2_X1 U107 ( .A1(n315), .A2(n397), .ZN(n46) );
  NAND2_X1 U108 ( .A1(n47), .A2(n46), .ZN(n427) );
  AOI21_X1 U109 ( .B1(n162), .B2(n466), .A(n48), .ZN(n49) );
  INV_X1 U110 ( .A(n49), .ZN(n109) );
  XNOR2_X1 U111 ( .A(n11), .B(\mult_x_1/n285 ), .ZN(n60) );
  OAI22_X1 U112 ( .A1(n236), .A2(n50), .B1(n237), .B2(n60), .ZN(n108) );
  NOR2_X1 U113 ( .A1(n473), .A2(n83), .ZN(n107) );
  INV_X1 U114 ( .A(n67), .ZN(n94) );
  XNOR2_X1 U115 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n53) );
  OAI22_X1 U116 ( .A1(n12), .A2(n51), .B1(n157), .B2(n53), .ZN(n75) );
  XNOR2_X1 U117 ( .A(n13), .B(\mult_x_1/n283 ), .ZN(n58) );
  OAI22_X1 U118 ( .A1(n8), .A2(n52), .B1(n15), .B2(n58), .ZN(n76) );
  NOR2_X1 U119 ( .A1(n472), .A2(n83), .ZN(n64) );
  NOR2_X1 U120 ( .A1(n65), .A2(n64), .ZN(n93) );
  NAND2_X1 U121 ( .A1(n64), .A2(n65), .ZN(n92) );
  OAI21_X1 U122 ( .B1(n94), .B2(n93), .A(n92), .ZN(n56) );
  XNOR2_X1 U123 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n59) );
  XNOR2_X1 U124 ( .A(n11), .B(\mult_x_1/n283 ), .ZN(n84) );
  OAI22_X1 U125 ( .A1(n236), .A2(n59), .B1(n237), .B2(n84), .ZN(n88) );
  XNOR2_X1 U126 ( .A(n182), .B(\mult_x_1/n312 ), .ZN(n54) );
  OAI22_X1 U127 ( .A1(n155), .A2(n53), .B1(n54), .B2(n157), .ZN(n87) );
  AOI21_X1 U128 ( .B1(n157), .B2(n12), .A(n54), .ZN(n55) );
  INV_X1 U129 ( .A(n55), .ZN(n86) );
  XNOR2_X1 U130 ( .A(n56), .B(n97), .ZN(n63) );
  CLKBUF_X1 U131 ( .A(n83), .Z(n239) );
  NOR2_X1 U132 ( .A1(n471), .A2(n239), .ZN(n91) );
  XNOR2_X1 U133 ( .A(n13), .B(\mult_x_1/n282 ), .ZN(n57) );
  XNOR2_X1 U134 ( .A(n13), .B(\mult_x_1/n281 ), .ZN(n85) );
  OAI22_X1 U135 ( .A1(n8), .A2(n57), .B1(n15), .B2(n85), .ZN(n90) );
  OAI22_X1 U136 ( .A1(n8), .A2(n58), .B1(n187), .B2(n57), .ZN(n68) );
  OAI22_X1 U137 ( .A1(n236), .A2(n60), .B1(n237), .B2(n59), .ZN(n69) );
  INV_X1 U138 ( .A(n87), .ZN(n70) );
  OAI21_X1 U139 ( .B1(n68), .B2(n69), .A(n70), .ZN(n62) );
  NAND2_X1 U140 ( .A1(n69), .A2(n68), .ZN(n61) );
  NAND2_X1 U141 ( .A1(n62), .A2(n61), .ZN(n89) );
  XNOR2_X1 U142 ( .A(n63), .B(n95), .ZN(n255) );
  XNOR2_X1 U143 ( .A(n65), .B(n64), .ZN(n66) );
  XNOR2_X1 U144 ( .A(n67), .B(n66), .ZN(n105) );
  XNOR2_X1 U145 ( .A(n69), .B(n68), .ZN(n71) );
  FA_X1 U146 ( .A(n74), .B(n73), .CI(n72), .CO(n114), .S(n267) );
  XNOR2_X1 U147 ( .A(n76), .B(n75), .ZN(n113) );
  NAND2_X1 U148 ( .A1(n255), .A2(n256), .ZN(n79) );
  NAND2_X1 U149 ( .A1(n79), .A2(n356), .ZN(n82) );
  INV_X1 U150 ( .A(n6), .ZN(n80) );
  NAND2_X1 U151 ( .A1(n80), .A2(n393), .ZN(n81) );
  NAND2_X1 U152 ( .A1(n82), .A2(n81), .ZN(n419) );
  NOR2_X1 U153 ( .A1(n470), .A2(n83), .ZN(n191) );
  XNOR2_X1 U154 ( .A(n11), .B(\mult_x_1/n282 ), .ZN(n184) );
  OAI22_X1 U155 ( .A1(n236), .A2(n84), .B1(n237), .B2(n184), .ZN(n190) );
  XNOR2_X1 U156 ( .A(n182), .B(\mult_x_1/n311 ), .ZN(n185) );
  OAI22_X1 U157 ( .A1(n9), .A2(n85), .B1(n185), .B2(n187), .ZN(n192) );
  INV_X1 U158 ( .A(n192), .ZN(n189) );
  FA_X1 U159 ( .A(n88), .B(n17), .CI(n86), .CO(n201), .S(n97) );
  FA_X1 U160 ( .A(n91), .B(n90), .CI(n89), .CO(n200), .S(n95) );
  NAND2_X1 U161 ( .A1(n95), .A2(n97), .ZN(n100) );
  OAI21_X1 U162 ( .B1(n94), .B2(n93), .A(n92), .ZN(n96) );
  NAND2_X1 U163 ( .A1(n95), .A2(n96), .ZN(n99) );
  NAND2_X1 U164 ( .A1(n97), .A2(n96), .ZN(n98) );
  NAND3_X1 U165 ( .A1(n100), .A2(n99), .A3(n98), .ZN(n251) );
  NAND2_X1 U166 ( .A1(n252), .A2(n251), .ZN(n101) );
  NAND2_X1 U167 ( .A1(n101), .A2(n356), .ZN(n103) );
  NAND2_X1 U168 ( .A1(n5), .A2(n391), .ZN(n102) );
  NAND2_X1 U169 ( .A1(n103), .A2(n102), .ZN(n415) );
  XNOR2_X1 U170 ( .A(n18), .B(n104), .ZN(n106) );
  XNOR2_X1 U171 ( .A(n106), .B(n105), .ZN(n181) );
  FA_X1 U172 ( .A(n109), .B(n108), .CI(n107), .CO(n67), .S(n263) );
  FA_X1 U173 ( .A(n112), .B(n111), .CI(n110), .CO(n262), .S(n265) );
  INV_X1 U174 ( .A(n113), .ZN(n115) );
  XNOR2_X1 U175 ( .A(n115), .B(n114), .ZN(n261) );
  NAND2_X1 U176 ( .A1(n181), .A2(n178), .ZN(n116) );
  NAND2_X1 U177 ( .A1(n116), .A2(n356), .ZN(n118) );
  NAND2_X1 U178 ( .A1(n315), .A2(n399), .ZN(n117) );
  NAND2_X1 U179 ( .A1(n118), .A2(n117), .ZN(n431) );
  OR2_X1 U180 ( .A1(\mult_x_1/n288 ), .A2(n461), .ZN(n119) );
  OAI22_X1 U181 ( .A1(n186), .A2(n461), .B1(n119), .B2(n187), .ZN(n129) );
  XNOR2_X1 U182 ( .A(n13), .B(\mult_x_1/n288 ), .ZN(n120) );
  XNOR2_X1 U183 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n122) );
  OAI22_X1 U184 ( .A1(n186), .A2(n120), .B1(n187), .B2(n122), .ZN(n128) );
  OAI22_X1 U185 ( .A1(n8), .A2(n122), .B1(n15), .B2(n121), .ZN(n210) );
  XNOR2_X1 U186 ( .A(n211), .B(n210), .ZN(n127) );
  XNOR2_X1 U187 ( .A(n124), .B(n123), .ZN(n125) );
  XNOR2_X1 U188 ( .A(n126), .B(n125), .ZN(n209) );
  XNOR2_X1 U189 ( .A(n127), .B(n209), .ZN(n175) );
  HA_X1 U190 ( .A(n129), .B(n128), .CO(n211), .S(n138) );
  XNOR2_X1 U191 ( .A(n7), .B(\mult_x_1/n286 ), .ZN(n139) );
  OAI22_X1 U192 ( .A1(n155), .A2(n139), .B1(n157), .B2(n130), .ZN(n136) );
  XNOR2_X1 U193 ( .A(n161), .B(\mult_x_1/n284 ), .ZN(n140) );
  OAI22_X1 U194 ( .A1(n162), .A2(n140), .B1(n131), .B2(n466), .ZN(n135) );
  OR2_X1 U195 ( .A1(n175), .A2(n174), .ZN(n275) );
  XNOR2_X1 U196 ( .A(n138), .B(n137), .ZN(n172) );
  XNOR2_X1 U197 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n149) );
  OAI22_X1 U198 ( .A1(n12), .A2(n149), .B1(n157), .B2(n139), .ZN(n147) );
  XNOR2_X1 U199 ( .A(n161), .B(\mult_x_1/n285 ), .ZN(n151) );
  OAI22_X1 U200 ( .A1(n162), .A2(n151), .B1(n140), .B2(n466), .ZN(n145) );
  NAND2_X1 U201 ( .A1(n14), .A2(\mult_x_1/n288 ), .ZN(n146) );
  XOR2_X1 U202 ( .A(n146), .B(n145), .Z(n148) );
  XNOR2_X1 U203 ( .A(n148), .B(n147), .ZN(n170) );
  XNOR2_X1 U204 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n150) );
  OAI22_X1 U205 ( .A1(n155), .A2(n150), .B1(n157), .B2(n149), .ZN(n153) );
  XNOR2_X1 U206 ( .A(n161), .B(\mult_x_1/n286 ), .ZN(n156) );
  OAI22_X1 U207 ( .A1(n162), .A2(n156), .B1(n151), .B2(n466), .ZN(n152) );
  NOR2_X1 U208 ( .A1(n170), .A2(n169), .ZN(n302) );
  HA_X1 U209 ( .A(n153), .B(n152), .CO(n169), .S(n167) );
  OR2_X1 U210 ( .A1(\mult_x_1/n288 ), .A2(n463), .ZN(n154) );
  OAI22_X1 U211 ( .A1(n12), .A2(n463), .B1(n154), .B2(n157), .ZN(n166) );
  OR2_X1 U212 ( .A1(n166), .A2(n167), .ZN(n297) );
  XNOR2_X1 U213 ( .A(n161), .B(\mult_x_1/n287 ), .ZN(n160) );
  OAI22_X1 U214 ( .A1(n162), .A2(n160), .B1(n156), .B2(n466), .ZN(n165) );
  INV_X1 U215 ( .A(n157), .ZN(n158) );
  AND2_X1 U216 ( .A1(\mult_x_1/n288 ), .A2(n158), .ZN(n164) );
  NOR2_X1 U217 ( .A1(n165), .A2(n164), .ZN(n289) );
  OAI22_X1 U218 ( .A1(n162), .A2(\mult_x_1/n288 ), .B1(n160), .B2(n466), .ZN(
        n285) );
  OR2_X1 U219 ( .A1(\mult_x_1/n288 ), .A2(n465), .ZN(n163) );
  NAND2_X1 U220 ( .A1(n163), .A2(n162), .ZN(n284) );
  NAND2_X1 U221 ( .A1(n285), .A2(n284), .ZN(n292) );
  NAND2_X1 U222 ( .A1(n165), .A2(n164), .ZN(n290) );
  OAI21_X1 U223 ( .B1(n289), .B2(n292), .A(n290), .ZN(n298) );
  NAND2_X1 U224 ( .A1(n167), .A2(n166), .ZN(n296) );
  INV_X1 U225 ( .A(n296), .ZN(n168) );
  AOI21_X1 U226 ( .B1(n297), .B2(n298), .A(n168), .ZN(n305) );
  NAND2_X1 U227 ( .A1(n170), .A2(n169), .ZN(n303) );
  OAI21_X1 U228 ( .B1(n302), .B2(n305), .A(n303), .ZN(n309) );
  NAND2_X1 U229 ( .A1(n10), .A2(n311), .ZN(n173) );
  NAND2_X1 U230 ( .A1(n173), .A2(n310), .ZN(n277) );
  NAND2_X1 U231 ( .A1(n175), .A2(n174), .ZN(n274) );
  INV_X1 U232 ( .A(n178), .ZN(n179) );
  NAND2_X1 U233 ( .A1(n179), .A2(n356), .ZN(n180) );
  OAI22_X1 U234 ( .A1(n181), .A2(n180), .B1(n383), .B2(n441), .ZN(n433) );
  NOR2_X1 U253 ( .A1(n468), .A2(n239), .ZN(n234) );
  XNOR2_X1 U254 ( .A(n11), .B(\mult_x_1/n281 ), .ZN(n183) );
  XNOR2_X1 U255 ( .A(n182), .B(n11), .ZN(n235) );
  OAI22_X1 U256 ( .A1(n236), .A2(n183), .B1(n235), .B2(n237), .ZN(n243) );
  INV_X1 U257 ( .A(n243), .ZN(n233) );
  OAI22_X1 U258 ( .A1(n236), .A2(n184), .B1(n237), .B2(n183), .ZN(n194) );
  AOI21_X1 U259 ( .B1(n15), .B2(n186), .A(n185), .ZN(n188) );
  INV_X1 U260 ( .A(n188), .ZN(n193) );
  FA_X1 U261 ( .A(n191), .B(n190), .CI(n189), .CO(n199), .S(n202) );
  NOR2_X1 U262 ( .A1(n469), .A2(n239), .ZN(n198) );
  FA_X1 U263 ( .A(n194), .B(n193), .CI(n192), .CO(n232), .S(n197) );
  OR2_X1 U264 ( .A1(n217), .A2(n216), .ZN(n195) );
  NAND2_X1 U265 ( .A1(n356), .A2(n195), .ZN(n196) );
  OAI21_X1 U266 ( .B1(n6), .B2(n454), .A(n196), .ZN(n403) );
  FA_X1 U267 ( .A(n199), .B(n198), .CI(n197), .CO(n216), .S(n229) );
  FA_X1 U268 ( .A(n202), .B(n201), .CI(n200), .CO(n228), .S(n252) );
  OR2_X1 U269 ( .A1(n229), .A2(n228), .ZN(n203) );
  NAND2_X1 U270 ( .A1(n6), .A2(n203), .ZN(n204) );
  OAI21_X1 U271 ( .B1(n383), .B2(n453), .A(n204), .ZN(n405) );
  FA_X1 U272 ( .A(n207), .B(n206), .CI(n205), .CO(n220), .S(n225) );
  OR2_X1 U273 ( .A1(n225), .A2(n224), .ZN(n214) );
  NAND2_X1 U274 ( .A1(n381), .A2(n214), .ZN(n215) );
  OAI21_X1 U275 ( .B1(n383), .B2(n451), .A(n215), .ZN(n409) );
  NAND2_X1 U276 ( .A1(n217), .A2(n216), .ZN(n218) );
  NAND2_X1 U277 ( .A1(n381), .A2(n218), .ZN(n219) );
  OAI21_X1 U278 ( .B1(n378), .B2(n449), .A(n219), .ZN(n413) );
  NOR2_X1 U279 ( .A1(n221), .A2(n220), .ZN(n222) );
  NAND2_X1 U280 ( .A1(n356), .A2(n222), .ZN(n223) );
  OAI21_X1 U281 ( .B1(n381), .B2(n443), .A(n223), .ZN(n425) );
  NAND2_X1 U282 ( .A1(n225), .A2(n224), .ZN(n226) );
  NAND2_X1 U283 ( .A1(n356), .A2(n226), .ZN(n227) );
  OAI21_X1 U284 ( .B1(n381), .B2(n442), .A(n227), .ZN(n429) );
  NAND2_X1 U285 ( .A1(n229), .A2(n228), .ZN(n230) );
  NAND2_X1 U286 ( .A1(n356), .A2(n230), .ZN(n231) );
  OAI21_X1 U287 ( .B1(n383), .B2(n440), .A(n231), .ZN(n435) );
  OR2_X1 U288 ( .A1(n6), .A2(n450), .ZN(n250) );
  FA_X1 U289 ( .A(n234), .B(n233), .CI(n232), .CO(n245), .S(n217) );
  AOI21_X1 U290 ( .B1(n237), .B2(n236), .A(n235), .ZN(n238) );
  INV_X1 U291 ( .A(n238), .ZN(n241) );
  NOR2_X1 U292 ( .A1(n467), .A2(n239), .ZN(n240) );
  XOR2_X1 U293 ( .A(n241), .B(n240), .Z(n242) );
  XOR2_X1 U294 ( .A(n243), .B(n242), .Z(n244) );
  OR2_X1 U295 ( .A1(n245), .A2(n244), .ZN(n247) );
  NAND2_X1 U296 ( .A1(n245), .A2(n244), .ZN(n246) );
  NAND2_X1 U297 ( .A1(n247), .A2(n246), .ZN(n248) );
  NAND2_X1 U298 ( .A1(n6), .A2(n248), .ZN(n249) );
  NAND2_X1 U299 ( .A1(n250), .A2(n249), .ZN(n411) );
  OR2_X1 U300 ( .A1(n381), .A2(n452), .ZN(n254) );
  OAI21_X1 U301 ( .B1(n252), .B2(n251), .A(n383), .ZN(n253) );
  NAND2_X1 U302 ( .A1(n254), .A2(n253), .ZN(n407) );
  OR2_X1 U303 ( .A1(n381), .A2(n447), .ZN(n260) );
  INV_X1 U304 ( .A(n255), .ZN(n258) );
  INV_X1 U305 ( .A(n256), .ZN(n257) );
  NAND3_X1 U306 ( .A1(n258), .A2(n257), .A3(n356), .ZN(n259) );
  NAND2_X1 U307 ( .A1(n260), .A2(n259), .ZN(n417) );
  FA_X1 U308 ( .A(n263), .B(n262), .CI(n261), .CO(n178), .S(n273) );
  OR2_X1 U309 ( .A1(n378), .A2(n444), .ZN(n271) );
  NAND2_X1 U310 ( .A1(n19), .A2(n356), .ZN(n270) );
  OAI211_X1 U311 ( .C1(n273), .C2(n5), .A(n271), .B(n270), .ZN(n423) );
  NAND2_X1 U312 ( .A1(n356), .A2(n19), .ZN(n272) );
  OAI22_X1 U313 ( .A1(n273), .A2(n272), .B1(n383), .B2(n445), .ZN(n421) );
  INV_X1 U314 ( .A(rst_n), .ZN(n643) );
  NAND2_X1 U315 ( .A1(n275), .A2(n274), .ZN(n276) );
  XNOR2_X1 U316 ( .A(n277), .B(n276), .ZN(n278) );
  INV_X2 U317 ( .A(n281), .ZN(n381) );
  NAND2_X1 U318 ( .A1(n278), .A2(n381), .ZN(n280) );
  INV_X2 U319 ( .A(n281), .ZN(n378) );
  NAND2_X1 U320 ( .A1(n5), .A2(n455), .ZN(n279) );
  NAND2_X1 U321 ( .A1(n280), .A2(n279), .ZN(n554) );
  BUF_X2 U322 ( .A(n281), .Z(n315) );
  AOI22_X1 U323 ( .A1(n356), .A2(n512), .B1(n513), .B2(n315), .ZN(n515) );
  AOI22_X1 U324 ( .A1(n356), .A2(n511), .B1(n512), .B2(n315), .ZN(n517) );
  INV_X4 U325 ( .A(n281), .ZN(n383) );
  AND2_X1 U326 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n282) );
  NAND2_X1 U327 ( .A1(n6), .A2(n282), .ZN(n283) );
  OAI21_X1 U328 ( .B1(n383), .B2(n511), .A(n283), .ZN(n519) );
  AOI22_X1 U329 ( .A1(n356), .A2(n509), .B1(n510), .B2(n315), .ZN(n521) );
  AOI22_X1 U330 ( .A1(n356), .A2(n508), .B1(n509), .B2(n315), .ZN(n523) );
  OR2_X1 U331 ( .A1(n285), .A2(n284), .ZN(n286) );
  AND2_X1 U332 ( .A1(n286), .A2(n292), .ZN(n287) );
  NAND2_X1 U333 ( .A1(n383), .A2(n287), .ZN(n288) );
  OAI21_X1 U334 ( .B1(n6), .B2(n508), .A(n288), .ZN(n525) );
  AOI22_X1 U335 ( .A1(n356), .A2(n506), .B1(n507), .B2(n315), .ZN(n527) );
  AOI22_X1 U336 ( .A1(n356), .A2(n505), .B1(n506), .B2(n315), .ZN(n529) );
  INV_X1 U337 ( .A(n289), .ZN(n291) );
  NAND2_X1 U338 ( .A1(n291), .A2(n290), .ZN(n293) );
  XOR2_X1 U339 ( .A(n293), .B(n292), .Z(n294) );
  NAND2_X1 U340 ( .A1(n383), .A2(n294), .ZN(n295) );
  OAI21_X1 U341 ( .B1(n378), .B2(n505), .A(n295), .ZN(n531) );
  AOI22_X1 U342 ( .A1(n356), .A2(n503), .B1(n504), .B2(n315), .ZN(n533) );
  AOI22_X1 U343 ( .A1(n356), .A2(n502), .B1(n503), .B2(n315), .ZN(n535) );
  NAND2_X1 U344 ( .A1(n297), .A2(n296), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  NAND2_X1 U346 ( .A1(n6), .A2(n300), .ZN(n301) );
  OAI21_X1 U347 ( .B1(n383), .B2(n502), .A(n301), .ZN(n537) );
  AOI22_X1 U348 ( .A1(n356), .A2(n500), .B1(n501), .B2(n315), .ZN(n539) );
  AOI22_X1 U349 ( .A1(n356), .A2(n499), .B1(n500), .B2(n315), .ZN(n541) );
  INV_X1 U350 ( .A(n302), .ZN(n304) );
  NAND2_X1 U351 ( .A1(n304), .A2(n303), .ZN(n306) );
  XOR2_X1 U352 ( .A(n306), .B(n305), .Z(n307) );
  NAND2_X1 U353 ( .A1(n383), .A2(n307), .ZN(n308) );
  OAI21_X1 U354 ( .B1(n381), .B2(n499), .A(n308), .ZN(n543) );
  AOI22_X1 U355 ( .A1(n356), .A2(n497), .B1(n498), .B2(n315), .ZN(n545) );
  AOI22_X1 U356 ( .A1(n356), .A2(n496), .B1(n497), .B2(n315), .ZN(n547) );
  NAND2_X1 U357 ( .A1(n311), .A2(n310), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n309), .B(n312), .ZN(n313) );
  NAND2_X1 U359 ( .A1(n378), .A2(n313), .ZN(n314) );
  OAI21_X1 U360 ( .B1(n6), .B2(n496), .A(n314), .ZN(n548) );
  AOI22_X1 U361 ( .A1(n356), .A2(n494), .B1(n495), .B2(n315), .ZN(n550) );
  AOI22_X1 U362 ( .A1(n378), .A2(n493), .B1(n494), .B2(n315), .ZN(n552) );
  AOI22_X1 U363 ( .A1(n378), .A2(n491), .B1(n492), .B2(n315), .ZN(n556) );
  NAND2_X1 U364 ( .A1(n388), .A2(n398), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n402), .B(n317), .ZN(n318) );
  NAND2_X1 U366 ( .A1(n381), .A2(n318), .ZN(n319) );
  OAI21_X1 U367 ( .B1(n378), .B2(n491), .A(n319), .ZN(n558) );
  AOI22_X1 U368 ( .A1(n381), .A2(n489), .B1(n490), .B2(n315), .ZN(n560) );
  AOI21_X1 U369 ( .B1(n402), .B2(n388), .A(n442), .ZN(n323) );
  NAND2_X1 U370 ( .A1(n443), .A2(n397), .ZN(n320) );
  XOR2_X1 U371 ( .A(n323), .B(n320), .Z(n321) );
  NAND2_X1 U372 ( .A1(n6), .A2(n321), .ZN(n322) );
  OAI21_X1 U373 ( .B1(n383), .B2(n489), .A(n322), .ZN(n562) );
  AOI22_X1 U374 ( .A1(n356), .A2(n487), .B1(n488), .B2(n315), .ZN(n564) );
  OAI21_X1 U375 ( .B1(n323), .B2(n396), .A(n397), .ZN(n333) );
  INV_X1 U376 ( .A(n333), .ZN(n327) );
  NAND2_X1 U377 ( .A1(n445), .A2(n395), .ZN(n324) );
  XOR2_X1 U378 ( .A(n327), .B(n324), .Z(n325) );
  NAND2_X1 U379 ( .A1(n383), .A2(n325), .ZN(n326) );
  OAI21_X1 U380 ( .B1(n381), .B2(n487), .A(n326), .ZN(n566) );
  AOI22_X1 U381 ( .A1(n378), .A2(n485), .B1(n486), .B2(n315), .ZN(n568) );
  OAI21_X1 U382 ( .B1(n327), .B2(n394), .A(n395), .ZN(n329) );
  NAND2_X1 U383 ( .A1(n441), .A2(n399), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  NAND2_X1 U385 ( .A1(n381), .A2(n330), .ZN(n331) );
  OAI21_X1 U386 ( .B1(n6), .B2(n485), .A(n331), .ZN(n570) );
  AOI22_X1 U387 ( .A1(n6), .A2(n483), .B1(n484), .B2(n315), .ZN(n572) );
  NOR2_X1 U388 ( .A1(n400), .A2(n394), .ZN(n334) );
  OAI21_X1 U389 ( .B1(n400), .B2(n395), .A(n399), .ZN(n332) );
  AOI21_X1 U390 ( .B1(n334), .B2(n333), .A(n332), .ZN(n361) );
  NAND2_X1 U391 ( .A1(n447), .A2(n393), .ZN(n335) );
  XOR2_X1 U392 ( .A(n361), .B(n335), .Z(n336) );
  NAND2_X1 U393 ( .A1(n383), .A2(n336), .ZN(n337) );
  OAI21_X1 U394 ( .B1(n383), .B2(n483), .A(n337), .ZN(n574) );
  AOI22_X1 U395 ( .A1(n356), .A2(n481), .B1(n482), .B2(n315), .ZN(n576) );
  OAI21_X1 U396 ( .B1(n361), .B2(n392), .A(n393), .ZN(n339) );
  NAND2_X1 U397 ( .A1(n387), .A2(n391), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  NAND2_X1 U399 ( .A1(n383), .A2(n340), .ZN(n341) );
  OAI21_X1 U400 ( .B1(n378), .B2(n481), .A(n341), .ZN(n578) );
  AOI22_X1 U401 ( .A1(n356), .A2(n479), .B1(n480), .B2(n315), .ZN(n580) );
  NAND2_X1 U402 ( .A1(n447), .A2(n387), .ZN(n343) );
  AOI21_X1 U403 ( .B1(n446), .B2(n387), .A(n448), .ZN(n342) );
  OAI21_X1 U404 ( .B1(n361), .B2(n343), .A(n342), .ZN(n345) );
  NAND2_X1 U405 ( .A1(n386), .A2(n401), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U407 ( .A1(n6), .A2(n346), .ZN(n347) );
  OAI21_X1 U408 ( .B1(n381), .B2(n479), .A(n347), .ZN(n582) );
  AOI22_X1 U409 ( .A1(n356), .A2(n477), .B1(n478), .B2(n315), .ZN(n584) );
  NAND2_X1 U410 ( .A1(n387), .A2(n386), .ZN(n349) );
  NOR2_X1 U411 ( .A1(n392), .A2(n349), .ZN(n357) );
  INV_X1 U412 ( .A(n357), .ZN(n351) );
  AOI21_X1 U413 ( .B1(n448), .B2(n386), .A(n440), .ZN(n348) );
  OAI21_X1 U414 ( .B1(n349), .B2(n393), .A(n348), .ZN(n358) );
  INV_X1 U415 ( .A(n358), .ZN(n350) );
  OAI21_X1 U416 ( .B1(n361), .B2(n351), .A(n350), .ZN(n353) );
  NAND2_X1 U417 ( .A1(n385), .A2(n390), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  NAND2_X1 U419 ( .A1(n383), .A2(n354), .ZN(n355) );
  OAI21_X1 U420 ( .B1(n6), .B2(n477), .A(n355), .ZN(n586) );
  AOI22_X1 U421 ( .A1(n356), .A2(n475), .B1(n476), .B2(n315), .ZN(n588) );
  NAND2_X1 U422 ( .A1(n357), .A2(n385), .ZN(n360) );
  AOI21_X1 U423 ( .B1(n358), .B2(n385), .A(n449), .ZN(n359) );
  OAI21_X1 U424 ( .B1(n361), .B2(n360), .A(n359), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n362), .B(n389), .ZN(n363) );
  NAND2_X1 U426 ( .A1(n378), .A2(n363), .ZN(n364) );
  OAI21_X1 U427 ( .B1(n6), .B2(n475), .A(n364), .ZN(n590) );
  NAND2_X1 U428 ( .A1(n6), .A2(B_extended[0]), .ZN(n365) );
  OAI21_X1 U429 ( .B1(n378), .B2(n474), .A(n365), .ZN(n592) );
  NAND2_X1 U430 ( .A1(n6), .A2(B_extended[1]), .ZN(n366) );
  OAI21_X1 U431 ( .B1(n383), .B2(n473), .A(n366), .ZN(n594) );
  NAND2_X1 U432 ( .A1(n378), .A2(B_extended[2]), .ZN(n367) );
  OAI21_X1 U433 ( .B1(n381), .B2(n472), .A(n367), .ZN(n596) );
  NAND2_X1 U434 ( .A1(n383), .A2(B_extended[3]), .ZN(n368) );
  OAI21_X1 U435 ( .B1(n378), .B2(n471), .A(n368), .ZN(n598) );
  NAND2_X1 U436 ( .A1(n383), .A2(B_extended[4]), .ZN(n369) );
  OAI21_X1 U437 ( .B1(n383), .B2(n470), .A(n369), .ZN(n600) );
  NAND2_X1 U438 ( .A1(n381), .A2(B_extended[5]), .ZN(n370) );
  OAI21_X1 U439 ( .B1(n381), .B2(n469), .A(n370), .ZN(n602) );
  NAND2_X1 U440 ( .A1(n381), .A2(B_extended[6]), .ZN(n371) );
  OAI21_X1 U441 ( .B1(n6), .B2(n468), .A(n371), .ZN(n604) );
  NAND2_X1 U442 ( .A1(n378), .A2(B_extended[7]), .ZN(n372) );
  OAI21_X1 U443 ( .B1(n378), .B2(n467), .A(n372), .ZN(n606) );
  NAND2_X1 U444 ( .A1(n6), .A2(A_extended[0]), .ZN(n373) );
  OAI21_X1 U445 ( .B1(n383), .B2(n466), .A(n373), .ZN(n608) );
  NAND2_X1 U446 ( .A1(n383), .A2(A_extended[1]), .ZN(n374) );
  OAI21_X1 U447 ( .B1(n381), .B2(n465), .A(n374), .ZN(n610) );
  NAND2_X1 U448 ( .A1(n378), .A2(A_extended[2]), .ZN(n375) );
  OAI21_X1 U449 ( .B1(n6), .B2(n464), .A(n375), .ZN(n612) );
  NAND2_X1 U450 ( .A1(n6), .A2(A_extended[3]), .ZN(n376) );
  OAI21_X1 U451 ( .B1(n378), .B2(n463), .A(n376), .ZN(n614) );
  NAND2_X1 U452 ( .A1(n378), .A2(A_extended[4]), .ZN(n377) );
  OAI21_X1 U453 ( .B1(n383), .B2(n462), .A(n377), .ZN(n616) );
  NAND2_X1 U454 ( .A1(n381), .A2(A_extended[5]), .ZN(n379) );
  OAI21_X1 U455 ( .B1(n381), .B2(n461), .A(n379), .ZN(n618) );
  NAND2_X1 U456 ( .A1(n381), .A2(A_extended[6]), .ZN(n380) );
  OAI21_X1 U457 ( .B1(n6), .B2(n460), .A(n380), .ZN(n620) );
  NAND2_X1 U458 ( .A1(n383), .A2(A_extended[7]), .ZN(n382) );
  OAI21_X1 U459 ( .B1(n383), .B2(n459), .A(n382), .ZN(n622) );
  NAND2_X1 U460 ( .A1(n458), .A2(n315), .ZN(n624) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_30 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n425,
         n427, n429, n431, n433, n435, n437, n439, n441, n443, n445, n447,
         n449, n451, n453, n455, n457, n459, n460, n461, n462, n463, n464,
         n465, n466, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n538, n540, n542, n544, n546, n548,
         n550, n552, n554, n556, n558, n560, n562, n564, n566, n568, n570,
         n572, n574, n576, n578, n580, n582, n584, n586, n588, n590, n592,
         n594, n596, n598, n600, n602, n604, n606, n608, n610, n612, n614,
         n616, n618, n620, n622, n624, n626, n628, n630, n632, n634, n636,
         n638, n640, n642, n644, n646, n648, n665, n666, n667;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n648), .CK(clk), .Q(n666), 
        .QN(n481) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n480), .SE(n644), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n483) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n480), .SE(n642), .CK(clk), .Q(n665), 
        .QN(n484) );
  SDFF_X1 clk_r_REG45_S1 ( .D(1'b0), .SI(n480), .SE(n640), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n485) );
  SDFF_X1 clk_r_REG53_S1 ( .D(1'b0), .SI(n480), .SE(n636), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n487) );
  SDFF_X1 clk_r_REG61_S1 ( .D(1'b0), .SI(n480), .SE(n632), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n489) );
  SDFF_X1 clk_r_REG65_S1 ( .D(1'b0), .SI(n480), .SE(n630), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n490) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n480), .SE(n628), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n491) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n480), .SE(n626), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n492) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n624), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n493) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n622), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n494) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n620), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n495) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n618), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n496) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n616), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n497) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n5), .SE(n614), .CK(clk), .QN(n498)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(rst_n), .SE(n612), .CK(clk), .Q(
        product[15]), .QN(n499) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n5), .SE(n610), .CK(clk), .QN(n500)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(rst_n), .SE(n608), .CK(clk), .Q(
        product[14]), .QN(n501) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(rst_n), .SE(n606), .CK(clk), .QN(n502) );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(rst_n), .SE(n604), .CK(clk), .Q(
        product[13]), .QN(n503) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n479), .SE(n602), .CK(clk), .QN(n504)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n479), .SE(n600), .CK(clk), .Q(
        product[12]), .QN(n505) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n479), .SE(n598), .CK(clk), .QN(n506)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n479), .SE(n596), .CK(clk), .Q(
        product[11]), .QN(n507) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n479), .SE(n594), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n479), .SE(n592), .CK(clk), .Q(
        product[10]), .QN(n509) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n479), .SE(n590), .CK(clk), .QN(n510)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n479), .SE(n588), .CK(clk), .Q(
        product[9]), .QN(n511) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n479), .SE(n586), .CK(clk), .QN(n512)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n479), .SE(n584), .CK(clk), .Q(
        product[8]), .QN(n513) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n479), .SE(n582), .CK(clk), .QN(n514)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n478), .SE(n580), .CK(clk), .Q(
        product[7]), .QN(n515) );
  SDFF_X1 clk_r_REG37_S2 ( .D(1'b0), .SI(n478), .SE(n578), .CK(clk), .QN(n516)
         );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n478), .SE(n576), .CK(clk), .QN(n517)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n478), .SE(n574), .CK(clk), .Q(
        product[6]), .QN(n518) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n478), .SE(n572), .CK(clk), .QN(n519)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n478), .SE(n570), .CK(clk), .QN(n520)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n478), .SE(n568), .CK(clk), .Q(
        product[5]), .QN(n521) );
  SDFF_X1 clk_r_REG46_S2 ( .D(1'b0), .SI(n478), .SE(n566), .CK(clk), .QN(n522)
         );
  SDFF_X1 clk_r_REG47_S3 ( .D(1'b0), .SI(n478), .SE(n564), .CK(clk), .QN(n523)
         );
  SDFF_X1 clk_r_REG48_S4 ( .D(1'b0), .SI(n478), .SE(n562), .CK(clk), .Q(
        product[4]), .QN(n524) );
  SDFF_X1 clk_r_REG50_S2 ( .D(1'b0), .SI(n478), .SE(n560), .CK(clk), .QN(n525)
         );
  SDFF_X1 clk_r_REG51_S3 ( .D(1'b0), .SI(n477), .SE(n558), .CK(clk), .QN(n526)
         );
  SDFF_X1 clk_r_REG52_S4 ( .D(1'b0), .SI(n477), .SE(n556), .CK(clk), .Q(
        product[3]), .QN(n527) );
  SDFF_X1 clk_r_REG54_S2 ( .D(1'b0), .SI(n477), .SE(n554), .CK(clk), .QN(n528)
         );
  SDFF_X1 clk_r_REG55_S3 ( .D(1'b0), .SI(n477), .SE(n552), .CK(clk), .QN(n529)
         );
  SDFF_X1 clk_r_REG56_S4 ( .D(1'b0), .SI(n477), .SE(n550), .CK(clk), .Q(
        product[2]), .QN(n530) );
  SDFF_X1 clk_r_REG58_S2 ( .D(1'b0), .SI(n477), .SE(n548), .CK(clk), .QN(n531)
         );
  SDFF_X1 clk_r_REG59_S3 ( .D(1'b0), .SI(n477), .SE(n546), .CK(clk), .QN(n532)
         );
  SDFF_X1 clk_r_REG60_S4 ( .D(1'b0), .SI(n477), .SE(n544), .CK(clk), .Q(
        product[1]), .QN(n533) );
  SDFF_X1 clk_r_REG62_S2 ( .D(1'b0), .SI(n477), .SE(n542), .CK(clk), .QN(n534)
         );
  SDFF_X1 clk_r_REG63_S3 ( .D(1'b0), .SI(n477), .SE(n540), .CK(clk), .QN(n535)
         );
  SDFF_X1 clk_r_REG64_S4 ( .D(1'b0), .SI(n477), .SE(n538), .CK(clk), .Q(
        product[0]), .QN(n536) );
  SDFF_X1 clk_r_REG57_S1 ( .D(1'b0), .SI(n480), .SE(n634), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n488) );
  SDFF_X1 clk_r_REG49_S1 ( .D(1'b0), .SI(n480), .SE(n638), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n486) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n667), .SI(1'b1), .SE(n437), .CK(clk), 
        .Q(n412), .QN(n469) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n667), .SI(1'b1), .SE(n457), .CK(clk), 
        .Q(n422), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n667), .SI(1'b1), .SE(n455), .CK(clk), 
        .Q(n421), .QN(n460) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n667), .SE(n453), .CK(
        clk), .Q(n461), .QN(n420) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n667), .SI(1'b1), .SE(n451), .CK(clk), 
        .Q(n419), .QN(n462) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n667), .SE(n449), .CK(
        clk), .Q(n463), .QN(n418) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n667), .SI(1'b1), .SE(n447), .CK(clk), 
        .Q(n417), .QN(n464) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n667), .SI(1'b1), .SE(n445), .CK(clk), 
        .Q(n416), .QN(n465) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n667), .SI(1'b1), .SE(n443), .CK(clk), 
        .Q(n415), .QN(n466) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n667), .SI(1'b1), .SE(n441), .CK(clk), 
        .Q(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n667), .SI(1'b1), .SE(n439), .CK(clk), 
        .Q(n413), .QN(n468) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n667), .SI(1'b1), .SE(n435), .CK(clk), 
        .Q(n411), .QN(n470) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n667), .SI(1'b1), .SE(n433), .CK(clk), 
        .Q(n410), .QN(n471) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n667), .SI(1'b1), .SE(n431), .CK(clk), 
        .Q(n409), .QN(n472) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n667), .SE(n429), .CK(
        clk), .Q(n473), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n667), .SE(n427), .CK(
        clk), .Q(n474), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n667), .SI(1'b1), .SE(n425), .CK(clk), 
        .Q(n406), .QN(n475) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n667), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n405), .QN(n476) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n480), .SE(n646), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n482) );
  BUF_X1 U2 ( .A(rst_n), .Z(n5) );
  INV_X1 U3 ( .A(rst_n), .ZN(n667) );
  BUF_X1 U4 ( .A(n93), .Z(n185) );
  NOR2_X2 U5 ( .A1(n481), .A2(n482), .ZN(n238) );
  XNOR2_X1 U6 ( .A(\mult_x_1/a[6] ), .B(n665), .ZN(n6) );
  XNOR2_X1 U7 ( .A(\mult_x_1/a[6] ), .B(n665), .ZN(n93) );
  BUF_X2 U8 ( .A(n138), .Z(n152) );
  BUF_X1 U9 ( .A(n78), .Z(n143) );
  INV_X1 U10 ( .A(n107), .ZN(n103) );
  OAI22_X1 U11 ( .A1(n92), .A2(n91), .B1(n90), .B2(n89), .ZN(n162) );
  INV_X1 U12 ( .A(n175), .ZN(n171) );
  XNOR2_X1 U13 ( .A(n97), .B(n160), .ZN(n173) );
  XNOR2_X1 U14 ( .A(n162), .B(n161), .ZN(n97) );
  CLKBUF_X1 U15 ( .A(n233), .Z(n19) );
  NAND2_X1 U16 ( .A1(n287), .A2(n286), .ZN(n291) );
  NAND2_X1 U17 ( .A1(n285), .A2(n284), .ZN(n286) );
  NAND2_X1 U18 ( .A1(n273), .A2(n272), .ZN(n277) );
  NAND2_X1 U19 ( .A1(n271), .A2(n270), .ZN(n272) );
  INV_X1 U20 ( .A(n274), .ZN(n271) );
  INV_X1 U21 ( .A(n275), .ZN(n270) );
  CLKBUF_X1 U22 ( .A(n184), .Z(n9) );
  NAND2_X1 U23 ( .A1(n263), .A2(n242), .ZN(n244) );
  NAND2_X1 U24 ( .A1(n110), .A2(n109), .ZN(n111) );
  NAND2_X1 U25 ( .A1(n104), .A2(n103), .ZN(n105) );
  AND2_X1 U26 ( .A1(n73), .A2(n72), .ZN(n74) );
  NAND2_X1 U27 ( .A1(n164), .A2(n163), .ZN(n207) );
  NAND2_X1 U28 ( .A1(n162), .A2(n161), .ZN(n163) );
  OAI21_X1 U29 ( .B1(n162), .B2(n161), .A(n160), .ZN(n164) );
  NAND2_X1 U30 ( .A1(n177), .A2(n176), .ZN(n217) );
  NAND2_X1 U31 ( .A1(n173), .A2(n172), .ZN(n177) );
  NAND2_X1 U32 ( .A1(n171), .A2(n170), .ZN(n172) );
  INV_X1 U33 ( .A(n10), .ZN(n312) );
  INV_X2 U34 ( .A(n318), .ZN(n403) );
  INV_X1 U35 ( .A(n53), .ZN(n54) );
  OAI21_X1 U36 ( .B1(n247), .B2(n246), .A(n255), .ZN(n245) );
  CLKBUF_X1 U37 ( .A(n292), .Z(n7) );
  NAND2_X1 U38 ( .A1(n277), .A2(n276), .ZN(n278) );
  NAND2_X1 U39 ( .A1(n275), .A2(n274), .ZN(n276) );
  BUF_X1 U40 ( .A(n5), .Z(n477) );
  BUF_X1 U41 ( .A(n5), .Z(n478) );
  BUF_X1 U42 ( .A(n5), .Z(n479) );
  BUF_X1 U43 ( .A(n5), .Z(n480) );
  NAND2_X1 U44 ( .A1(n215), .A2(n54), .ZN(n55) );
  NAND2_X1 U45 ( .A1(n404), .A2(n414), .ZN(n8) );
  NAND2_X1 U46 ( .A1(n8), .A2(n216), .ZN(n441) );
  AND2_X1 U47 ( .A1(n68), .A2(n67), .ZN(n10) );
  INV_X1 U48 ( .A(n29), .ZN(n11) );
  XNOR2_X1 U49 ( .A(n485), .B(n665), .ZN(n21) );
  XNOR2_X1 U50 ( .A(n173), .B(n102), .ZN(n112) );
  BUF_X2 U51 ( .A(n138), .Z(n60) );
  INV_X1 U52 ( .A(n89), .ZN(n12) );
  OAI22_X1 U53 ( .A1(n76), .A2(n141), .B1(n78), .B2(n484), .ZN(n101) );
  AND2_X1 U54 ( .A1(n13), .A2(n29), .ZN(n261) );
  XOR2_X1 U55 ( .A(n238), .B(\mult_x_1/n286 ), .Z(n13) );
  NAND2_X1 U56 ( .A1(n106), .A2(n105), .ZN(n110) );
  XNOR2_X1 U57 ( .A(n106), .B(n82), .ZN(n87) );
  OR2_X1 U58 ( .A1(n295), .A2(n462), .ZN(n14) );
  NAND2_X1 U59 ( .A1(n14), .A2(n249), .ZN(n451) );
  OAI22_X1 U60 ( .A1(n56), .A2(n55), .B1(n293), .B2(n470), .ZN(n435) );
  XNOR2_X1 U61 ( .A(n108), .B(n107), .ZN(n82) );
  INV_X1 U62 ( .A(n108), .ZN(n104) );
  NAND2_X1 U63 ( .A1(n108), .A2(n107), .ZN(n109) );
  NAND2_X1 U64 ( .A1(n244), .A2(n243), .ZN(n280) );
  OR2_X1 U65 ( .A1(n241), .A2(n240), .ZN(n260) );
  AND2_X1 U66 ( .A1(n15), .A2(n26), .ZN(n157) );
  XOR2_X1 U67 ( .A(n238), .B(\mult_x_1/n284 ), .Z(n15) );
  INV_X1 U68 ( .A(n26), .ZN(n239) );
  NAND2_X2 U69 ( .A1(n89), .A2(n17), .ZN(n92) );
  BUF_X1 U70 ( .A(\mult_x_1/n310 ), .Z(n16) );
  INV_X1 U71 ( .A(n488), .ZN(n17) );
  INV_X1 U72 ( .A(n62), .ZN(n18) );
  INV_X1 U73 ( .A(n62), .ZN(n153) );
  OAI22_X1 U74 ( .A1(n152), .A2(n96), .B1(n18), .B2(n95), .ZN(n160) );
  XNOR2_X1 U75 ( .A(n175), .B(n174), .ZN(n102) );
  INV_X1 U76 ( .A(n174), .ZN(n170) );
  NAND2_X1 U77 ( .A1(n175), .A2(n174), .ZN(n176) );
  AND2_X1 U78 ( .A1(n20), .A2(n29), .ZN(n229) );
  XOR2_X1 U79 ( .A(n238), .B(\mult_x_1/n285 ), .Z(n20) );
  OAI21_X1 U80 ( .B1(n285), .B2(n284), .A(n283), .ZN(n287) );
  OR2_X1 U81 ( .A1(n261), .A2(n260), .ZN(n242) );
  NAND2_X1 U82 ( .A1(n261), .A2(n260), .ZN(n243) );
  INV_X1 U83 ( .A(n318), .ZN(n399) );
  XNOR2_X1 U84 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n22) );
  NAND2_X1 U85 ( .A1(n21), .A2(n22), .ZN(n78) );
  BUF_X2 U86 ( .A(n665), .Z(n134) );
  XNOR2_X1 U87 ( .A(n134), .B(\mult_x_1/n284 ), .ZN(n34) );
  INV_X1 U88 ( .A(n22), .ZN(n70) );
  INV_X2 U89 ( .A(n70), .ZN(n141) );
  XNOR2_X1 U90 ( .A(n134), .B(\mult_x_1/n283 ), .ZN(n135) );
  OAI22_X1 U91 ( .A1(n78), .A2(n34), .B1(n141), .B2(n135), .ZN(n241) );
  XOR2_X1 U92 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n23) );
  XNOR2_X1 U93 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n24) );
  NAND2_X1 U94 ( .A1(n23), .A2(n24), .ZN(n138) );
  BUF_X2 U95 ( .A(\mult_x_1/n312 ), .Z(n136) );
  XNOR2_X1 U96 ( .A(n136), .B(\mult_x_1/n282 ), .ZN(n35) );
  INV_X1 U97 ( .A(n24), .ZN(n62) );
  XNOR2_X1 U98 ( .A(n136), .B(\mult_x_1/n281 ), .ZN(n139) );
  OAI22_X1 U99 ( .A1(n60), .A2(n35), .B1(n153), .B2(n139), .ZN(n240) );
  XNOR2_X1 U100 ( .A(n241), .B(n240), .ZN(n259) );
  INV_X1 U101 ( .A(n238), .ZN(n25) );
  OR2_X1 U102 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n27) );
  INV_X1 U103 ( .A(\mult_x_1/n310 ), .ZN(n37) );
  XNOR2_X1 U104 ( .A(n238), .B(n37), .ZN(n26) );
  NOR2_X1 U105 ( .A1(n27), .A2(n11), .ZN(n258) );
  XOR2_X1 U106 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n28) );
  NAND2_X2 U107 ( .A1(n28), .A2(n6), .ZN(n184) );
  XNOR2_X1 U108 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n38) );
  XNOR2_X1 U109 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n32) );
  OAI22_X1 U110 ( .A1(n184), .A2(n38), .B1(n185), .B2(n32), .ZN(n43) );
  INV_X2 U111 ( .A(\mult_x_1/n180 ), .ZN(n89) );
  BUF_X2 U112 ( .A(\mult_x_1/n313 ), .Z(n80) );
  XNOR2_X1 U113 ( .A(n80), .B(\mult_x_1/n281 ), .ZN(n45) );
  AND2_X1 U114 ( .A1(n666), .A2(\mult_x_1/n281 ), .ZN(n137) );
  XNOR2_X1 U115 ( .A(n137), .B(n80), .ZN(n30) );
  OAI22_X1 U116 ( .A1(n92), .A2(n45), .B1(n30), .B2(n89), .ZN(n42) );
  XNOR2_X1 U117 ( .A(n238), .B(n37), .ZN(n29) );
  AND2_X1 U118 ( .A1(n29), .A2(\mult_x_1/n288 ), .ZN(n41) );
  AOI21_X1 U119 ( .B1(n92), .B2(n89), .A(n30), .ZN(n31) );
  INV_X1 U120 ( .A(n31), .ZN(n237) );
  XNOR2_X1 U121 ( .A(n16), .B(\mult_x_1/n285 ), .ZN(n133) );
  OAI22_X1 U122 ( .A1(n184), .A2(n32), .B1(n185), .B2(n133), .ZN(n236) );
  XNOR2_X1 U123 ( .A(n238), .B(\mult_x_1/n287 ), .ZN(n33) );
  NOR2_X1 U124 ( .A1(n33), .A2(n239), .ZN(n235) );
  XNOR2_X1 U125 ( .A(n134), .B(\mult_x_1/n285 ), .ZN(n44) );
  OAI22_X1 U126 ( .A1(n143), .A2(n44), .B1(n141), .B2(n34), .ZN(n49) );
  XNOR2_X1 U127 ( .A(n136), .B(\mult_x_1/n283 ), .ZN(n46) );
  OAI22_X1 U128 ( .A1(n60), .A2(n46), .B1(n18), .B2(n35), .ZN(n48) );
  OR2_X1 U129 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n36) );
  OAI22_X1 U130 ( .A1(n184), .A2(n37), .B1(n36), .B2(n185), .ZN(n166) );
  XNOR2_X1 U131 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n39) );
  OAI22_X1 U132 ( .A1(n184), .A2(n39), .B1(n185), .B2(n38), .ZN(n165) );
  XNOR2_X1 U133 ( .A(n275), .B(n274), .ZN(n40) );
  XNOR2_X1 U134 ( .A(n273), .B(n40), .ZN(n56) );
  FA_X1 U135 ( .A(n43), .B(n42), .CI(n41), .CO(n257), .S(n204) );
  XNOR2_X1 U136 ( .A(n134), .B(\mult_x_1/n286 ), .ZN(n98) );
  OAI22_X1 U137 ( .A1(n143), .A2(n98), .B1(n141), .B2(n44), .ZN(n169) );
  XNOR2_X1 U138 ( .A(n80), .B(\mult_x_1/n282 ), .ZN(n90) );
  OAI22_X1 U139 ( .A1(n92), .A2(n90), .B1(n45), .B2(n89), .ZN(n168) );
  XNOR2_X1 U140 ( .A(n136), .B(\mult_x_1/n284 ), .ZN(n95) );
  OAI22_X1 U141 ( .A1(n60), .A2(n95), .B1(n18), .B2(n46), .ZN(n167) );
  FA_X1 U142 ( .A(n49), .B(n48), .CI(n47), .CO(n274), .S(n202) );
  NAND2_X1 U143 ( .A1(n56), .A2(n53), .ZN(n50) );
  INV_X1 U144 ( .A(en), .ZN(n116) );
  INV_X4 U145 ( .A(n116), .ZN(n374) );
  BUF_X1 U146 ( .A(n374), .Z(n215) );
  NAND2_X1 U147 ( .A1(n50), .A2(n215), .ZN(n52) );
  BUF_X2 U148 ( .A(n374), .Z(n293) );
  OR2_X1 U149 ( .A1(n293), .A2(n469), .ZN(n51) );
  NAND2_X1 U150 ( .A1(n52), .A2(n51), .ZN(n437) );
  XNOR2_X1 U151 ( .A(n136), .B(\mult_x_1/n288 ), .ZN(n57) );
  XNOR2_X1 U152 ( .A(n136), .B(\mult_x_1/n287 ), .ZN(n71) );
  OAI22_X1 U153 ( .A1(n60), .A2(n57), .B1(n153), .B2(n71), .ZN(n73) );
  XNOR2_X1 U154 ( .A(n80), .B(\mult_x_1/n286 ), .ZN(n61) );
  XNOR2_X1 U155 ( .A(n80), .B(\mult_x_1/n285 ), .ZN(n69) );
  OAI22_X1 U156 ( .A1(n92), .A2(n61), .B1(n69), .B2(n89), .ZN(n72) );
  INV_X1 U157 ( .A(n72), .ZN(n58) );
  XNOR2_X1 U158 ( .A(n73), .B(n58), .ZN(n68) );
  OR2_X1 U159 ( .A1(\mult_x_1/n288 ), .A2(n486), .ZN(n59) );
  OAI22_X1 U160 ( .A1(n60), .A2(n486), .B1(n59), .B2(n18), .ZN(n67) );
  OR2_X1 U161 ( .A1(n68), .A2(n67), .ZN(n313) );
  XNOR2_X1 U162 ( .A(n80), .B(\mult_x_1/n287 ), .ZN(n63) );
  OAI22_X1 U163 ( .A1(n92), .A2(n63), .B1(n61), .B2(n89), .ZN(n66) );
  AND2_X1 U164 ( .A1(\mult_x_1/n288 ), .A2(n62), .ZN(n65) );
  NOR2_X1 U165 ( .A1(n66), .A2(n65), .ZN(n305) );
  OAI22_X1 U166 ( .A1(n92), .A2(\mult_x_1/n288 ), .B1(n63), .B2(n89), .ZN(n301) );
  OR2_X1 U167 ( .A1(\mult_x_1/n288 ), .A2(n488), .ZN(n64) );
  NAND2_X1 U168 ( .A1(n64), .A2(n92), .ZN(n300) );
  NAND2_X1 U169 ( .A1(n301), .A2(n300), .ZN(n308) );
  NAND2_X1 U170 ( .A1(n66), .A2(n65), .ZN(n306) );
  OAI21_X1 U171 ( .B1(n305), .B2(n308), .A(n306), .ZN(n314) );
  AOI21_X1 U172 ( .B1(n313), .B2(n314), .A(n10), .ZN(n322) );
  XNOR2_X1 U173 ( .A(n80), .B(\mult_x_1/n284 ), .ZN(n81) );
  OAI22_X1 U174 ( .A1(n92), .A2(n69), .B1(n81), .B2(n89), .ZN(n85) );
  AND2_X1 U175 ( .A1(n70), .A2(\mult_x_1/n288 ), .ZN(n84) );
  XNOR2_X1 U176 ( .A(n136), .B(\mult_x_1/n286 ), .ZN(n79) );
  OAI22_X1 U177 ( .A1(n152), .A2(n71), .B1(n153), .B2(n79), .ZN(n83) );
  NOR2_X1 U178 ( .A1(n75), .A2(n74), .ZN(n319) );
  NAND2_X1 U179 ( .A1(n75), .A2(n74), .ZN(n320) );
  OAI21_X1 U180 ( .B1(n322), .B2(n319), .A(n320), .ZN(n328) );
  OR2_X1 U181 ( .A1(\mult_x_1/n288 ), .A2(n484), .ZN(n76) );
  XNOR2_X1 U182 ( .A(n134), .B(\mult_x_1/n288 ), .ZN(n77) );
  XNOR2_X1 U183 ( .A(n134), .B(\mult_x_1/n287 ), .ZN(n99) );
  OAI22_X1 U184 ( .A1(n78), .A2(n77), .B1(n141), .B2(n99), .ZN(n100) );
  XNOR2_X1 U185 ( .A(n136), .B(\mult_x_1/n285 ), .ZN(n96) );
  OAI22_X1 U186 ( .A1(n152), .A2(n79), .B1(n153), .B2(n96), .ZN(n108) );
  XNOR2_X1 U187 ( .A(n80), .B(\mult_x_1/n283 ), .ZN(n91) );
  OAI22_X1 U188 ( .A1(n92), .A2(n81), .B1(n91), .B2(n89), .ZN(n107) );
  FA_X1 U189 ( .A(n85), .B(n84), .CI(n83), .CO(n86), .S(n75) );
  OR2_X1 U190 ( .A1(n87), .A2(n86), .ZN(n327) );
  NAND2_X1 U191 ( .A1(n87), .A2(n86), .ZN(n326) );
  INV_X1 U192 ( .A(n326), .ZN(n88) );
  AOI21_X1 U193 ( .B1(n328), .B2(n327), .A(n88), .ZN(n252) );
  INV_X1 U194 ( .A(n252), .ZN(n114) );
  INV_X1 U195 ( .A(n6), .ZN(n94) );
  AND2_X1 U196 ( .A1(\mult_x_1/n288 ), .A2(n94), .ZN(n161) );
  OAI22_X1 U197 ( .A1(n143), .A2(n99), .B1(n141), .B2(n98), .ZN(n175) );
  HA_X1 U198 ( .A(n101), .B(n100), .CO(n174), .S(n106) );
  OR2_X1 U199 ( .A1(n112), .A2(n111), .ZN(n250) );
  NAND2_X1 U200 ( .A1(n112), .A2(n111), .ZN(n251) );
  NAND2_X1 U201 ( .A1(n250), .A2(n251), .ZN(n113) );
  XNOR2_X1 U202 ( .A(n114), .B(n113), .ZN(n115) );
  INV_X2 U203 ( .A(n318), .ZN(n401) );
  NAND2_X1 U204 ( .A1(n115), .A2(n401), .ZN(n118) );
  BUF_X2 U205 ( .A(n116), .Z(n318) );
  INV_X2 U206 ( .A(n318), .ZN(n390) );
  OR2_X1 U207 ( .A1(n390), .A2(n516), .ZN(n117) );
  NAND2_X1 U208 ( .A1(n118), .A2(n117), .ZN(n578) );
  BUF_X2 U227 ( .A(n374), .Z(n295) );
  XNOR2_X1 U228 ( .A(n238), .B(\mult_x_1/n282 ), .ZN(n119) );
  NOR2_X1 U229 ( .A1(n119), .A2(n11), .ZN(n182) );
  XNOR2_X1 U230 ( .A(n16), .B(\mult_x_1/n281 ), .ZN(n120) );
  XNOR2_X1 U231 ( .A(n137), .B(n16), .ZN(n183) );
  OAI22_X1 U232 ( .A1(n9), .A2(n120), .B1(n183), .B2(n185), .ZN(n191) );
  INV_X1 U233 ( .A(n191), .ZN(n181) );
  XNOR2_X1 U234 ( .A(n16), .B(\mult_x_1/n282 ), .ZN(n123) );
  OAI22_X1 U235 ( .A1(n184), .A2(n123), .B1(n185), .B2(n120), .ZN(n127) );
  XNOR2_X1 U236 ( .A(n137), .B(n134), .ZN(n122) );
  AOI21_X1 U237 ( .B1(n141), .B2(n78), .A(n122), .ZN(n121) );
  INV_X1 U238 ( .A(n121), .ZN(n126) );
  XNOR2_X1 U239 ( .A(n134), .B(\mult_x_1/n281 ), .ZN(n140) );
  OAI22_X1 U240 ( .A1(n78), .A2(n140), .B1(n122), .B2(n141), .ZN(n125) );
  XNOR2_X1 U241 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n149) );
  OAI22_X1 U242 ( .A1(n184), .A2(n149), .B1(n185), .B2(n123), .ZN(n156) );
  INV_X1 U243 ( .A(n125), .ZN(n155) );
  XNOR2_X1 U244 ( .A(n238), .B(\mult_x_1/n283 ), .ZN(n124) );
  NOR2_X1 U245 ( .A1(n124), .A2(n11), .ZN(n131) );
  FA_X1 U246 ( .A(n127), .B(n126), .CI(n125), .CO(n180), .S(n130) );
  OR2_X1 U247 ( .A1(n199), .A2(n198), .ZN(n128) );
  NAND2_X1 U248 ( .A1(n399), .A2(n128), .ZN(n129) );
  OAI21_X1 U249 ( .B1(n295), .B2(n476), .A(n129), .ZN(n423) );
  FA_X1 U250 ( .A(n132), .B(n131), .CI(n130), .CO(n198), .S(n222) );
  XNOR2_X1 U251 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n150) );
  OAI22_X1 U252 ( .A1(n184), .A2(n133), .B1(n185), .B2(n150), .ZN(n266) );
  XNOR2_X1 U253 ( .A(n134), .B(\mult_x_1/n282 ), .ZN(n142) );
  OAI22_X1 U254 ( .A1(n78), .A2(n135), .B1(n141), .B2(n142), .ZN(n265) );
  XNOR2_X1 U255 ( .A(n137), .B(n136), .ZN(n151) );
  OAI22_X1 U256 ( .A1(n139), .A2(n138), .B1(n151), .B2(n153), .ZN(n233) );
  INV_X1 U257 ( .A(n233), .ZN(n264) );
  INV_X1 U258 ( .A(n229), .ZN(n145) );
  OAI22_X1 U259 ( .A1(n143), .A2(n142), .B1(n141), .B2(n140), .ZN(n228) );
  INV_X1 U260 ( .A(n228), .ZN(n144) );
  NAND2_X1 U261 ( .A1(n145), .A2(n144), .ZN(n146) );
  NAND2_X1 U262 ( .A1(n231), .A2(n146), .ZN(n148) );
  NAND2_X1 U263 ( .A1(n229), .A2(n228), .ZN(n147) );
  NAND2_X1 U264 ( .A1(n148), .A2(n147), .ZN(n227) );
  OAI22_X1 U265 ( .A1(n184), .A2(n150), .B1(n185), .B2(n149), .ZN(n234) );
  AOI21_X1 U266 ( .B1(n18), .B2(n152), .A(n151), .ZN(n154) );
  INV_X1 U267 ( .A(n154), .ZN(n232) );
  FA_X1 U268 ( .A(n157), .B(n156), .CI(n155), .CO(n132), .S(n225) );
  OR2_X1 U269 ( .A1(n222), .A2(n221), .ZN(n158) );
  NAND2_X1 U270 ( .A1(n293), .A2(n158), .ZN(n159) );
  OAI21_X1 U271 ( .B1(n295), .B2(n475), .A(n159), .ZN(n425) );
  HA_X1 U272 ( .A(n165), .B(n166), .CO(n47), .S(n206) );
  FA_X1 U273 ( .A(n169), .B(n168), .CI(n167), .CO(n203), .S(n205) );
  OR2_X1 U274 ( .A1(n218), .A2(n217), .ZN(n178) );
  NAND2_X1 U275 ( .A1(n293), .A2(n178), .ZN(n179) );
  OAI21_X1 U276 ( .B1(n295), .B2(n474), .A(n179), .ZN(n427) );
  FA_X1 U277 ( .A(n182), .B(n181), .CI(n180), .CO(n193), .S(n199) );
  AOI21_X1 U278 ( .B1(n185), .B2(n184), .A(n183), .ZN(n186) );
  INV_X1 U279 ( .A(n186), .ZN(n189) );
  XNOR2_X1 U280 ( .A(n238), .B(\mult_x_1/n281 ), .ZN(n187) );
  NOR2_X1 U281 ( .A1(n187), .A2(n11), .ZN(n188) );
  XOR2_X1 U282 ( .A(n189), .B(n188), .Z(n190) );
  XOR2_X1 U283 ( .A(n191), .B(n190), .Z(n192) );
  OR2_X1 U284 ( .A1(n193), .A2(n192), .ZN(n195) );
  NAND2_X1 U285 ( .A1(n193), .A2(n192), .ZN(n194) );
  NAND2_X1 U286 ( .A1(n195), .A2(n194), .ZN(n196) );
  NAND2_X1 U287 ( .A1(n293), .A2(n196), .ZN(n197) );
  OAI21_X1 U288 ( .B1(n293), .B2(n473), .A(n197), .ZN(n429) );
  NAND2_X1 U289 ( .A1(n199), .A2(n198), .ZN(n200) );
  NAND2_X1 U290 ( .A1(n293), .A2(n200), .ZN(n201) );
  OAI21_X1 U291 ( .B1(n293), .B2(n472), .A(n201), .ZN(n431) );
  FA_X1 U292 ( .A(n204), .B(n203), .CI(n202), .CO(n53), .S(n213) );
  INV_X1 U293 ( .A(n213), .ZN(n210) );
  FA_X1 U294 ( .A(n207), .B(n206), .CI(n205), .CO(n212), .S(n218) );
  INV_X1 U295 ( .A(n212), .ZN(n208) );
  AND2_X1 U296 ( .A1(n215), .A2(n208), .ZN(n209) );
  NAND2_X1 U297 ( .A1(n210), .A2(n209), .ZN(n211) );
  OAI21_X1 U298 ( .B1(n293), .B2(n468), .A(n211), .ZN(n439) );
  NAND2_X1 U299 ( .A1(n213), .A2(n212), .ZN(n214) );
  NAND2_X1 U300 ( .A1(n215), .A2(n214), .ZN(n216) );
  BUF_X1 U301 ( .A(n374), .Z(n255) );
  NAND2_X1 U302 ( .A1(n218), .A2(n217), .ZN(n219) );
  NAND2_X1 U303 ( .A1(n255), .A2(n219), .ZN(n220) );
  OAI21_X1 U304 ( .B1(n295), .B2(n466), .A(n220), .ZN(n443) );
  NAND2_X1 U305 ( .A1(n222), .A2(n221), .ZN(n223) );
  NAND2_X1 U306 ( .A1(n255), .A2(n223), .ZN(n224) );
  OAI21_X1 U307 ( .B1(n295), .B2(n465), .A(n224), .ZN(n445) );
  FA_X1 U308 ( .A(n227), .B(n226), .CI(n225), .CO(n221), .S(n247) );
  XNOR2_X1 U309 ( .A(n229), .B(n228), .ZN(n230) );
  XNOR2_X1 U310 ( .A(n231), .B(n230), .ZN(n282) );
  FA_X1 U311 ( .A(n234), .B(n19), .CI(n232), .CO(n226), .S(n281) );
  FA_X1 U312 ( .A(n237), .B(n236), .CI(n235), .CO(n263), .S(n275) );
  OAI21_X1 U313 ( .B1(n295), .B2(n464), .A(n245), .ZN(n447) );
  NAND2_X1 U314 ( .A1(n247), .A2(n246), .ZN(n248) );
  NAND2_X1 U315 ( .A1(n399), .A2(n248), .ZN(n249) );
  INV_X1 U316 ( .A(n250), .ZN(n253) );
  OAI21_X1 U317 ( .B1(n253), .B2(n252), .A(n251), .ZN(n254) );
  NAND2_X1 U318 ( .A1(n255), .A2(n254), .ZN(n256) );
  OAI21_X1 U319 ( .B1(n295), .B2(n461), .A(n256), .ZN(n453) );
  FA_X1 U320 ( .A(n259), .B(n258), .CI(n257), .CO(n285), .S(n273) );
  XNOR2_X1 U321 ( .A(n261), .B(n260), .ZN(n262) );
  XNOR2_X1 U322 ( .A(n263), .B(n262), .ZN(n283) );
  FA_X1 U323 ( .A(n265), .B(n266), .CI(n264), .CO(n231), .S(n284) );
  XNOR2_X1 U324 ( .A(n283), .B(n284), .ZN(n267) );
  XNOR2_X1 U325 ( .A(n285), .B(n267), .ZN(n268) );
  NAND2_X1 U326 ( .A1(n399), .A2(n268), .ZN(n269) );
  OAI21_X1 U327 ( .B1(n295), .B2(n460), .A(n269), .ZN(n455) );
  NAND2_X1 U328 ( .A1(n293), .A2(n278), .ZN(n279) );
  OAI21_X1 U329 ( .B1(n295), .B2(n459), .A(n279), .ZN(n457) );
  FA_X1 U330 ( .A(n282), .B(n281), .CI(n280), .CO(n246), .S(n292) );
  INV_X1 U331 ( .A(n291), .ZN(n288) );
  NAND2_X1 U332 ( .A1(n288), .A2(n399), .ZN(n290) );
  OR2_X1 U333 ( .A1(n295), .A2(n463), .ZN(n289) );
  OAI21_X1 U334 ( .B1(n7), .B2(n290), .A(n289), .ZN(n449) );
  NAND2_X1 U335 ( .A1(n292), .A2(n291), .ZN(n294) );
  NAND2_X1 U336 ( .A1(n294), .A2(n293), .ZN(n297) );
  OR2_X1 U337 ( .A1(n295), .A2(n471), .ZN(n296) );
  NAND2_X1 U338 ( .A1(n297), .A2(n296), .ZN(n433) );
  AOI22_X1 U339 ( .A1(n374), .A2(n535), .B1(n536), .B2(n318), .ZN(n538) );
  AOI22_X1 U340 ( .A1(n374), .A2(n534), .B1(n535), .B2(n318), .ZN(n540) );
  AND2_X1 U341 ( .A1(\mult_x_1/n288 ), .A2(n12), .ZN(n298) );
  NAND2_X1 U342 ( .A1(n399), .A2(n298), .ZN(n299) );
  OAI21_X1 U343 ( .B1(n403), .B2(n534), .A(n299), .ZN(n542) );
  AOI22_X1 U344 ( .A1(n374), .A2(n532), .B1(n533), .B2(n318), .ZN(n544) );
  AOI22_X1 U345 ( .A1(n374), .A2(n531), .B1(n532), .B2(n318), .ZN(n546) );
  OR2_X1 U346 ( .A1(n301), .A2(n300), .ZN(n302) );
  AND2_X1 U347 ( .A1(n302), .A2(n308), .ZN(n303) );
  NAND2_X1 U348 ( .A1(n399), .A2(n303), .ZN(n304) );
  OAI21_X1 U349 ( .B1(n390), .B2(n531), .A(n304), .ZN(n548) );
  AOI22_X1 U350 ( .A1(n374), .A2(n529), .B1(n530), .B2(n404), .ZN(n550) );
  AOI22_X1 U351 ( .A1(n374), .A2(n528), .B1(n529), .B2(n404), .ZN(n552) );
  INV_X1 U352 ( .A(n305), .ZN(n307) );
  NAND2_X1 U353 ( .A1(n307), .A2(n306), .ZN(n309) );
  XOR2_X1 U354 ( .A(n309), .B(n308), .Z(n310) );
  NAND2_X1 U355 ( .A1(n399), .A2(n310), .ZN(n311) );
  OAI21_X1 U356 ( .B1(n390), .B2(n528), .A(n311), .ZN(n554) );
  AOI22_X1 U357 ( .A1(n374), .A2(n526), .B1(n527), .B2(n404), .ZN(n556) );
  AOI22_X1 U358 ( .A1(n374), .A2(n525), .B1(n526), .B2(n404), .ZN(n558) );
  NAND2_X1 U359 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  NAND2_X1 U361 ( .A1(n401), .A2(n316), .ZN(n317) );
  OAI21_X1 U362 ( .B1(n390), .B2(n525), .A(n317), .ZN(n560) );
  AOI22_X1 U363 ( .A1(n374), .A2(n523), .B1(n524), .B2(n404), .ZN(n562) );
  BUF_X2 U364 ( .A(n318), .Z(n404) );
  AOI22_X1 U365 ( .A1(n374), .A2(n522), .B1(n523), .B2(n404), .ZN(n564) );
  INV_X1 U366 ( .A(n319), .ZN(n321) );
  NAND2_X1 U367 ( .A1(n321), .A2(n320), .ZN(n323) );
  XOR2_X1 U368 ( .A(n323), .B(n322), .Z(n324) );
  NAND2_X1 U369 ( .A1(n401), .A2(n324), .ZN(n325) );
  OAI21_X1 U370 ( .B1(n390), .B2(n522), .A(n325), .ZN(n566) );
  AOI22_X1 U371 ( .A1(n374), .A2(n520), .B1(n521), .B2(n404), .ZN(n568) );
  AOI22_X1 U372 ( .A1(n374), .A2(n519), .B1(n520), .B2(n404), .ZN(n570) );
  NAND2_X1 U373 ( .A1(n327), .A2(n326), .ZN(n329) );
  XNOR2_X1 U374 ( .A(n329), .B(n328), .ZN(n330) );
  NAND2_X1 U375 ( .A1(n401), .A2(n330), .ZN(n331) );
  OAI21_X1 U376 ( .B1(n390), .B2(n519), .A(n331), .ZN(n572) );
  AOI22_X1 U377 ( .A1(n374), .A2(n517), .B1(n518), .B2(n404), .ZN(n574) );
  AOI22_X1 U378 ( .A1(n403), .A2(n516), .B1(n517), .B2(n404), .ZN(n576) );
  AOI22_X1 U379 ( .A1(n403), .A2(n514), .B1(n515), .B2(n404), .ZN(n580) );
  NAND2_X1 U380 ( .A1(n407), .A2(n415), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n420), .B(n332), .ZN(n333) );
  NAND2_X1 U382 ( .A1(n401), .A2(n333), .ZN(n334) );
  OAI21_X1 U383 ( .B1(n390), .B2(n514), .A(n334), .ZN(n582) );
  AOI22_X1 U384 ( .A1(n403), .A2(n512), .B1(n513), .B2(n404), .ZN(n584) );
  AOI21_X1 U385 ( .B1(n420), .B2(n407), .A(n466), .ZN(n338) );
  NAND2_X1 U386 ( .A1(n468), .A2(n414), .ZN(n335) );
  XOR2_X1 U387 ( .A(n338), .B(n335), .Z(n336) );
  NAND2_X1 U388 ( .A1(n401), .A2(n336), .ZN(n337) );
  OAI21_X1 U389 ( .B1(n390), .B2(n512), .A(n337), .ZN(n586) );
  AOI22_X1 U390 ( .A1(n374), .A2(n510), .B1(n511), .B2(n404), .ZN(n588) );
  OAI21_X1 U391 ( .B1(n338), .B2(n413), .A(n414), .ZN(n351) );
  INV_X1 U392 ( .A(n351), .ZN(n342) );
  NAND2_X1 U393 ( .A1(n470), .A2(n412), .ZN(n339) );
  XOR2_X1 U394 ( .A(n342), .B(n339), .Z(n340) );
  NAND2_X1 U395 ( .A1(n401), .A2(n340), .ZN(n341) );
  OAI21_X1 U396 ( .B1(n390), .B2(n510), .A(n341), .ZN(n590) );
  AOI22_X1 U397 ( .A1(n403), .A2(n508), .B1(n509), .B2(n404), .ZN(n592) );
  OAI21_X1 U398 ( .B1(n342), .B2(n411), .A(n412), .ZN(n345) );
  OR2_X1 U399 ( .A1(n421), .A2(n422), .ZN(n343) );
  NAND2_X1 U400 ( .A1(n421), .A2(n422), .ZN(n348) );
  NAND2_X1 U401 ( .A1(n343), .A2(n348), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U403 ( .A1(n401), .A2(n346), .ZN(n347) );
  OAI21_X1 U404 ( .B1(n390), .B2(n508), .A(n347), .ZN(n594) );
  AOI22_X1 U405 ( .A1(n403), .A2(n506), .B1(n507), .B2(n404), .ZN(n596) );
  NOR2_X1 U406 ( .A1(n421), .A2(n422), .ZN(n349) );
  NOR2_X1 U407 ( .A1(n349), .A2(n411), .ZN(n352) );
  OAI21_X1 U408 ( .B1(n349), .B2(n412), .A(n348), .ZN(n350) );
  AOI21_X1 U409 ( .B1(n352), .B2(n351), .A(n350), .ZN(n380) );
  NAND2_X1 U410 ( .A1(n463), .A2(n410), .ZN(n353) );
  XOR2_X1 U411 ( .A(n380), .B(n353), .Z(n354) );
  NAND2_X1 U412 ( .A1(n390), .A2(n354), .ZN(n355) );
  OAI21_X1 U413 ( .B1(n390), .B2(n506), .A(n355), .ZN(n598) );
  AOI22_X1 U414 ( .A1(n374), .A2(n504), .B1(n505), .B2(n404), .ZN(n600) );
  OAI21_X1 U415 ( .B1(n380), .B2(n418), .A(n410), .ZN(n357) );
  NAND2_X1 U416 ( .A1(n417), .A2(n419), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  NAND2_X1 U418 ( .A1(n390), .A2(n358), .ZN(n359) );
  OAI21_X1 U419 ( .B1(n390), .B2(n504), .A(n359), .ZN(n602) );
  AOI22_X1 U420 ( .A1(n374), .A2(n502), .B1(n503), .B2(n404), .ZN(n604) );
  NAND2_X1 U421 ( .A1(n463), .A2(n417), .ZN(n361) );
  AOI21_X1 U422 ( .B1(n471), .B2(n417), .A(n462), .ZN(n360) );
  OAI21_X1 U423 ( .B1(n380), .B2(n361), .A(n360), .ZN(n363) );
  NAND2_X1 U424 ( .A1(n406), .A2(n416), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  NAND2_X1 U426 ( .A1(n390), .A2(n364), .ZN(n365) );
  OAI21_X1 U427 ( .B1(n390), .B2(n502), .A(n365), .ZN(n606) );
  AOI22_X1 U428 ( .A1(n374), .A2(n500), .B1(n501), .B2(n404), .ZN(n608) );
  NAND2_X1 U429 ( .A1(n417), .A2(n406), .ZN(n367) );
  INV_X1 U430 ( .A(n367), .ZN(n375) );
  NAND2_X1 U431 ( .A1(n463), .A2(n375), .ZN(n369) );
  AOI21_X1 U432 ( .B1(n462), .B2(n406), .A(n465), .ZN(n366) );
  OAI21_X1 U433 ( .B1(n367), .B2(n410), .A(n366), .ZN(n377) );
  INV_X1 U434 ( .A(n377), .ZN(n368) );
  OAI21_X1 U435 ( .B1(n380), .B2(n369), .A(n368), .ZN(n371) );
  NAND2_X1 U436 ( .A1(n405), .A2(n409), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U438 ( .A1(n401), .A2(n372), .ZN(n373) );
  OAI21_X1 U439 ( .B1(n403), .B2(n500), .A(n373), .ZN(n610) );
  AOI22_X1 U440 ( .A1(n374), .A2(n498), .B1(n499), .B2(n404), .ZN(n612) );
  AND2_X1 U441 ( .A1(n405), .A2(n375), .ZN(n376) );
  NAND2_X1 U442 ( .A1(n376), .A2(n463), .ZN(n379) );
  AOI21_X1 U443 ( .B1(n377), .B2(n405), .A(n472), .ZN(n378) );
  OAI21_X1 U444 ( .B1(n380), .B2(n379), .A(n378), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n381), .B(n408), .ZN(n382) );
  NAND2_X1 U446 ( .A1(n401), .A2(n382), .ZN(n383) );
  OAI21_X1 U447 ( .B1(n390), .B2(n498), .A(n383), .ZN(n614) );
  NAND2_X1 U448 ( .A1(n401), .A2(B_extended[0]), .ZN(n384) );
  OAI21_X1 U449 ( .B1(n403), .B2(n497), .A(n384), .ZN(n616) );
  NAND2_X1 U450 ( .A1(n401), .A2(B_extended[1]), .ZN(n385) );
  OAI21_X1 U451 ( .B1(n390), .B2(n496), .A(n385), .ZN(n618) );
  NAND2_X1 U452 ( .A1(n401), .A2(B_extended[2]), .ZN(n386) );
  OAI21_X1 U453 ( .B1(n403), .B2(n495), .A(n386), .ZN(n620) );
  NAND2_X1 U454 ( .A1(n401), .A2(B_extended[3]), .ZN(n387) );
  OAI21_X1 U455 ( .B1(n390), .B2(n494), .A(n387), .ZN(n622) );
  NAND2_X1 U456 ( .A1(n401), .A2(B_extended[4]), .ZN(n388) );
  OAI21_X1 U457 ( .B1(n403), .B2(n493), .A(n388), .ZN(n624) );
  NAND2_X1 U458 ( .A1(n401), .A2(B_extended[5]), .ZN(n389) );
  OAI21_X1 U459 ( .B1(n390), .B2(n492), .A(n389), .ZN(n626) );
  NAND2_X1 U460 ( .A1(n401), .A2(B_extended[6]), .ZN(n391) );
  OAI21_X1 U461 ( .B1(n403), .B2(n491), .A(n391), .ZN(n628) );
  NAND2_X1 U462 ( .A1(n401), .A2(B_extended[7]), .ZN(n392) );
  OAI21_X1 U463 ( .B1(n403), .B2(n490), .A(n392), .ZN(n630) );
  NAND2_X1 U464 ( .A1(n401), .A2(A_extended[0]), .ZN(n393) );
  OAI21_X1 U465 ( .B1(n403), .B2(n489), .A(n393), .ZN(n632) );
  NAND2_X1 U466 ( .A1(n399), .A2(A_extended[1]), .ZN(n394) );
  OAI21_X1 U467 ( .B1(n403), .B2(n488), .A(n394), .ZN(n634) );
  NAND2_X1 U468 ( .A1(n401), .A2(A_extended[2]), .ZN(n395) );
  OAI21_X1 U469 ( .B1(n403), .B2(n487), .A(n395), .ZN(n636) );
  NAND2_X1 U470 ( .A1(n399), .A2(A_extended[3]), .ZN(n396) );
  OAI21_X1 U471 ( .B1(n403), .B2(n486), .A(n396), .ZN(n638) );
  NAND2_X1 U472 ( .A1(n399), .A2(A_extended[4]), .ZN(n397) );
  OAI21_X1 U473 ( .B1(n403), .B2(n485), .A(n397), .ZN(n640) );
  NAND2_X1 U474 ( .A1(n399), .A2(A_extended[5]), .ZN(n398) );
  OAI21_X1 U475 ( .B1(n403), .B2(n484), .A(n398), .ZN(n642) );
  NAND2_X1 U476 ( .A1(n399), .A2(A_extended[6]), .ZN(n400) );
  OAI21_X1 U477 ( .B1(n403), .B2(n483), .A(n400), .ZN(n644) );
  NAND2_X1 U478 ( .A1(n401), .A2(A_extended[7]), .ZN(n402) );
  OAI21_X1 U479 ( .B1(n403), .B2(n482), .A(n402), .ZN(n646) );
  NAND2_X1 U480 ( .A1(n481), .A2(n404), .ZN(n648) );
endmodule


module conv_128_32_opt_DW_mult_pipe_J1_31 ( clk, rst_n, en, tc, a, b, product
 );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n407, n409, n411, n413, n415, n417, n419, n421,
         n423, n425, n427, n429, n431, n433, n435, n437, n439, n441, n443,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n526, n528, n530, n532, n534, n536, n538, n540,
         n542, n544, n546, n548, n550, n552, n554, n556, n558, n560, n562,
         n564, n566, n568, n570, n572, n574, n576, n578, n580, n582, n584,
         n586, n588, n590, n592, n594, n596, n598, n600, n602, n604, n606,
         n608, n610, n612, n614, n616, n618, n620, n622, n624, n626, n628,
         n630, n632, n634, n651, n652;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n469), .SE(n634), .CK(clk), .Q(n651), 
        .QN(n470) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n469), .SE(n630), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n472) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n469), .SE(n628), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n473) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n469), .SE(n626), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n474) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n469), .SE(n624), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n475) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n469), .SE(n622), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n476) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n469), .SE(n618), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n478) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n469), .SE(n616), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n479) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n469), .SE(n614), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n480) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n468), .SE(n612), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n481) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n468), .SE(n610), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n482) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n468), .SE(n608), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n483) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n468), .SE(n606), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n484) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n468), .SE(n604), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n485) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n468), .SE(n602), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n486) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n468), .SE(n600), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n468), .SE(n598), .CK(clk), .Q(
        product[15]), .QN(n488) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n468), .SE(n596), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n468), .SE(n594), .CK(clk), .Q(
        product[14]), .QN(n490) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n468), .SE(n592), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n467), .SE(n590), .CK(clk), .Q(
        product[13]), .QN(n492) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n467), .SE(n588), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n467), .SE(n586), .CK(clk), .Q(
        product[12]), .QN(n494) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n467), .SE(n584), .CK(clk), .QN(n495)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n467), .SE(n582), .CK(clk), .Q(
        product[11]), .QN(n496) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n467), .SE(n580), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n467), .SE(n578), .CK(clk), .Q(
        product[10]), .QN(n498) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n467), .SE(n576), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n467), .SE(n574), .CK(clk), .Q(
        product[9]), .QN(n500) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n467), .SE(n572), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n467), .SE(n570), .CK(clk), .Q(
        product[8]), .QN(n502) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n466), .SE(n568), .CK(clk), .QN(n503)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n466), .SE(n566), .CK(clk), .Q(
        product[7]), .QN(n504) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n466), .SE(n564), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n466), .SE(n562), .CK(clk), .Q(
        product[6]), .QN(n506) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n466), .SE(n560), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n466), .SE(n558), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n466), .SE(n556), .CK(clk), .Q(
        product[5]), .QN(n509) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n466), .SE(n554), .CK(clk), .QN(n510)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n466), .SE(n552), .CK(clk), .QN(n511)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n466), .SE(n550), .CK(clk), .Q(
        product[4]), .QN(n512) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n466), .SE(n548), .CK(clk), .QN(n513)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n465), .SE(n546), .CK(clk), .QN(n514)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n465), .SE(n544), .CK(clk), .Q(
        product[3]), .QN(n515) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n465), .SE(n542), .CK(clk), .QN(n516)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n465), .SE(n540), .CK(clk), .QN(n517)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n465), .SE(n538), .CK(clk), .Q(
        product[2]), .QN(n518) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n465), .SE(n536), .CK(clk), .QN(n519)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n465), .SE(n534), .CK(clk), .QN(n520)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n465), .SE(n532), .CK(clk), .Q(
        product[1]), .QN(n521) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n465), .SE(n530), .CK(clk), .QN(n522)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n465), .SE(n528), .CK(clk), .QN(n523)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n465), .SE(n526), .CK(clk), .Q(
        product[0]), .QN(n524) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n469), .SE(n620), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n477) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n652), .SE(n439), .CK(
        clk), .Q(n447), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n652), .SI(1'b1), .SE(n443), .CK(clk), 
        .Q(n404), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2_IP  ( .D(1'b1), .SI(n652), .SE(n441), .CK(
        clk), .Q(n446), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n652), .SI(1'b1), .SE(n437), .CK(clk), 
        .Q(n401), .QN(n448) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n652), .SI(1'b1), .SE(n435), .CK(clk), 
        .Q(n400), .QN(n449) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n652), .SE(n433), .CK(
        clk), .Q(n450), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n652), .SE(n431), .CK(
        clk), .Q(n451), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n652), .SI(1'b1), .SE(n429), .CK(clk), 
        .Q(n397), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n652), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n396), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n652), .SI(1'b1), .SE(n425), .CK(clk), 
        .Q(n395), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n652), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n394), .QN(n455) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n652), .SI(1'b1), .SE(n421), .CK(clk), 
        .Q(n393), .QN(n456) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n652), .SI(1'b1), .SE(n419), .CK(clk), 
        .Q(n392), .QN(n457) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n652), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n391), .QN(n458) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n652), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n390), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n652), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n389), .QN(n460) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n652), .SE(n411), .CK(
        clk), .Q(n461), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n652), .SE(n409), .CK(
        clk), .Q(n462), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n652), .SI(1'b1), .SE(n407), .CK(clk), 
        .Q(n386), .QN(n463) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n652), .SI(1'b1), .SE(n405), .CK(clk), 
        .Q(n385), .QN(n464) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n469), .SE(n632), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n471) );
  OR2_X1 U2 ( .A1(n189), .A2(n11), .ZN(n187) );
  NAND2_X1 U3 ( .A1(n12), .A2(n348), .ZN(n11) );
  INV_X1 U4 ( .A(n188), .ZN(n12) );
  NAND2_X1 U5 ( .A1(n6), .A2(n5), .ZN(n266) );
  OAI21_X1 U6 ( .B1(n110), .B2(n109), .A(n7), .ZN(n6) );
  INV_X1 U7 ( .A(n10), .ZN(n7) );
  BUF_X1 U8 ( .A(\mult_x_1/n312 ), .Z(n225) );
  BUF_X1 U9 ( .A(\mult_x_1/n313 ), .Z(n236) );
  XOR2_X1 U10 ( .A(n142), .B(n141), .Z(n184) );
  NAND2_X2 U11 ( .A1(n110), .A2(n109), .ZN(n5) );
  XNOR2_X1 U12 ( .A(n9), .B(n8), .ZN(n180) );
  INV_X1 U13 ( .A(n110), .ZN(n8) );
  XNOR2_X1 U14 ( .A(n10), .B(n109), .ZN(n9) );
  NAND2_X1 U15 ( .A1(n142), .A2(n141), .ZN(n10) );
  OAI21_X1 U16 ( .B1(n14), .B2(n13), .A(n348), .ZN(n209) );
  INV_X1 U17 ( .A(n249), .ZN(n13) );
  INV_X1 U18 ( .A(n19), .ZN(n14) );
  AND2_X1 U19 ( .A1(n651), .A2(\mult_x_1/n281 ), .ZN(n116) );
  BUF_X1 U20 ( .A(n357), .Z(n384) );
  INV_X1 U21 ( .A(n357), .ZN(n253) );
  INV_X2 U22 ( .A(n280), .ZN(n348) );
  CLKBUF_X1 U23 ( .A(n279), .Z(n466) );
  CLKBUF_X1 U24 ( .A(n279), .Z(n467) );
  CLKBUF_X1 U25 ( .A(n279), .Z(n468) );
  CLKBUF_X1 U26 ( .A(n279), .Z(n469) );
  CLKBUF_X1 U27 ( .A(n279), .Z(n465) );
  INV_X1 U28 ( .A(rst_n), .ZN(n652) );
  INV_X1 U29 ( .A(n30), .ZN(n40) );
  BUF_X2 U30 ( .A(n38), .Z(n15) );
  INV_X1 U31 ( .A(n471), .ZN(n16) );
  INV_X1 U32 ( .A(n471), .ZN(n115) );
  OR2_X1 U33 ( .A1(n253), .A2(n454), .ZN(n17) );
  NAND2_X1 U34 ( .A1(n17), .A2(n191), .ZN(n425) );
  XNOR2_X1 U35 ( .A(n215), .B(n214), .ZN(n216) );
  XNOR2_X1 U36 ( .A(n265), .B(n101), .ZN(n278) );
  XNOR2_X1 U37 ( .A(n267), .B(n266), .ZN(n101) );
  NAND2_X1 U38 ( .A1(n267), .A2(n266), .ZN(n268) );
  NAND2_X1 U39 ( .A1(n265), .A2(n264), .ZN(n269) );
  OR2_X1 U40 ( .A1(n266), .A2(n267), .ZN(n264) );
  OAI21_X1 U41 ( .B1(n21), .B2(n83), .A(n82), .ZN(n133) );
  NAND2_X1 U42 ( .A1(n215), .A2(n214), .ZN(n204) );
  NAND2_X1 U43 ( .A1(n217), .A2(n203), .ZN(n205) );
  OR2_X1 U44 ( .A1(n215), .A2(n214), .ZN(n203) );
  INV_X1 U45 ( .A(n652), .ZN(n279) );
  CLKBUF_X1 U46 ( .A(n77), .Z(n18) );
  OR2_X1 U47 ( .A1(n207), .A2(n206), .ZN(n19) );
  NAND2_X1 U48 ( .A1(n205), .A2(n204), .ZN(n206) );
  OR2_X1 U49 ( .A1(n477), .A2(\mult_x_1/n180 ), .ZN(n237) );
  INV_X1 U50 ( .A(n479), .ZN(n20) );
  AND3_X1 U51 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n21) );
  INV_X1 U52 ( .A(n225), .ZN(n22) );
  XNOR2_X1 U53 ( .A(n217), .B(n216), .ZN(n247) );
  NAND2_X1 U54 ( .A1(n81), .A2(n80), .ZN(n82) );
  NOR2_X1 U55 ( .A1(n81), .A2(n80), .ZN(n83) );
  XOR2_X1 U56 ( .A(n53), .B(n54), .Z(n23) );
  XOR2_X1 U57 ( .A(n55), .B(n23), .Z(n262) );
  NAND2_X1 U58 ( .A1(n53), .A2(n55), .ZN(n24) );
  NAND2_X1 U59 ( .A1(n55), .A2(n54), .ZN(n25) );
  NAND2_X1 U60 ( .A1(n53), .A2(n54), .ZN(n26) );
  NAND3_X1 U61 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n79) );
  BUF_X2 U62 ( .A(n51), .Z(n151) );
  BUF_X4 U63 ( .A(n348), .Z(n27) );
  INV_X1 U64 ( .A(n295), .ZN(n28) );
  INV_X1 U65 ( .A(n295), .ZN(n29) );
  XNOR2_X1 U66 ( .A(n476), .B(\mult_x_1/n313 ), .ZN(n30) );
  BUF_X1 U67 ( .A(n280), .Z(n295) );
  AND2_X1 U68 ( .A1(n269), .A2(n268), .ZN(n31) );
  INV_X1 U69 ( .A(n295), .ZN(n381) );
  INV_X1 U70 ( .A(en), .ZN(n280) );
  XOR2_X1 U71 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n32) );
  XNOR2_X1 U72 ( .A(n474), .B(n475), .ZN(n33) );
  NAND2_X1 U73 ( .A1(n32), .A2(n33), .ZN(n51) );
  BUF_X2 U74 ( .A(\mult_x_1/n311 ), .Z(n147) );
  XNOR2_X1 U75 ( .A(n147), .B(\mult_x_1/n284 ), .ZN(n96) );
  BUF_X2 U76 ( .A(n33), .Z(n219) );
  XNOR2_X1 U77 ( .A(n147), .B(\mult_x_1/n283 ), .ZN(n39) );
  OAI22_X1 U78 ( .A1(n151), .A2(n96), .B1(n219), .B2(n39), .ZN(n43) );
  XNOR2_X1 U79 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n34) );
  OR2_X2 U80 ( .A1(n34), .A2(n30), .ZN(n232) );
  XNOR2_X1 U81 ( .A(n225), .B(\mult_x_1/n282 ), .ZN(n97) );
  XNOR2_X1 U82 ( .A(n225), .B(\mult_x_1/n281 ), .ZN(n41) );
  OAI22_X1 U83 ( .A1(n232), .A2(n97), .B1(n40), .B2(n41), .ZN(n42) );
  XNOR2_X1 U84 ( .A(n43), .B(n42), .ZN(n92) );
  AND2_X2 U85 ( .A1(n651), .A2(\mult_x_1/n310 ), .ZN(n163) );
  XNOR2_X1 U86 ( .A(n163), .B(n115), .ZN(n74) );
  CLKBUF_X1 U87 ( .A(n74), .Z(n164) );
  INV_X1 U88 ( .A(n163), .ZN(n35) );
  OR2_X1 U89 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n36) );
  NOR2_X1 U90 ( .A1(n164), .A2(n36), .ZN(n91) );
  XNOR2_X1 U91 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n38) );
  XNOR2_X1 U92 ( .A(n472), .B(\mult_x_1/n310 ), .ZN(n37) );
  NAND2_X2 U93 ( .A1(n38), .A2(n37), .ZN(n161) );
  XNOR2_X1 U94 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n99) );
  XNOR2_X1 U95 ( .A(n115), .B(\mult_x_1/n286 ), .ZN(n48) );
  OAI22_X1 U96 ( .A1(n161), .A2(n99), .B1(n15), .B2(n48), .ZN(n104) );
  XNOR2_X1 U97 ( .A(n236), .B(n20), .ZN(n106) );
  XNOR2_X1 U98 ( .A(n116), .B(\mult_x_1/n313 ), .ZN(n45) );
  OAI22_X1 U99 ( .A1(n237), .A2(n106), .B1(n45), .B2(n478), .ZN(n103) );
  NOR2_X1 U100 ( .A1(n74), .A2(n486), .ZN(n102) );
  XNOR2_X1 U101 ( .A(n147), .B(\mult_x_1/n282 ), .ZN(n52) );
  OAI22_X1 U102 ( .A1(n151), .A2(n39), .B1(n219), .B2(n52), .ZN(n55) );
  XNOR2_X1 U103 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n57) );
  XNOR2_X1 U104 ( .A(n115), .B(\mult_x_1/n285 ), .ZN(n47) );
  OAI22_X1 U105 ( .A1(n15), .A2(n57), .B1(n47), .B2(n161), .ZN(n54) );
  XNOR2_X1 U106 ( .A(n116), .B(n225), .ZN(n58) );
  OAI22_X1 U107 ( .A1(n232), .A2(n41), .B1(n58), .B2(n40), .ZN(n77) );
  INV_X1 U108 ( .A(n77), .ZN(n53) );
  OR2_X1 U109 ( .A1(n43), .A2(n42), .ZN(n62) );
  XNOR2_X1 U110 ( .A(n163), .B(\mult_x_1/n286 ), .ZN(n44) );
  NOR2_X1 U111 ( .A1(n164), .A2(n44), .ZN(n61) );
  AOI21_X1 U112 ( .B1(n237), .B2(n478), .A(n45), .ZN(n46) );
  INV_X1 U113 ( .A(n46), .ZN(n95) );
  OAI22_X1 U114 ( .A1(n161), .A2(n48), .B1(n15), .B2(n47), .ZN(n94) );
  XNOR2_X1 U115 ( .A(n163), .B(\mult_x_1/n287 ), .ZN(n49) );
  NOR2_X1 U116 ( .A1(n74), .A2(n49), .ZN(n93) );
  NOR2_X1 U117 ( .A1(n357), .A2(n67), .ZN(n64) );
  XNOR2_X1 U118 ( .A(n163), .B(\mult_x_1/n285 ), .ZN(n50) );
  NOR2_X1 U119 ( .A1(n50), .A2(n74), .ZN(n81) );
  XNOR2_X1 U120 ( .A(n147), .B(\mult_x_1/n281 ), .ZN(n72) );
  OAI22_X1 U121 ( .A1(n151), .A2(n52), .B1(n219), .B2(n72), .ZN(n80) );
  XNOR2_X1 U122 ( .A(n81), .B(n80), .ZN(n56) );
  XNOR2_X1 U123 ( .A(n56), .B(n79), .ZN(n86) );
  XNOR2_X1 U124 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n73) );
  OAI22_X1 U125 ( .A1(n161), .A2(n57), .B1(n15), .B2(n73), .ZN(n78) );
  AOI21_X1 U126 ( .B1(n40), .B2(n232), .A(n58), .ZN(n59) );
  INV_X1 U127 ( .A(n59), .ZN(n76) );
  FA_X1 U128 ( .A(n62), .B(n61), .CI(n60), .CO(n84), .S(n261) );
  INV_X1 U129 ( .A(n68), .ZN(n63) );
  NAND2_X1 U130 ( .A1(n64), .A2(n63), .ZN(n66) );
  OR2_X1 U131 ( .A1(n29), .A2(n447), .ZN(n65) );
  NAND2_X1 U132 ( .A1(n66), .A2(n65), .ZN(n439) );
  NAND2_X1 U133 ( .A1(n68), .A2(n67), .ZN(n69) );
  BUF_X2 U134 ( .A(n280), .Z(n357) );
  NAND2_X1 U135 ( .A1(n69), .A2(n253), .ZN(n71) );
  OR2_X1 U136 ( .A1(n27), .A2(n458), .ZN(n70) );
  NAND2_X1 U137 ( .A1(n71), .A2(n70), .ZN(n417) );
  XNOR2_X1 U138 ( .A(n116), .B(n147), .ZN(n119) );
  OAI22_X1 U139 ( .A1(n51), .A2(n72), .B1(n119), .B2(n219), .ZN(n126) );
  INV_X1 U140 ( .A(n126), .ZN(n123) );
  XNOR2_X1 U141 ( .A(n115), .B(\mult_x_1/n282 ), .ZN(n118) );
  OAI22_X1 U142 ( .A1(n161), .A2(n73), .B1(n15), .B2(n118), .ZN(n122) );
  XNOR2_X1 U143 ( .A(n163), .B(\mult_x_1/n284 ), .ZN(n75) );
  NOR2_X1 U144 ( .A1(n75), .A2(n74), .ZN(n121) );
  FA_X1 U145 ( .A(n78), .B(n76), .CI(n18), .CO(n134), .S(n85) );
  FA_X1 U146 ( .A(n86), .B(n85), .CI(n84), .CO(n256), .S(n68) );
  OR2_X1 U147 ( .A1(n257), .A2(n256), .ZN(n87) );
  NAND2_X1 U148 ( .A1(n87), .A2(n27), .ZN(n89) );
  OR2_X1 U149 ( .A1(n28), .A2(n448), .ZN(n88) );
  NAND2_X1 U150 ( .A1(n89), .A2(n88), .ZN(n437) );
  FA_X1 U151 ( .A(n92), .B(n91), .CI(n90), .CO(n263), .S(n265) );
  FA_X1 U152 ( .A(n95), .B(n94), .CI(n93), .CO(n60), .S(n267) );
  XNOR2_X1 U153 ( .A(n147), .B(\mult_x_1/n285 ), .ZN(n105) );
  OAI22_X1 U154 ( .A1(n151), .A2(n105), .B1(n219), .B2(n96), .ZN(n110) );
  XNOR2_X1 U155 ( .A(n225), .B(\mult_x_1/n283 ), .ZN(n107) );
  OAI22_X1 U156 ( .A1(n232), .A2(n107), .B1(n40), .B2(n97), .ZN(n109) );
  OR2_X1 U157 ( .A1(\mult_x_1/n288 ), .A2(n471), .ZN(n98) );
  OAI22_X1 U158 ( .A1(n161), .A2(n471), .B1(n98), .B2(n15), .ZN(n142) );
  XNOR2_X1 U159 ( .A(n115), .B(\mult_x_1/n288 ), .ZN(n100) );
  OAI22_X1 U160 ( .A1(n161), .A2(n100), .B1(n15), .B2(n99), .ZN(n141) );
  FA_X1 U161 ( .A(n104), .B(n103), .CI(n102), .CO(n90), .S(n182) );
  XNOR2_X1 U162 ( .A(n147), .B(\mult_x_1/n286 ), .ZN(n149) );
  OAI22_X1 U163 ( .A1(n51), .A2(n149), .B1(n219), .B2(n105), .ZN(n145) );
  XNOR2_X1 U164 ( .A(n236), .B(\mult_x_1/n282 ), .ZN(n138) );
  OAI22_X1 U165 ( .A1(n237), .A2(n138), .B1(n106), .B2(n478), .ZN(n144) );
  XNOR2_X1 U166 ( .A(n225), .B(\mult_x_1/n284 ), .ZN(n140) );
  OAI22_X1 U167 ( .A1(n232), .A2(n140), .B1(n40), .B2(n107), .ZN(n143) );
  NAND2_X1 U168 ( .A1(n278), .A2(n274), .ZN(n111) );
  NAND2_X1 U169 ( .A1(n111), .A2(n253), .ZN(n113) );
  OR2_X1 U170 ( .A1(n29), .A2(n456), .ZN(n112) );
  NAND2_X1 U171 ( .A1(n113), .A2(n112), .ZN(n421) );
  XNOR2_X1 U192 ( .A(n163), .B(\mult_x_1/n282 ), .ZN(n114) );
  NOR2_X1 U193 ( .A1(n164), .A2(n114), .ZN(n159) );
  XNOR2_X1 U194 ( .A(n16), .B(n20), .ZN(n117) );
  XNOR2_X1 U195 ( .A(n116), .B(n16), .ZN(n160) );
  OAI22_X1 U196 ( .A1(n161), .A2(n117), .B1(n160), .B2(n15), .ZN(n169) );
  INV_X1 U197 ( .A(n169), .ZN(n158) );
  OAI22_X1 U198 ( .A1(n161), .A2(n118), .B1(n15), .B2(n117), .ZN(n127) );
  AOI21_X1 U199 ( .B1(n219), .B2(n51), .A(n119), .ZN(n120) );
  INV_X1 U200 ( .A(n120), .ZN(n125) );
  FA_X1 U201 ( .A(n123), .B(n122), .CI(n121), .CO(n132), .S(n135) );
  XNOR2_X1 U202 ( .A(n163), .B(\mult_x_1/n283 ), .ZN(n124) );
  NOR2_X1 U203 ( .A1(n124), .A2(n164), .ZN(n131) );
  FA_X1 U204 ( .A(n127), .B(n126), .CI(n125), .CO(n157), .S(n130) );
  OR2_X1 U205 ( .A1(n177), .A2(n176), .ZN(n128) );
  NAND2_X1 U206 ( .A1(n253), .A2(n128), .ZN(n129) );
  OAI21_X1 U207 ( .B1(n27), .B2(n464), .A(n129), .ZN(n405) );
  FA_X1 U208 ( .A(n132), .B(n131), .CI(n130), .CO(n176), .S(n211) );
  FA_X1 U209 ( .A(n135), .B(n134), .CI(n133), .CO(n210), .S(n257) );
  OR2_X1 U210 ( .A1(n211), .A2(n210), .ZN(n136) );
  NAND2_X1 U211 ( .A1(n253), .A2(n136), .ZN(n137) );
  OAI21_X1 U212 ( .B1(n29), .B2(n463), .A(n137), .ZN(n407) );
  XNOR2_X1 U213 ( .A(n236), .B(\mult_x_1/n283 ), .ZN(n202) );
  OAI22_X1 U214 ( .A1(n237), .A2(n202), .B1(n138), .B2(n478), .ZN(n154) );
  INV_X1 U215 ( .A(n38), .ZN(n139) );
  AND2_X1 U216 ( .A1(\mult_x_1/n288 ), .A2(n139), .ZN(n153) );
  XNOR2_X1 U217 ( .A(n225), .B(\mult_x_1/n285 ), .ZN(n201) );
  OAI22_X1 U218 ( .A1(n232), .A2(n201), .B1(n40), .B2(n140), .ZN(n152) );
  FA_X1 U219 ( .A(n145), .B(n144), .CI(n143), .CO(n181), .S(n183) );
  OR2_X1 U220 ( .A1(\mult_x_1/n288 ), .A2(n473), .ZN(n146) );
  OAI22_X1 U221 ( .A1(n151), .A2(n473), .B1(n146), .B2(n219), .ZN(n200) );
  XNOR2_X1 U222 ( .A(n147), .B(\mult_x_1/n288 ), .ZN(n148) );
  XNOR2_X1 U223 ( .A(n147), .B(\mult_x_1/n287 ), .ZN(n150) );
  OAI22_X1 U224 ( .A1(n51), .A2(n148), .B1(n219), .B2(n150), .ZN(n199) );
  OAI22_X1 U225 ( .A1(n151), .A2(n150), .B1(n219), .B2(n149), .ZN(n197) );
  FA_X1 U226 ( .A(n154), .B(n153), .CI(n152), .CO(n185), .S(n196) );
  OR2_X1 U227 ( .A1(n193), .A2(n192), .ZN(n155) );
  NAND2_X1 U228 ( .A1(n253), .A2(n155), .ZN(n156) );
  OAI21_X1 U229 ( .B1(n253), .B2(n462), .A(n156), .ZN(n409) );
  FA_X1 U230 ( .A(n159), .B(n158), .CI(n157), .CO(n171), .S(n177) );
  AOI21_X1 U231 ( .B1(n15), .B2(n161), .A(n160), .ZN(n162) );
  INV_X1 U232 ( .A(n162), .ZN(n167) );
  XNOR2_X1 U233 ( .A(n163), .B(n20), .ZN(n165) );
  NOR2_X1 U234 ( .A1(n165), .A2(n164), .ZN(n166) );
  XOR2_X1 U235 ( .A(n167), .B(n166), .Z(n168) );
  XOR2_X1 U236 ( .A(n169), .B(n168), .Z(n170) );
  OR2_X1 U237 ( .A1(n171), .A2(n170), .ZN(n173) );
  NAND2_X1 U238 ( .A1(n171), .A2(n170), .ZN(n172) );
  NAND2_X1 U239 ( .A1(n173), .A2(n172), .ZN(n174) );
  NAND2_X1 U240 ( .A1(n348), .A2(n174), .ZN(n175) );
  OAI21_X1 U241 ( .B1(n253), .B2(n461), .A(n175), .ZN(n411) );
  NAND2_X1 U242 ( .A1(n177), .A2(n176), .ZN(n178) );
  NAND2_X1 U243 ( .A1(n348), .A2(n178), .ZN(n179) );
  OAI21_X1 U244 ( .B1(n381), .B2(n460), .A(n179), .ZN(n413) );
  FA_X1 U245 ( .A(n182), .B(n181), .CI(n180), .CO(n274), .S(n189) );
  FA_X1 U246 ( .A(n185), .B(n184), .CI(n183), .CO(n188), .S(n193) );
  OAI21_X1 U247 ( .B1(n253), .B2(n455), .A(n187), .ZN(n423) );
  NAND2_X1 U248 ( .A1(n189), .A2(n188), .ZN(n190) );
  NAND2_X1 U249 ( .A1(n253), .A2(n190), .ZN(n191) );
  NAND2_X1 U250 ( .A1(n193), .A2(n192), .ZN(n194) );
  NAND2_X1 U251 ( .A1(n383), .A2(n194), .ZN(n195) );
  OAI21_X1 U252 ( .B1(n253), .B2(n453), .A(n195), .ZN(n427) );
  FA_X1 U253 ( .A(n198), .B(n197), .CI(n196), .CO(n192), .S(n207) );
  HA_X1 U254 ( .A(n200), .B(n199), .CO(n198), .S(n217) );
  XNOR2_X1 U255 ( .A(n225), .B(\mult_x_1/n286 ), .ZN(n221) );
  OAI22_X1 U256 ( .A1(n232), .A2(n221), .B1(n40), .B2(n201), .ZN(n215) );
  XNOR2_X1 U257 ( .A(n236), .B(\mult_x_1/n284 ), .ZN(n218) );
  OAI22_X1 U258 ( .A1(n237), .A2(n218), .B1(n202), .B2(n478), .ZN(n214) );
  NOR2_X1 U259 ( .A1(n207), .A2(n206), .ZN(n250) );
  NAND2_X1 U260 ( .A1(n207), .A2(n206), .ZN(n249) );
  OAI21_X1 U261 ( .B1(n253), .B2(n452), .A(n209), .ZN(n429) );
  NAND2_X1 U262 ( .A1(n211), .A2(n210), .ZN(n212) );
  NAND2_X1 U263 ( .A1(n348), .A2(n212), .ZN(n213) );
  OAI21_X1 U264 ( .B1(n253), .B2(n449), .A(n213), .ZN(n435) );
  XNOR2_X1 U265 ( .A(n236), .B(\mult_x_1/n285 ), .ZN(n228) );
  OAI22_X1 U266 ( .A1(n237), .A2(n228), .B1(n218), .B2(n478), .ZN(n224) );
  INV_X1 U267 ( .A(n219), .ZN(n220) );
  AND2_X1 U268 ( .A1(\mult_x_1/n288 ), .A2(n220), .ZN(n223) );
  XNOR2_X1 U269 ( .A(n225), .B(\mult_x_1/n287 ), .ZN(n226) );
  OAI22_X1 U270 ( .A1(n232), .A2(n226), .B1(n40), .B2(n221), .ZN(n222) );
  OR2_X1 U271 ( .A1(n247), .A2(n246), .ZN(n310) );
  FA_X1 U272 ( .A(n224), .B(n223), .CI(n222), .CO(n246), .S(n245) );
  XNOR2_X1 U273 ( .A(n225), .B(\mult_x_1/n288 ), .ZN(n227) );
  OAI22_X1 U274 ( .A1(n232), .A2(n227), .B1(n40), .B2(n226), .ZN(n230) );
  XNOR2_X1 U275 ( .A(n236), .B(\mult_x_1/n286 ), .ZN(n233) );
  OAI22_X1 U276 ( .A1(n237), .A2(n233), .B1(n228), .B2(n478), .ZN(n229) );
  NOR2_X1 U277 ( .A1(n245), .A2(n244), .ZN(n302) );
  HA_X1 U278 ( .A(n230), .B(n229), .CO(n244), .S(n242) );
  OR2_X1 U279 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n231) );
  OAI22_X1 U280 ( .A1(n232), .A2(n22), .B1(n231), .B2(n40), .ZN(n241) );
  OR2_X1 U281 ( .A1(n242), .A2(n241), .ZN(n297) );
  XNOR2_X1 U282 ( .A(n236), .B(\mult_x_1/n287 ), .ZN(n235) );
  OAI22_X1 U283 ( .A1(n237), .A2(n235), .B1(n233), .B2(n478), .ZN(n240) );
  INV_X1 U284 ( .A(n40), .ZN(n234) );
  AND2_X1 U285 ( .A1(\mult_x_1/n288 ), .A2(n234), .ZN(n239) );
  NOR2_X1 U286 ( .A1(n240), .A2(n239), .ZN(n288) );
  OAI22_X1 U287 ( .A1(n237), .A2(\mult_x_1/n288 ), .B1(n235), .B2(n478), .ZN(
        n284) );
  OR2_X1 U288 ( .A1(\mult_x_1/n288 ), .A2(n477), .ZN(n238) );
  NAND2_X1 U289 ( .A1(n238), .A2(n237), .ZN(n283) );
  NAND2_X1 U290 ( .A1(n284), .A2(n283), .ZN(n291) );
  NAND2_X1 U291 ( .A1(n240), .A2(n239), .ZN(n289) );
  OAI21_X1 U292 ( .B1(n288), .B2(n291), .A(n289), .ZN(n298) );
  NAND2_X1 U293 ( .A1(n242), .A2(n241), .ZN(n296) );
  INV_X1 U294 ( .A(n296), .ZN(n243) );
  AOI21_X1 U295 ( .B1(n297), .B2(n298), .A(n243), .ZN(n305) );
  NAND2_X1 U296 ( .A1(n245), .A2(n244), .ZN(n303) );
  OAI21_X1 U297 ( .B1(n302), .B2(n305), .A(n303), .ZN(n311) );
  NAND2_X1 U298 ( .A1(n247), .A2(n246), .ZN(n309) );
  INV_X1 U299 ( .A(n309), .ZN(n248) );
  AOI21_X1 U300 ( .B1(n310), .B2(n311), .A(n248), .ZN(n254) );
  OAI21_X1 U301 ( .B1(n254), .B2(n250), .A(n249), .ZN(n251) );
  NAND2_X1 U302 ( .A1(n251), .A2(n348), .ZN(n252) );
  OAI21_X1 U303 ( .B1(n253), .B2(n446), .A(n252), .ZN(n441) );
  NAND2_X1 U304 ( .A1(n28), .A2(n254), .ZN(n255) );
  OAI21_X1 U305 ( .B1(n381), .B2(n445), .A(n255), .ZN(n443) );
  OR2_X1 U306 ( .A1(n27), .A2(n459), .ZN(n260) );
  NAND2_X1 U307 ( .A1(n257), .A2(n256), .ZN(n258) );
  NAND2_X1 U308 ( .A1(n27), .A2(n258), .ZN(n259) );
  NAND2_X1 U309 ( .A1(n260), .A2(n259), .ZN(n415) );
  FA_X1 U310 ( .A(n263), .B(n262), .CI(n261), .CO(n67), .S(n273) );
  NAND2_X1 U311 ( .A1(n31), .A2(n348), .ZN(n270) );
  OAI22_X1 U312 ( .A1(n273), .A2(n270), .B1(n27), .B2(n451), .ZN(n431) );
  OR2_X1 U313 ( .A1(n381), .A2(n450), .ZN(n272) );
  NAND2_X1 U314 ( .A1(n31), .A2(n348), .ZN(n271) );
  OAI211_X1 U315 ( .C1(n273), .C2(n295), .A(n272), .B(n271), .ZN(n433) );
  INV_X1 U316 ( .A(n274), .ZN(n275) );
  NAND2_X1 U317 ( .A1(n348), .A2(n275), .ZN(n277) );
  OR2_X1 U318 ( .A1(n28), .A2(n457), .ZN(n276) );
  OAI21_X1 U319 ( .B1(n278), .B2(n277), .A(n276), .ZN(n419) );
  AOI22_X1 U320 ( .A1(n27), .A2(n523), .B1(n524), .B2(n384), .ZN(n526) );
  AOI22_X1 U321 ( .A1(n27), .A2(n522), .B1(n523), .B2(n384), .ZN(n528) );
  INV_X2 U322 ( .A(n295), .ZN(n383) );
  AND2_X1 U323 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n281) );
  NAND2_X1 U324 ( .A1(n28), .A2(n281), .ZN(n282) );
  OAI21_X1 U325 ( .B1(n383), .B2(n522), .A(n282), .ZN(n530) );
  AOI22_X1 U326 ( .A1(n27), .A2(n520), .B1(n521), .B2(n384), .ZN(n532) );
  AOI22_X1 U327 ( .A1(n27), .A2(n519), .B1(n520), .B2(n384), .ZN(n534) );
  OR2_X1 U328 ( .A1(n284), .A2(n283), .ZN(n285) );
  AND2_X1 U329 ( .A1(n285), .A2(n291), .ZN(n286) );
  NAND2_X1 U330 ( .A1(n29), .A2(n286), .ZN(n287) );
  OAI21_X1 U331 ( .B1(n28), .B2(n519), .A(n287), .ZN(n536) );
  AOI22_X1 U332 ( .A1(n27), .A2(n517), .B1(n518), .B2(n384), .ZN(n538) );
  AOI22_X1 U333 ( .A1(n27), .A2(n516), .B1(n517), .B2(n384), .ZN(n540) );
  INV_X1 U334 ( .A(n288), .ZN(n290) );
  NAND2_X1 U335 ( .A1(n290), .A2(n289), .ZN(n292) );
  XOR2_X1 U336 ( .A(n292), .B(n291), .Z(n293) );
  NAND2_X1 U337 ( .A1(n383), .A2(n293), .ZN(n294) );
  OAI21_X1 U338 ( .B1(n383), .B2(n516), .A(n294), .ZN(n542) );
  AOI22_X1 U339 ( .A1(n27), .A2(n514), .B1(n515), .B2(n384), .ZN(n544) );
  AOI22_X1 U340 ( .A1(n27), .A2(n513), .B1(n514), .B2(n384), .ZN(n546) );
  NAND2_X1 U341 ( .A1(n297), .A2(n296), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  NAND2_X1 U343 ( .A1(n28), .A2(n300), .ZN(n301) );
  OAI21_X1 U344 ( .B1(n27), .B2(n513), .A(n301), .ZN(n548) );
  AOI22_X1 U345 ( .A1(n27), .A2(n511), .B1(n512), .B2(n384), .ZN(n550) );
  AOI22_X1 U346 ( .A1(n27), .A2(n510), .B1(n511), .B2(n384), .ZN(n552) );
  INV_X1 U347 ( .A(n302), .ZN(n304) );
  NAND2_X1 U348 ( .A1(n304), .A2(n303), .ZN(n306) );
  XOR2_X1 U349 ( .A(n306), .B(n305), .Z(n307) );
  NAND2_X1 U350 ( .A1(n381), .A2(n307), .ZN(n308) );
  OAI21_X1 U351 ( .B1(n27), .B2(n510), .A(n308), .ZN(n554) );
  AOI22_X1 U352 ( .A1(n27), .A2(n508), .B1(n509), .B2(n384), .ZN(n556) );
  AOI22_X1 U353 ( .A1(n29), .A2(n507), .B1(n508), .B2(n357), .ZN(n558) );
  NAND2_X1 U354 ( .A1(n310), .A2(n309), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n313) );
  NAND2_X1 U356 ( .A1(n28), .A2(n313), .ZN(n314) );
  OAI21_X1 U357 ( .B1(n29), .B2(n507), .A(n314), .ZN(n560) );
  AOI22_X1 U358 ( .A1(n29), .A2(n505), .B1(n506), .B2(n357), .ZN(n562) );
  XOR2_X1 U359 ( .A(n397), .B(n404), .Z(n315) );
  NAND2_X1 U360 ( .A1(n29), .A2(n315), .ZN(n316) );
  OAI21_X1 U361 ( .B1(n27), .B2(n505), .A(n316), .ZN(n564) );
  AOI22_X1 U362 ( .A1(n381), .A2(n503), .B1(n504), .B2(n357), .ZN(n566) );
  NAND2_X1 U363 ( .A1(n387), .A2(n396), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n403), .B(n317), .ZN(n318) );
  NAND2_X1 U365 ( .A1(n383), .A2(n318), .ZN(n319) );
  OAI21_X1 U366 ( .B1(n381), .B2(n503), .A(n319), .ZN(n568) );
  AOI22_X1 U367 ( .A1(n29), .A2(n501), .B1(n502), .B2(n357), .ZN(n570) );
  AOI21_X1 U368 ( .B1(n403), .B2(n387), .A(n453), .ZN(n323) );
  NAND2_X1 U369 ( .A1(n455), .A2(n395), .ZN(n320) );
  XOR2_X1 U370 ( .A(n323), .B(n320), .Z(n321) );
  NAND2_X1 U371 ( .A1(n383), .A2(n321), .ZN(n322) );
  OAI21_X1 U372 ( .B1(n28), .B2(n501), .A(n322), .ZN(n572) );
  AOI22_X1 U373 ( .A1(n28), .A2(n499), .B1(n500), .B2(n357), .ZN(n574) );
  OAI21_X1 U374 ( .B1(n323), .B2(n394), .A(n395), .ZN(n333) );
  INV_X1 U375 ( .A(n333), .ZN(n327) );
  NAND2_X1 U376 ( .A1(n457), .A2(n393), .ZN(n324) );
  XOR2_X1 U377 ( .A(n327), .B(n324), .Z(n325) );
  NAND2_X1 U378 ( .A1(n383), .A2(n325), .ZN(n326) );
  OAI21_X1 U379 ( .B1(n383), .B2(n499), .A(n326), .ZN(n576) );
  AOI22_X1 U380 ( .A1(n383), .A2(n497), .B1(n498), .B2(n357), .ZN(n578) );
  OAI21_X1 U381 ( .B1(n327), .B2(n392), .A(n393), .ZN(n329) );
  NAND2_X1 U382 ( .A1(n451), .A2(n399), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  NAND2_X1 U384 ( .A1(n383), .A2(n330), .ZN(n331) );
  OAI21_X1 U385 ( .B1(n27), .B2(n497), .A(n331), .ZN(n580) );
  AOI22_X1 U386 ( .A1(n383), .A2(n495), .B1(n496), .B2(n357), .ZN(n582) );
  NOR2_X1 U387 ( .A1(n398), .A2(n392), .ZN(n334) );
  OAI21_X1 U388 ( .B1(n398), .B2(n393), .A(n399), .ZN(n332) );
  AOI21_X1 U389 ( .B1(n334), .B2(n333), .A(n332), .ZN(n362) );
  NAND2_X1 U390 ( .A1(n447), .A2(n391), .ZN(n335) );
  XOR2_X1 U391 ( .A(n362), .B(n335), .Z(n336) );
  NAND2_X1 U392 ( .A1(n29), .A2(n336), .ZN(n337) );
  OAI21_X1 U393 ( .B1(n27), .B2(n495), .A(n337), .ZN(n584) );
  AOI22_X1 U394 ( .A1(n27), .A2(n493), .B1(n494), .B2(n357), .ZN(n586) );
  OAI21_X1 U395 ( .B1(n362), .B2(n402), .A(n391), .ZN(n339) );
  NAND2_X1 U396 ( .A1(n401), .A2(n390), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  NAND2_X1 U398 ( .A1(n383), .A2(n340), .ZN(n341) );
  OAI21_X1 U399 ( .B1(n29), .B2(n493), .A(n341), .ZN(n588) );
  AOI22_X1 U400 ( .A1(n27), .A2(n491), .B1(n492), .B2(n384), .ZN(n590) );
  NAND2_X1 U401 ( .A1(n447), .A2(n401), .ZN(n343) );
  AOI21_X1 U402 ( .B1(n458), .B2(n401), .A(n459), .ZN(n342) );
  OAI21_X1 U403 ( .B1(n362), .B2(n343), .A(n342), .ZN(n345) );
  NAND2_X1 U404 ( .A1(n386), .A2(n400), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U406 ( .A1(n29), .A2(n346), .ZN(n347) );
  OAI21_X1 U407 ( .B1(n28), .B2(n491), .A(n347), .ZN(n592) );
  AOI22_X1 U408 ( .A1(n27), .A2(n489), .B1(n490), .B2(n384), .ZN(n594) );
  NAND2_X1 U409 ( .A1(n401), .A2(n386), .ZN(n350) );
  NOR2_X1 U410 ( .A1(n402), .A2(n350), .ZN(n358) );
  INV_X1 U411 ( .A(n358), .ZN(n352) );
  AOI21_X1 U412 ( .B1(n459), .B2(n386), .A(n449), .ZN(n349) );
  OAI21_X1 U413 ( .B1(n350), .B2(n391), .A(n349), .ZN(n359) );
  INV_X1 U414 ( .A(n359), .ZN(n351) );
  OAI21_X1 U415 ( .B1(n362), .B2(n352), .A(n351), .ZN(n354) );
  NAND2_X1 U416 ( .A1(n385), .A2(n389), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  NAND2_X1 U418 ( .A1(n383), .A2(n355), .ZN(n356) );
  OAI21_X1 U419 ( .B1(n27), .B2(n489), .A(n356), .ZN(n596) );
  AOI22_X1 U420 ( .A1(n27), .A2(n487), .B1(n488), .B2(n357), .ZN(n598) );
  NAND2_X1 U421 ( .A1(n358), .A2(n385), .ZN(n361) );
  AOI21_X1 U422 ( .B1(n359), .B2(n385), .A(n460), .ZN(n360) );
  OAI21_X1 U423 ( .B1(n362), .B2(n361), .A(n360), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n363), .B(n388), .ZN(n364) );
  NAND2_X1 U425 ( .A1(n383), .A2(n364), .ZN(n365) );
  OAI21_X1 U426 ( .B1(n28), .B2(n487), .A(n365), .ZN(n600) );
  NAND2_X1 U427 ( .A1(n381), .A2(B_extended[0]), .ZN(n366) );
  OAI21_X1 U428 ( .B1(n29), .B2(n486), .A(n366), .ZN(n602) );
  NAND2_X1 U429 ( .A1(n29), .A2(B_extended[1]), .ZN(n367) );
  OAI21_X1 U430 ( .B1(n28), .B2(n485), .A(n367), .ZN(n604) );
  NAND2_X1 U431 ( .A1(n381), .A2(B_extended[2]), .ZN(n368) );
  OAI21_X1 U432 ( .B1(n27), .B2(n484), .A(n368), .ZN(n606) );
  NAND2_X1 U433 ( .A1(n383), .A2(B_extended[3]), .ZN(n369) );
  OAI21_X1 U434 ( .B1(n381), .B2(n483), .A(n369), .ZN(n608) );
  NAND2_X1 U435 ( .A1(n383), .A2(B_extended[4]), .ZN(n370) );
  OAI21_X1 U436 ( .B1(n381), .B2(n482), .A(n370), .ZN(n610) );
  NAND2_X1 U437 ( .A1(n383), .A2(B_extended[5]), .ZN(n371) );
  OAI21_X1 U438 ( .B1(n27), .B2(n481), .A(n371), .ZN(n612) );
  NAND2_X1 U439 ( .A1(n381), .A2(B_extended[6]), .ZN(n372) );
  OAI21_X1 U440 ( .B1(n383), .B2(n480), .A(n372), .ZN(n614) );
  NAND2_X1 U441 ( .A1(n383), .A2(B_extended[7]), .ZN(n373) );
  OAI21_X1 U442 ( .B1(n381), .B2(n479), .A(n373), .ZN(n616) );
  NAND2_X1 U443 ( .A1(n383), .A2(A_extended[0]), .ZN(n374) );
  OAI21_X1 U444 ( .B1(n28), .B2(n478), .A(n374), .ZN(n618) );
  NAND2_X1 U445 ( .A1(n381), .A2(A_extended[1]), .ZN(n375) );
  OAI21_X1 U446 ( .B1(n29), .B2(n477), .A(n375), .ZN(n620) );
  NAND2_X1 U447 ( .A1(n28), .A2(A_extended[2]), .ZN(n376) );
  OAI21_X1 U448 ( .B1(n381), .B2(n476), .A(n376), .ZN(n622) );
  NAND2_X1 U449 ( .A1(n383), .A2(A_extended[3]), .ZN(n377) );
  OAI21_X1 U450 ( .B1(n27), .B2(n22), .A(n377), .ZN(n624) );
  NAND2_X1 U451 ( .A1(n253), .A2(A_extended[4]), .ZN(n378) );
  OAI21_X1 U452 ( .B1(n383), .B2(n474), .A(n378), .ZN(n626) );
  NAND2_X1 U453 ( .A1(n29), .A2(A_extended[5]), .ZN(n379) );
  OAI21_X1 U454 ( .B1(n27), .B2(n473), .A(n379), .ZN(n628) );
  NAND2_X1 U455 ( .A1(n348), .A2(A_extended[6]), .ZN(n380) );
  OAI21_X1 U456 ( .B1(n381), .B2(n472), .A(n380), .ZN(n630) );
  NAND2_X1 U457 ( .A1(n383), .A2(A_extended[7]), .ZN(n382) );
  OAI21_X1 U458 ( .B1(n28), .B2(n471), .A(n382), .ZN(n632) );
  NAND2_X1 U459 ( .A1(n470), .A2(n384), .ZN(n634) );
endmodule


module conv_128_32_opt ( clk, reset, s_valid_x, s_valid_f, m_ready_y, 
        s_data_in_x, s_data_in_f, s_ready_f, s_ready_x, m_valid_y, 
        m_data_out_y );
  input [7:0] s_data_in_x;
  input [7:0] s_data_in_f;
  output [20:0] m_data_out_y;
  input clk, reset, s_valid_x, s_valid_f, m_ready_y;
  output s_ready_f, s_ready_x, m_valid_y;
  wire   conv_done, xmem_full, \xmem_data[31][7] , \xmem_data[31][6] ,
         \xmem_data[31][5] , \xmem_data[31][4] , \xmem_data[31][3] ,
         \xmem_data[31][2] , \xmem_data[31][1] , \xmem_data[31][0] ,
         \xmem_data[30][7] , \xmem_data[30][6] , \xmem_data[30][5] ,
         \xmem_data[30][4] , \xmem_data[30][3] , \xmem_data[30][2] ,
         \xmem_data[30][1] , \xmem_data[30][0] , \xmem_data[29][7] ,
         \xmem_data[29][6] , \xmem_data[29][5] , \xmem_data[29][4] ,
         \xmem_data[29][3] , \xmem_data[29][2] , \xmem_data[29][1] ,
         \xmem_data[29][0] , \xmem_data[28][7] , \xmem_data[28][6] ,
         \xmem_data[28][5] , \xmem_data[28][4] , \xmem_data[28][3] ,
         \xmem_data[28][2] , \xmem_data[28][1] , \xmem_data[28][0] ,
         \xmem_data[27][7] , \xmem_data[27][6] , \xmem_data[27][5] ,
         \xmem_data[27][4] , \xmem_data[27][3] , \xmem_data[27][2] ,
         \xmem_data[27][1] , \xmem_data[27][0] , \xmem_data[26][7] ,
         \xmem_data[26][6] , \xmem_data[26][5] , \xmem_data[26][4] ,
         \xmem_data[26][3] , \xmem_data[26][2] , \xmem_data[26][1] ,
         \xmem_data[26][0] , \xmem_data[25][7] , \xmem_data[25][6] ,
         \xmem_data[25][5] , \xmem_data[25][4] , \xmem_data[25][3] ,
         \xmem_data[25][2] , \xmem_data[25][1] , \xmem_data[25][0] ,
         \xmem_data[24][7] , \xmem_data[24][6] , \xmem_data[24][5] ,
         \xmem_data[24][4] , \xmem_data[24][3] , \xmem_data[24][2] ,
         \xmem_data[24][1] , \xmem_data[24][0] , \xmem_data[23][7] ,
         \xmem_data[23][6] , \xmem_data[23][5] , \xmem_data[23][4] ,
         \xmem_data[23][3] , \xmem_data[23][2] , \xmem_data[23][1] ,
         \xmem_data[23][0] , \xmem_data[22][7] , \xmem_data[22][6] ,
         \xmem_data[22][5] , \xmem_data[22][4] , \xmem_data[22][3] ,
         \xmem_data[22][2] , \xmem_data[22][1] , \xmem_data[22][0] ,
         \xmem_data[21][7] , \xmem_data[21][6] , \xmem_data[21][5] ,
         \xmem_data[21][4] , \xmem_data[21][3] , \xmem_data[21][2] ,
         \xmem_data[21][1] , \xmem_data[21][0] , \xmem_data[20][7] ,
         \xmem_data[20][6] , \xmem_data[20][5] , \xmem_data[20][4] ,
         \xmem_data[20][3] , \xmem_data[20][2] , \xmem_data[20][1] ,
         \xmem_data[20][0] , \xmem_data[19][7] , \xmem_data[19][6] ,
         \xmem_data[19][5] , \xmem_data[19][4] , \xmem_data[19][3] ,
         \xmem_data[19][2] , \xmem_data[19][1] , \xmem_data[19][0] ,
         \xmem_data[18][7] , \xmem_data[18][6] , \xmem_data[18][5] ,
         \xmem_data[18][4] , \xmem_data[18][3] , \xmem_data[18][2] ,
         \xmem_data[18][1] , \xmem_data[18][0] , \xmem_data[17][7] ,
         \xmem_data[17][6] , \xmem_data[17][5] , \xmem_data[17][4] ,
         \xmem_data[17][3] , \xmem_data[17][2] , \xmem_data[17][1] ,
         \xmem_data[17][0] , \xmem_data[16][7] , \xmem_data[16][6] ,
         \xmem_data[16][5] , \xmem_data[16][4] , \xmem_data[16][3] ,
         \xmem_data[16][2] , \xmem_data[16][1] , \xmem_data[16][0] ,
         \xmem_data[15][7] , \xmem_data[15][6] , \xmem_data[15][5] ,
         \xmem_data[15][4] , \xmem_data[15][3] , \xmem_data[15][2] ,
         \xmem_data[15][1] , \xmem_data[15][0] , \xmem_data[14][7] ,
         \xmem_data[14][6] , \xmem_data[14][5] , \xmem_data[14][4] ,
         \xmem_data[14][3] , \xmem_data[14][2] , \xmem_data[14][1] ,
         \xmem_data[14][0] , \xmem_data[13][7] , \xmem_data[13][6] ,
         \xmem_data[13][5] , \xmem_data[13][4] , \xmem_data[13][3] ,
         \xmem_data[13][2] , \xmem_data[13][1] , \xmem_data[13][0] ,
         \xmem_data[12][7] , \xmem_data[12][6] , \xmem_data[12][5] ,
         \xmem_data[12][4] , \xmem_data[12][3] , \xmem_data[12][2] ,
         \xmem_data[12][1] , \xmem_data[12][0] , \xmem_data[11][7] ,
         \xmem_data[11][6] , \xmem_data[11][5] , \xmem_data[11][4] ,
         \xmem_data[11][3] , \xmem_data[11][2] , \xmem_data[11][1] ,
         \xmem_data[11][0] , \xmem_data[10][7] , \xmem_data[10][6] ,
         \xmem_data[10][5] , \xmem_data[10][4] , \xmem_data[10][3] ,
         \xmem_data[10][2] , \xmem_data[10][1] , \xmem_data[10][0] ,
         \xmem_data[9][7] , \xmem_data[9][6] , \xmem_data[9][5] ,
         \xmem_data[9][4] , \xmem_data[9][3] , \xmem_data[9][2] ,
         \xmem_data[9][1] , \xmem_data[9][0] , \xmem_data[8][7] ,
         \xmem_data[8][6] , \xmem_data[8][5] , \xmem_data[8][4] ,
         \xmem_data[8][3] , \xmem_data[8][2] , \xmem_data[8][1] ,
         \xmem_data[8][0] , \xmem_data[7][7] , \xmem_data[7][6] ,
         \xmem_data[7][5] , \xmem_data[7][4] , \xmem_data[7][3] ,
         \xmem_data[7][2] , \xmem_data[7][1] , \xmem_data[7][0] ,
         \xmem_data[6][7] , \xmem_data[6][6] , \xmem_data[6][5] ,
         \xmem_data[6][4] , \xmem_data[6][3] , \xmem_data[6][2] ,
         \xmem_data[6][1] , \xmem_data[6][0] , \xmem_data[5][7] ,
         \xmem_data[5][6] , \xmem_data[5][5] , \xmem_data[5][4] ,
         \xmem_data[5][3] , \xmem_data[5][2] , \xmem_data[5][1] ,
         \xmem_data[5][0] , \xmem_data[4][7] , \xmem_data[4][6] ,
         \xmem_data[4][5] , \xmem_data[4][4] , \xmem_data[4][3] ,
         \xmem_data[4][2] , \xmem_data[4][1] , \xmem_data[4][0] ,
         \xmem_data[3][7] , \xmem_data[3][6] , \xmem_data[3][5] ,
         \xmem_data[3][4] , \xmem_data[3][3] , \xmem_data[3][2] ,
         \xmem_data[3][1] , \xmem_data[3][0] , \xmem_data[2][7] ,
         \xmem_data[2][6] , \xmem_data[2][5] , \xmem_data[2][4] ,
         \xmem_data[2][3] , \xmem_data[2][2] , \xmem_data[2][1] ,
         \xmem_data[2][0] , \xmem_data[1][7] , \xmem_data[1][6] ,
         \xmem_data[1][5] , \xmem_data[1][4] , \xmem_data[1][3] ,
         \xmem_data[1][2] , \xmem_data[1][1] , \xmem_data[1][0] ,
         \xmem_data[0][7] , \xmem_data[0][6] , \xmem_data[0][5] ,
         \xmem_data[0][4] , \xmem_data[0][3] , \xmem_data[0][2] ,
         \xmem_data[0][1] , \xmem_data[0][0] , \fmem_data[31][7] ,
         \fmem_data[31][6] , \fmem_data[31][5] , \fmem_data[31][4] ,
         \fmem_data[31][3] , \fmem_data[31][2] , \fmem_data[31][1] ,
         \fmem_data[31][0] , \fmem_data[30][7] , \fmem_data[30][6] ,
         \fmem_data[30][5] , \fmem_data[30][4] , \fmem_data[30][3] ,
         \fmem_data[30][2] , \fmem_data[30][1] , \fmem_data[30][0] ,
         \fmem_data[29][7] , \fmem_data[29][6] , \fmem_data[29][5] ,
         \fmem_data[29][4] , \fmem_data[29][3] , \fmem_data[29][2] ,
         \fmem_data[29][1] , \fmem_data[29][0] , \fmem_data[28][7] ,
         \fmem_data[28][6] , \fmem_data[28][5] , \fmem_data[28][4] ,
         \fmem_data[28][3] , \fmem_data[28][2] , \fmem_data[28][1] ,
         \fmem_data[28][0] , \fmem_data[27][7] , \fmem_data[27][6] ,
         \fmem_data[27][5] , \fmem_data[27][4] , \fmem_data[27][3] ,
         \fmem_data[27][2] , \fmem_data[27][1] , \fmem_data[27][0] ,
         \fmem_data[26][7] , \fmem_data[26][6] , \fmem_data[26][5] ,
         \fmem_data[26][4] , \fmem_data[26][3] , \fmem_data[26][2] ,
         \fmem_data[26][1] , \fmem_data[26][0] , \fmem_data[25][7] ,
         \fmem_data[25][6] , \fmem_data[25][5] , \fmem_data[25][4] ,
         \fmem_data[25][3] , \fmem_data[25][2] , \fmem_data[25][1] ,
         \fmem_data[25][0] , \fmem_data[24][7] , \fmem_data[24][6] ,
         \fmem_data[24][5] , \fmem_data[24][4] , \fmem_data[24][3] ,
         \fmem_data[24][2] , \fmem_data[24][1] , \fmem_data[24][0] ,
         \fmem_data[23][7] , \fmem_data[23][6] , \fmem_data[23][5] ,
         \fmem_data[23][4] , \fmem_data[23][3] , \fmem_data[23][2] ,
         \fmem_data[23][1] , \fmem_data[23][0] , \fmem_data[22][7] ,
         \fmem_data[22][6] , \fmem_data[22][5] , \fmem_data[22][4] ,
         \fmem_data[22][3] , \fmem_data[22][2] , \fmem_data[22][1] ,
         \fmem_data[22][0] , \fmem_data[21][7] , \fmem_data[21][6] ,
         \fmem_data[21][5] , \fmem_data[21][4] , \fmem_data[21][3] ,
         \fmem_data[21][2] , \fmem_data[21][1] , \fmem_data[21][0] ,
         \fmem_data[20][7] , \fmem_data[20][6] , \fmem_data[20][5] ,
         \fmem_data[20][4] , \fmem_data[20][3] , \fmem_data[20][2] ,
         \fmem_data[20][1] , \fmem_data[20][0] , \fmem_data[19][7] ,
         \fmem_data[19][6] , \fmem_data[19][5] , \fmem_data[19][4] ,
         \fmem_data[19][3] , \fmem_data[19][2] , \fmem_data[19][1] ,
         \fmem_data[19][0] , \fmem_data[18][7] , \fmem_data[18][6] ,
         \fmem_data[18][5] , \fmem_data[18][4] , \fmem_data[18][3] ,
         \fmem_data[18][2] , \fmem_data[18][1] , \fmem_data[18][0] ,
         \fmem_data[17][7] , \fmem_data[17][6] , \fmem_data[17][5] ,
         \fmem_data[17][4] , \fmem_data[17][3] , \fmem_data[17][2] ,
         \fmem_data[17][1] , \fmem_data[17][0] , \fmem_data[16][7] ,
         \fmem_data[16][6] , \fmem_data[16][5] , \fmem_data[16][4] ,
         \fmem_data[16][3] , \fmem_data[16][2] , \fmem_data[16][1] ,
         \fmem_data[16][0] , \fmem_data[15][7] , \fmem_data[15][6] ,
         \fmem_data[15][5] , \fmem_data[15][4] , \fmem_data[15][3] ,
         \fmem_data[15][2] , \fmem_data[15][1] , \fmem_data[15][0] ,
         \fmem_data[14][7] , \fmem_data[14][6] , \fmem_data[14][5] ,
         \fmem_data[14][4] , \fmem_data[14][3] , \fmem_data[14][2] ,
         \fmem_data[14][1] , \fmem_data[14][0] , \fmem_data[13][7] ,
         \fmem_data[13][6] , \fmem_data[13][5] , \fmem_data[13][4] ,
         \fmem_data[13][3] , \fmem_data[13][2] , \fmem_data[13][1] ,
         \fmem_data[13][0] , \fmem_data[12][7] , \fmem_data[12][6] ,
         \fmem_data[12][5] , \fmem_data[12][4] , \fmem_data[12][3] ,
         \fmem_data[12][2] , \fmem_data[12][1] , \fmem_data[12][0] ,
         \fmem_data[11][7] , \fmem_data[11][6] , \fmem_data[11][5] ,
         \fmem_data[11][4] , \fmem_data[11][3] , \fmem_data[11][2] ,
         \fmem_data[11][1] , \fmem_data[11][0] , \fmem_data[10][7] ,
         \fmem_data[10][6] , \fmem_data[10][5] , \fmem_data[10][4] ,
         \fmem_data[10][3] , \fmem_data[10][2] , \fmem_data[10][1] ,
         \fmem_data[10][0] , \fmem_data[9][7] , \fmem_data[9][6] ,
         \fmem_data[9][5] , \fmem_data[9][4] , \fmem_data[9][3] ,
         \fmem_data[9][2] , \fmem_data[9][1] , \fmem_data[9][0] ,
         \fmem_data[8][7] , \fmem_data[8][6] , \fmem_data[8][5] ,
         \fmem_data[8][4] , \fmem_data[8][3] , \fmem_data[8][2] ,
         \fmem_data[8][1] , \fmem_data[8][0] , \fmem_data[7][7] ,
         \fmem_data[7][6] , \fmem_data[7][5] , \fmem_data[7][4] ,
         \fmem_data[7][3] , \fmem_data[7][2] , \fmem_data[7][1] ,
         \fmem_data[7][0] , \fmem_data[6][7] , \fmem_data[6][6] ,
         \fmem_data[6][5] , \fmem_data[6][4] , \fmem_data[6][3] ,
         \fmem_data[6][2] , \fmem_data[6][1] , \fmem_data[6][0] ,
         \fmem_data[5][7] , \fmem_data[5][6] , \fmem_data[5][5] ,
         \fmem_data[5][4] , \fmem_data[5][3] , \fmem_data[5][2] ,
         \fmem_data[5][1] , \fmem_data[5][0] , \fmem_data[4][7] ,
         \fmem_data[4][6] , \fmem_data[4][5] , \fmem_data[4][4] ,
         \fmem_data[4][3] , \fmem_data[4][2] , \fmem_data[4][1] ,
         \fmem_data[4][0] , \fmem_data[3][7] , \fmem_data[3][6] ,
         \fmem_data[3][5] , \fmem_data[3][4] , \fmem_data[3][3] ,
         \fmem_data[3][2] , \fmem_data[3][1] , \fmem_data[3][0] ,
         \fmem_data[2][7] , \fmem_data[2][6] , \fmem_data[2][5] ,
         \fmem_data[2][4] , \fmem_data[2][3] , \fmem_data[2][2] ,
         \fmem_data[2][1] , \fmem_data[2][0] , \fmem_data[1][7] ,
         \fmem_data[1][6] , \fmem_data[1][5] , \fmem_data[1][4] ,
         \fmem_data[1][3] , \fmem_data[1][2] , \fmem_data[1][1] ,
         \fmem_data[1][0] , \fmem_data[0][7] , \fmem_data[0][6] ,
         \fmem_data[0][5] , \fmem_data[0][4] , \fmem_data[0][3] ,
         \fmem_data[0][2] , \fmem_data[0][1] , \fmem_data[0][0] ,
         \x_mult_f_int[31][15] , \x_mult_f_int[31][14] ,
         \x_mult_f_int[31][13] , \x_mult_f_int[31][12] ,
         \x_mult_f_int[31][11] , \x_mult_f_int[31][10] , \x_mult_f_int[31][9] ,
         \x_mult_f_int[31][8] , \x_mult_f_int[31][7] , \x_mult_f_int[31][6] ,
         \x_mult_f_int[31][5] , \x_mult_f_int[31][4] , \x_mult_f_int[31][3] ,
         \x_mult_f_int[31][2] , \x_mult_f_int[31][1] , \x_mult_f_int[31][0] ,
         \x_mult_f_int[30][15] , \x_mult_f_int[30][14] ,
         \x_mult_f_int[30][13] , \x_mult_f_int[30][12] ,
         \x_mult_f_int[30][11] , \x_mult_f_int[30][10] , \x_mult_f_int[30][9] ,
         \x_mult_f_int[30][8] , \x_mult_f_int[30][7] , \x_mult_f_int[30][6] ,
         \x_mult_f_int[30][5] , \x_mult_f_int[30][4] , \x_mult_f_int[30][3] ,
         \x_mult_f_int[30][2] , \x_mult_f_int[30][1] , \x_mult_f_int[30][0] ,
         \x_mult_f_int[29][15] , \x_mult_f_int[29][14] ,
         \x_mult_f_int[29][13] , \x_mult_f_int[29][12] ,
         \x_mult_f_int[29][11] , \x_mult_f_int[29][10] , \x_mult_f_int[29][9] ,
         \x_mult_f_int[29][8] , \x_mult_f_int[29][7] , \x_mult_f_int[29][6] ,
         \x_mult_f_int[29][5] , \x_mult_f_int[29][4] , \x_mult_f_int[29][3] ,
         \x_mult_f_int[29][2] , \x_mult_f_int[29][1] , \x_mult_f_int[29][0] ,
         \x_mult_f_int[28][15] , \x_mult_f_int[28][14] ,
         \x_mult_f_int[28][13] , \x_mult_f_int[28][12] ,
         \x_mult_f_int[28][11] , \x_mult_f_int[28][10] , \x_mult_f_int[28][9] ,
         \x_mult_f_int[28][8] , \x_mult_f_int[28][7] , \x_mult_f_int[28][6] ,
         \x_mult_f_int[28][5] , \x_mult_f_int[28][4] , \x_mult_f_int[28][3] ,
         \x_mult_f_int[28][2] , \x_mult_f_int[28][1] , \x_mult_f_int[28][0] ,
         \x_mult_f_int[27][15] , \x_mult_f_int[27][14] ,
         \x_mult_f_int[27][13] , \x_mult_f_int[27][12] ,
         \x_mult_f_int[27][11] , \x_mult_f_int[27][10] , \x_mult_f_int[27][9] ,
         \x_mult_f_int[27][8] , \x_mult_f_int[27][7] , \x_mult_f_int[27][6] ,
         \x_mult_f_int[27][5] , \x_mult_f_int[27][4] , \x_mult_f_int[27][3] ,
         \x_mult_f_int[27][2] , \x_mult_f_int[27][1] , \x_mult_f_int[27][0] ,
         \x_mult_f_int[26][15] , \x_mult_f_int[26][14] ,
         \x_mult_f_int[26][13] , \x_mult_f_int[26][12] ,
         \x_mult_f_int[26][11] , \x_mult_f_int[26][10] , \x_mult_f_int[26][9] ,
         \x_mult_f_int[26][8] , \x_mult_f_int[26][7] , \x_mult_f_int[26][6] ,
         \x_mult_f_int[26][5] , \x_mult_f_int[26][4] , \x_mult_f_int[26][3] ,
         \x_mult_f_int[26][2] , \x_mult_f_int[26][1] , \x_mult_f_int[26][0] ,
         \x_mult_f_int[25][15] , \x_mult_f_int[25][14] ,
         \x_mult_f_int[25][13] , \x_mult_f_int[25][12] ,
         \x_mult_f_int[25][11] , \x_mult_f_int[25][10] , \x_mult_f_int[25][9] ,
         \x_mult_f_int[25][8] , \x_mult_f_int[25][7] , \x_mult_f_int[25][6] ,
         \x_mult_f_int[25][5] , \x_mult_f_int[25][4] , \x_mult_f_int[25][3] ,
         \x_mult_f_int[25][2] , \x_mult_f_int[25][1] , \x_mult_f_int[25][0] ,
         \x_mult_f_int[24][15] , \x_mult_f_int[24][14] ,
         \x_mult_f_int[24][13] , \x_mult_f_int[24][12] ,
         \x_mult_f_int[24][11] , \x_mult_f_int[24][10] , \x_mult_f_int[24][9] ,
         \x_mult_f_int[24][8] , \x_mult_f_int[24][7] , \x_mult_f_int[24][6] ,
         \x_mult_f_int[24][5] , \x_mult_f_int[24][4] , \x_mult_f_int[24][3] ,
         \x_mult_f_int[24][2] , \x_mult_f_int[24][1] , \x_mult_f_int[24][0] ,
         \x_mult_f_int[23][15] , \x_mult_f_int[23][14] ,
         \x_mult_f_int[23][13] , \x_mult_f_int[23][12] ,
         \x_mult_f_int[23][11] , \x_mult_f_int[23][10] , \x_mult_f_int[23][9] ,
         \x_mult_f_int[23][8] , \x_mult_f_int[23][7] , \x_mult_f_int[23][6] ,
         \x_mult_f_int[23][5] , \x_mult_f_int[23][4] , \x_mult_f_int[23][3] ,
         \x_mult_f_int[23][2] , \x_mult_f_int[23][1] , \x_mult_f_int[23][0] ,
         \x_mult_f_int[22][15] , \x_mult_f_int[22][14] ,
         \x_mult_f_int[22][13] , \x_mult_f_int[22][12] ,
         \x_mult_f_int[22][11] , \x_mult_f_int[22][10] , \x_mult_f_int[22][9] ,
         \x_mult_f_int[22][8] , \x_mult_f_int[22][7] , \x_mult_f_int[22][6] ,
         \x_mult_f_int[22][5] , \x_mult_f_int[22][4] , \x_mult_f_int[22][3] ,
         \x_mult_f_int[22][2] , \x_mult_f_int[22][1] , \x_mult_f_int[22][0] ,
         \x_mult_f_int[21][15] , \x_mult_f_int[21][14] ,
         \x_mult_f_int[21][13] , \x_mult_f_int[21][12] ,
         \x_mult_f_int[21][11] , \x_mult_f_int[21][10] , \x_mult_f_int[21][9] ,
         \x_mult_f_int[21][8] , \x_mult_f_int[21][7] , \x_mult_f_int[21][6] ,
         \x_mult_f_int[21][5] , \x_mult_f_int[21][4] , \x_mult_f_int[21][3] ,
         \x_mult_f_int[21][2] , \x_mult_f_int[21][1] , \x_mult_f_int[21][0] ,
         \x_mult_f_int[20][15] , \x_mult_f_int[20][14] ,
         \x_mult_f_int[20][13] , \x_mult_f_int[20][12] ,
         \x_mult_f_int[20][11] , \x_mult_f_int[20][10] , \x_mult_f_int[20][9] ,
         \x_mult_f_int[20][8] , \x_mult_f_int[20][7] , \x_mult_f_int[20][6] ,
         \x_mult_f_int[20][5] , \x_mult_f_int[20][4] , \x_mult_f_int[20][3] ,
         \x_mult_f_int[20][2] , \x_mult_f_int[20][1] , \x_mult_f_int[20][0] ,
         \x_mult_f_int[19][15] , \x_mult_f_int[19][14] ,
         \x_mult_f_int[19][13] , \x_mult_f_int[19][12] ,
         \x_mult_f_int[19][11] , \x_mult_f_int[19][10] , \x_mult_f_int[19][9] ,
         \x_mult_f_int[19][8] , \x_mult_f_int[19][7] , \x_mult_f_int[19][6] ,
         \x_mult_f_int[19][5] , \x_mult_f_int[19][4] , \x_mult_f_int[19][3] ,
         \x_mult_f_int[19][2] , \x_mult_f_int[19][1] , \x_mult_f_int[19][0] ,
         \x_mult_f_int[18][15] , \x_mult_f_int[18][14] ,
         \x_mult_f_int[18][13] , \x_mult_f_int[18][12] ,
         \x_mult_f_int[18][11] , \x_mult_f_int[18][10] , \x_mult_f_int[18][9] ,
         \x_mult_f_int[18][8] , \x_mult_f_int[18][7] , \x_mult_f_int[18][6] ,
         \x_mult_f_int[18][5] , \x_mult_f_int[18][4] , \x_mult_f_int[18][3] ,
         \x_mult_f_int[18][2] , \x_mult_f_int[18][1] , \x_mult_f_int[18][0] ,
         \x_mult_f_int[17][15] , \x_mult_f_int[17][14] ,
         \x_mult_f_int[17][13] , \x_mult_f_int[17][12] ,
         \x_mult_f_int[17][11] , \x_mult_f_int[17][10] , \x_mult_f_int[17][9] ,
         \x_mult_f_int[17][8] , \x_mult_f_int[17][7] , \x_mult_f_int[17][6] ,
         \x_mult_f_int[17][5] , \x_mult_f_int[17][4] , \x_mult_f_int[17][3] ,
         \x_mult_f_int[17][2] , \x_mult_f_int[17][1] , \x_mult_f_int[17][0] ,
         \x_mult_f_int[16][15] , \x_mult_f_int[16][14] ,
         \x_mult_f_int[16][13] , \x_mult_f_int[16][12] ,
         \x_mult_f_int[16][11] , \x_mult_f_int[16][10] , \x_mult_f_int[16][9] ,
         \x_mult_f_int[16][8] , \x_mult_f_int[16][7] , \x_mult_f_int[16][6] ,
         \x_mult_f_int[16][5] , \x_mult_f_int[16][4] , \x_mult_f_int[16][3] ,
         \x_mult_f_int[16][2] , \x_mult_f_int[16][1] , \x_mult_f_int[16][0] ,
         \x_mult_f_int[15][15] , \x_mult_f_int[15][14] ,
         \x_mult_f_int[15][13] , \x_mult_f_int[15][12] ,
         \x_mult_f_int[15][11] , \x_mult_f_int[15][10] , \x_mult_f_int[15][9] ,
         \x_mult_f_int[15][8] , \x_mult_f_int[15][7] , \x_mult_f_int[15][6] ,
         \x_mult_f_int[15][5] , \x_mult_f_int[15][4] , \x_mult_f_int[15][3] ,
         \x_mult_f_int[15][2] , \x_mult_f_int[15][1] , \x_mult_f_int[15][0] ,
         \x_mult_f_int[14][15] , \x_mult_f_int[14][14] ,
         \x_mult_f_int[14][13] , \x_mult_f_int[14][12] ,
         \x_mult_f_int[14][11] , \x_mult_f_int[14][10] , \x_mult_f_int[14][9] ,
         \x_mult_f_int[14][8] , \x_mult_f_int[14][7] , \x_mult_f_int[14][6] ,
         \x_mult_f_int[14][5] , \x_mult_f_int[14][4] , \x_mult_f_int[14][3] ,
         \x_mult_f_int[14][2] , \x_mult_f_int[14][1] , \x_mult_f_int[14][0] ,
         \x_mult_f_int[13][15] , \x_mult_f_int[13][14] ,
         \x_mult_f_int[13][13] , \x_mult_f_int[13][12] ,
         \x_mult_f_int[13][11] , \x_mult_f_int[13][10] , \x_mult_f_int[13][9] ,
         \x_mult_f_int[13][8] , \x_mult_f_int[13][7] , \x_mult_f_int[13][6] ,
         \x_mult_f_int[13][5] , \x_mult_f_int[13][4] , \x_mult_f_int[13][3] ,
         \x_mult_f_int[13][2] , \x_mult_f_int[13][1] , \x_mult_f_int[13][0] ,
         \x_mult_f_int[12][15] , \x_mult_f_int[12][14] ,
         \x_mult_f_int[12][13] , \x_mult_f_int[12][12] ,
         \x_mult_f_int[12][11] , \x_mult_f_int[12][10] , \x_mult_f_int[12][9] ,
         \x_mult_f_int[12][8] , \x_mult_f_int[12][7] , \x_mult_f_int[12][6] ,
         \x_mult_f_int[12][5] , \x_mult_f_int[12][4] , \x_mult_f_int[12][3] ,
         \x_mult_f_int[12][2] , \x_mult_f_int[12][1] , \x_mult_f_int[12][0] ,
         \x_mult_f_int[11][15] , \x_mult_f_int[11][14] ,
         \x_mult_f_int[11][13] , \x_mult_f_int[11][12] ,
         \x_mult_f_int[11][11] , \x_mult_f_int[11][10] , \x_mult_f_int[11][9] ,
         \x_mult_f_int[11][8] , \x_mult_f_int[11][7] , \x_mult_f_int[11][6] ,
         \x_mult_f_int[11][5] , \x_mult_f_int[11][4] , \x_mult_f_int[11][3] ,
         \x_mult_f_int[11][2] , \x_mult_f_int[11][1] , \x_mult_f_int[11][0] ,
         \x_mult_f_int[10][15] , \x_mult_f_int[10][14] ,
         \x_mult_f_int[10][13] , \x_mult_f_int[10][12] ,
         \x_mult_f_int[10][11] , \x_mult_f_int[10][10] , \x_mult_f_int[10][9] ,
         \x_mult_f_int[10][8] , \x_mult_f_int[10][7] , \x_mult_f_int[10][6] ,
         \x_mult_f_int[10][5] , \x_mult_f_int[10][4] , \x_mult_f_int[10][3] ,
         \x_mult_f_int[10][2] , \x_mult_f_int[10][1] , \x_mult_f_int[10][0] ,
         \x_mult_f_int[9][15] , \x_mult_f_int[9][14] , \x_mult_f_int[9][13] ,
         \x_mult_f_int[9][12] , \x_mult_f_int[9][11] , \x_mult_f_int[9][10] ,
         \x_mult_f_int[9][9] , \x_mult_f_int[9][8] , \x_mult_f_int[9][7] ,
         \x_mult_f_int[9][6] , \x_mult_f_int[9][5] , \x_mult_f_int[9][4] ,
         \x_mult_f_int[9][3] , \x_mult_f_int[9][2] , \x_mult_f_int[9][1] ,
         \x_mult_f_int[9][0] , \x_mult_f_int[8][15] , \x_mult_f_int[8][14] ,
         \x_mult_f_int[8][13] , \x_mult_f_int[8][12] , \x_mult_f_int[8][11] ,
         \x_mult_f_int[8][10] , \x_mult_f_int[8][9] , \x_mult_f_int[8][8] ,
         \x_mult_f_int[8][7] , \x_mult_f_int[8][6] , \x_mult_f_int[8][5] ,
         \x_mult_f_int[8][4] , \x_mult_f_int[8][3] , \x_mult_f_int[8][2] ,
         \x_mult_f_int[8][1] , \x_mult_f_int[8][0] , \x_mult_f_int[7][15] ,
         \x_mult_f_int[7][14] , \x_mult_f_int[7][13] , \x_mult_f_int[7][12] ,
         \x_mult_f_int[7][11] , \x_mult_f_int[7][10] , \x_mult_f_int[7][9] ,
         \x_mult_f_int[7][8] , \x_mult_f_int[7][7] , \x_mult_f_int[7][6] ,
         \x_mult_f_int[7][5] , \x_mult_f_int[7][4] , \x_mult_f_int[7][3] ,
         \x_mult_f_int[7][2] , \x_mult_f_int[7][1] , \x_mult_f_int[7][0] ,
         \x_mult_f_int[6][15] , \x_mult_f_int[6][14] , \x_mult_f_int[6][13] ,
         \x_mult_f_int[6][12] , \x_mult_f_int[6][11] , \x_mult_f_int[6][10] ,
         \x_mult_f_int[6][9] , \x_mult_f_int[6][8] , \x_mult_f_int[6][7] ,
         \x_mult_f_int[6][6] , \x_mult_f_int[6][5] , \x_mult_f_int[6][4] ,
         \x_mult_f_int[6][3] , \x_mult_f_int[6][2] , \x_mult_f_int[6][1] ,
         \x_mult_f_int[6][0] , \x_mult_f_int[5][15] , \x_mult_f_int[5][14] ,
         \x_mult_f_int[5][13] , \x_mult_f_int[5][12] , \x_mult_f_int[5][11] ,
         \x_mult_f_int[5][10] , \x_mult_f_int[5][9] , \x_mult_f_int[5][8] ,
         \x_mult_f_int[5][7] , \x_mult_f_int[5][6] , \x_mult_f_int[5][5] ,
         \x_mult_f_int[5][4] , \x_mult_f_int[5][3] , \x_mult_f_int[5][2] ,
         \x_mult_f_int[5][1] , \x_mult_f_int[5][0] , \x_mult_f_int[4][15] ,
         \x_mult_f_int[4][14] , \x_mult_f_int[4][13] , \x_mult_f_int[4][12] ,
         \x_mult_f_int[4][11] , \x_mult_f_int[4][10] , \x_mult_f_int[4][9] ,
         \x_mult_f_int[4][8] , \x_mult_f_int[4][7] , \x_mult_f_int[4][6] ,
         \x_mult_f_int[4][5] , \x_mult_f_int[4][4] , \x_mult_f_int[4][3] ,
         \x_mult_f_int[4][2] , \x_mult_f_int[4][1] , \x_mult_f_int[4][0] ,
         \x_mult_f_int[3][15] , \x_mult_f_int[3][14] , \x_mult_f_int[3][13] ,
         \x_mult_f_int[3][12] , \x_mult_f_int[3][11] , \x_mult_f_int[3][10] ,
         \x_mult_f_int[3][9] , \x_mult_f_int[3][8] , \x_mult_f_int[3][7] ,
         \x_mult_f_int[3][6] , \x_mult_f_int[3][5] , \x_mult_f_int[3][4] ,
         \x_mult_f_int[3][3] , \x_mult_f_int[3][2] , \x_mult_f_int[3][1] ,
         \x_mult_f_int[3][0] , \x_mult_f_int[2][15] , \x_mult_f_int[2][14] ,
         \x_mult_f_int[2][13] , \x_mult_f_int[2][12] , \x_mult_f_int[2][11] ,
         \x_mult_f_int[2][10] , \x_mult_f_int[2][9] , \x_mult_f_int[2][8] ,
         \x_mult_f_int[2][7] , \x_mult_f_int[2][6] , \x_mult_f_int[2][5] ,
         \x_mult_f_int[2][4] , \x_mult_f_int[2][3] , \x_mult_f_int[2][2] ,
         \x_mult_f_int[2][1] , \x_mult_f_int[2][0] , \x_mult_f_int[1][15] ,
         \x_mult_f_int[1][14] , \x_mult_f_int[1][13] , \x_mult_f_int[1][12] ,
         \x_mult_f_int[1][11] , \x_mult_f_int[1][10] , \x_mult_f_int[1][9] ,
         \x_mult_f_int[1][8] , \x_mult_f_int[1][7] , \x_mult_f_int[1][6] ,
         \x_mult_f_int[1][5] , \x_mult_f_int[1][4] , \x_mult_f_int[1][3] ,
         \x_mult_f_int[1][2] , \x_mult_f_int[1][1] , \x_mult_f_int[1][0] ,
         \x_mult_f_int[0][15] , \x_mult_f_int[0][14] , \x_mult_f_int[0][13] ,
         \x_mult_f_int[0][12] , \x_mult_f_int[0][11] , \x_mult_f_int[0][10] ,
         \x_mult_f_int[0][9] , \x_mult_f_int[0][8] , \x_mult_f_int[0][7] ,
         \x_mult_f_int[0][6] , \x_mult_f_int[0][5] , \x_mult_f_int[0][4] ,
         \x_mult_f_int[0][3] , \x_mult_f_int[0][2] , \x_mult_f_int[0][1] ,
         \x_mult_f_int[0][0] , \x_mult_f[31][15] , \x_mult_f[31][14] ,
         \x_mult_f[31][13] , \x_mult_f[31][12] , \x_mult_f[31][11] ,
         \x_mult_f[31][10] , \x_mult_f[31][9] , \x_mult_f[31][8] ,
         \x_mult_f[31][7] , \x_mult_f[31][6] , \x_mult_f[31][5] ,
         \x_mult_f[31][4] , \x_mult_f[31][3] , \x_mult_f[31][2] ,
         \x_mult_f[31][1] , \x_mult_f[31][0] , \x_mult_f[30][15] ,
         \x_mult_f[30][14] , \x_mult_f[30][13] , \x_mult_f[30][12] ,
         \x_mult_f[30][11] , \x_mult_f[30][10] , \x_mult_f[30][9] ,
         \x_mult_f[30][8] , \x_mult_f[30][7] , \x_mult_f[30][6] ,
         \x_mult_f[30][5] , \x_mult_f[30][4] , \x_mult_f[30][3] ,
         \x_mult_f[30][2] , \x_mult_f[30][1] , \x_mult_f[30][0] ,
         \x_mult_f[29][15] , \x_mult_f[29][14] , \x_mult_f[29][13] ,
         \x_mult_f[29][12] , \x_mult_f[29][11] , \x_mult_f[29][10] ,
         \x_mult_f[29][9] , \x_mult_f[29][8] , \x_mult_f[29][7] ,
         \x_mult_f[29][6] , \x_mult_f[29][5] , \x_mult_f[29][4] ,
         \x_mult_f[29][3] , \x_mult_f[29][2] , \x_mult_f[29][1] ,
         \x_mult_f[29][0] , \x_mult_f[28][15] , \x_mult_f[28][14] ,
         \x_mult_f[28][13] , \x_mult_f[28][12] , \x_mult_f[28][11] ,
         \x_mult_f[28][10] , \x_mult_f[28][9] , \x_mult_f[28][8] ,
         \x_mult_f[28][7] , \x_mult_f[28][6] , \x_mult_f[28][5] ,
         \x_mult_f[28][4] , \x_mult_f[28][3] , \x_mult_f[28][2] ,
         \x_mult_f[28][1] , \x_mult_f[28][0] , \x_mult_f[27][15] ,
         \x_mult_f[27][14] , \x_mult_f[27][13] , \x_mult_f[27][12] ,
         \x_mult_f[27][11] , \x_mult_f[27][10] , \x_mult_f[27][9] ,
         \x_mult_f[27][8] , \x_mult_f[27][7] , \x_mult_f[27][6] ,
         \x_mult_f[27][5] , \x_mult_f[27][4] , \x_mult_f[27][3] ,
         \x_mult_f[27][2] , \x_mult_f[27][1] , \x_mult_f[27][0] ,
         \x_mult_f[26][15] , \x_mult_f[26][14] , \x_mult_f[26][13] ,
         \x_mult_f[26][12] , \x_mult_f[26][11] , \x_mult_f[26][10] ,
         \x_mult_f[26][9] , \x_mult_f[26][8] , \x_mult_f[26][7] ,
         \x_mult_f[26][6] , \x_mult_f[26][5] , \x_mult_f[26][4] ,
         \x_mult_f[26][3] , \x_mult_f[26][2] , \x_mult_f[26][1] ,
         \x_mult_f[26][0] , \x_mult_f[25][15] , \x_mult_f[25][14] ,
         \x_mult_f[25][13] , \x_mult_f[25][12] , \x_mult_f[25][11] ,
         \x_mult_f[25][10] , \x_mult_f[25][9] , \x_mult_f[25][8] ,
         \x_mult_f[25][7] , \x_mult_f[25][6] , \x_mult_f[25][5] ,
         \x_mult_f[25][4] , \x_mult_f[25][3] , \x_mult_f[25][2] ,
         \x_mult_f[25][1] , \x_mult_f[25][0] , \x_mult_f[24][15] ,
         \x_mult_f[24][14] , \x_mult_f[24][13] , \x_mult_f[24][12] ,
         \x_mult_f[24][11] , \x_mult_f[24][10] , \x_mult_f[24][9] ,
         \x_mult_f[24][8] , \x_mult_f[24][7] , \x_mult_f[24][6] ,
         \x_mult_f[24][5] , \x_mult_f[24][4] , \x_mult_f[24][3] ,
         \x_mult_f[24][2] , \x_mult_f[24][1] , \x_mult_f[24][0] ,
         \x_mult_f[23][15] , \x_mult_f[23][14] , \x_mult_f[23][13] ,
         \x_mult_f[23][12] , \x_mult_f[23][11] , \x_mult_f[23][10] ,
         \x_mult_f[23][9] , \x_mult_f[23][8] , \x_mult_f[23][7] ,
         \x_mult_f[23][6] , \x_mult_f[23][5] , \x_mult_f[23][4] ,
         \x_mult_f[23][3] , \x_mult_f[23][2] , \x_mult_f[23][1] ,
         \x_mult_f[23][0] , \x_mult_f[22][15] , \x_mult_f[22][14] ,
         \x_mult_f[22][13] , \x_mult_f[22][12] , \x_mult_f[22][11] ,
         \x_mult_f[22][10] , \x_mult_f[22][9] , \x_mult_f[22][8] ,
         \x_mult_f[22][7] , \x_mult_f[22][6] , \x_mult_f[22][5] ,
         \x_mult_f[22][4] , \x_mult_f[22][3] , \x_mult_f[22][2] ,
         \x_mult_f[22][1] , \x_mult_f[22][0] , \x_mult_f[21][15] ,
         \x_mult_f[21][14] , \x_mult_f[21][13] , \x_mult_f[21][12] ,
         \x_mult_f[21][11] , \x_mult_f[21][10] , \x_mult_f[21][9] ,
         \x_mult_f[21][8] , \x_mult_f[21][7] , \x_mult_f[21][6] ,
         \x_mult_f[21][5] , \x_mult_f[21][4] , \x_mult_f[21][3] ,
         \x_mult_f[21][2] , \x_mult_f[21][1] , \x_mult_f[21][0] ,
         \x_mult_f[20][15] , \x_mult_f[20][14] , \x_mult_f[20][13] ,
         \x_mult_f[20][12] , \x_mult_f[20][11] , \x_mult_f[20][10] ,
         \x_mult_f[20][9] , \x_mult_f[20][8] , \x_mult_f[20][7] ,
         \x_mult_f[20][6] , \x_mult_f[20][5] , \x_mult_f[20][4] ,
         \x_mult_f[20][3] , \x_mult_f[20][2] , \x_mult_f[20][1] ,
         \x_mult_f[20][0] , \x_mult_f[19][15] , \x_mult_f[19][14] ,
         \x_mult_f[19][13] , \x_mult_f[19][12] , \x_mult_f[19][11] ,
         \x_mult_f[19][10] , \x_mult_f[19][9] , \x_mult_f[19][8] ,
         \x_mult_f[19][7] , \x_mult_f[19][6] , \x_mult_f[19][5] ,
         \x_mult_f[19][4] , \x_mult_f[19][3] , \x_mult_f[19][2] ,
         \x_mult_f[19][1] , \x_mult_f[19][0] , \x_mult_f[18][15] ,
         \x_mult_f[18][14] , \x_mult_f[18][13] , \x_mult_f[18][12] ,
         \x_mult_f[18][11] , \x_mult_f[18][10] , \x_mult_f[18][9] ,
         \x_mult_f[18][8] , \x_mult_f[18][7] , \x_mult_f[18][6] ,
         \x_mult_f[18][5] , \x_mult_f[18][4] , \x_mult_f[18][3] ,
         \x_mult_f[18][2] , \x_mult_f[18][1] , \x_mult_f[18][0] ,
         \x_mult_f[17][15] , \x_mult_f[17][14] , \x_mult_f[17][13] ,
         \x_mult_f[17][12] , \x_mult_f[17][11] , \x_mult_f[17][10] ,
         \x_mult_f[17][9] , \x_mult_f[17][8] , \x_mult_f[17][7] ,
         \x_mult_f[17][6] , \x_mult_f[17][5] , \x_mult_f[17][4] ,
         \x_mult_f[17][3] , \x_mult_f[17][2] , \x_mult_f[17][1] ,
         \x_mult_f[17][0] , \x_mult_f[16][15] , \x_mult_f[16][14] ,
         \x_mult_f[16][13] , \x_mult_f[16][12] , \x_mult_f[16][11] ,
         \x_mult_f[16][10] , \x_mult_f[16][9] , \x_mult_f[16][8] ,
         \x_mult_f[16][7] , \x_mult_f[16][6] , \x_mult_f[16][5] ,
         \x_mult_f[16][4] , \x_mult_f[16][3] , \x_mult_f[16][2] ,
         \x_mult_f[16][1] , \x_mult_f[16][0] , \x_mult_f[15][15] ,
         \x_mult_f[15][14] , \x_mult_f[15][13] , \x_mult_f[15][12] ,
         \x_mult_f[15][11] , \x_mult_f[15][10] , \x_mult_f[15][9] ,
         \x_mult_f[15][8] , \x_mult_f[15][7] , \x_mult_f[15][6] ,
         \x_mult_f[15][5] , \x_mult_f[15][4] , \x_mult_f[15][3] ,
         \x_mult_f[15][2] , \x_mult_f[15][1] , \x_mult_f[15][0] ,
         \x_mult_f[14][15] , \x_mult_f[14][14] , \x_mult_f[14][13] ,
         \x_mult_f[14][12] , \x_mult_f[14][11] , \x_mult_f[14][10] ,
         \x_mult_f[14][9] , \x_mult_f[14][8] , \x_mult_f[14][7] ,
         \x_mult_f[14][6] , \x_mult_f[14][5] , \x_mult_f[14][4] ,
         \x_mult_f[14][3] , \x_mult_f[14][2] , \x_mult_f[14][1] ,
         \x_mult_f[14][0] , \x_mult_f[13][15] , \x_mult_f[13][14] ,
         \x_mult_f[13][13] , \x_mult_f[13][12] , \x_mult_f[13][11] ,
         \x_mult_f[13][10] , \x_mult_f[13][9] , \x_mult_f[13][8] ,
         \x_mult_f[13][7] , \x_mult_f[13][6] , \x_mult_f[13][5] ,
         \x_mult_f[13][4] , \x_mult_f[13][3] , \x_mult_f[13][2] ,
         \x_mult_f[13][1] , \x_mult_f[13][0] , \x_mult_f[12][15] ,
         \x_mult_f[12][14] , \x_mult_f[12][13] , \x_mult_f[12][12] ,
         \x_mult_f[12][11] , \x_mult_f[12][10] , \x_mult_f[12][9] ,
         \x_mult_f[12][8] , \x_mult_f[12][7] , \x_mult_f[12][6] ,
         \x_mult_f[12][5] , \x_mult_f[12][4] , \x_mult_f[12][3] ,
         \x_mult_f[12][2] , \x_mult_f[12][1] , \x_mult_f[12][0] ,
         \x_mult_f[11][15] , \x_mult_f[11][14] , \x_mult_f[11][13] ,
         \x_mult_f[11][12] , \x_mult_f[11][11] , \x_mult_f[11][10] ,
         \x_mult_f[11][9] , \x_mult_f[11][8] , \x_mult_f[11][7] ,
         \x_mult_f[11][6] , \x_mult_f[11][5] , \x_mult_f[11][4] ,
         \x_mult_f[11][3] , \x_mult_f[11][2] , \x_mult_f[11][1] ,
         \x_mult_f[11][0] , \x_mult_f[10][15] , \x_mult_f[10][14] ,
         \x_mult_f[10][13] , \x_mult_f[10][12] , \x_mult_f[10][11] ,
         \x_mult_f[10][10] , \x_mult_f[10][9] , \x_mult_f[10][8] ,
         \x_mult_f[10][7] , \x_mult_f[10][6] , \x_mult_f[10][5] ,
         \x_mult_f[10][4] , \x_mult_f[10][3] , \x_mult_f[10][2] ,
         \x_mult_f[10][1] , \x_mult_f[10][0] , \x_mult_f[9][15] ,
         \x_mult_f[9][14] , \x_mult_f[9][13] , \x_mult_f[9][12] ,
         \x_mult_f[9][11] , \x_mult_f[9][10] , \x_mult_f[9][9] ,
         \x_mult_f[9][8] , \x_mult_f[9][7] , \x_mult_f[9][6] ,
         \x_mult_f[9][5] , \x_mult_f[9][4] , \x_mult_f[9][3] ,
         \x_mult_f[9][2] , \x_mult_f[9][1] , \x_mult_f[9][0] ,
         \x_mult_f[8][15] , \x_mult_f[8][14] , \x_mult_f[8][13] ,
         \x_mult_f[8][12] , \x_mult_f[8][11] , \x_mult_f[8][10] ,
         \x_mult_f[8][9] , \x_mult_f[8][8] , \x_mult_f[8][7] ,
         \x_mult_f[8][6] , \x_mult_f[8][5] , \x_mult_f[8][4] ,
         \x_mult_f[8][3] , \x_mult_f[8][2] , \x_mult_f[8][1] ,
         \x_mult_f[8][0] , \x_mult_f[7][15] , \x_mult_f[7][14] ,
         \x_mult_f[7][13] , \x_mult_f[7][12] , \x_mult_f[7][11] ,
         \x_mult_f[7][10] , \x_mult_f[7][9] , \x_mult_f[7][8] ,
         \x_mult_f[7][7] , \x_mult_f[7][6] , \x_mult_f[7][5] ,
         \x_mult_f[7][4] , \x_mult_f[7][3] , \x_mult_f[7][2] ,
         \x_mult_f[7][1] , \x_mult_f[7][0] , \x_mult_f[6][15] ,
         \x_mult_f[6][14] , \x_mult_f[6][13] , \x_mult_f[6][12] ,
         \x_mult_f[6][11] , \x_mult_f[6][10] , \x_mult_f[6][9] ,
         \x_mult_f[6][8] , \x_mult_f[6][7] , \x_mult_f[6][6] ,
         \x_mult_f[6][5] , \x_mult_f[6][4] , \x_mult_f[6][3] ,
         \x_mult_f[6][2] , \x_mult_f[6][1] , \x_mult_f[6][0] ,
         \x_mult_f[5][15] , \x_mult_f[5][14] , \x_mult_f[5][13] ,
         \x_mult_f[5][12] , \x_mult_f[5][11] , \x_mult_f[5][10] ,
         \x_mult_f[5][9] , \x_mult_f[5][8] , \x_mult_f[5][7] ,
         \x_mult_f[5][6] , \x_mult_f[5][5] , \x_mult_f[5][4] ,
         \x_mult_f[5][3] , \x_mult_f[5][2] , \x_mult_f[5][1] ,
         \x_mult_f[5][0] , \x_mult_f[4][15] , \x_mult_f[4][14] ,
         \x_mult_f[4][13] , \x_mult_f[4][12] , \x_mult_f[4][11] ,
         \x_mult_f[4][10] , \x_mult_f[4][9] , \x_mult_f[4][8] ,
         \x_mult_f[4][7] , \x_mult_f[4][6] , \x_mult_f[4][5] ,
         \x_mult_f[4][4] , \x_mult_f[4][3] , \x_mult_f[4][2] ,
         \x_mult_f[4][1] , \x_mult_f[4][0] , \x_mult_f[3][15] ,
         \x_mult_f[3][14] , \x_mult_f[3][13] , \x_mult_f[3][12] ,
         \x_mult_f[3][11] , \x_mult_f[3][10] , \x_mult_f[3][9] ,
         \x_mult_f[3][8] , \x_mult_f[3][7] , \x_mult_f[3][6] ,
         \x_mult_f[3][5] , \x_mult_f[3][4] , \x_mult_f[3][3] ,
         \x_mult_f[3][2] , \x_mult_f[3][1] , \x_mult_f[3][0] ,
         \x_mult_f[2][15] , \x_mult_f[2][14] , \x_mult_f[2][13] ,
         \x_mult_f[2][12] , \x_mult_f[2][11] , \x_mult_f[2][10] ,
         \x_mult_f[2][9] , \x_mult_f[2][8] , \x_mult_f[2][7] ,
         \x_mult_f[2][6] , \x_mult_f[2][5] , \x_mult_f[2][4] ,
         \x_mult_f[2][3] , \x_mult_f[2][2] , \x_mult_f[2][1] ,
         \x_mult_f[2][0] , \x_mult_f[1][15] , \x_mult_f[1][14] ,
         \x_mult_f[1][13] , \x_mult_f[1][12] , \x_mult_f[1][11] ,
         \x_mult_f[1][10] , \x_mult_f[1][9] , \x_mult_f[1][8] ,
         \x_mult_f[1][7] , \x_mult_f[1][6] , \x_mult_f[1][5] ,
         \x_mult_f[1][4] , \x_mult_f[1][3] , \x_mult_f[1][2] ,
         \x_mult_f[1][1] , \x_mult_f[1][0] , \x_mult_f[0][15] ,
         \x_mult_f[0][14] , \x_mult_f[0][13] , \x_mult_f[0][12] ,
         \x_mult_f[0][11] , \x_mult_f[0][10] , \x_mult_f[0][9] ,
         \x_mult_f[0][8] , \x_mult_f[0][7] , \x_mult_f[0][6] ,
         \x_mult_f[0][5] , \x_mult_f[0][4] , \x_mult_f[0][3] ,
         \x_mult_f[0][2] , \x_mult_f[0][1] , \x_mult_f[0][0] ,
         \adder_stage1[15][20] , \adder_stage1[15][15] ,
         \adder_stage1[15][14] , \adder_stage1[15][13] ,
         \adder_stage1[15][12] , \adder_stage1[15][11] ,
         \adder_stage1[15][10] , \adder_stage1[15][9] , \adder_stage1[15][8] ,
         \adder_stage1[15][7] , \adder_stage1[15][6] , \adder_stage1[15][5] ,
         \adder_stage1[15][4] , \adder_stage1[15][3] , \adder_stage1[15][2] ,
         \adder_stage1[15][1] , \adder_stage1[15][0] , \adder_stage1[14][20] ,
         \adder_stage1[14][15] , \adder_stage1[14][14] ,
         \adder_stage1[14][13] , \adder_stage1[14][12] ,
         \adder_stage1[14][11] , \adder_stage1[14][10] , \adder_stage1[14][9] ,
         \adder_stage1[14][8] , \adder_stage1[14][7] , \adder_stage1[14][6] ,
         \adder_stage1[14][5] , \adder_stage1[14][4] , \adder_stage1[14][3] ,
         \adder_stage1[14][2] , \adder_stage1[14][1] , \adder_stage1[14][0] ,
         \adder_stage1[13][20] , \adder_stage1[13][15] ,
         \adder_stage1[13][14] , \adder_stage1[13][13] ,
         \adder_stage1[13][12] , \adder_stage1[13][11] ,
         \adder_stage1[13][10] , \adder_stage1[13][9] , \adder_stage1[13][8] ,
         \adder_stage1[13][7] , \adder_stage1[13][6] , \adder_stage1[13][5] ,
         \adder_stage1[13][4] , \adder_stage1[13][3] , \adder_stage1[13][2] ,
         \adder_stage1[13][1] , \adder_stage1[13][0] , \adder_stage1[12][20] ,
         \adder_stage1[12][15] , \adder_stage1[12][14] ,
         \adder_stage1[12][13] , \adder_stage1[12][12] ,
         \adder_stage1[12][11] , \adder_stage1[12][10] , \adder_stage1[12][9] ,
         \adder_stage1[12][8] , \adder_stage1[12][7] , \adder_stage1[12][6] ,
         \adder_stage1[12][5] , \adder_stage1[12][4] , \adder_stage1[12][3] ,
         \adder_stage1[12][2] , \adder_stage1[12][1] , \adder_stage1[12][0] ,
         \adder_stage1[11][20] , \adder_stage1[11][15] ,
         \adder_stage1[11][14] , \adder_stage1[11][13] ,
         \adder_stage1[11][12] , \adder_stage1[11][11] ,
         \adder_stage1[11][10] , \adder_stage1[11][9] , \adder_stage1[11][8] ,
         \adder_stage1[11][7] , \adder_stage1[11][6] , \adder_stage1[11][5] ,
         \adder_stage1[11][4] , \adder_stage1[11][3] , \adder_stage1[11][2] ,
         \adder_stage1[11][1] , \adder_stage1[11][0] , \adder_stage1[10][20] ,
         \adder_stage1[10][15] , \adder_stage1[10][14] ,
         \adder_stage1[10][13] , \adder_stage1[10][12] ,
         \adder_stage1[10][11] , \adder_stage1[10][10] , \adder_stage1[10][9] ,
         \adder_stage1[10][8] , \adder_stage1[10][7] , \adder_stage1[10][6] ,
         \adder_stage1[10][5] , \adder_stage1[10][4] , \adder_stage1[10][3] ,
         \adder_stage1[10][2] , \adder_stage1[10][1] , \adder_stage1[10][0] ,
         \adder_stage1[9][20] , \adder_stage1[9][15] , \adder_stage1[9][14] ,
         \adder_stage1[9][13] , \adder_stage1[9][12] , \adder_stage1[9][11] ,
         \adder_stage1[9][10] , \adder_stage1[9][9] , \adder_stage1[9][8] ,
         \adder_stage1[9][7] , \adder_stage1[9][6] , \adder_stage1[9][5] ,
         \adder_stage1[9][4] , \adder_stage1[9][3] , \adder_stage1[9][2] ,
         \adder_stage1[9][1] , \adder_stage1[9][0] , \adder_stage1[8][20] ,
         \adder_stage1[8][15] , \adder_stage1[8][14] , \adder_stage1[8][13] ,
         \adder_stage1[8][12] , \adder_stage1[8][11] , \adder_stage1[8][10] ,
         \adder_stage1[8][9] , \adder_stage1[8][8] , \adder_stage1[8][7] ,
         \adder_stage1[8][6] , \adder_stage1[8][5] , \adder_stage1[8][4] ,
         \adder_stage1[8][3] , \adder_stage1[8][2] , \adder_stage1[8][1] ,
         \adder_stage1[8][0] , \adder_stage1[7][20] , \adder_stage1[7][15] ,
         \adder_stage1[7][14] , \adder_stage1[7][13] , \adder_stage1[7][12] ,
         \adder_stage1[7][11] , \adder_stage1[7][10] , \adder_stage1[7][9] ,
         \adder_stage1[7][8] , \adder_stage1[7][7] , \adder_stage1[7][6] ,
         \adder_stage1[7][5] , \adder_stage1[7][4] , \adder_stage1[7][3] ,
         \adder_stage1[7][2] , \adder_stage1[7][1] , \adder_stage1[7][0] ,
         \adder_stage1[6][20] , \adder_stage1[6][15] , \adder_stage1[6][14] ,
         \adder_stage1[6][13] , \adder_stage1[6][12] , \adder_stage1[6][11] ,
         \adder_stage1[6][10] , \adder_stage1[6][9] , \adder_stage1[6][8] ,
         \adder_stage1[6][7] , \adder_stage1[6][6] , \adder_stage1[6][5] ,
         \adder_stage1[6][4] , \adder_stage1[6][3] , \adder_stage1[6][2] ,
         \adder_stage1[6][1] , \adder_stage1[6][0] , \adder_stage1[5][20] ,
         \adder_stage1[5][15] , \adder_stage1[5][14] , \adder_stage1[5][13] ,
         \adder_stage1[5][12] , \adder_stage1[5][11] , \adder_stage1[5][10] ,
         \adder_stage1[5][9] , \adder_stage1[5][8] , \adder_stage1[5][7] ,
         \adder_stage1[5][6] , \adder_stage1[5][5] , \adder_stage1[5][4] ,
         \adder_stage1[5][3] , \adder_stage1[5][2] , \adder_stage1[5][1] ,
         \adder_stage1[5][0] , \adder_stage1[4][20] , \adder_stage1[4][15] ,
         \adder_stage1[4][14] , \adder_stage1[4][13] , \adder_stage1[4][12] ,
         \adder_stage1[4][11] , \adder_stage1[4][10] , \adder_stage1[4][9] ,
         \adder_stage1[4][8] , \adder_stage1[4][7] , \adder_stage1[4][6] ,
         \adder_stage1[4][5] , \adder_stage1[4][4] , \adder_stage1[4][3] ,
         \adder_stage1[4][2] , \adder_stage1[4][1] , \adder_stage1[4][0] ,
         \adder_stage1[3][20] , \adder_stage1[3][15] , \adder_stage1[3][14] ,
         \adder_stage1[3][13] , \adder_stage1[3][12] , \adder_stage1[3][11] ,
         \adder_stage1[3][10] , \adder_stage1[3][9] , \adder_stage1[3][8] ,
         \adder_stage1[3][7] , \adder_stage1[3][6] , \adder_stage1[3][5] ,
         \adder_stage1[3][4] , \adder_stage1[3][3] , \adder_stage1[3][2] ,
         \adder_stage1[3][1] , \adder_stage1[3][0] , \adder_stage1[2][20] ,
         \adder_stage1[2][15] , \adder_stage1[2][14] , \adder_stage1[2][13] ,
         \adder_stage1[2][12] , \adder_stage1[2][11] , \adder_stage1[2][10] ,
         \adder_stage1[2][9] , \adder_stage1[2][8] , \adder_stage1[2][7] ,
         \adder_stage1[2][6] , \adder_stage1[2][5] , \adder_stage1[2][4] ,
         \adder_stage1[2][3] , \adder_stage1[2][2] , \adder_stage1[2][1] ,
         \adder_stage1[2][0] , \adder_stage1[1][20] , \adder_stage1[1][15] ,
         \adder_stage1[1][14] , \adder_stage1[1][13] , \adder_stage1[1][12] ,
         \adder_stage1[1][11] , \adder_stage1[1][10] , \adder_stage1[1][9] ,
         \adder_stage1[1][8] , \adder_stage1[1][7] , \adder_stage1[1][6] ,
         \adder_stage1[1][5] , \adder_stage1[1][4] , \adder_stage1[1][3] ,
         \adder_stage1[1][2] , \adder_stage1[1][1] , \adder_stage1[1][0] ,
         \adder_stage1[0][20] , \adder_stage1[0][15] , \adder_stage1[0][14] ,
         \adder_stage1[0][13] , \adder_stage1[0][12] , \adder_stage1[0][11] ,
         \adder_stage1[0][10] , \adder_stage1[0][9] , \adder_stage1[0][8] ,
         \adder_stage1[0][7] , \adder_stage1[0][6] , \adder_stage1[0][5] ,
         \adder_stage1[0][4] , \adder_stage1[0][3] , \adder_stage1[0][2] ,
         \adder_stage1[0][1] , \adder_stage1[0][0] , \adder_stage2[7][20] ,
         \adder_stage2[7][19] , \adder_stage2[7][18] , \adder_stage2[7][17] ,
         \adder_stage2[7][16] , \adder_stage2[7][15] , \adder_stage2[7][14] ,
         \adder_stage2[7][13] , \adder_stage2[7][12] , \adder_stage2[7][11] ,
         \adder_stage2[7][10] , \adder_stage2[7][9] , \adder_stage2[7][8] ,
         \adder_stage2[7][7] , \adder_stage2[7][6] , \adder_stage2[7][5] ,
         \adder_stage2[7][4] , \adder_stage2[7][3] , \adder_stage2[7][2] ,
         \adder_stage2[7][1] , \adder_stage2[7][0] , \adder_stage2[6][20] ,
         \adder_stage2[6][19] , \adder_stage2[6][18] , \adder_stage2[6][17] ,
         \adder_stage2[6][16] , \adder_stage2[6][15] , \adder_stage2[6][14] ,
         \adder_stage2[6][13] , \adder_stage2[6][12] , \adder_stage2[6][11] ,
         \adder_stage2[6][10] , \adder_stage2[6][9] , \adder_stage2[6][8] ,
         \adder_stage2[6][7] , \adder_stage2[6][6] , \adder_stage2[6][5] ,
         \adder_stage2[6][4] , \adder_stage2[6][3] , \adder_stage2[6][2] ,
         \adder_stage2[6][1] , \adder_stage2[6][0] , \adder_stage2[5][20] ,
         \adder_stage2[5][19] , \adder_stage2[5][18] , \adder_stage2[5][17] ,
         \adder_stage2[5][16] , \adder_stage2[5][15] , \adder_stage2[5][14] ,
         \adder_stage2[5][13] , \adder_stage2[5][12] , \adder_stage2[5][11] ,
         \adder_stage2[5][10] , \adder_stage2[5][9] , \adder_stage2[5][8] ,
         \adder_stage2[5][7] , \adder_stage2[5][6] , \adder_stage2[5][5] ,
         \adder_stage2[5][4] , \adder_stage2[5][3] , \adder_stage2[5][2] ,
         \adder_stage2[5][1] , \adder_stage2[5][0] , \adder_stage2[4][20] ,
         \adder_stage2[4][19] , \adder_stage2[4][18] , \adder_stage2[4][17] ,
         \adder_stage2[4][16] , \adder_stage2[4][15] , \adder_stage2[4][14] ,
         \adder_stage2[4][13] , \adder_stage2[4][12] , \adder_stage2[4][11] ,
         \adder_stage2[4][10] , \adder_stage2[4][9] , \adder_stage2[4][8] ,
         \adder_stage2[4][7] , \adder_stage2[4][6] , \adder_stage2[4][5] ,
         \adder_stage2[4][4] , \adder_stage2[4][3] , \adder_stage2[4][2] ,
         \adder_stage2[4][1] , \adder_stage2[4][0] , \adder_stage2[3][20] ,
         \adder_stage2[3][19] , \adder_stage2[3][18] , \adder_stage2[3][17] ,
         \adder_stage2[3][16] , \adder_stage2[3][15] , \adder_stage2[3][14] ,
         \adder_stage2[3][13] , \adder_stage2[3][12] , \adder_stage2[3][11] ,
         \adder_stage2[3][10] , \adder_stage2[3][9] , \adder_stage2[3][8] ,
         \adder_stage2[3][7] , \adder_stage2[3][6] , \adder_stage2[3][5] ,
         \adder_stage2[3][4] , \adder_stage2[3][3] , \adder_stage2[3][2] ,
         \adder_stage2[3][1] , \adder_stage2[3][0] , \adder_stage2[2][20] ,
         \adder_stage2[2][19] , \adder_stage2[2][18] , \adder_stage2[2][17] ,
         \adder_stage2[2][16] , \adder_stage2[2][15] , \adder_stage2[2][14] ,
         \adder_stage2[2][13] , \adder_stage2[2][12] , \adder_stage2[2][11] ,
         \adder_stage2[2][10] , \adder_stage2[2][9] , \adder_stage2[2][8] ,
         \adder_stage2[2][7] , \adder_stage2[2][6] , \adder_stage2[2][5] ,
         \adder_stage2[2][4] , \adder_stage2[2][3] , \adder_stage2[2][2] ,
         \adder_stage2[2][1] , \adder_stage2[2][0] , \adder_stage2[1][20] ,
         \adder_stage2[1][19] , \adder_stage2[1][18] , \adder_stage2[1][17] ,
         \adder_stage2[1][16] , \adder_stage2[1][15] , \adder_stage2[1][14] ,
         \adder_stage2[1][13] , \adder_stage2[1][12] , \adder_stage2[1][11] ,
         \adder_stage2[1][10] , \adder_stage2[1][9] , \adder_stage2[1][8] ,
         \adder_stage2[1][7] , \adder_stage2[1][6] , \adder_stage2[1][5] ,
         \adder_stage2[1][4] , \adder_stage2[1][3] , \adder_stage2[1][2] ,
         \adder_stage2[1][1] , \adder_stage2[1][0] , \adder_stage2[0][20] ,
         \adder_stage2[0][19] , \adder_stage2[0][18] , \adder_stage2[0][17] ,
         \adder_stage2[0][16] , \adder_stage2[0][15] , \adder_stage2[0][14] ,
         \adder_stage2[0][13] , \adder_stage2[0][12] , \adder_stage2[0][11] ,
         \adder_stage2[0][10] , \adder_stage2[0][9] , \adder_stage2[0][8] ,
         \adder_stage2[0][7] , \adder_stage2[0][6] , \adder_stage2[0][5] ,
         \adder_stage2[0][4] , \adder_stage2[0][3] , \adder_stage2[0][2] ,
         \adder_stage2[0][1] , \adder_stage2[0][0] , \adder_stage3[3][20] ,
         \adder_stage3[3][19] , \adder_stage3[3][18] , \adder_stage3[3][17] ,
         \adder_stage3[3][16] , \adder_stage3[3][15] , \adder_stage3[3][14] ,
         \adder_stage3[3][13] , \adder_stage3[3][12] , \adder_stage3[3][11] ,
         \adder_stage3[3][10] , \adder_stage3[3][9] , \adder_stage3[3][8] ,
         \adder_stage3[3][7] , \adder_stage3[3][6] , \adder_stage3[3][5] ,
         \adder_stage3[3][4] , \adder_stage3[3][3] , \adder_stage3[3][2] ,
         \adder_stage3[3][1] , \adder_stage3[3][0] , \adder_stage3[2][20] ,
         \adder_stage3[2][19] , \adder_stage3[2][18] , \adder_stage3[2][17] ,
         \adder_stage3[2][16] , \adder_stage3[2][15] , \adder_stage3[2][14] ,
         \adder_stage3[2][13] , \adder_stage3[2][12] , \adder_stage3[2][11] ,
         \adder_stage3[2][10] , \adder_stage3[2][9] , \adder_stage3[2][8] ,
         \adder_stage3[2][7] , \adder_stage3[2][6] , \adder_stage3[2][5] ,
         \adder_stage3[2][4] , \adder_stage3[2][3] , \adder_stage3[2][2] ,
         \adder_stage3[2][1] , \adder_stage3[2][0] , \adder_stage3[1][20] ,
         \adder_stage3[1][19] , \adder_stage3[1][18] , \adder_stage3[1][17] ,
         \adder_stage3[1][16] , \adder_stage3[1][15] , \adder_stage3[1][14] ,
         \adder_stage3[1][13] , \adder_stage3[1][12] , \adder_stage3[1][11] ,
         \adder_stage3[1][10] , \adder_stage3[1][9] , \adder_stage3[1][8] ,
         \adder_stage3[1][7] , \adder_stage3[1][6] , \adder_stage3[1][5] ,
         \adder_stage3[1][4] , \adder_stage3[1][3] , \adder_stage3[1][2] ,
         \adder_stage3[1][1] , \adder_stage3[1][0] , \adder_stage3[0][20] ,
         \adder_stage3[0][19] , \adder_stage3[0][18] , \adder_stage3[0][17] ,
         \adder_stage3[0][16] , \adder_stage3[0][15] , \adder_stage3[0][14] ,
         \adder_stage3[0][13] , \adder_stage3[0][12] , \adder_stage3[0][11] ,
         \adder_stage3[0][10] , \adder_stage3[0][9] , \adder_stage3[0][8] ,
         \adder_stage3[0][7] , \adder_stage3[0][6] , \adder_stage3[0][5] ,
         \adder_stage3[0][4] , \adder_stage3[0][3] , \adder_stage3[0][2] ,
         \adder_stage3[0][1] , \adder_stage3[0][0] , \adder_stage4[1][20] ,
         \adder_stage4[1][19] , \adder_stage4[1][18] , \adder_stage4[1][17] ,
         \adder_stage4[1][16] , \adder_stage4[1][15] , \adder_stage4[1][14] ,
         \adder_stage4[1][13] , \adder_stage4[1][12] , \adder_stage4[1][11] ,
         \adder_stage4[1][10] , \adder_stage4[1][9] , \adder_stage4[1][8] ,
         \adder_stage4[1][7] , \adder_stage4[1][6] , \adder_stage4[1][5] ,
         \adder_stage4[1][4] , \adder_stage4[1][3] , \adder_stage4[1][2] ,
         \adder_stage4[1][1] , \adder_stage4[1][0] , \adder_stage4[0][20] ,
         \adder_stage4[0][19] , \adder_stage4[0][18] , \adder_stage4[0][17] ,
         \adder_stage4[0][16] , \adder_stage4[0][15] , \adder_stage4[0][14] ,
         \adder_stage4[0][13] , \adder_stage4[0][12] , \adder_stage4[0][11] ,
         \adder_stage4[0][10] , \adder_stage4[0][9] , \adder_stage4[0][8] ,
         \adder_stage4[0][7] , \adder_stage4[0][6] , \adder_stage4[0][5] ,
         \adder_stage4[0][4] , \adder_stage4[0][3] , \adder_stage4[0][2] ,
         \adder_stage4[0][1] , \adder_stage4[0][0] , \ctrl_inst/s_ready_fsm ,
         n1909, n1910, n1911, n1912, n1930, n1931, n1932, n1933, n1951, n1952,
         n1953, n1954, n1972, n1973, n1974, n1975, n1993, n1994, n1995, n1996,
         n2014, n2015, n2016, n2017, n2035, n2036, n2037, n2038, n2056, n2057,
         n2058, n2059, n3118, n3119, n3120, n3121, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3383, n3385, n3386, n3387, n3388,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8322, n8323, n8324, n8325, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421;
  wire   [4:0] fmem_addr;
  wire   [6:0] \ctrl_inst/xmem_tracker ;
  wire   [3:0] \ctrl_inst/pline_cntr ;
  wire   [2:0] \ctrl_inst/state ;

  DFF_X1 \ctrl_inst/s_ready_fsm_reg  ( .D(n3385), .CK(clk), .Q(
        \ctrl_inst/s_ready_fsm ), .QN(n8812) );
  DFF_X1 \xmem_inst/mem_reg[31][7]  ( .D(n3377), .CK(clk), .Q(
        \xmem_data[31][7] ) );
  DFF_X1 \xmem_inst/mem_reg[31][6]  ( .D(n3376), .CK(clk), .Q(
        \xmem_data[31][6] ) );
  DFF_X1 \xmem_inst/mem_reg[31][5]  ( .D(n3375), .CK(clk), .Q(
        \xmem_data[31][5] ) );
  DFF_X1 \xmem_inst/mem_reg[31][4]  ( .D(n3374), .CK(clk), .Q(
        \xmem_data[31][4] ) );
  DFF_X1 \xmem_inst/mem_reg[31][3]  ( .D(n3373), .CK(clk), .Q(
        \xmem_data[31][3] ) );
  DFF_X1 \xmem_inst/mem_reg[31][2]  ( .D(n3372), .CK(clk), .Q(
        \xmem_data[31][2] ) );
  DFF_X1 \xmem_inst/mem_reg[31][1]  ( .D(n3371), .CK(clk), .Q(
        \xmem_data[31][1] ) );
  DFF_X1 \xmem_inst/mem_reg[31][0]  ( .D(n3370), .CK(clk), .Q(
        \xmem_data[31][0] ) );
  DFF_X1 \xmem_inst/mem_reg[30][7]  ( .D(n10417), .CK(clk), .Q(
        \xmem_data[30][7] ) );
  DFF_X1 \xmem_inst/mem_reg[30][6]  ( .D(n10416), .CK(clk), .Q(
        \xmem_data[30][6] ) );
  DFF_X1 \xmem_inst/mem_reg[30][5]  ( .D(n10415), .CK(clk), .Q(
        \xmem_data[30][5] ) );
  DFF_X1 \xmem_inst/mem_reg[30][4]  ( .D(n10414), .CK(clk), .Q(
        \xmem_data[30][4] ) );
  DFF_X1 \xmem_inst/mem_reg[30][3]  ( .D(n10413), .CK(clk), .Q(
        \xmem_data[30][3] ) );
  DFF_X1 \xmem_inst/mem_reg[30][2]  ( .D(n10412), .CK(clk), .Q(
        \xmem_data[30][2] ) );
  DFF_X1 \xmem_inst/mem_reg[30][1]  ( .D(n10411), .CK(clk), .Q(
        \xmem_data[30][1] ) );
  DFF_X1 \xmem_inst/mem_reg[30][0]  ( .D(n10410), .CK(clk), .Q(
        \xmem_data[30][0] ) );
  DFF_X1 \xmem_inst/mem_reg[29][7]  ( .D(n10409), .CK(clk), .Q(
        \xmem_data[29][7] ) );
  DFF_X1 \xmem_inst/mem_reg[29][6]  ( .D(n10408), .CK(clk), .Q(
        \xmem_data[29][6] ) );
  DFF_X1 \xmem_inst/mem_reg[29][5]  ( .D(n10407), .CK(clk), .Q(
        \xmem_data[29][5] ) );
  DFF_X1 \xmem_inst/mem_reg[29][4]  ( .D(n10406), .CK(clk), .Q(
        \xmem_data[29][4] ) );
  DFF_X1 \xmem_inst/mem_reg[29][3]  ( .D(n10405), .CK(clk), .Q(
        \xmem_data[29][3] ) );
  DFF_X1 \xmem_inst/mem_reg[29][2]  ( .D(n10404), .CK(clk), .Q(
        \xmem_data[29][2] ) );
  DFF_X1 \xmem_inst/mem_reg[29][1]  ( .D(n10403), .CK(clk), .Q(
        \xmem_data[29][1] ) );
  DFF_X1 \xmem_inst/mem_reg[29][0]  ( .D(n10402), .CK(clk), .Q(
        \xmem_data[29][0] ) );
  DFF_X1 \xmem_inst/mem_reg[28][7]  ( .D(n10401), .CK(clk), .Q(
        \xmem_data[28][7] ) );
  DFF_X1 \xmem_inst/mem_reg[28][6]  ( .D(n10400), .CK(clk), .Q(
        \xmem_data[28][6] ) );
  DFF_X1 \xmem_inst/mem_reg[28][5]  ( .D(n10399), .CK(clk), .Q(
        \xmem_data[28][5] ) );
  DFF_X1 \xmem_inst/mem_reg[28][4]  ( .D(n10398), .CK(clk), .Q(
        \xmem_data[28][4] ) );
  DFF_X1 \xmem_inst/mem_reg[28][3]  ( .D(n10397), .CK(clk), .Q(
        \xmem_data[28][3] ) );
  DFF_X1 \xmem_inst/mem_reg[28][2]  ( .D(n10396), .CK(clk), .Q(
        \xmem_data[28][2] ) );
  DFF_X1 \xmem_inst/mem_reg[28][1]  ( .D(n10395), .CK(clk), .Q(
        \xmem_data[28][1] ) );
  DFF_X1 \xmem_inst/mem_reg[28][0]  ( .D(n10394), .CK(clk), .Q(
        \xmem_data[28][0] ) );
  DFF_X1 \xmem_inst/mem_reg[27][7]  ( .D(n10393), .CK(clk), .Q(
        \xmem_data[27][7] ) );
  DFF_X1 \xmem_inst/mem_reg[27][6]  ( .D(n10392), .CK(clk), .Q(
        \xmem_data[27][6] ) );
  DFF_X1 \xmem_inst/mem_reg[27][5]  ( .D(n10391), .CK(clk), .Q(
        \xmem_data[27][5] ) );
  DFF_X1 \xmem_inst/mem_reg[27][4]  ( .D(n10390), .CK(clk), .Q(
        \xmem_data[27][4] ) );
  DFF_X1 \xmem_inst/mem_reg[27][3]  ( .D(n10389), .CK(clk), .Q(
        \xmem_data[27][3] ) );
  DFF_X1 \xmem_inst/mem_reg[27][2]  ( .D(n10388), .CK(clk), .Q(
        \xmem_data[27][2] ) );
  DFF_X1 \xmem_inst/mem_reg[27][1]  ( .D(n10387), .CK(clk), .Q(
        \xmem_data[27][1] ) );
  DFF_X1 \xmem_inst/mem_reg[27][0]  ( .D(n10386), .CK(clk), .Q(
        \xmem_data[27][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][7]  ( .D(n10385), .CK(clk), .Q(
        \xmem_data[26][7] ) );
  DFF_X1 \xmem_inst/mem_reg[26][6]  ( .D(n10384), .CK(clk), .Q(
        \xmem_data[26][6] ) );
  DFF_X1 \xmem_inst/mem_reg[26][5]  ( .D(n10383), .CK(clk), .Q(
        \xmem_data[26][5] ) );
  DFF_X1 \xmem_inst/mem_reg[26][4]  ( .D(n10382), .CK(clk), .Q(
        \xmem_data[26][4] ) );
  DFF_X1 \xmem_inst/mem_reg[26][3]  ( .D(n10381), .CK(clk), .Q(
        \xmem_data[26][3] ) );
  DFF_X1 \xmem_inst/mem_reg[26][2]  ( .D(n10380), .CK(clk), .Q(
        \xmem_data[26][2] ) );
  DFF_X1 \xmem_inst/mem_reg[26][1]  ( .D(n10379), .CK(clk), .Q(
        \xmem_data[26][1] ) );
  DFF_X1 \xmem_inst/mem_reg[26][0]  ( .D(n10378), .CK(clk), .Q(
        \xmem_data[26][0] ) );
  DFF_X1 \xmem_inst/mem_reg[25][7]  ( .D(n10377), .CK(clk), .Q(
        \xmem_data[25][7] ) );
  DFF_X1 \xmem_inst/mem_reg[25][6]  ( .D(n10376), .CK(clk), .Q(
        \xmem_data[25][6] ) );
  DFF_X1 \xmem_inst/mem_reg[25][5]  ( .D(n10375), .CK(clk), .Q(
        \xmem_data[25][5] ) );
  DFF_X1 \xmem_inst/mem_reg[24][5]  ( .D(n10374), .CK(clk), .Q(
        \xmem_data[24][5] ) );
  DFF_X1 \xmem_inst/mem_reg[23][5]  ( .D(n10373), .CK(clk), .Q(
        \xmem_data[23][5] ) );
  DFF_X1 \xmem_inst/mem_reg[22][5]  ( .D(n10372), .CK(clk), .Q(
        \xmem_data[22][5] ) );
  DFF_X1 \xmem_inst/mem_reg[21][5]  ( .D(n10371), .CK(clk), .Q(
        \xmem_data[21][5] ) );
  DFF_X1 \xmem_inst/mem_reg[20][5]  ( .D(n10370), .CK(clk), .Q(
        \xmem_data[20][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n10369), .CK(clk), .Q(
        \xmem_data[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n10368), .CK(clk), .Q(
        \xmem_data[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n10367), .CK(clk), .Q(
        \xmem_data[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n10366), .CK(clk), .Q(
        \xmem_data[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n10365), .CK(clk), .Q(
        \xmem_data[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n10364), .CK(clk), .Q(
        \xmem_data[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n10363), .CK(clk), .Q(
        \xmem_data[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n10362), .CK(clk), .Q(
        \xmem_data[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n10361), .CK(clk), .Q(
        \xmem_data[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n10360), .CK(clk), .Q(
        \xmem_data[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n10359), .CK(clk), .Q(
        \xmem_data[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n10358), .CK(clk), .Q(
        \xmem_data[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n10357), .CK(clk), .Q(
        \xmem_data[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n10356), .CK(clk), .Q(
        \xmem_data[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n10355), .CK(clk), .Q(
        \xmem_data[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n10354), .CK(clk), .Q(
        \xmem_data[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n10353), .CK(clk), .Q(
        \xmem_data[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n10352), .CK(clk), .Q(
        \xmem_data[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n10351), .CK(clk), .Q(
        \xmem_data[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n10350), .CK(clk), .Q(
        \xmem_data[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[25][4]  ( .D(n10349), .CK(clk), .Q(
        \xmem_data[25][4] ) );
  DFF_X1 \xmem_inst/mem_reg[24][4]  ( .D(n10348), .CK(clk), .Q(
        \xmem_data[24][4] ) );
  DFF_X1 \xmem_inst/mem_reg[23][4]  ( .D(n10347), .CK(clk), .Q(
        \xmem_data[23][4] ) );
  DFF_X1 \xmem_inst/mem_reg[22][4]  ( .D(n10346), .CK(clk), .Q(
        \xmem_data[22][4] ) );
  DFF_X1 \xmem_inst/mem_reg[21][4]  ( .D(n10345), .CK(clk), .Q(
        \xmem_data[21][4] ) );
  DFF_X1 \xmem_inst/mem_reg[20][4]  ( .D(n10344), .CK(clk), .Q(
        \xmem_data[20][4] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n10343), .CK(clk), .Q(
        \xmem_data[19][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n10342), .CK(clk), .Q(
        \xmem_data[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n10341), .CK(clk), .Q(
        \xmem_data[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n10340), .CK(clk), .Q(
        \xmem_data[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n10339), .CK(clk), .Q(
        \xmem_data[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n10338), .CK(clk), .Q(
        \xmem_data[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n10337), .CK(clk), .Q(
        \xmem_data[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n10336), .CK(clk), .Q(
        \xmem_data[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n10335), .CK(clk), .Q(
        \xmem_data[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n10334), .CK(clk), .Q(
        \xmem_data[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n10333), .CK(clk), .Q(
        \xmem_data[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n10332), .CK(clk), .Q(
        \xmem_data[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n10331), .CK(clk), .Q(
        \xmem_data[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n10330), .CK(clk), .Q(
        \xmem_data[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n10329), .CK(clk), .Q(
        \xmem_data[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n10328), .CK(clk), .Q(
        \xmem_data[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n10327), .CK(clk), .Q(
        \xmem_data[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n10326), .CK(clk), .Q(
        \xmem_data[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n10325), .CK(clk), .Q(
        \xmem_data[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n10324), .CK(clk), .Q(
        \xmem_data[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[25][3]  ( .D(n10323), .CK(clk), .Q(
        \xmem_data[25][3] ) );
  DFF_X1 \xmem_inst/mem_reg[24][3]  ( .D(n10322), .CK(clk), .Q(
        \xmem_data[24][3] ) );
  DFF_X1 \xmem_inst/mem_reg[23][3]  ( .D(n10321), .CK(clk), .Q(
        \xmem_data[23][3] ) );
  DFF_X1 \xmem_inst/mem_reg[22][3]  ( .D(n10320), .CK(clk), .Q(
        \xmem_data[22][3] ) );
  DFF_X1 \xmem_inst/mem_reg[21][3]  ( .D(n10319), .CK(clk), .Q(
        \xmem_data[21][3] ) );
  DFF_X1 \xmem_inst/mem_reg[20][3]  ( .D(n10318), .CK(clk), .Q(
        \xmem_data[20][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n10317), .CK(clk), .Q(
        \xmem_data[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n10316), .CK(clk), .Q(
        \xmem_data[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n10315), .CK(clk), .Q(
        \xmem_data[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n10314), .CK(clk), .Q(
        \xmem_data[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n10313), .CK(clk), .Q(
        \xmem_data[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n10312), .CK(clk), .Q(
        \xmem_data[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n10311), .CK(clk), .Q(
        \xmem_data[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n10310), .CK(clk), .Q(
        \xmem_data[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n10309), .CK(clk), .Q(
        \xmem_data[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n10308), .CK(clk), .Q(
        \xmem_data[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n10307), .CK(clk), .Q(
        \xmem_data[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n10306), .CK(clk), .Q(
        \xmem_data[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n10305), .CK(clk), .Q(
        \xmem_data[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n10304), .CK(clk), .Q(
        \xmem_data[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n10303), .CK(clk), .Q(
        \xmem_data[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n10302), .CK(clk), .Q(
        \xmem_data[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n10301), .CK(clk), .Q(
        \xmem_data[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n10300), .CK(clk), .Q(
        \xmem_data[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n10299), .CK(clk), .Q(
        \xmem_data[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n10298), .CK(clk), .Q(
        \xmem_data[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[25][2]  ( .D(n10297), .CK(clk), .Q(
        \xmem_data[25][2] ) );
  DFF_X1 \xmem_inst/mem_reg[24][2]  ( .D(n10296), .CK(clk), .Q(
        \xmem_data[24][2] ) );
  DFF_X1 \xmem_inst/mem_reg[23][2]  ( .D(n10295), .CK(clk), .Q(
        \xmem_data[23][2] ) );
  DFF_X1 \xmem_inst/mem_reg[22][2]  ( .D(n10294), .CK(clk), .Q(
        \xmem_data[22][2] ) );
  DFF_X1 \xmem_inst/mem_reg[21][2]  ( .D(n10293), .CK(clk), .Q(
        \xmem_data[21][2] ) );
  DFF_X1 \xmem_inst/mem_reg[20][2]  ( .D(n10292), .CK(clk), .Q(
        \xmem_data[20][2] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n10291), .CK(clk), .Q(
        \xmem_data[19][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n10290), .CK(clk), .Q(
        \xmem_data[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n10289), .CK(clk), .Q(
        \xmem_data[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n10288), .CK(clk), .Q(
        \xmem_data[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n10287), .CK(clk), .Q(
        \xmem_data[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n10286), .CK(clk), .Q(
        \xmem_data[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n10285), .CK(clk), .Q(
        \xmem_data[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n10284), .CK(clk), .Q(
        \xmem_data[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n10283), .CK(clk), .Q(
        \xmem_data[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n10282), .CK(clk), .Q(
        \xmem_data[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n10281), .CK(clk), .Q(
        \xmem_data[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n10280), .CK(clk), .Q(
        \xmem_data[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n10279), .CK(clk), .Q(
        \xmem_data[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n10278), .CK(clk), .Q(
        \xmem_data[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n10277), .CK(clk), .Q(
        \xmem_data[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n10276), .CK(clk), .Q(
        \xmem_data[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n10275), .CK(clk), .Q(
        \xmem_data[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n10274), .CK(clk), .Q(
        \xmem_data[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n10273), .CK(clk), .Q(
        \xmem_data[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n10272), .CK(clk), .Q(
        \xmem_data[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[25][1]  ( .D(n10271), .CK(clk), .Q(
        \xmem_data[25][1] ) );
  DFF_X1 \xmem_inst/mem_reg[24][1]  ( .D(n10270), .CK(clk), .Q(
        \xmem_data[24][1] ) );
  DFF_X1 \xmem_inst/mem_reg[23][1]  ( .D(n10269), .CK(clk), .Q(
        \xmem_data[23][1] ) );
  DFF_X1 \xmem_inst/mem_reg[22][1]  ( .D(n10268), .CK(clk), .Q(
        \xmem_data[22][1] ) );
  DFF_X1 \xmem_inst/mem_reg[21][1]  ( .D(n10267), .CK(clk), .Q(
        \xmem_data[21][1] ) );
  DFF_X1 \xmem_inst/mem_reg[20][1]  ( .D(n10266), .CK(clk), .Q(
        \xmem_data[20][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n10265), .CK(clk), .Q(
        \xmem_data[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n10264), .CK(clk), .Q(
        \xmem_data[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n10263), .CK(clk), .Q(
        \xmem_data[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n10262), .CK(clk), .Q(
        \xmem_data[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n10261), .CK(clk), .Q(
        \xmem_data[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n10260), .CK(clk), .Q(
        \xmem_data[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n10259), .CK(clk), .Q(
        \xmem_data[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n10258), .CK(clk), .Q(
        \xmem_data[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n10257), .CK(clk), .Q(
        \xmem_data[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n10256), .CK(clk), .Q(
        \xmem_data[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n10255), .CK(clk), .Q(
        \xmem_data[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n10254), .CK(clk), .Q(
        \xmem_data[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n10253), .CK(clk), .Q(
        \xmem_data[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n10252), .CK(clk), .Q(
        \xmem_data[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n10251), .CK(clk), .Q(
        \xmem_data[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n10250), .CK(clk), .Q(
        \xmem_data[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n10249), .CK(clk), .Q(
        \xmem_data[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n10248), .CK(clk), .Q(
        \xmem_data[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n10247), .CK(clk), .Q(
        \xmem_data[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n10246), .CK(clk), .Q(
        \xmem_data[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[25][0]  ( .D(n10245), .CK(clk), .Q(
        \xmem_data[25][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][0]  ( .D(n10244), .CK(clk), .Q(
        \xmem_data[24][0] ) );
  DFF_X1 \xmem_inst/mem_reg[23][0]  ( .D(n10243), .CK(clk), .Q(
        \xmem_data[23][0] ) );
  DFF_X1 \xmem_inst/mem_reg[22][0]  ( .D(n10242), .CK(clk), .Q(
        \xmem_data[22][0] ) );
  DFF_X1 \xmem_inst/mem_reg[21][0]  ( .D(n10241), .CK(clk), .Q(
        \xmem_data[21][0] ) );
  DFF_X1 \xmem_inst/mem_reg[20][0]  ( .D(n10240), .CK(clk), .Q(
        \xmem_data[20][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n10239), .CK(clk), .Q(
        \xmem_data[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n10238), .CK(clk), .Q(
        \xmem_data[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n10237), .CK(clk), .Q(
        \xmem_data[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n10236), .CK(clk), .Q(
        \xmem_data[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n10235), .CK(clk), .Q(
        \xmem_data[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n10234), .CK(clk), .Q(
        \xmem_data[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n10233), .CK(clk), .Q(
        \xmem_data[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n10232), .CK(clk), .Q(
        \xmem_data[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n10231), .CK(clk), .Q(
        \xmem_data[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n10230), .CK(clk), .Q(
        \xmem_data[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n10229), .CK(clk), .Q(
        \xmem_data[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n10228), .CK(clk), .Q(
        \xmem_data[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n10227), .CK(clk), .Q(
        \xmem_data[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n10226), .CK(clk), .Q(
        \xmem_data[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n10225), .CK(clk), .Q(
        \xmem_data[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n10224), .CK(clk), .Q(
        \xmem_data[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n10223), .CK(clk), .Q(
        \xmem_data[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n10222), .CK(clk), .Q(
        \xmem_data[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n10221), .CK(clk), .Q(
        \xmem_data[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n10220), .CK(clk), .Q(
        \xmem_data[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][7]  ( .D(n10219), .CK(clk), .Q(
        \xmem_data[24][7] ) );
  DFF_X1 \xmem_inst/mem_reg[23][7]  ( .D(n10218), .CK(clk), .Q(
        \xmem_data[23][7] ) );
  DFF_X1 \xmem_inst/mem_reg[22][7]  ( .D(n10217), .CK(clk), .Q(
        \xmem_data[22][7] ) );
  DFF_X1 \xmem_inst/mem_reg[21][7]  ( .D(n10216), .CK(clk), .Q(
        \xmem_data[21][7] ) );
  DFF_X1 \xmem_inst/mem_reg[20][7]  ( .D(n10215), .CK(clk), .Q(
        \xmem_data[20][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n10214), .CK(clk), .Q(
        \xmem_data[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n10213), .CK(clk), .Q(
        \xmem_data[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n10212), .CK(clk), .Q(
        \xmem_data[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n10211), .CK(clk), .Q(
        \xmem_data[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n10210), .CK(clk), .Q(
        \xmem_data[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n10209), .CK(clk), .Q(
        \xmem_data[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n10208), .CK(clk), .Q(
        \xmem_data[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n10207), .CK(clk), .Q(
        \xmem_data[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n10206), .CK(clk), .Q(
        \xmem_data[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n10205), .CK(clk), .Q(
        \xmem_data[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n10204), .CK(clk), .Q(
        \xmem_data[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n10203), .CK(clk), .Q(
        \xmem_data[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n10202), .CK(clk), .Q(
        \xmem_data[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n10201), .CK(clk), .Q(
        \xmem_data[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n10200), .CK(clk), .Q(
        \xmem_data[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n10199), .CK(clk), .Q(
        \xmem_data[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n10198), .CK(clk), .Q(
        \xmem_data[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n10197), .CK(clk), .Q(
        \xmem_data[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n10196), .CK(clk), .Q(
        \xmem_data[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n10195), .CK(clk), .Q(
        \xmem_data[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[24][6]  ( .D(n10194), .CK(clk), .Q(
        \xmem_data[24][6] ) );
  DFF_X1 \xmem_inst/mem_reg[23][6]  ( .D(n10193), .CK(clk), .Q(
        \xmem_data[23][6] ) );
  DFF_X1 \xmem_inst/mem_reg[22][6]  ( .D(n10192), .CK(clk), .Q(
        \xmem_data[22][6] ) );
  DFF_X1 \xmem_inst/mem_reg[21][6]  ( .D(n10191), .CK(clk), .Q(
        \xmem_data[21][6] ) );
  DFF_X1 \xmem_inst/mem_reg[20][6]  ( .D(n10190), .CK(clk), .Q(
        \xmem_data[20][6] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n10189), .CK(clk), .Q(
        \xmem_data[19][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n10188), .CK(clk), .Q(
        \xmem_data[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n10187), .CK(clk), .Q(
        \xmem_data[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n10186), .CK(clk), .Q(
        \xmem_data[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n10185), .CK(clk), .Q(
        \xmem_data[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n10184), .CK(clk), .Q(
        \xmem_data[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n10183), .CK(clk), .Q(
        \xmem_data[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n10182), .CK(clk), .Q(
        \xmem_data[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n10181), .CK(clk), .Q(
        \xmem_data[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n10180), .CK(clk), .Q(
        \xmem_data[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n10179), .CK(clk), .Q(
        \xmem_data[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n10178), .CK(clk), .Q(
        \xmem_data[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n10177), .CK(clk), .Q(
        \xmem_data[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n10176), .CK(clk), .Q(
        \xmem_data[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n10175), .CK(clk), .Q(
        \xmem_data[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n10174), .CK(clk), .Q(
        \xmem_data[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n10173), .CK(clk), .Q(
        \xmem_data[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n10172), .CK(clk), .Q(
        \xmem_data[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n10171), .CK(clk), .Q(
        \xmem_data[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n10170), .CK(clk), .Q(
        \xmem_data[0][6] ) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[3]  ( .D(n3118), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [3]), .QN(n8841) );
  DFF_X1 \ctrl_inst/state_reg[2]  ( .D(n3386), .CK(clk), .Q(
        \ctrl_inst/state [2]), .QN(n8806) );
  DFF_X1 \ctrl_inst/conv_done_reg  ( .D(n3390), .CK(clk), .Q(conv_done), .QN(
        n8844) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[0]  ( .D(n3383), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [0]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[1]  ( .D(n10421), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [1]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[2]  ( .D(n10420), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [2]), .QN(n8843) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[3]  ( .D(n10419), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [3]), .QN(n3483) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[4]  ( .D(n10418), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [4]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[5]  ( .D(n3378), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [5]), .QN(n8807) );
  DFF_X1 \ctrl_inst/state_reg[0]  ( .D(n3388), .CK(clk), .Q(
        \ctrl_inst/state [0]), .QN(n8813) );
  DFF_X1 \ctrl_inst/xmem_full_reg  ( .D(n3391), .CK(clk), .Q(xmem_full) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[3]  ( .D(n3396), .CK(clk), .Q(
        fmem_addr[3]), .QN(n8809) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[2]  ( .D(n3393), .CK(clk), .Q(
        fmem_addr[2]), .QN(n8804) );
  DFF_X1 \fmem_inst/mem_reg[0][0]  ( .D(n9645), .CK(clk), .Q(\fmem_data[0][0] ) );
  DFF_X1 \fmem_inst/mem_reg[0][1]  ( .D(n9644), .CK(clk), .Q(\fmem_data[0][1] ) );
  DFF_X1 \fmem_inst/mem_reg[0][2]  ( .D(n9643), .CK(clk), .Q(\fmem_data[0][2] ) );
  DFF_X1 \fmem_inst/mem_reg[0][3]  ( .D(n9642), .CK(clk), .Q(\fmem_data[0][3] ) );
  DFF_X1 \fmem_inst/mem_reg[0][4]  ( .D(n9641), .CK(clk), .Q(\fmem_data[0][4] ) );
  DFF_X1 \fmem_inst/mem_reg[0][5]  ( .D(n9640), .CK(clk), .Q(\fmem_data[0][5] ) );
  DFF_X1 \fmem_inst/mem_reg[0][6]  ( .D(n9639), .CK(clk), .Q(\fmem_data[0][6] ) );
  DFF_X1 \fmem_inst/mem_reg[0][7]  ( .D(n9638), .CK(clk), .Q(\fmem_data[0][7] ) );
  DFF_X1 \fmem_inst/mem_reg[1][0]  ( .D(n9637), .CK(clk), .Q(\fmem_data[1][0] ) );
  DFF_X1 \fmem_inst/mem_reg[1][1]  ( .D(n9636), .CK(clk), .Q(\fmem_data[1][1] ) );
  DFF_X1 \fmem_inst/mem_reg[1][2]  ( .D(n9635), .CK(clk), .Q(\fmem_data[1][2] ) );
  DFF_X1 \fmem_inst/mem_reg[1][3]  ( .D(n9634), .CK(clk), .Q(\fmem_data[1][3] ) );
  DFF_X1 \fmem_inst/mem_reg[1][4]  ( .D(n9633), .CK(clk), .Q(\fmem_data[1][4] ) );
  DFF_X1 \fmem_inst/mem_reg[1][5]  ( .D(n9632), .CK(clk), .Q(\fmem_data[1][5] ) );
  DFF_X1 \fmem_inst/mem_reg[1][6]  ( .D(n9631), .CK(clk), .Q(\fmem_data[1][6] ) );
  DFF_X1 \fmem_inst/mem_reg[1][7]  ( .D(n9630), .CK(clk), .Q(\fmem_data[1][7] ) );
  DFF_X1 \fmem_inst/mem_reg[2][0]  ( .D(n9629), .CK(clk), .Q(\fmem_data[2][0] ) );
  DFF_X1 \fmem_inst/mem_reg[2][1]  ( .D(n9628), .CK(clk), .Q(\fmem_data[2][1] ) );
  DFF_X1 \fmem_inst/mem_reg[2][2]  ( .D(n9627), .CK(clk), .Q(\fmem_data[2][2] ) );
  DFF_X1 \fmem_inst/mem_reg[2][3]  ( .D(n9626), .CK(clk), .Q(\fmem_data[2][3] ) );
  DFF_X1 \fmem_inst/mem_reg[2][4]  ( .D(n9625), .CK(clk), .Q(\fmem_data[2][4] ) );
  DFF_X1 \fmem_inst/mem_reg[2][5]  ( .D(n9624), .CK(clk), .Q(\fmem_data[2][5] ) );
  DFF_X1 \fmem_inst/mem_reg[2][6]  ( .D(n9623), .CK(clk), .Q(\fmem_data[2][6] ) );
  DFF_X1 \fmem_inst/mem_reg[2][7]  ( .D(n9622), .CK(clk), .Q(\fmem_data[2][7] ) );
  DFF_X1 \fmem_inst/mem_reg[3][0]  ( .D(n9621), .CK(clk), .Q(\fmem_data[3][0] ) );
  DFF_X1 \fmem_inst/mem_reg[3][1]  ( .D(n9620), .CK(clk), .Q(\fmem_data[3][1] ) );
  DFF_X1 \fmem_inst/mem_reg[3][2]  ( .D(n9619), .CK(clk), .Q(\fmem_data[3][2] ) );
  DFF_X1 \fmem_inst/mem_reg[3][3]  ( .D(n9618), .CK(clk), .Q(\fmem_data[3][3] ) );
  DFF_X1 \fmem_inst/mem_reg[3][4]  ( .D(n9617), .CK(clk), .Q(\fmem_data[3][4] ) );
  DFF_X1 \fmem_inst/mem_reg[3][5]  ( .D(n9616), .CK(clk), .Q(\fmem_data[3][5] ) );
  DFF_X1 \fmem_inst/mem_reg[3][6]  ( .D(n9615), .CK(clk), .Q(\fmem_data[3][6] ) );
  DFF_X1 \fmem_inst/mem_reg[3][7]  ( .D(n9614), .CK(clk), .Q(\fmem_data[3][7] ) );
  DFF_X1 \fmem_inst/mem_reg[4][0]  ( .D(n9613), .CK(clk), .Q(\fmem_data[4][0] ) );
  DFF_X1 \fmem_inst/mem_reg[4][1]  ( .D(n9612), .CK(clk), .Q(\fmem_data[4][1] ) );
  DFF_X1 \fmem_inst/mem_reg[4][2]  ( .D(n9611), .CK(clk), .Q(\fmem_data[4][2] ) );
  DFF_X1 \fmem_inst/mem_reg[4][3]  ( .D(n9610), .CK(clk), .Q(\fmem_data[4][3] ) );
  DFF_X1 \fmem_inst/mem_reg[4][4]  ( .D(n9609), .CK(clk), .Q(\fmem_data[4][4] ) );
  DFF_X1 \fmem_inst/mem_reg[4][5]  ( .D(n9608), .CK(clk), .Q(\fmem_data[4][5] ) );
  DFF_X1 \fmem_inst/mem_reg[4][6]  ( .D(n9607), .CK(clk), .Q(\fmem_data[4][6] ) );
  DFF_X1 \fmem_inst/mem_reg[4][7]  ( .D(n9606), .CK(clk), .Q(\fmem_data[4][7] ) );
  DFF_X1 \fmem_inst/mem_reg[5][0]  ( .D(n9605), .CK(clk), .Q(\fmem_data[5][0] ) );
  DFF_X1 \fmem_inst/mem_reg[5][1]  ( .D(n9604), .CK(clk), .Q(\fmem_data[5][1] ) );
  DFF_X1 \fmem_inst/mem_reg[5][2]  ( .D(n9603), .CK(clk), .Q(\fmem_data[5][2] ) );
  DFF_X1 \fmem_inst/mem_reg[5][3]  ( .D(n9602), .CK(clk), .Q(\fmem_data[5][3] ) );
  DFF_X1 \fmem_inst/mem_reg[5][4]  ( .D(n9601), .CK(clk), .Q(\fmem_data[5][4] ) );
  DFF_X1 \fmem_inst/mem_reg[5][5]  ( .D(n9600), .CK(clk), .Q(\fmem_data[5][5] ) );
  DFF_X1 \fmem_inst/mem_reg[5][6]  ( .D(n9599), .CK(clk), .Q(\fmem_data[5][6] ) );
  DFF_X1 \fmem_inst/mem_reg[5][7]  ( .D(n9598), .CK(clk), .Q(\fmem_data[5][7] ) );
  DFF_X1 \fmem_inst/mem_reg[6][0]  ( .D(n9597), .CK(clk), .Q(\fmem_data[6][0] ) );
  DFF_X1 \fmem_inst/mem_reg[6][1]  ( .D(n9596), .CK(clk), .Q(\fmem_data[6][1] ) );
  DFF_X1 \fmem_inst/mem_reg[6][2]  ( .D(n9595), .CK(clk), .Q(\fmem_data[6][2] ) );
  DFF_X1 \fmem_inst/mem_reg[6][3]  ( .D(n9594), .CK(clk), .Q(\fmem_data[6][3] ) );
  DFF_X1 \fmem_inst/mem_reg[6][4]  ( .D(n9593), .CK(clk), .Q(\fmem_data[6][4] ) );
  DFF_X1 \fmem_inst/mem_reg[6][5]  ( .D(n9592), .CK(clk), .Q(\fmem_data[6][5] ) );
  DFF_X1 \fmem_inst/mem_reg[6][6]  ( .D(n9591), .CK(clk), .Q(\fmem_data[6][6] ) );
  DFF_X1 \fmem_inst/mem_reg[6][7]  ( .D(n9590), .CK(clk), .Q(\fmem_data[6][7] ) );
  DFF_X1 \fmem_inst/mem_reg[7][0]  ( .D(n9589), .CK(clk), .Q(\fmem_data[7][0] ) );
  DFF_X1 \fmem_inst/mem_reg[7][1]  ( .D(n9588), .CK(clk), .Q(\fmem_data[7][1] ) );
  DFF_X1 \fmem_inst/mem_reg[7][2]  ( .D(n9587), .CK(clk), .Q(\fmem_data[7][2] ) );
  DFF_X1 \fmem_inst/mem_reg[7][3]  ( .D(n9586), .CK(clk), .Q(\fmem_data[7][3] ) );
  DFF_X1 \fmem_inst/mem_reg[7][4]  ( .D(n9585), .CK(clk), .Q(\fmem_data[7][4] ) );
  DFF_X1 \fmem_inst/mem_reg[7][5]  ( .D(n9584), .CK(clk), .Q(\fmem_data[7][5] ) );
  DFF_X1 \fmem_inst/mem_reg[7][6]  ( .D(n9583), .CK(clk), .Q(\fmem_data[7][6] ) );
  DFF_X1 \fmem_inst/mem_reg[7][7]  ( .D(n9582), .CK(clk), .Q(\fmem_data[7][7] ) );
  DFF_X1 \fmem_inst/mem_reg[8][0]  ( .D(n9581), .CK(clk), .Q(\fmem_data[8][0] ) );
  DFF_X1 \fmem_inst/mem_reg[8][1]  ( .D(n9580), .CK(clk), .Q(\fmem_data[8][1] ) );
  DFF_X1 \fmem_inst/mem_reg[8][2]  ( .D(n9579), .CK(clk), .Q(\fmem_data[8][2] ) );
  DFF_X1 \fmem_inst/mem_reg[8][3]  ( .D(n9578), .CK(clk), .Q(\fmem_data[8][3] ) );
  DFF_X1 \fmem_inst/mem_reg[8][4]  ( .D(n9577), .CK(clk), .Q(\fmem_data[8][4] ) );
  DFF_X1 \fmem_inst/mem_reg[8][5]  ( .D(n9576), .CK(clk), .Q(\fmem_data[8][5] ) );
  DFF_X1 \fmem_inst/mem_reg[8][6]  ( .D(n9575), .CK(clk), .Q(\fmem_data[8][6] ) );
  DFF_X1 \fmem_inst/mem_reg[8][7]  ( .D(n9574), .CK(clk), .Q(\fmem_data[8][7] ) );
  DFF_X1 \fmem_inst/mem_reg[9][0]  ( .D(n9573), .CK(clk), .Q(\fmem_data[9][0] ) );
  DFF_X1 \fmem_inst/mem_reg[9][1]  ( .D(n9572), .CK(clk), .Q(\fmem_data[9][1] ) );
  DFF_X1 \fmem_inst/mem_reg[9][2]  ( .D(n9571), .CK(clk), .Q(\fmem_data[9][2] ) );
  DFF_X1 \fmem_inst/mem_reg[9][3]  ( .D(n9570), .CK(clk), .Q(\fmem_data[9][3] ) );
  DFF_X1 \fmem_inst/mem_reg[9][4]  ( .D(n9569), .CK(clk), .Q(\fmem_data[9][4] ) );
  DFF_X1 \fmem_inst/mem_reg[9][5]  ( .D(n9568), .CK(clk), .Q(\fmem_data[9][5] ) );
  DFF_X1 \fmem_inst/mem_reg[9][6]  ( .D(n9567), .CK(clk), .Q(\fmem_data[9][6] ) );
  DFF_X1 \fmem_inst/mem_reg[9][7]  ( .D(n9566), .CK(clk), .Q(\fmem_data[9][7] ) );
  DFF_X1 \fmem_inst/mem_reg[10][0]  ( .D(n9565), .CK(clk), .Q(
        \fmem_data[10][0] ) );
  DFF_X1 \fmem_inst/mem_reg[10][1]  ( .D(n9564), .CK(clk), .Q(
        \fmem_data[10][1] ) );
  DFF_X1 \fmem_inst/mem_reg[10][2]  ( .D(n9563), .CK(clk), .Q(
        \fmem_data[10][2] ) );
  DFF_X1 \fmem_inst/mem_reg[10][3]  ( .D(n9562), .CK(clk), .Q(
        \fmem_data[10][3] ) );
  DFF_X1 \fmem_inst/mem_reg[10][4]  ( .D(n9561), .CK(clk), .Q(
        \fmem_data[10][4] ) );
  DFF_X1 \fmem_inst/mem_reg[10][5]  ( .D(n9560), .CK(clk), .Q(
        \fmem_data[10][5] ) );
  DFF_X1 \fmem_inst/mem_reg[10][6]  ( .D(n9559), .CK(clk), .Q(
        \fmem_data[10][6] ) );
  DFF_X1 \fmem_inst/mem_reg[10][7]  ( .D(n9558), .CK(clk), .Q(
        \fmem_data[10][7] ) );
  DFF_X1 \fmem_inst/mem_reg[11][0]  ( .D(n9557), .CK(clk), .Q(
        \fmem_data[11][0] ) );
  DFF_X1 \fmem_inst/mem_reg[11][1]  ( .D(n9556), .CK(clk), .Q(
        \fmem_data[11][1] ) );
  DFF_X1 \fmem_inst/mem_reg[11][2]  ( .D(n9555), .CK(clk), .Q(
        \fmem_data[11][2] ) );
  DFF_X1 \fmem_inst/mem_reg[11][3]  ( .D(n9554), .CK(clk), .Q(
        \fmem_data[11][3] ) );
  DFF_X1 \fmem_inst/mem_reg[11][4]  ( .D(n9553), .CK(clk), .Q(
        \fmem_data[11][4] ) );
  DFF_X1 \fmem_inst/mem_reg[11][5]  ( .D(n9552), .CK(clk), .Q(
        \fmem_data[11][5] ) );
  DFF_X1 \fmem_inst/mem_reg[11][6]  ( .D(n9551), .CK(clk), .Q(
        \fmem_data[11][6] ) );
  DFF_X1 \fmem_inst/mem_reg[11][7]  ( .D(n9550), .CK(clk), .Q(
        \fmem_data[11][7] ) );
  DFF_X1 \fmem_inst/mem_reg[12][0]  ( .D(n9549), .CK(clk), .Q(
        \fmem_data[12][0] ) );
  DFF_X1 \fmem_inst/mem_reg[12][1]  ( .D(n9548), .CK(clk), .Q(
        \fmem_data[12][1] ) );
  DFF_X1 \fmem_inst/mem_reg[12][2]  ( .D(n9547), .CK(clk), .Q(
        \fmem_data[12][2] ) );
  DFF_X1 \fmem_inst/mem_reg[12][3]  ( .D(n9546), .CK(clk), .Q(
        \fmem_data[12][3] ) );
  DFF_X1 \fmem_inst/mem_reg[12][4]  ( .D(n9545), .CK(clk), .Q(
        \fmem_data[12][4] ) );
  DFF_X1 \fmem_inst/mem_reg[12][5]  ( .D(n9544), .CK(clk), .Q(
        \fmem_data[12][5] ) );
  DFF_X1 \fmem_inst/mem_reg[12][6]  ( .D(n9543), .CK(clk), .Q(
        \fmem_data[12][6] ) );
  DFF_X1 \fmem_inst/mem_reg[12][7]  ( .D(n9542), .CK(clk), .Q(
        \fmem_data[12][7] ) );
  DFF_X1 \fmem_inst/mem_reg[13][0]  ( .D(n9541), .CK(clk), .Q(
        \fmem_data[13][0] ) );
  DFF_X1 \fmem_inst/mem_reg[13][1]  ( .D(n9540), .CK(clk), .Q(
        \fmem_data[13][1] ) );
  DFF_X1 \fmem_inst/mem_reg[13][2]  ( .D(n9539), .CK(clk), .Q(
        \fmem_data[13][2] ) );
  DFF_X1 \fmem_inst/mem_reg[13][3]  ( .D(n9538), .CK(clk), .Q(
        \fmem_data[13][3] ) );
  DFF_X1 \fmem_inst/mem_reg[13][4]  ( .D(n9537), .CK(clk), .Q(
        \fmem_data[13][4] ) );
  DFF_X1 \fmem_inst/mem_reg[13][5]  ( .D(n9536), .CK(clk), .Q(
        \fmem_data[13][5] ) );
  DFF_X1 \fmem_inst/mem_reg[13][6]  ( .D(n9535), .CK(clk), .Q(
        \fmem_data[13][6] ) );
  DFF_X1 \fmem_inst/mem_reg[13][7]  ( .D(n9534), .CK(clk), .Q(
        \fmem_data[13][7] ) );
  DFF_X1 \fmem_inst/mem_reg[14][0]  ( .D(n9533), .CK(clk), .Q(
        \fmem_data[14][0] ) );
  DFF_X1 \fmem_inst/mem_reg[14][1]  ( .D(n9532), .CK(clk), .Q(
        \fmem_data[14][1] ) );
  DFF_X1 \fmem_inst/mem_reg[14][2]  ( .D(n9531), .CK(clk), .Q(
        \fmem_data[14][2] ) );
  DFF_X1 \fmem_inst/mem_reg[14][3]  ( .D(n9530), .CK(clk), .Q(
        \fmem_data[14][3] ) );
  DFF_X1 \fmem_inst/mem_reg[14][4]  ( .D(n9529), .CK(clk), .Q(
        \fmem_data[14][4] ) );
  DFF_X1 \fmem_inst/mem_reg[14][5]  ( .D(n9528), .CK(clk), .Q(
        \fmem_data[14][5] ) );
  DFF_X1 \fmem_inst/mem_reg[14][6]  ( .D(n9527), .CK(clk), .Q(
        \fmem_data[14][6] ) );
  DFF_X1 \fmem_inst/mem_reg[14][7]  ( .D(n9526), .CK(clk), .Q(
        \fmem_data[14][7] ) );
  DFF_X1 \fmem_inst/mem_reg[15][0]  ( .D(n9525), .CK(clk), .Q(
        \fmem_data[15][0] ) );
  DFF_X1 \fmem_inst/mem_reg[15][1]  ( .D(n9524), .CK(clk), .Q(
        \fmem_data[15][1] ) );
  DFF_X1 \fmem_inst/mem_reg[15][2]  ( .D(n9523), .CK(clk), .Q(
        \fmem_data[15][2] ) );
  DFF_X1 \fmem_inst/mem_reg[15][3]  ( .D(n9522), .CK(clk), .Q(
        \fmem_data[15][3] ) );
  DFF_X1 \fmem_inst/mem_reg[15][4]  ( .D(n9521), .CK(clk), .Q(
        \fmem_data[15][4] ) );
  DFF_X1 \fmem_inst/mem_reg[15][5]  ( .D(n9520), .CK(clk), .Q(
        \fmem_data[15][5] ) );
  DFF_X1 \fmem_inst/mem_reg[15][6]  ( .D(n9519), .CK(clk), .Q(
        \fmem_data[15][6] ) );
  DFF_X1 \fmem_inst/mem_reg[15][7]  ( .D(n9518), .CK(clk), .Q(
        \fmem_data[15][7] ) );
  DFF_X1 \fmem_inst/mem_reg[16][0]  ( .D(n9517), .CK(clk), .Q(
        \fmem_data[16][0] ) );
  DFF_X1 \fmem_inst/mem_reg[16][1]  ( .D(n9516), .CK(clk), .Q(
        \fmem_data[16][1] ) );
  DFF_X1 \fmem_inst/mem_reg[16][2]  ( .D(n9515), .CK(clk), .Q(
        \fmem_data[16][2] ) );
  DFF_X1 \fmem_inst/mem_reg[16][3]  ( .D(n9514), .CK(clk), .Q(
        \fmem_data[16][3] ) );
  DFF_X1 \fmem_inst/mem_reg[16][4]  ( .D(n9513), .CK(clk), .Q(
        \fmem_data[16][4] ) );
  DFF_X1 \fmem_inst/mem_reg[16][5]  ( .D(n9512), .CK(clk), .Q(
        \fmem_data[16][5] ) );
  DFF_X1 \fmem_inst/mem_reg[16][6]  ( .D(n9511), .CK(clk), .Q(
        \fmem_data[16][6] ) );
  DFF_X1 \fmem_inst/mem_reg[16][7]  ( .D(n9510), .CK(clk), .Q(
        \fmem_data[16][7] ) );
  DFF_X1 \fmem_inst/mem_reg[17][0]  ( .D(n9509), .CK(clk), .Q(
        \fmem_data[17][0] ) );
  DFF_X1 \fmem_inst/mem_reg[17][1]  ( .D(n9508), .CK(clk), .Q(
        \fmem_data[17][1] ) );
  DFF_X1 \fmem_inst/mem_reg[17][2]  ( .D(n9507), .CK(clk), .Q(
        \fmem_data[17][2] ) );
  DFF_X1 \fmem_inst/mem_reg[17][3]  ( .D(n9506), .CK(clk), .Q(
        \fmem_data[17][3] ) );
  DFF_X1 \fmem_inst/mem_reg[17][4]  ( .D(n9505), .CK(clk), .Q(
        \fmem_data[17][4] ) );
  DFF_X1 \fmem_inst/mem_reg[17][5]  ( .D(n9504), .CK(clk), .Q(
        \fmem_data[17][5] ) );
  DFF_X1 \fmem_inst/mem_reg[17][6]  ( .D(n9503), .CK(clk), .Q(
        \fmem_data[17][6] ) );
  DFF_X1 \fmem_inst/mem_reg[17][7]  ( .D(n9502), .CK(clk), .Q(
        \fmem_data[17][7] ) );
  DFF_X1 \fmem_inst/mem_reg[18][0]  ( .D(n9501), .CK(clk), .Q(
        \fmem_data[18][0] ) );
  DFF_X1 \fmem_inst/mem_reg[18][1]  ( .D(n9500), .CK(clk), .Q(
        \fmem_data[18][1] ) );
  DFF_X1 \fmem_inst/mem_reg[18][2]  ( .D(n9499), .CK(clk), .Q(
        \fmem_data[18][2] ) );
  DFF_X1 \fmem_inst/mem_reg[18][3]  ( .D(n9498), .CK(clk), .Q(
        \fmem_data[18][3] ) );
  DFF_X1 \fmem_inst/mem_reg[18][4]  ( .D(n9497), .CK(clk), .Q(
        \fmem_data[18][4] ) );
  DFF_X1 \fmem_inst/mem_reg[18][5]  ( .D(n9496), .CK(clk), .Q(
        \fmem_data[18][5] ) );
  DFF_X1 \fmem_inst/mem_reg[18][6]  ( .D(n9495), .CK(clk), .Q(
        \fmem_data[18][6] ) );
  DFF_X1 \fmem_inst/mem_reg[18][7]  ( .D(n9494), .CK(clk), .Q(
        \fmem_data[18][7] ) );
  DFF_X1 \fmem_inst/mem_reg[19][0]  ( .D(n9493), .CK(clk), .Q(
        \fmem_data[19][0] ) );
  DFF_X1 \fmem_inst/mem_reg[19][1]  ( .D(n9492), .CK(clk), .Q(
        \fmem_data[19][1] ) );
  DFF_X1 \fmem_inst/mem_reg[19][2]  ( .D(n9491), .CK(clk), .Q(
        \fmem_data[19][2] ) );
  DFF_X1 \fmem_inst/mem_reg[19][3]  ( .D(n9490), .CK(clk), .Q(
        \fmem_data[19][3] ) );
  DFF_X1 \fmem_inst/mem_reg[19][4]  ( .D(n9489), .CK(clk), .Q(
        \fmem_data[19][4] ) );
  DFF_X1 \fmem_inst/mem_reg[19][5]  ( .D(n9488), .CK(clk), .Q(
        \fmem_data[19][5] ) );
  DFF_X1 \fmem_inst/mem_reg[19][6]  ( .D(n9487), .CK(clk), .Q(
        \fmem_data[19][6] ) );
  DFF_X1 \fmem_inst/mem_reg[19][7]  ( .D(n9486), .CK(clk), .Q(
        \fmem_data[19][7] ) );
  DFF_X1 \fmem_inst/mem_reg[20][0]  ( .D(n9485), .CK(clk), .Q(
        \fmem_data[20][0] ) );
  DFF_X1 \fmem_inst/mem_reg[20][1]  ( .D(n9484), .CK(clk), .Q(
        \fmem_data[20][1] ) );
  DFF_X1 \fmem_inst/mem_reg[20][2]  ( .D(n9483), .CK(clk), .Q(
        \fmem_data[20][2] ) );
  DFF_X1 \fmem_inst/mem_reg[20][3]  ( .D(n9482), .CK(clk), .Q(
        \fmem_data[20][3] ) );
  DFF_X1 \fmem_inst/mem_reg[20][4]  ( .D(n9481), .CK(clk), .Q(
        \fmem_data[20][4] ) );
  DFF_X1 \fmem_inst/mem_reg[20][5]  ( .D(n9480), .CK(clk), .Q(
        \fmem_data[20][5] ) );
  DFF_X1 \fmem_inst/mem_reg[20][6]  ( .D(n9479), .CK(clk), .Q(
        \fmem_data[20][6] ) );
  DFF_X1 \fmem_inst/mem_reg[20][7]  ( .D(n9478), .CK(clk), .Q(
        \fmem_data[20][7] ) );
  DFF_X1 \fmem_inst/mem_reg[21][0]  ( .D(n9477), .CK(clk), .Q(
        \fmem_data[21][0] ) );
  DFF_X1 \fmem_inst/mem_reg[21][1]  ( .D(n9476), .CK(clk), .Q(
        \fmem_data[21][1] ) );
  DFF_X1 \fmem_inst/mem_reg[21][2]  ( .D(n9475), .CK(clk), .Q(
        \fmem_data[21][2] ) );
  DFF_X1 \fmem_inst/mem_reg[21][3]  ( .D(n9474), .CK(clk), .Q(
        \fmem_data[21][3] ) );
  DFF_X1 \fmem_inst/mem_reg[21][4]  ( .D(n9473), .CK(clk), .Q(
        \fmem_data[21][4] ) );
  DFF_X1 \fmem_inst/mem_reg[21][5]  ( .D(n9472), .CK(clk), .Q(
        \fmem_data[21][5] ) );
  DFF_X1 \fmem_inst/mem_reg[21][6]  ( .D(n9471), .CK(clk), .Q(
        \fmem_data[21][6] ) );
  DFF_X1 \fmem_inst/mem_reg[21][7]  ( .D(n9470), .CK(clk), .Q(
        \fmem_data[21][7] ) );
  DFF_X1 \fmem_inst/mem_reg[22][0]  ( .D(n9469), .CK(clk), .Q(
        \fmem_data[22][0] ) );
  DFF_X1 \fmem_inst/mem_reg[22][1]  ( .D(n9468), .CK(clk), .Q(
        \fmem_data[22][1] ) );
  DFF_X1 \fmem_inst/mem_reg[22][2]  ( .D(n9467), .CK(clk), .Q(
        \fmem_data[22][2] ) );
  DFF_X1 \fmem_inst/mem_reg[22][3]  ( .D(n9466), .CK(clk), .Q(
        \fmem_data[22][3] ) );
  DFF_X1 \fmem_inst/mem_reg[22][4]  ( .D(n9465), .CK(clk), .Q(
        \fmem_data[22][4] ) );
  DFF_X1 \fmem_inst/mem_reg[22][5]  ( .D(n9464), .CK(clk), .Q(
        \fmem_data[22][5] ) );
  DFF_X1 \fmem_inst/mem_reg[22][6]  ( .D(n9463), .CK(clk), .Q(
        \fmem_data[22][6] ) );
  DFF_X1 \fmem_inst/mem_reg[22][7]  ( .D(n9462), .CK(clk), .Q(
        \fmem_data[22][7] ) );
  DFF_X1 \fmem_inst/mem_reg[23][0]  ( .D(n9461), .CK(clk), .Q(
        \fmem_data[23][0] ) );
  DFF_X1 \fmem_inst/mem_reg[23][1]  ( .D(n9460), .CK(clk), .Q(
        \fmem_data[23][1] ) );
  DFF_X1 \fmem_inst/mem_reg[23][2]  ( .D(n9459), .CK(clk), .Q(
        \fmem_data[23][2] ) );
  DFF_X1 \fmem_inst/mem_reg[23][3]  ( .D(n9458), .CK(clk), .Q(
        \fmem_data[23][3] ) );
  DFF_X1 \fmem_inst/mem_reg[23][4]  ( .D(n9457), .CK(clk), .Q(
        \fmem_data[23][4] ) );
  DFF_X1 \fmem_inst/mem_reg[23][5]  ( .D(n9456), .CK(clk), .Q(
        \fmem_data[23][5] ) );
  DFF_X1 \fmem_inst/mem_reg[23][6]  ( .D(n9455), .CK(clk), .Q(
        \fmem_data[23][6] ) );
  DFF_X1 \fmem_inst/mem_reg[23][7]  ( .D(n9454), .CK(clk), .Q(
        \fmem_data[23][7] ) );
  DFF_X1 \fmem_inst/mem_reg[24][0]  ( .D(n9453), .CK(clk), .Q(
        \fmem_data[24][0] ) );
  DFF_X1 \fmem_inst/mem_reg[24][1]  ( .D(n9452), .CK(clk), .Q(
        \fmem_data[24][1] ) );
  DFF_X1 \fmem_inst/mem_reg[24][2]  ( .D(n9451), .CK(clk), .Q(
        \fmem_data[24][2] ) );
  DFF_X1 \fmem_inst/mem_reg[24][3]  ( .D(n9450), .CK(clk), .Q(
        \fmem_data[24][3] ) );
  DFF_X1 \fmem_inst/mem_reg[24][4]  ( .D(n9449), .CK(clk), .Q(
        \fmem_data[24][4] ) );
  DFF_X1 \fmem_inst/mem_reg[24][5]  ( .D(n9448), .CK(clk), .Q(
        \fmem_data[24][5] ) );
  DFF_X1 \fmem_inst/mem_reg[24][6]  ( .D(n9447), .CK(clk), .Q(
        \fmem_data[24][6] ) );
  DFF_X1 \fmem_inst/mem_reg[24][7]  ( .D(n9446), .CK(clk), .Q(
        \fmem_data[24][7] ) );
  DFF_X1 \fmem_inst/mem_reg[25][0]  ( .D(n9445), .CK(clk), .Q(
        \fmem_data[25][0] ) );
  DFF_X1 \fmem_inst/mem_reg[25][1]  ( .D(n9444), .CK(clk), .Q(
        \fmem_data[25][1] ) );
  DFF_X1 \fmem_inst/mem_reg[25][2]  ( .D(n9443), .CK(clk), .Q(
        \fmem_data[25][2] ) );
  DFF_X1 \fmem_inst/mem_reg[25][3]  ( .D(n9442), .CK(clk), .Q(
        \fmem_data[25][3] ) );
  DFF_X1 \fmem_inst/mem_reg[25][4]  ( .D(n9441), .CK(clk), .Q(
        \fmem_data[25][4] ) );
  DFF_X1 \fmem_inst/mem_reg[25][5]  ( .D(n9440), .CK(clk), .Q(
        \fmem_data[25][5] ) );
  DFF_X1 \fmem_inst/mem_reg[25][6]  ( .D(n9439), .CK(clk), .Q(
        \fmem_data[25][6] ) );
  DFF_X1 \fmem_inst/mem_reg[25][7]  ( .D(n9438), .CK(clk), .Q(
        \fmem_data[25][7] ) );
  DFF_X1 \fmem_inst/mem_reg[26][0]  ( .D(n9437), .CK(clk), .Q(
        \fmem_data[26][0] ) );
  DFF_X1 \fmem_inst/mem_reg[26][1]  ( .D(n9436), .CK(clk), .Q(
        \fmem_data[26][1] ) );
  DFF_X1 \fmem_inst/mem_reg[26][2]  ( .D(n9435), .CK(clk), .Q(
        \fmem_data[26][2] ) );
  DFF_X1 \fmem_inst/mem_reg[26][3]  ( .D(n9434), .CK(clk), .Q(
        \fmem_data[26][3] ) );
  DFF_X1 \fmem_inst/mem_reg[26][4]  ( .D(n9433), .CK(clk), .Q(
        \fmem_data[26][4] ) );
  DFF_X1 \fmem_inst/mem_reg[26][5]  ( .D(n9432), .CK(clk), .Q(
        \fmem_data[26][5] ) );
  DFF_X1 \fmem_inst/mem_reg[26][6]  ( .D(n9431), .CK(clk), .Q(
        \fmem_data[26][6] ) );
  DFF_X1 \fmem_inst/mem_reg[26][7]  ( .D(n9430), .CK(clk), .Q(
        \fmem_data[26][7] ) );
  DFF_X1 \fmem_inst/mem_reg[27][0]  ( .D(n9429), .CK(clk), .Q(
        \fmem_data[27][0] ) );
  DFF_X1 \fmem_inst/mem_reg[27][1]  ( .D(n9428), .CK(clk), .Q(
        \fmem_data[27][1] ) );
  DFF_X1 \fmem_inst/mem_reg[27][2]  ( .D(n9427), .CK(clk), .Q(
        \fmem_data[27][2] ) );
  DFF_X1 \fmem_inst/mem_reg[27][3]  ( .D(n9426), .CK(clk), .Q(
        \fmem_data[27][3] ) );
  DFF_X1 \fmem_inst/mem_reg[27][4]  ( .D(n9425), .CK(clk), .Q(
        \fmem_data[27][4] ) );
  DFF_X1 \fmem_inst/mem_reg[27][5]  ( .D(n9424), .CK(clk), .Q(
        \fmem_data[27][5] ) );
  DFF_X1 \fmem_inst/mem_reg[27][6]  ( .D(n9423), .CK(clk), .Q(
        \fmem_data[27][6] ) );
  DFF_X1 \fmem_inst/mem_reg[27][7]  ( .D(n9422), .CK(clk), .Q(
        \fmem_data[27][7] ) );
  DFF_X1 \fmem_inst/mem_reg[28][0]  ( .D(n9421), .CK(clk), .Q(
        \fmem_data[28][0] ) );
  DFF_X1 \fmem_inst/mem_reg[28][1]  ( .D(n9420), .CK(clk), .Q(
        \fmem_data[28][1] ) );
  DFF_X1 \fmem_inst/mem_reg[28][2]  ( .D(n9419), .CK(clk), .Q(
        \fmem_data[28][2] ) );
  DFF_X1 \fmem_inst/mem_reg[28][3]  ( .D(n9418), .CK(clk), .Q(
        \fmem_data[28][3] ) );
  DFF_X1 \fmem_inst/mem_reg[28][4]  ( .D(n9417), .CK(clk), .Q(
        \fmem_data[28][4] ) );
  DFF_X1 \fmem_inst/mem_reg[28][5]  ( .D(n9416), .CK(clk), .Q(
        \fmem_data[28][5] ) );
  DFF_X1 \fmem_inst/mem_reg[28][6]  ( .D(n9415), .CK(clk), .Q(
        \fmem_data[28][6] ) );
  DFF_X1 \fmem_inst/mem_reg[28][7]  ( .D(n9414), .CK(clk), .Q(
        \fmem_data[28][7] ) );
  DFF_X1 \fmem_inst/mem_reg[29][0]  ( .D(n9413), .CK(clk), .Q(
        \fmem_data[29][0] ) );
  DFF_X1 \fmem_inst/mem_reg[29][1]  ( .D(n9412), .CK(clk), .Q(
        \fmem_data[29][1] ) );
  DFF_X1 \fmem_inst/mem_reg[29][2]  ( .D(n9411), .CK(clk), .Q(
        \fmem_data[29][2] ) );
  DFF_X1 \fmem_inst/mem_reg[29][3]  ( .D(n9410), .CK(clk), .Q(
        \fmem_data[29][3] ) );
  DFF_X1 \fmem_inst/mem_reg[29][4]  ( .D(n9409), .CK(clk), .Q(
        \fmem_data[29][4] ) );
  DFF_X1 \fmem_inst/mem_reg[29][5]  ( .D(n9408), .CK(clk), .Q(
        \fmem_data[29][5] ) );
  DFF_X1 \fmem_inst/mem_reg[29][6]  ( .D(n9407), .CK(clk), .Q(
        \fmem_data[29][6] ) );
  DFF_X1 \fmem_inst/mem_reg[29][7]  ( .D(n9406), .CK(clk), .Q(
        \fmem_data[29][7] ) );
  DFF_X1 \fmem_inst/mem_reg[30][0]  ( .D(n9405), .CK(clk), .Q(
        \fmem_data[30][0] ) );
  DFF_X1 \fmem_inst/mem_reg[30][1]  ( .D(n9404), .CK(clk), .Q(
        \fmem_data[30][1] ) );
  DFF_X1 \fmem_inst/mem_reg[30][2]  ( .D(n9403), .CK(clk), .Q(
        \fmem_data[30][2] ) );
  DFF_X1 \fmem_inst/mem_reg[30][3]  ( .D(n9402), .CK(clk), .Q(
        \fmem_data[30][3] ) );
  DFF_X1 \fmem_inst/mem_reg[30][4]  ( .D(n9401), .CK(clk), .Q(
        \fmem_data[30][4] ) );
  DFF_X1 \fmem_inst/mem_reg[30][5]  ( .D(n9400), .CK(clk), .Q(
        \fmem_data[30][5] ) );
  DFF_X1 \fmem_inst/mem_reg[30][6]  ( .D(n9399), .CK(clk), .Q(
        \fmem_data[30][6] ) );
  DFF_X1 \fmem_inst/mem_reg[30][7]  ( .D(n9398), .CK(clk), .Q(
        \fmem_data[30][7] ) );
  DFF_X1 \fmem_inst/mem_reg[31][0]  ( .D(n9397), .CK(clk), .Q(
        \fmem_data[31][0] ) );
  DFF_X1 \fmem_inst/mem_reg[31][1]  ( .D(n9396), .CK(clk), .Q(
        \fmem_data[31][1] ) );
  DFF_X1 \fmem_inst/mem_reg[31][2]  ( .D(n9395), .CK(clk), .Q(
        \fmem_data[31][2] ) );
  DFF_X1 \fmem_inst/mem_reg[31][3]  ( .D(n9394), .CK(clk), .Q(
        \fmem_data[31][3] ) );
  DFF_X1 \fmem_inst/mem_reg[31][4]  ( .D(n9393), .CK(clk), .Q(
        \fmem_data[31][4] ) );
  DFF_X1 \fmem_inst/mem_reg[31][5]  ( .D(n9392), .CK(clk), .Q(
        \fmem_data[31][5] ) );
  DFF_X1 \fmem_inst/mem_reg[31][6]  ( .D(n9391), .CK(clk), .Q(
        \fmem_data[31][6] ) );
  DFF_X1 \fmem_inst/mem_reg[31][7]  ( .D(n9390), .CK(clk), .Q(
        \fmem_data[31][7] ) );
  DFF_X1 \x_mult_f_reg[0][0]  ( .D(n9327), .CK(clk), .Q(\x_mult_f[0][0] ) );
  DFF_X1 \x_mult_f_reg[0][1]  ( .D(n9326), .CK(clk), .Q(\x_mult_f[0][1] ) );
  DFF_X1 \x_mult_f_reg[0][2]  ( .D(n8926), .CK(clk), .Q(\x_mult_f[0][2] ) );
  DFF_X1 \x_mult_f_reg[0][3]  ( .D(n8925), .CK(clk), .Q(\x_mult_f[0][3] ) );
  DFF_X1 \x_mult_f_reg[0][4]  ( .D(n8924), .CK(clk), .Q(\x_mult_f[0][4] ) );
  DFF_X1 \x_mult_f_reg[0][5]  ( .D(n8923), .CK(clk), .Q(\x_mult_f[0][5] ) );
  DFF_X1 \x_mult_f_reg[0][6]  ( .D(n8922), .CK(clk), .Q(\x_mult_f[0][6] ) );
  DFF_X1 \x_mult_f_reg[0][7]  ( .D(n8921), .CK(clk), .Q(\x_mult_f[0][7] ) );
  DFF_X1 \x_mult_f_reg[0][8]  ( .D(n8920), .CK(clk), .Q(\x_mult_f[0][8] ) );
  DFF_X1 \x_mult_f_reg[0][9]  ( .D(n8919), .CK(clk), .Q(\x_mult_f[0][9] ) );
  DFF_X1 \x_mult_f_reg[0][10]  ( .D(n8918), .CK(clk), .Q(\x_mult_f[0][10] ) );
  DFF_X1 \x_mult_f_reg[0][11]  ( .D(n8917), .CK(clk), .Q(\x_mult_f[0][11] ) );
  DFF_X1 \x_mult_f_reg[0][12]  ( .D(n8916), .CK(clk), .Q(\x_mult_f[0][12] ) );
  DFF_X1 \x_mult_f_reg[0][13]  ( .D(n8915), .CK(clk), .Q(\x_mult_f[0][13] ) );
  DFF_X1 \x_mult_f_reg[0][14]  ( .D(n8914), .CK(clk), .Q(\x_mult_f[0][14] ) );
  DFF_X1 \x_mult_f_reg[0][15]  ( .D(n8913), .CK(clk), .Q(\x_mult_f[0][15] ), 
        .QN(n8788) );
  DFF_X1 \x_mult_f_reg[1][0]  ( .D(n9329), .CK(clk), .Q(\x_mult_f[1][0] ) );
  DFF_X1 \x_mult_f_reg[1][1]  ( .D(n9328), .CK(clk), .Q(\x_mult_f[1][1] ) );
  DFF_X1 \x_mult_f_reg[1][2]  ( .D(n8940), .CK(clk), .Q(\x_mult_f[1][2] ) );
  DFF_X1 \x_mult_f_reg[1][3]  ( .D(n8939), .CK(clk), .Q(\x_mult_f[1][3] ) );
  DFF_X1 \x_mult_f_reg[1][4]  ( .D(n8938), .CK(clk), .Q(\x_mult_f[1][4] ) );
  DFF_X1 \x_mult_f_reg[1][5]  ( .D(n8937), .CK(clk), .Q(\x_mult_f[1][5] ) );
  DFF_X1 \x_mult_f_reg[1][6]  ( .D(n8936), .CK(clk), .Q(\x_mult_f[1][6] ) );
  DFF_X1 \x_mult_f_reg[1][7]  ( .D(n8935), .CK(clk), .Q(\x_mult_f[1][7] ) );
  DFF_X1 \x_mult_f_reg[1][8]  ( .D(n8934), .CK(clk), .Q(\x_mult_f[1][8] ) );
  DFF_X1 \x_mult_f_reg[1][9]  ( .D(n8933), .CK(clk), .Q(\x_mult_f[1][9] ) );
  DFF_X1 \x_mult_f_reg[1][10]  ( .D(n8932), .CK(clk), .Q(\x_mult_f[1][10] ) );
  DFF_X1 \x_mult_f_reg[1][11]  ( .D(n8931), .CK(clk), .Q(\x_mult_f[1][11] ) );
  DFF_X1 \x_mult_f_reg[1][12]  ( .D(n8930), .CK(clk), .Q(\x_mult_f[1][12] ) );
  DFF_X1 \x_mult_f_reg[1][13]  ( .D(n8929), .CK(clk), .Q(\x_mult_f[1][13] ) );
  DFF_X1 \x_mult_f_reg[1][14]  ( .D(n8928), .CK(clk), .Q(\x_mult_f[1][14] ) );
  DFF_X1 \x_mult_f_reg[1][15]  ( .D(n8927), .CK(clk), .Q(\x_mult_f[1][15] ), 
        .QN(n3476) );
  DFF_X1 \x_mult_f_reg[2][0]  ( .D(n9331), .CK(clk), .Q(\x_mult_f[2][0] ) );
  DFF_X1 \x_mult_f_reg[2][1]  ( .D(n9330), .CK(clk), .Q(\x_mult_f[2][1] ) );
  DFF_X1 \x_mult_f_reg[2][2]  ( .D(n8954), .CK(clk), .Q(\x_mult_f[2][2] ) );
  DFF_X1 \x_mult_f_reg[2][3]  ( .D(n8953), .CK(clk), .Q(\x_mult_f[2][3] ) );
  DFF_X1 \x_mult_f_reg[2][4]  ( .D(n8952), .CK(clk), .Q(\x_mult_f[2][4] ) );
  DFF_X1 \x_mult_f_reg[2][5]  ( .D(n8951), .CK(clk), .Q(\x_mult_f[2][5] ) );
  DFF_X1 \x_mult_f_reg[2][6]  ( .D(n8950), .CK(clk), .Q(\x_mult_f[2][6] ) );
  DFF_X1 \x_mult_f_reg[2][7]  ( .D(n8949), .CK(clk), .Q(\x_mult_f[2][7] ) );
  DFF_X1 \x_mult_f_reg[2][8]  ( .D(n8948), .CK(clk), .Q(\x_mult_f[2][8] ) );
  DFF_X1 \x_mult_f_reg[2][9]  ( .D(n8947), .CK(clk), .Q(\x_mult_f[2][9] ) );
  DFF_X1 \x_mult_f_reg[2][10]  ( .D(n8946), .CK(clk), .Q(\x_mult_f[2][10] ) );
  DFF_X1 \x_mult_f_reg[2][11]  ( .D(n8945), .CK(clk), .Q(\x_mult_f[2][11] ) );
  DFF_X1 \x_mult_f_reg[2][12]  ( .D(n8944), .CK(clk), .Q(\x_mult_f[2][12] ) );
  DFF_X1 \x_mult_f_reg[2][13]  ( .D(n8943), .CK(clk), .Q(\x_mult_f[2][13] ) );
  DFF_X1 \x_mult_f_reg[2][14]  ( .D(n8942), .CK(clk), .Q(\x_mult_f[2][14] ) );
  DFF_X1 \x_mult_f_reg[2][15]  ( .D(n8941), .CK(clk), .Q(\x_mult_f[2][15] ), 
        .QN(n8789) );
  DFF_X1 \x_mult_f_reg[3][2]  ( .D(n8968), .CK(clk), .Q(\x_mult_f[3][2] ) );
  DFF_X1 \x_mult_f_reg[3][3]  ( .D(n8967), .CK(clk), .Q(\x_mult_f[3][3] ) );
  DFF_X1 \x_mult_f_reg[3][4]  ( .D(n8966), .CK(clk), .Q(\x_mult_f[3][4] ) );
  DFF_X1 \x_mult_f_reg[3][5]  ( .D(n8965), .CK(clk), .Q(\x_mult_f[3][5] ) );
  DFF_X1 \x_mult_f_reg[3][6]  ( .D(n8964), .CK(clk), .Q(\x_mult_f[3][6] ) );
  DFF_X1 \x_mult_f_reg[3][7]  ( .D(n8963), .CK(clk), .Q(\x_mult_f[3][7] ) );
  DFF_X1 \x_mult_f_reg[3][8]  ( .D(n8962), .CK(clk), .Q(\x_mult_f[3][8] ) );
  DFF_X1 \x_mult_f_reg[3][9]  ( .D(n8961), .CK(clk), .Q(\x_mult_f[3][9] ) );
  DFF_X1 \x_mult_f_reg[3][10]  ( .D(n8960), .CK(clk), .Q(\x_mult_f[3][10] ) );
  DFF_X1 \x_mult_f_reg[3][11]  ( .D(n8959), .CK(clk), .Q(\x_mult_f[3][11] ) );
  DFF_X1 \x_mult_f_reg[3][12]  ( .D(n8958), .CK(clk), .Q(\x_mult_f[3][12] ) );
  DFF_X1 \x_mult_f_reg[3][13]  ( .D(n8957), .CK(clk), .Q(\x_mult_f[3][13] ) );
  DFF_X1 \x_mult_f_reg[3][14]  ( .D(n8956), .CK(clk), .Q(\x_mult_f[3][14] ) );
  DFF_X1 \x_mult_f_reg[3][15]  ( .D(n8955), .CK(clk), .Q(\x_mult_f[3][15] ), 
        .QN(n3471) );
  DFF_X1 \x_mult_f_reg[4][0]  ( .D(n9335), .CK(clk), .Q(\x_mult_f[4][0] ) );
  DFF_X1 \x_mult_f_reg[4][1]  ( .D(n9334), .CK(clk), .Q(\x_mult_f[4][1] ) );
  DFF_X1 \x_mult_f_reg[4][2]  ( .D(n8978), .CK(clk), .Q(\x_mult_f[4][2] ) );
  DFF_X1 \x_mult_f_reg[4][3]  ( .D(n8977), .CK(clk), .Q(\x_mult_f[4][3] ) );
  DFF_X1 \x_mult_f_reg[4][4]  ( .D(n8976), .CK(clk), .Q(\x_mult_f[4][4] ) );
  DFF_X1 \x_mult_f_reg[4][5]  ( .D(n8975), .CK(clk), .Q(\x_mult_f[4][5] ) );
  DFF_X1 \x_mult_f_reg[4][10]  ( .D(n8974), .CK(clk), .Q(\x_mult_f[4][10] ) );
  DFF_X1 \x_mult_f_reg[4][11]  ( .D(n8973), .CK(clk), .Q(\x_mult_f[4][11] ) );
  DFF_X1 \x_mult_f_reg[4][12]  ( .D(n8972), .CK(clk), .Q(\x_mult_f[4][12] ) );
  DFF_X1 \x_mult_f_reg[4][13]  ( .D(n8971), .CK(clk), .Q(\x_mult_f[4][13] ) );
  DFF_X1 \x_mult_f_reg[4][14]  ( .D(n8970), .CK(clk), .Q(\x_mult_f[4][14] ) );
  DFF_X1 \x_mult_f_reg[4][15]  ( .D(n8969), .CK(clk), .Q(\x_mult_f[4][15] ), 
        .QN(n3465) );
  DFF_X1 \x_mult_f_reg[5][0]  ( .D(n9337), .CK(clk), .Q(\x_mult_f[5][0] ) );
  DFF_X1 \x_mult_f_reg[5][1]  ( .D(n9336), .CK(clk), .Q(\x_mult_f[5][1] ) );
  DFF_X1 \x_mult_f_reg[5][2]  ( .D(n8983), .CK(clk), .Q(\x_mult_f[5][2] ) );
  DFF_X1 \x_mult_f_reg[5][3]  ( .D(n8982), .CK(clk), .Q(\x_mult_f[5][3] ) );
  DFF_X1 \x_mult_f_reg[5][4]  ( .D(n8981), .CK(clk), .Q(\x_mult_f[5][4] ) );
  DFF_X1 \x_mult_f_reg[5][5]  ( .D(n8980), .CK(clk), .Q(\x_mult_f[5][5] ) );
  DFF_X1 \x_mult_f_reg[5][13]  ( .D(n8979), .CK(clk), .Q(\x_mult_f[5][13] ) );
  DFF_X1 \x_mult_f_reg[6][0]  ( .D(n9339), .CK(clk), .Q(\x_mult_f[6][0] ) );
  DFF_X1 \x_mult_f_reg[6][1]  ( .D(n9338), .CK(clk), .Q(\x_mult_f[6][1] ) );
  DFF_X1 \x_mult_f_reg[6][2]  ( .D(n8997), .CK(clk), .Q(\x_mult_f[6][2] ) );
  DFF_X1 \x_mult_f_reg[6][3]  ( .D(n8996), .CK(clk), .Q(\x_mult_f[6][3] ) );
  DFF_X1 \x_mult_f_reg[6][4]  ( .D(n8995), .CK(clk), .Q(\x_mult_f[6][4] ) );
  DFF_X1 \x_mult_f_reg[6][5]  ( .D(n8994), .CK(clk), .Q(\x_mult_f[6][5] ) );
  DFF_X1 \x_mult_f_reg[6][6]  ( .D(n8993), .CK(clk), .Q(\x_mult_f[6][6] ) );
  DFF_X1 \x_mult_f_reg[6][7]  ( .D(n8992), .CK(clk), .Q(\x_mult_f[6][7] ) );
  DFF_X1 \x_mult_f_reg[6][8]  ( .D(n8991), .CK(clk), .Q(\x_mult_f[6][8] ) );
  DFF_X1 \x_mult_f_reg[6][9]  ( .D(n8990), .CK(clk), .Q(\x_mult_f[6][9] ) );
  DFF_X1 \x_mult_f_reg[6][10]  ( .D(n8989), .CK(clk), .Q(\x_mult_f[6][10] ) );
  DFF_X1 \x_mult_f_reg[6][11]  ( .D(n8988), .CK(clk), .Q(\x_mult_f[6][11] ) );
  DFF_X1 \x_mult_f_reg[6][12]  ( .D(n8987), .CK(clk), .Q(\x_mult_f[6][12] ) );
  DFF_X1 \x_mult_f_reg[6][13]  ( .D(n8986), .CK(clk), .Q(\x_mult_f[6][13] ) );
  DFF_X1 \x_mult_f_reg[6][14]  ( .D(n8985), .CK(clk), .Q(\x_mult_f[6][14] ) );
  DFF_X1 \x_mult_f_reg[6][15]  ( .D(n8984), .CK(clk), .Q(\x_mult_f[6][15] ), 
        .QN(n3455) );
  DFF_X1 \x_mult_f_reg[7][0]  ( .D(n9341), .CK(clk), .Q(\x_mult_f[7][0] ) );
  DFF_X1 \x_mult_f_reg[7][1]  ( .D(n9340), .CK(clk), .Q(\x_mult_f[7][1] ) );
  DFF_X1 \x_mult_f_reg[7][2]  ( .D(n9011), .CK(clk), .Q(\x_mult_f[7][2] ) );
  DFF_X1 \x_mult_f_reg[7][3]  ( .D(n9010), .CK(clk), .Q(\x_mult_f[7][3] ) );
  DFF_X1 \x_mult_f_reg[7][4]  ( .D(n9009), .CK(clk), .Q(\x_mult_f[7][4] ) );
  DFF_X1 \x_mult_f_reg[7][5]  ( .D(n9008), .CK(clk), .Q(\x_mult_f[7][5] ) );
  DFF_X1 \x_mult_f_reg[7][6]  ( .D(n9007), .CK(clk), .Q(\x_mult_f[7][6] ) );
  DFF_X1 \x_mult_f_reg[7][7]  ( .D(n9006), .CK(clk), .Q(\x_mult_f[7][7] ) );
  DFF_X1 \x_mult_f_reg[7][8]  ( .D(n9005), .CK(clk), .Q(\x_mult_f[7][8] ) );
  DFF_X1 \x_mult_f_reg[7][9]  ( .D(n9004), .CK(clk), .Q(\x_mult_f[7][9] ) );
  DFF_X1 \x_mult_f_reg[7][10]  ( .D(n9003), .CK(clk), .Q(\x_mult_f[7][10] ) );
  DFF_X1 \x_mult_f_reg[7][11]  ( .D(n9002), .CK(clk), .Q(\x_mult_f[7][11] ) );
  DFF_X1 \x_mult_f_reg[7][12]  ( .D(n9001), .CK(clk), .Q(\x_mult_f[7][12] ) );
  DFF_X1 \x_mult_f_reg[7][13]  ( .D(n9000), .CK(clk), .Q(\x_mult_f[7][13] ) );
  DFF_X1 \x_mult_f_reg[7][14]  ( .D(n8999), .CK(clk), .Q(\x_mult_f[7][14] ) );
  DFF_X1 \x_mult_f_reg[7][15]  ( .D(n8998), .CK(clk), .Q(\x_mult_f[7][15] ), 
        .QN(n3478) );
  DFF_X1 \x_mult_f_reg[8][0]  ( .D(n9343), .CK(clk), .Q(\x_mult_f[8][0] ) );
  DFF_X1 \x_mult_f_reg[8][1]  ( .D(n9342), .CK(clk), .Q(\x_mult_f[8][1] ) );
  DFF_X1 \x_mult_f_reg[8][2]  ( .D(n9025), .CK(clk), .Q(\x_mult_f[8][2] ) );
  DFF_X1 \x_mult_f_reg[8][3]  ( .D(n9024), .CK(clk), .Q(\x_mult_f[8][3] ) );
  DFF_X1 \x_mult_f_reg[8][4]  ( .D(n9023), .CK(clk), .Q(\x_mult_f[8][4] ) );
  DFF_X1 \x_mult_f_reg[8][5]  ( .D(n9022), .CK(clk), .Q(\x_mult_f[8][5] ) );
  DFF_X1 \x_mult_f_reg[8][6]  ( .D(n9021), .CK(clk), .Q(\x_mult_f[8][6] ) );
  DFF_X1 \x_mult_f_reg[8][7]  ( .D(n9020), .CK(clk), .Q(\x_mult_f[8][7] ) );
  DFF_X1 \x_mult_f_reg[8][8]  ( .D(n9019), .CK(clk), .Q(\x_mult_f[8][8] ) );
  DFF_X1 \x_mult_f_reg[8][9]  ( .D(n9018), .CK(clk), .Q(\x_mult_f[8][9] ) );
  DFF_X1 \x_mult_f_reg[8][10]  ( .D(n9017), .CK(clk), .Q(\x_mult_f[8][10] ) );
  DFF_X1 \x_mult_f_reg[8][11]  ( .D(n9016), .CK(clk), .Q(\x_mult_f[8][11] ) );
  DFF_X1 \x_mult_f_reg[8][12]  ( .D(n9015), .CK(clk), .Q(\x_mult_f[8][12] ) );
  DFF_X1 \x_mult_f_reg[8][13]  ( .D(n9014), .CK(clk), .Q(\x_mult_f[8][13] ) );
  DFF_X1 \x_mult_f_reg[8][14]  ( .D(n9013), .CK(clk), .Q(\x_mult_f[8][14] ) );
  DFF_X1 \x_mult_f_reg[8][15]  ( .D(n9012), .CK(clk), .Q(\x_mult_f[8][15] ), 
        .QN(n8791) );
  DFF_X1 \x_mult_f_reg[9][0]  ( .D(n9345), .CK(clk), .Q(\x_mult_f[9][0] ) );
  DFF_X1 \x_mult_f_reg[9][1]  ( .D(n9344), .CK(clk), .Q(\x_mult_f[9][1] ) );
  DFF_X1 \x_mult_f_reg[9][2]  ( .D(n9039), .CK(clk), .Q(\x_mult_f[9][2] ) );
  DFF_X1 \x_mult_f_reg[9][3]  ( .D(n9038), .CK(clk), .Q(\x_mult_f[9][3] ) );
  DFF_X1 \x_mult_f_reg[9][4]  ( .D(n9037), .CK(clk), .Q(\x_mult_f[9][4] ) );
  DFF_X1 \x_mult_f_reg[9][5]  ( .D(n9036), .CK(clk), .Q(\x_mult_f[9][5] ) );
  DFF_X1 \x_mult_f_reg[9][6]  ( .D(n9035), .CK(clk), .Q(\x_mult_f[9][6] ) );
  DFF_X1 \x_mult_f_reg[9][7]  ( .D(n9034), .CK(clk), .Q(\x_mult_f[9][7] ) );
  DFF_X1 \x_mult_f_reg[9][8]  ( .D(n9033), .CK(clk), .Q(\x_mult_f[9][8] ) );
  DFF_X1 \x_mult_f_reg[9][9]  ( .D(n9032), .CK(clk), .Q(\x_mult_f[9][9] ) );
  DFF_X1 \x_mult_f_reg[9][10]  ( .D(n9031), .CK(clk), .Q(\x_mult_f[9][10] ) );
  DFF_X1 \x_mult_f_reg[9][11]  ( .D(n9030), .CK(clk), .Q(\x_mult_f[9][11] ) );
  DFF_X1 \x_mult_f_reg[9][12]  ( .D(n9029), .CK(clk), .Q(\x_mult_f[9][12] ) );
  DFF_X1 \x_mult_f_reg[9][13]  ( .D(n9028), .CK(clk), .Q(\x_mult_f[9][13] ) );
  DFF_X1 \x_mult_f_reg[9][14]  ( .D(n9027), .CK(clk), .Q(\x_mult_f[9][14] ) );
  DFF_X1 \x_mult_f_reg[9][15]  ( .D(n9026), .CK(clk), .Q(\x_mult_f[9][15] ), 
        .QN(n8792) );
  DFF_X1 \x_mult_f_reg[10][0]  ( .D(n9347), .CK(clk), .Q(\x_mult_f[10][0] ) );
  DFF_X1 \x_mult_f_reg[10][1]  ( .D(n9346), .CK(clk), .Q(\x_mult_f[10][1] ) );
  DFF_X1 \x_mult_f_reg[10][2]  ( .D(n9053), .CK(clk), .Q(\x_mult_f[10][2] ) );
  DFF_X1 \x_mult_f_reg[10][3]  ( .D(n9052), .CK(clk), .Q(\x_mult_f[10][3] ) );
  DFF_X1 \x_mult_f_reg[10][4]  ( .D(n9051), .CK(clk), .Q(\x_mult_f[10][4] ) );
  DFF_X1 \x_mult_f_reg[10][5]  ( .D(n9050), .CK(clk), .Q(\x_mult_f[10][5] ) );
  DFF_X1 \x_mult_f_reg[10][6]  ( .D(n9049), .CK(clk), .Q(\x_mult_f[10][6] ) );
  DFF_X1 \x_mult_f_reg[10][7]  ( .D(n9048), .CK(clk), .Q(\x_mult_f[10][7] ) );
  DFF_X1 \x_mult_f_reg[10][8]  ( .D(n9047), .CK(clk), .Q(\x_mult_f[10][8] ) );
  DFF_X1 \x_mult_f_reg[10][9]  ( .D(n9046), .CK(clk), .Q(\x_mult_f[10][9] ) );
  DFF_X1 \x_mult_f_reg[10][10]  ( .D(n9045), .CK(clk), .Q(\x_mult_f[10][10] )
         );
  DFF_X1 \x_mult_f_reg[10][11]  ( .D(n9044), .CK(clk), .Q(\x_mult_f[10][11] )
         );
  DFF_X1 \x_mult_f_reg[10][12]  ( .D(n9043), .CK(clk), .Q(\x_mult_f[10][12] )
         );
  DFF_X1 \x_mult_f_reg[10][13]  ( .D(n9042), .CK(clk), .Q(\x_mult_f[10][13] )
         );
  DFF_X1 \x_mult_f_reg[10][14]  ( .D(n9041), .CK(clk), .Q(\x_mult_f[10][14] )
         );
  DFF_X1 \x_mult_f_reg[10][15]  ( .D(n9040), .CK(clk), .Q(\x_mult_f[10][15] ), 
        .QN(n3462) );
  DFF_X1 \x_mult_f_reg[11][0]  ( .D(n9349), .CK(clk), .Q(\x_mult_f[11][0] ) );
  DFF_X1 \x_mult_f_reg[11][1]  ( .D(n9348), .CK(clk), .Q(\x_mult_f[11][1] ) );
  DFF_X1 \x_mult_f_reg[11][2]  ( .D(n9066), .CK(clk), .Q(\x_mult_f[11][2] ) );
  DFF_X1 \x_mult_f_reg[11][3]  ( .D(n9065), .CK(clk), .Q(\x_mult_f[11][3] ) );
  DFF_X1 \x_mult_f_reg[11][4]  ( .D(n9064), .CK(clk), .Q(\x_mult_f[11][4] ) );
  DFF_X1 \x_mult_f_reg[11][5]  ( .D(n9063), .CK(clk), .Q(\x_mult_f[11][5] ) );
  DFF_X1 \x_mult_f_reg[11][6]  ( .D(n9062), .CK(clk), .Q(\x_mult_f[11][6] ) );
  DFF_X1 \x_mult_f_reg[11][7]  ( .D(n9061), .CK(clk), .Q(\x_mult_f[11][7] ) );
  DFF_X1 \x_mult_f_reg[11][8]  ( .D(n9060), .CK(clk), .Q(\x_mult_f[11][8] ) );
  DFF_X1 \x_mult_f_reg[11][9]  ( .D(n9059), .CK(clk), .Q(\x_mult_f[11][9] ) );
  DFF_X1 \x_mult_f_reg[11][10]  ( .D(n9058), .CK(clk), .Q(\x_mult_f[11][10] )
         );
  DFF_X1 \x_mult_f_reg[11][11]  ( .D(n9057), .CK(clk), .Q(\x_mult_f[11][11] )
         );
  DFF_X1 \x_mult_f_reg[11][12]  ( .D(n9056), .CK(clk), .Q(\x_mult_f[11][12] )
         );
  DFF_X1 \x_mult_f_reg[11][13]  ( .D(n9055), .CK(clk), .Q(\x_mult_f[11][13] )
         );
  DFF_X1 \x_mult_f_reg[11][14]  ( .D(n9054), .CK(clk), .Q(\x_mult_f[11][14] )
         );
  DFF_X1 \x_mult_f_reg[12][0]  ( .D(n9351), .CK(clk), .Q(\x_mult_f[12][0] ) );
  DFF_X1 \x_mult_f_reg[12][1]  ( .D(n9350), .CK(clk), .Q(\x_mult_f[12][1] ) );
  DFF_X1 \x_mult_f_reg[12][2]  ( .D(n9080), .CK(clk), .Q(\x_mult_f[12][2] ) );
  DFF_X1 \x_mult_f_reg[12][3]  ( .D(n9079), .CK(clk), .Q(\x_mult_f[12][3] ) );
  DFF_X1 \x_mult_f_reg[12][4]  ( .D(n9078), .CK(clk), .Q(\x_mult_f[12][4] ) );
  DFF_X1 \x_mult_f_reg[12][5]  ( .D(n9077), .CK(clk), .Q(\x_mult_f[12][5] ) );
  DFF_X1 \x_mult_f_reg[12][6]  ( .D(n9076), .CK(clk), .Q(\x_mult_f[12][6] ) );
  DFF_X1 \x_mult_f_reg[12][7]  ( .D(n9075), .CK(clk), .Q(\x_mult_f[12][7] ) );
  DFF_X1 \x_mult_f_reg[12][8]  ( .D(n9074), .CK(clk), .Q(\x_mult_f[12][8] ) );
  DFF_X1 \x_mult_f_reg[12][9]  ( .D(n9073), .CK(clk), .Q(\x_mult_f[12][9] ) );
  DFF_X1 \x_mult_f_reg[12][10]  ( .D(n9072), .CK(clk), .Q(\x_mult_f[12][10] )
         );
  DFF_X1 \x_mult_f_reg[12][11]  ( .D(n9071), .CK(clk), .Q(\x_mult_f[12][11] )
         );
  DFF_X1 \x_mult_f_reg[12][12]  ( .D(n9070), .CK(clk), .Q(\x_mult_f[12][12] )
         );
  DFF_X1 \x_mult_f_reg[12][13]  ( .D(n9069), .CK(clk), .Q(\x_mult_f[12][13] )
         );
  DFF_X1 \x_mult_f_reg[12][14]  ( .D(n9068), .CK(clk), .Q(\x_mult_f[12][14] )
         );
  DFF_X1 \x_mult_f_reg[12][15]  ( .D(n9067), .CK(clk), .Q(\x_mult_f[12][15] ), 
        .QN(n3447) );
  DFF_X1 \x_mult_f_reg[13][0]  ( .D(n9353), .CK(clk), .Q(\x_mult_f[13][0] ) );
  DFF_X1 \x_mult_f_reg[13][1]  ( .D(n9352), .CK(clk), .Q(\x_mult_f[13][1] ) );
  DFF_X1 \x_mult_f_reg[13][2]  ( .D(n9094), .CK(clk), .Q(\x_mult_f[13][2] ) );
  DFF_X1 \x_mult_f_reg[13][3]  ( .D(n9093), .CK(clk), .Q(\x_mult_f[13][3] ) );
  DFF_X1 \x_mult_f_reg[13][4]  ( .D(n9092), .CK(clk), .Q(\x_mult_f[13][4] ) );
  DFF_X1 \x_mult_f_reg[13][5]  ( .D(n9091), .CK(clk), .Q(\x_mult_f[13][5] ) );
  DFF_X1 \x_mult_f_reg[13][6]  ( .D(n9090), .CK(clk), .Q(\x_mult_f[13][6] ) );
  DFF_X1 \x_mult_f_reg[13][7]  ( .D(n9089), .CK(clk), .Q(\x_mult_f[13][7] ) );
  DFF_X1 \x_mult_f_reg[13][8]  ( .D(n9088), .CK(clk), .Q(\x_mult_f[13][8] ) );
  DFF_X1 \x_mult_f_reg[13][9]  ( .D(n9087), .CK(clk), .Q(\x_mult_f[13][9] ) );
  DFF_X1 \x_mult_f_reg[13][10]  ( .D(n9086), .CK(clk), .Q(\x_mult_f[13][10] )
         );
  DFF_X1 \x_mult_f_reg[13][11]  ( .D(n9085), .CK(clk), .Q(\x_mult_f[13][11] )
         );
  DFF_X1 \x_mult_f_reg[13][12]  ( .D(n9084), .CK(clk), .Q(\x_mult_f[13][12] )
         );
  DFF_X1 \x_mult_f_reg[13][13]  ( .D(n9083), .CK(clk), .Q(\x_mult_f[13][13] )
         );
  DFF_X1 \x_mult_f_reg[13][14]  ( .D(n9082), .CK(clk), .Q(\x_mult_f[13][14] )
         );
  DFF_X1 \x_mult_f_reg[13][15]  ( .D(n9081), .CK(clk), .Q(\x_mult_f[13][15] ), 
        .QN(n3466) );
  DFF_X1 \x_mult_f_reg[14][0]  ( .D(n9355), .CK(clk), .Q(\x_mult_f[14][0] ) );
  DFF_X1 \x_mult_f_reg[14][1]  ( .D(n9354), .CK(clk), .Q(\x_mult_f[14][1] ) );
  DFF_X1 \x_mult_f_reg[14][2]  ( .D(n9108), .CK(clk), .Q(\x_mult_f[14][2] ) );
  DFF_X1 \x_mult_f_reg[14][3]  ( .D(n9107), .CK(clk), .Q(\x_mult_f[14][3] ) );
  DFF_X1 \x_mult_f_reg[14][4]  ( .D(n9106), .CK(clk), .Q(\x_mult_f[14][4] ) );
  DFF_X1 \x_mult_f_reg[14][5]  ( .D(n9105), .CK(clk), .Q(\x_mult_f[14][5] ) );
  DFF_X1 \x_mult_f_reg[14][6]  ( .D(n9104), .CK(clk), .Q(\x_mult_f[14][6] ) );
  DFF_X1 \x_mult_f_reg[14][8]  ( .D(n9102), .CK(clk), .Q(\x_mult_f[14][8] ) );
  DFF_X1 \x_mult_f_reg[14][9]  ( .D(n9101), .CK(clk), .Q(\x_mult_f[14][9] ) );
  DFF_X1 \x_mult_f_reg[14][10]  ( .D(n9100), .CK(clk), .Q(\x_mult_f[14][10] )
         );
  DFF_X1 \x_mult_f_reg[14][11]  ( .D(n9099), .CK(clk), .Q(\x_mult_f[14][11] )
         );
  DFF_X1 \x_mult_f_reg[14][12]  ( .D(n9098), .CK(clk), .Q(\x_mult_f[14][12] )
         );
  DFF_X1 \x_mult_f_reg[14][13]  ( .D(n9097), .CK(clk), .Q(\x_mult_f[14][13] )
         );
  DFF_X1 \x_mult_f_reg[14][14]  ( .D(n9096), .CK(clk), .Q(\x_mult_f[14][14] )
         );
  DFF_X1 \x_mult_f_reg[14][15]  ( .D(n9095), .CK(clk), .Q(\x_mult_f[14][15] ), 
        .QN(n3450) );
  DFF_X1 \x_mult_f_reg[15][0]  ( .D(n9357), .CK(clk), .Q(\x_mult_f[15][0] ) );
  DFF_X1 \x_mult_f_reg[15][1]  ( .D(n9356), .CK(clk), .Q(\x_mult_f[15][1] ) );
  DFF_X1 \x_mult_f_reg[15][2]  ( .D(n9122), .CK(clk), .Q(\x_mult_f[15][2] ) );
  DFF_X1 \x_mult_f_reg[15][3]  ( .D(n9121), .CK(clk), .Q(\x_mult_f[15][3] ) );
  DFF_X1 \x_mult_f_reg[15][4]  ( .D(n9120), .CK(clk), .Q(\x_mult_f[15][4] ) );
  DFF_X1 \x_mult_f_reg[15][5]  ( .D(n9119), .CK(clk), .Q(\x_mult_f[15][5] ) );
  DFF_X1 \x_mult_f_reg[15][6]  ( .D(n9118), .CK(clk), .Q(\x_mult_f[15][6] ) );
  DFF_X1 \x_mult_f_reg[15][7]  ( .D(n9117), .CK(clk), .Q(\x_mult_f[15][7] ) );
  DFF_X1 \x_mult_f_reg[15][8]  ( .D(n9116), .CK(clk), .Q(\x_mult_f[15][8] ) );
  DFF_X1 \x_mult_f_reg[15][9]  ( .D(n9115), .CK(clk), .Q(\x_mult_f[15][9] ) );
  DFF_X1 \x_mult_f_reg[15][10]  ( .D(n9114), .CK(clk), .Q(\x_mult_f[15][10] )
         );
  DFF_X1 \x_mult_f_reg[15][11]  ( .D(n9113), .CK(clk), .Q(\x_mult_f[15][11] )
         );
  DFF_X1 \x_mult_f_reg[15][12]  ( .D(n9112), .CK(clk), .Q(\x_mult_f[15][12] )
         );
  DFF_X1 \x_mult_f_reg[15][13]  ( .D(n9111), .CK(clk), .Q(\x_mult_f[15][13] )
         );
  DFF_X1 \x_mult_f_reg[15][14]  ( .D(n9110), .CK(clk), .Q(\x_mult_f[15][14] )
         );
  DFF_X1 \x_mult_f_reg[15][15]  ( .D(n9109), .CK(clk), .Q(\x_mult_f[15][15] ), 
        .QN(n3469) );
  DFF_X1 \x_mult_f_reg[16][0]  ( .D(n9359), .CK(clk), .Q(\x_mult_f[16][0] ) );
  DFF_X1 \x_mult_f_reg[16][1]  ( .D(n9358), .CK(clk), .Q(\x_mult_f[16][1] ) );
  DFF_X1 \x_mult_f_reg[16][2]  ( .D(n9129), .CK(clk), .Q(\x_mult_f[16][2] ) );
  DFF_X1 \x_mult_f_reg[16][3]  ( .D(n9128), .CK(clk), .Q(\x_mult_f[16][3] ) );
  DFF_X1 \x_mult_f_reg[16][4]  ( .D(n9127), .CK(clk), .Q(\x_mult_f[16][4] ) );
  DFF_X1 \x_mult_f_reg[16][5]  ( .D(n9126), .CK(clk), .Q(\x_mult_f[16][5] ) );
  DFF_X1 \x_mult_f_reg[16][13]  ( .D(n9125), .CK(clk), .Q(\x_mult_f[16][13] )
         );
  DFF_X1 \x_mult_f_reg[16][14]  ( .D(n9124), .CK(clk), .Q(\x_mult_f[16][14] )
         );
  DFF_X1 \x_mult_f_reg[16][15]  ( .D(n9123), .CK(clk), .Q(\x_mult_f[16][15] ), 
        .QN(n3464) );
  DFF_X1 \x_mult_f_reg[17][0]  ( .D(n9361), .CK(clk), .Q(\x_mult_f[17][0] ) );
  DFF_X1 \x_mult_f_reg[17][1]  ( .D(n9360), .CK(clk), .Q(\x_mult_f[17][1] ) );
  DFF_X1 \x_mult_f_reg[17][2]  ( .D(n9139), .CK(clk), .Q(\x_mult_f[17][2] ) );
  DFF_X1 \x_mult_f_reg[17][3]  ( .D(n9138), .CK(clk), .Q(\x_mult_f[17][3] ) );
  DFF_X1 \x_mult_f_reg[17][4]  ( .D(n9137), .CK(clk), .Q(\x_mult_f[17][4] ) );
  DFF_X1 \x_mult_f_reg[17][6]  ( .D(n9135), .CK(clk), .Q(\x_mult_f[17][6] ) );
  DFF_X1 \x_mult_f_reg[17][7]  ( .D(n9134), .CK(clk), .Q(\x_mult_f[17][7] ) );
  DFF_X1 \x_mult_f_reg[17][8]  ( .D(n9133), .CK(clk), .Q(\x_mult_f[17][8] ) );
  DFF_X1 \x_mult_f_reg[17][9]  ( .D(n9132), .CK(clk), .Q(\x_mult_f[17][9] ) );
  DFF_X1 \x_mult_f_reg[17][10]  ( .D(n9131), .CK(clk), .Q(\x_mult_f[17][10] )
         );
  DFF_X1 \x_mult_f_reg[17][11]  ( .D(n9130), .CK(clk), .Q(\x_mult_f[17][11] )
         );
  DFF_X1 \x_mult_f_reg[18][0]  ( .D(n9363), .CK(clk), .Q(\x_mult_f[18][0] ) );
  DFF_X1 \x_mult_f_reg[18][1]  ( .D(n9362), .CK(clk), .Q(\x_mult_f[18][1] ) );
  DFF_X1 \x_mult_f_reg[18][2]  ( .D(n9153), .CK(clk), .Q(\x_mult_f[18][2] ) );
  DFF_X1 \x_mult_f_reg[18][3]  ( .D(n9152), .CK(clk), .Q(\x_mult_f[18][3] ), 
        .QN(n3415) );
  DFF_X1 \x_mult_f_reg[18][4]  ( .D(n9151), .CK(clk), .Q(\x_mult_f[18][4] ) );
  DFF_X1 \x_mult_f_reg[18][5]  ( .D(n9150), .CK(clk), .Q(\x_mult_f[18][5] ) );
  DFF_X1 \x_mult_f_reg[18][6]  ( .D(n9149), .CK(clk), .Q(\x_mult_f[18][6] ) );
  DFF_X1 \x_mult_f_reg[18][7]  ( .D(n9148), .CK(clk), .Q(\x_mult_f[18][7] ) );
  DFF_X1 \x_mult_f_reg[18][8]  ( .D(n9147), .CK(clk), .Q(\x_mult_f[18][8] ) );
  DFF_X1 \x_mult_f_reg[18][9]  ( .D(n9146), .CK(clk), .Q(\x_mult_f[18][9] ) );
  DFF_X1 \x_mult_f_reg[18][10]  ( .D(n9145), .CK(clk), .Q(\x_mult_f[18][10] )
         );
  DFF_X1 \x_mult_f_reg[18][11]  ( .D(n9144), .CK(clk), .Q(\x_mult_f[18][11] )
         );
  DFF_X1 \x_mult_f_reg[18][12]  ( .D(n9143), .CK(clk), .Q(\x_mult_f[18][12] )
         );
  DFF_X1 \x_mult_f_reg[18][13]  ( .D(n9142), .CK(clk), .Q(\x_mult_f[18][13] )
         );
  DFF_X1 \x_mult_f_reg[18][14]  ( .D(n9141), .CK(clk), .Q(\x_mult_f[18][14] )
         );
  DFF_X1 \x_mult_f_reg[18][15]  ( .D(n9140), .CK(clk), .Q(\x_mult_f[18][15] ), 
        .QN(n3461) );
  DFF_X1 \x_mult_f_reg[19][0]  ( .D(n9365), .CK(clk), .Q(\x_mult_f[19][0] ) );
  DFF_X1 \x_mult_f_reg[19][1]  ( .D(n9364), .CK(clk), .Q(\x_mult_f[19][1] ) );
  DFF_X1 \x_mult_f_reg[19][2]  ( .D(n9167), .CK(clk), .Q(\x_mult_f[19][2] ) );
  DFF_X1 \x_mult_f_reg[19][3]  ( .D(n9166), .CK(clk), .Q(\x_mult_f[19][3] ), 
        .QN(n3416) );
  DFF_X1 \x_mult_f_reg[19][4]  ( .D(n9165), .CK(clk), .Q(\x_mult_f[19][4] ) );
  DFF_X1 \x_mult_f_reg[19][5]  ( .D(n9164), .CK(clk), .Q(\x_mult_f[19][5] ) );
  DFF_X1 \x_mult_f_reg[19][6]  ( .D(n9163), .CK(clk), .Q(\x_mult_f[19][6] ) );
  DFF_X1 \x_mult_f_reg[19][7]  ( .D(n9162), .CK(clk), .Q(\x_mult_f[19][7] ) );
  DFF_X1 \x_mult_f_reg[19][8]  ( .D(n9161), .CK(clk), .Q(\x_mult_f[19][8] ) );
  DFF_X1 \x_mult_f_reg[19][9]  ( .D(n9160), .CK(clk), .Q(\x_mult_f[19][9] ) );
  DFF_X1 \x_mult_f_reg[19][10]  ( .D(n9159), .CK(clk), .Q(\x_mult_f[19][10] )
         );
  DFF_X1 \x_mult_f_reg[19][11]  ( .D(n9158), .CK(clk), .Q(\x_mult_f[19][11] )
         );
  DFF_X1 \x_mult_f_reg[19][12]  ( .D(n9157), .CK(clk), .Q(\x_mult_f[19][12] )
         );
  DFF_X1 \x_mult_f_reg[19][13]  ( .D(n9156), .CK(clk), .Q(\x_mult_f[19][13] )
         );
  DFF_X1 \x_mult_f_reg[19][14]  ( .D(n9155), .CK(clk), .Q(\x_mult_f[19][14] )
         );
  DFF_X1 \x_mult_f_reg[19][15]  ( .D(n9154), .CK(clk), .Q(\x_mult_f[19][15] ), 
        .QN(n8795) );
  DFF_X1 \x_mult_f_reg[20][0]  ( .D(n9367), .CK(clk), .Q(\x_mult_f[20][0] ) );
  DFF_X1 \x_mult_f_reg[20][1]  ( .D(n9366), .CK(clk), .Q(\x_mult_f[20][1] ) );
  DFF_X1 \x_mult_f_reg[20][2]  ( .D(n9181), .CK(clk), .Q(\x_mult_f[20][2] ) );
  DFF_X1 \x_mult_f_reg[20][3]  ( .D(n9180), .CK(clk), .Q(\x_mult_f[20][3] ) );
  DFF_X1 \x_mult_f_reg[20][4]  ( .D(n9179), .CK(clk), .Q(\x_mult_f[20][4] ) );
  DFF_X1 \x_mult_f_reg[20][5]  ( .D(n9178), .CK(clk), .Q(\x_mult_f[20][5] ) );
  DFF_X1 \x_mult_f_reg[20][6]  ( .D(n9177), .CK(clk), .Q(\x_mult_f[20][6] ) );
  DFF_X1 \x_mult_f_reg[20][7]  ( .D(n9176), .CK(clk), .Q(\x_mult_f[20][7] ) );
  DFF_X1 \x_mult_f_reg[20][8]  ( .D(n9175), .CK(clk), .Q(\x_mult_f[20][8] ) );
  DFF_X1 \x_mult_f_reg[20][9]  ( .D(n9174), .CK(clk), .Q(\x_mult_f[20][9] ) );
  DFF_X1 \x_mult_f_reg[20][10]  ( .D(n9173), .CK(clk), .Q(\x_mult_f[20][10] )
         );
  DFF_X1 \x_mult_f_reg[20][11]  ( .D(n9172), .CK(clk), .Q(\x_mult_f[20][11] )
         );
  DFF_X1 \x_mult_f_reg[20][12]  ( .D(n9171), .CK(clk), .Q(\x_mult_f[20][12] )
         );
  DFF_X1 \x_mult_f_reg[20][13]  ( .D(n9170), .CK(clk), .Q(\x_mult_f[20][13] )
         );
  DFF_X1 \x_mult_f_reg[20][14]  ( .D(n9169), .CK(clk), .Q(\x_mult_f[20][14] )
         );
  DFF_X1 \x_mult_f_reg[20][15]  ( .D(n9168), .CK(clk), .Q(\x_mult_f[20][15] ), 
        .QN(n8796) );
  DFF_X1 \x_mult_f_reg[21][0]  ( .D(n9369), .CK(clk), .Q(\x_mult_f[21][0] ) );
  DFF_X1 \x_mult_f_reg[21][1]  ( .D(n9368), .CK(clk), .Q(\x_mult_f[21][1] ) );
  DFF_X1 \x_mult_f_reg[21][2]  ( .D(n9195), .CK(clk), .Q(\x_mult_f[21][2] ) );
  DFF_X1 \x_mult_f_reg[21][3]  ( .D(n9194), .CK(clk), .Q(\x_mult_f[21][3] ) );
  DFF_X1 \x_mult_f_reg[21][4]  ( .D(n9193), .CK(clk), .Q(\x_mult_f[21][4] ) );
  DFF_X1 \x_mult_f_reg[21][5]  ( .D(n9192), .CK(clk), .Q(\x_mult_f[21][5] ) );
  DFF_X1 \x_mult_f_reg[21][6]  ( .D(n9191), .CK(clk), .Q(\x_mult_f[21][6] ) );
  DFF_X1 \x_mult_f_reg[21][7]  ( .D(n9190), .CK(clk), .Q(\x_mult_f[21][7] ) );
  DFF_X1 \x_mult_f_reg[21][8]  ( .D(n9189), .CK(clk), .Q(\x_mult_f[21][8] ) );
  DFF_X1 \x_mult_f_reg[21][9]  ( .D(n9188), .CK(clk), .Q(\x_mult_f[21][9] ) );
  DFF_X1 \x_mult_f_reg[21][10]  ( .D(n9187), .CK(clk), .Q(\x_mult_f[21][10] )
         );
  DFF_X1 \x_mult_f_reg[21][11]  ( .D(n9186), .CK(clk), .Q(\x_mult_f[21][11] )
         );
  DFF_X1 \x_mult_f_reg[21][12]  ( .D(n9185), .CK(clk), .Q(\x_mult_f[21][12] )
         );
  DFF_X1 \x_mult_f_reg[21][13]  ( .D(n9184), .CK(clk), .Q(\x_mult_f[21][13] )
         );
  DFF_X1 \x_mult_f_reg[21][14]  ( .D(n9183), .CK(clk), .Q(\x_mult_f[21][14] )
         );
  DFF_X1 \x_mult_f_reg[21][15]  ( .D(n9182), .CK(clk), .Q(\x_mult_f[21][15] ), 
        .QN(n3470) );
  DFF_X1 \x_mult_f_reg[22][0]  ( .D(n9371), .CK(clk), .Q(\x_mult_f[22][0] ) );
  DFF_X1 \x_mult_f_reg[22][1]  ( .D(n9370), .CK(clk), .Q(\x_mult_f[22][1] ) );
  DFF_X1 \x_mult_f_reg[22][2]  ( .D(n9209), .CK(clk), .Q(\x_mult_f[22][2] ) );
  DFF_X1 \x_mult_f_reg[22][3]  ( .D(n9208), .CK(clk), .Q(\x_mult_f[22][3] ) );
  DFF_X1 \x_mult_f_reg[22][4]  ( .D(n9207), .CK(clk), .Q(\x_mult_f[22][4] ) );
  DFF_X1 \x_mult_f_reg[22][5]  ( .D(n9206), .CK(clk), .Q(\x_mult_f[22][5] ) );
  DFF_X1 \x_mult_f_reg[22][6]  ( .D(n9205), .CK(clk), .Q(\x_mult_f[22][6] ) );
  DFF_X1 \x_mult_f_reg[22][7]  ( .D(n9204), .CK(clk), .Q(\x_mult_f[22][7] ) );
  DFF_X1 \x_mult_f_reg[22][8]  ( .D(n9203), .CK(clk), .Q(\x_mult_f[22][8] ) );
  DFF_X1 \x_mult_f_reg[22][9]  ( .D(n9202), .CK(clk), .Q(\x_mult_f[22][9] ) );
  DFF_X1 \x_mult_f_reg[22][10]  ( .D(n9201), .CK(clk), .Q(\x_mult_f[22][10] )
         );
  DFF_X1 \x_mult_f_reg[22][11]  ( .D(n9200), .CK(clk), .Q(\x_mult_f[22][11] )
         );
  DFF_X1 \x_mult_f_reg[22][12]  ( .D(n9199), .CK(clk), .Q(\x_mult_f[22][12] )
         );
  DFF_X1 \x_mult_f_reg[22][13]  ( .D(n9198), .CK(clk), .Q(\x_mult_f[22][13] )
         );
  DFF_X1 \x_mult_f_reg[22][14]  ( .D(n9197), .CK(clk), .Q(\x_mult_f[22][14] )
         );
  DFF_X1 \x_mult_f_reg[22][15]  ( .D(n9196), .CK(clk), .Q(\x_mult_f[22][15] ), 
        .QN(n3454) );
  DFF_X1 \x_mult_f_reg[23][0]  ( .D(n9373), .CK(clk), .Q(\x_mult_f[23][0] ) );
  DFF_X1 \x_mult_f_reg[23][1]  ( .D(n9372), .CK(clk), .Q(\x_mult_f[23][1] ) );
  DFF_X1 \x_mult_f_reg[23][2]  ( .D(n9223), .CK(clk), .Q(\x_mult_f[23][2] ) );
  DFF_X1 \x_mult_f_reg[23][4]  ( .D(n9221), .CK(clk), .Q(\x_mult_f[23][4] ) );
  DFF_X1 \x_mult_f_reg[23][5]  ( .D(n9220), .CK(clk), .Q(\x_mult_f[23][5] ) );
  DFF_X1 \x_mult_f_reg[23][6]  ( .D(n9219), .CK(clk), .Q(\x_mult_f[23][6] ) );
  DFF_X1 \x_mult_f_reg[23][7]  ( .D(n9218), .CK(clk), .Q(\x_mult_f[23][7] ) );
  DFF_X1 \x_mult_f_reg[23][8]  ( .D(n9217), .CK(clk), .Q(\x_mult_f[23][8] ) );
  DFF_X1 \x_mult_f_reg[23][9]  ( .D(n9216), .CK(clk), .Q(\x_mult_f[23][9] ) );
  DFF_X1 \x_mult_f_reg[23][10]  ( .D(n9215), .CK(clk), .Q(\x_mult_f[23][10] )
         );
  DFF_X1 \x_mult_f_reg[23][11]  ( .D(n9214), .CK(clk), .Q(\x_mult_f[23][11] )
         );
  DFF_X1 \x_mult_f_reg[23][12]  ( .D(n9213), .CK(clk), .Q(\x_mult_f[23][12] )
         );
  DFF_X1 \x_mult_f_reg[23][13]  ( .D(n9212), .CK(clk), .Q(\x_mult_f[23][13] )
         );
  DFF_X1 \x_mult_f_reg[23][14]  ( .D(n9211), .CK(clk), .Q(\x_mult_f[23][14] )
         );
  DFF_X1 \x_mult_f_reg[23][15]  ( .D(n9210), .CK(clk), .Q(\x_mult_f[23][15] ), 
        .QN(n3475) );
  DFF_X1 \x_mult_f_reg[24][0]  ( .D(n9375), .CK(clk), .Q(\x_mult_f[24][0] ) );
  DFF_X1 \x_mult_f_reg[24][1]  ( .D(n9374), .CK(clk), .Q(\x_mult_f[24][1] ) );
  DFF_X1 \x_mult_f_reg[24][2]  ( .D(n9229), .CK(clk), .Q(\x_mult_f[24][2] ) );
  DFF_X1 \x_mult_f_reg[24][3]  ( .D(n9228), .CK(clk), .Q(\x_mult_f[24][3] ) );
  DFF_X1 \x_mult_f_reg[24][4]  ( .D(n9227), .CK(clk), .Q(\x_mult_f[24][4] ) );
  DFF_X1 \x_mult_f_reg[24][5]  ( .D(n9226), .CK(clk), .Q(\x_mult_f[24][5] ) );
  DFF_X1 \x_mult_f_reg[24][6]  ( .D(n9225), .CK(clk), .Q(\x_mult_f[24][6] ) );
  DFF_X1 \x_mult_f_reg[24][12]  ( .D(n9224), .CK(clk), .Q(\x_mult_f[24][12] )
         );
  DFF_X1 \x_mult_f_reg[25][0]  ( .D(n9377), .CK(clk), .Q(\x_mult_f[25][0] ) );
  DFF_X1 \x_mult_f_reg[25][1]  ( .D(n9376), .CK(clk), .Q(\x_mult_f[25][1] ) );
  DFF_X1 \x_mult_f_reg[25][2]  ( .D(n9243), .CK(clk), .Q(\x_mult_f[25][2] ) );
  DFF_X1 \x_mult_f_reg[25][3]  ( .D(n9242), .CK(clk), .Q(\x_mult_f[25][3] ) );
  DFF_X1 \x_mult_f_reg[25][4]  ( .D(n9241), .CK(clk), .Q(\x_mult_f[25][4] ) );
  DFF_X1 \x_mult_f_reg[25][6]  ( .D(n9239), .CK(clk), .Q(\x_mult_f[25][6] ) );
  DFF_X1 \x_mult_f_reg[25][7]  ( .D(n9238), .CK(clk), .Q(\x_mult_f[25][7] ) );
  DFF_X1 \x_mult_f_reg[25][8]  ( .D(n9237), .CK(clk), .Q(\x_mult_f[25][8] ) );
  DFF_X1 \x_mult_f_reg[25][9]  ( .D(n9236), .CK(clk), .Q(\x_mult_f[25][9] ) );
  DFF_X1 \x_mult_f_reg[25][10]  ( .D(n9235), .CK(clk), .Q(\x_mult_f[25][10] )
         );
  DFF_X1 \x_mult_f_reg[25][11]  ( .D(n9234), .CK(clk), .Q(\x_mult_f[25][11] )
         );
  DFF_X1 \x_mult_f_reg[25][12]  ( .D(n9233), .CK(clk), .Q(\x_mult_f[25][12] )
         );
  DFF_X1 \x_mult_f_reg[25][13]  ( .D(n9232), .CK(clk), .Q(\x_mult_f[25][13] )
         );
  DFF_X1 \x_mult_f_reg[25][14]  ( .D(n9231), .CK(clk), .Q(\x_mult_f[25][14] )
         );
  DFF_X1 \x_mult_f_reg[25][15]  ( .D(n9230), .CK(clk), .Q(\x_mult_f[25][15] ), 
        .QN(n3479) );
  DFF_X1 \x_mult_f_reg[26][0]  ( .D(n9379), .CK(clk), .Q(\x_mult_f[26][0] ) );
  DFF_X1 \x_mult_f_reg[26][1]  ( .D(n9378), .CK(clk), .Q(\x_mult_f[26][1] ) );
  DFF_X1 \x_mult_f_reg[26][2]  ( .D(n9257), .CK(clk), .Q(\x_mult_f[26][2] ) );
  DFF_X1 \x_mult_f_reg[26][3]  ( .D(n9256), .CK(clk), .Q(\x_mult_f[26][3] ) );
  DFF_X1 \x_mult_f_reg[26][4]  ( .D(n9255), .CK(clk), .Q(\x_mult_f[26][4] ) );
  DFF_X1 \x_mult_f_reg[26][5]  ( .D(n9254), .CK(clk), .Q(\x_mult_f[26][5] ) );
  DFF_X1 \x_mult_f_reg[26][6]  ( .D(n9253), .CK(clk), .Q(\x_mult_f[26][6] ) );
  DFF_X1 \x_mult_f_reg[26][7]  ( .D(n9252), .CK(clk), .Q(\x_mult_f[26][7] ) );
  DFF_X1 \x_mult_f_reg[26][8]  ( .D(n9251), .CK(clk), .Q(\x_mult_f[26][8] ) );
  DFF_X1 \x_mult_f_reg[26][9]  ( .D(n9250), .CK(clk), .Q(\x_mult_f[26][9] ) );
  DFF_X1 \x_mult_f_reg[26][10]  ( .D(n9249), .CK(clk), .Q(\x_mult_f[26][10] )
         );
  DFF_X1 \x_mult_f_reg[26][11]  ( .D(n9248), .CK(clk), .Q(\x_mult_f[26][11] )
         );
  DFF_X1 \x_mult_f_reg[26][12]  ( .D(n9247), .CK(clk), .Q(\x_mult_f[26][12] )
         );
  DFF_X1 \x_mult_f_reg[26][13]  ( .D(n9246), .CK(clk), .Q(\x_mult_f[26][13] )
         );
  DFF_X1 \x_mult_f_reg[26][14]  ( .D(n9245), .CK(clk), .Q(\x_mult_f[26][14] )
         );
  DFF_X1 \x_mult_f_reg[26][15]  ( .D(n9244), .CK(clk), .Q(\x_mult_f[26][15] ), 
        .QN(n3448) );
  DFF_X1 \x_mult_f_reg[27][0]  ( .D(n9381), .CK(clk), .Q(\x_mult_f[27][0] ) );
  DFF_X1 \x_mult_f_reg[27][1]  ( .D(n9380), .CK(clk), .Q(\x_mult_f[27][1] ) );
  DFF_X1 \x_mult_f_reg[27][2]  ( .D(n9271), .CK(clk), .Q(\x_mult_f[27][2] ) );
  DFF_X1 \x_mult_f_reg[27][3]  ( .D(n9270), .CK(clk), .Q(\x_mult_f[27][3] ) );
  DFF_X1 \x_mult_f_reg[27][4]  ( .D(n9269), .CK(clk), .Q(\x_mult_f[27][4] ) );
  DFF_X1 \x_mult_f_reg[27][5]  ( .D(n9268), .CK(clk), .Q(\x_mult_f[27][5] ) );
  DFF_X1 \x_mult_f_reg[27][6]  ( .D(n9267), .CK(clk), .Q(\x_mult_f[27][6] ) );
  DFF_X1 \x_mult_f_reg[27][7]  ( .D(n9266), .CK(clk), .Q(\x_mult_f[27][7] ) );
  DFF_X1 \x_mult_f_reg[27][8]  ( .D(n9265), .CK(clk), .Q(\x_mult_f[27][8] ) );
  DFF_X1 \x_mult_f_reg[27][9]  ( .D(n9264), .CK(clk), .Q(\x_mult_f[27][9] ) );
  DFF_X1 \x_mult_f_reg[27][10]  ( .D(n9263), .CK(clk), .Q(\x_mult_f[27][10] )
         );
  DFF_X1 \x_mult_f_reg[27][11]  ( .D(n9262), .CK(clk), .Q(\x_mult_f[27][11] )
         );
  DFF_X1 \x_mult_f_reg[27][12]  ( .D(n9261), .CK(clk), .Q(\x_mult_f[27][12] )
         );
  DFF_X1 \x_mult_f_reg[27][13]  ( .D(n9260), .CK(clk), .Q(\x_mult_f[27][13] )
         );
  DFF_X1 \x_mult_f_reg[27][14]  ( .D(n9259), .CK(clk), .Q(\x_mult_f[27][14] )
         );
  DFF_X1 \x_mult_f_reg[27][15]  ( .D(n9258), .CK(clk), .Q(\x_mult_f[27][15] ), 
        .QN(n3467) );
  DFF_X1 \x_mult_f_reg[28][1]  ( .D(n9382), .CK(clk), .Q(\x_mult_f[28][1] ) );
  DFF_X1 \x_mult_f_reg[28][2]  ( .D(n9285), .CK(clk), .Q(\x_mult_f[28][2] ) );
  DFF_X1 \x_mult_f_reg[28][3]  ( .D(n9284), .CK(clk), .Q(\x_mult_f[28][3] ) );
  DFF_X1 \x_mult_f_reg[28][4]  ( .D(n9283), .CK(clk), .Q(\x_mult_f[28][4] ) );
  DFF_X1 \x_mult_f_reg[28][5]  ( .D(n9282), .CK(clk), .Q(\x_mult_f[28][5] ) );
  DFF_X1 \x_mult_f_reg[28][6]  ( .D(n9281), .CK(clk), .Q(\x_mult_f[28][6] ) );
  DFF_X1 \x_mult_f_reg[28][7]  ( .D(n9280), .CK(clk), .Q(\x_mult_f[28][7] ) );
  DFF_X1 \x_mult_f_reg[28][8]  ( .D(n9279), .CK(clk), .Q(\x_mult_f[28][8] ) );
  DFF_X1 \x_mult_f_reg[28][9]  ( .D(n9278), .CK(clk), .Q(\x_mult_f[28][9] ) );
  DFF_X1 \x_mult_f_reg[28][10]  ( .D(n9277), .CK(clk), .Q(\x_mult_f[28][10] )
         );
  DFF_X1 \x_mult_f_reg[28][11]  ( .D(n9276), .CK(clk), .Q(\x_mult_f[28][11] )
         );
  DFF_X1 \x_mult_f_reg[28][12]  ( .D(n9275), .CK(clk), .Q(\x_mult_f[28][12] )
         );
  DFF_X1 \x_mult_f_reg[28][13]  ( .D(n9274), .CK(clk), .Q(\x_mult_f[28][13] )
         );
  DFF_X1 \x_mult_f_reg[28][14]  ( .D(n9273), .CK(clk), .Q(\x_mult_f[28][14] )
         );
  DFF_X1 \x_mult_f_reg[28][15]  ( .D(n9272), .CK(clk), .Q(\x_mult_f[28][15] ), 
        .QN(n8798) );
  DFF_X1 \x_mult_f_reg[29][0]  ( .D(n9385), .CK(clk), .Q(\x_mult_f[29][0] ) );
  DFF_X1 \x_mult_f_reg[29][1]  ( .D(n9384), .CK(clk), .Q(\x_mult_f[29][1] ) );
  DFF_X1 \x_mult_f_reg[29][2]  ( .D(n9299), .CK(clk), .Q(\x_mult_f[29][2] ) );
  DFF_X1 \x_mult_f_reg[29][3]  ( .D(n9298), .CK(clk), .Q(\x_mult_f[29][3] ) );
  DFF_X1 \x_mult_f_reg[29][4]  ( .D(n9297), .CK(clk), .Q(\x_mult_f[29][4] ) );
  DFF_X1 \x_mult_f_reg[29][5]  ( .D(n9296), .CK(clk), .Q(\x_mult_f[29][5] ) );
  DFF_X1 \x_mult_f_reg[29][6]  ( .D(n9295), .CK(clk), .Q(\x_mult_f[29][6] ) );
  DFF_X1 \x_mult_f_reg[29][7]  ( .D(n9294), .CK(clk), .Q(\x_mult_f[29][7] ) );
  DFF_X1 \x_mult_f_reg[29][8]  ( .D(n9293), .CK(clk), .Q(\x_mult_f[29][8] ) );
  DFF_X1 \x_mult_f_reg[29][9]  ( .D(n9292), .CK(clk), .Q(\x_mult_f[29][9] ) );
  DFF_X1 \x_mult_f_reg[29][10]  ( .D(n9291), .CK(clk), .Q(\x_mult_f[29][10] )
         );
  DFF_X1 \x_mult_f_reg[29][11]  ( .D(n9290), .CK(clk), .Q(\x_mult_f[29][11] )
         );
  DFF_X1 \x_mult_f_reg[29][12]  ( .D(n9289), .CK(clk), .Q(\x_mult_f[29][12] )
         );
  DFF_X1 \x_mult_f_reg[29][13]  ( .D(n9288), .CK(clk), .Q(\x_mult_f[29][13] )
         );
  DFF_X1 \x_mult_f_reg[29][14]  ( .D(n9287), .CK(clk), .Q(\x_mult_f[29][14] )
         );
  DFF_X1 \x_mult_f_reg[29][15]  ( .D(n9286), .CK(clk), .Q(\x_mult_f[29][15] ), 
        .QN(n3477) );
  DFF_X1 \x_mult_f_reg[30][0]  ( .D(n9387), .CK(clk), .Q(\x_mult_f[30][0] ) );
  DFF_X1 \x_mult_f_reg[30][1]  ( .D(n9386), .CK(clk), .Q(\x_mult_f[30][1] ) );
  DFF_X1 \x_mult_f_reg[30][2]  ( .D(n9313), .CK(clk), .Q(\x_mult_f[30][2] ) );
  DFF_X1 \x_mult_f_reg[30][3]  ( .D(n9312), .CK(clk), .Q(\x_mult_f[30][3] ) );
  DFF_X1 \x_mult_f_reg[30][4]  ( .D(n9311), .CK(clk), .Q(\x_mult_f[30][4] ) );
  DFF_X1 \x_mult_f_reg[30][5]  ( .D(n9310), .CK(clk), .Q(\x_mult_f[30][5] ) );
  DFF_X1 \x_mult_f_reg[30][6]  ( .D(n9309), .CK(clk), .Q(\x_mult_f[30][6] ) );
  DFF_X1 \x_mult_f_reg[30][7]  ( .D(n9308), .CK(clk), .Q(\x_mult_f[30][7] ) );
  DFF_X1 \x_mult_f_reg[30][8]  ( .D(n9307), .CK(clk), .Q(\x_mult_f[30][8] ) );
  DFF_X1 \x_mult_f_reg[30][9]  ( .D(n9306), .CK(clk), .Q(\x_mult_f[30][9] ) );
  DFF_X1 \x_mult_f_reg[30][10]  ( .D(n9305), .CK(clk), .Q(\x_mult_f[30][10] )
         );
  DFF_X1 \x_mult_f_reg[30][11]  ( .D(n9304), .CK(clk), .Q(\x_mult_f[30][11] )
         );
  DFF_X1 \x_mult_f_reg[30][12]  ( .D(n9303), .CK(clk), .Q(\x_mult_f[30][12] )
         );
  DFF_X1 \x_mult_f_reg[30][13]  ( .D(n9302), .CK(clk), .Q(\x_mult_f[30][13] )
         );
  DFF_X1 \x_mult_f_reg[30][14]  ( .D(n9301), .CK(clk), .Q(\x_mult_f[30][14] )
         );
  DFF_X1 \x_mult_f_reg[30][15]  ( .D(n9300), .CK(clk), .Q(\x_mult_f[30][15] ), 
        .QN(n3449) );
  DFF_X1 \x_mult_f_reg[31][0]  ( .D(n9389), .CK(clk), .Q(\x_mult_f[31][0] ) );
  DFF_X1 \x_mult_f_reg[31][1]  ( .D(n9388), .CK(clk), .Q(\x_mult_f[31][1] ) );
  DFF_X1 \x_mult_f_reg[31][2]  ( .D(n9325), .CK(clk), .Q(\x_mult_f[31][2] ) );
  DFF_X1 \x_mult_f_reg[31][3]  ( .D(n9324), .CK(clk), .Q(\x_mult_f[31][3] ) );
  DFF_X1 \x_mult_f_reg[31][4]  ( .D(n9323), .CK(clk), .Q(\x_mult_f[31][4] ) );
  DFF_X1 \x_mult_f_reg[31][5]  ( .D(n9322), .CK(clk), .Q(\x_mult_f[31][5] ) );
  DFF_X1 \x_mult_f_reg[31][8]  ( .D(n9321), .CK(clk), .Q(\x_mult_f[31][8] ) );
  DFF_X1 \x_mult_f_reg[31][9]  ( .D(n9320), .CK(clk), .Q(\x_mult_f[31][9] ) );
  DFF_X1 \x_mult_f_reg[31][10]  ( .D(n9319), .CK(clk), .Q(\x_mult_f[31][10] )
         );
  DFF_X1 \x_mult_f_reg[31][11]  ( .D(n9318), .CK(clk), .Q(\x_mult_f[31][11] )
         );
  DFF_X1 \x_mult_f_reg[31][12]  ( .D(n9317), .CK(clk), .Q(\x_mult_f[31][12] )
         );
  DFF_X1 \x_mult_f_reg[31][13]  ( .D(n9316), .CK(clk), .Q(\x_mult_f[31][13] )
         );
  DFF_X1 \x_mult_f_reg[31][14]  ( .D(n9315), .CK(clk), .Q(\x_mult_f[31][14] )
         );
  DFF_X1 \x_mult_f_reg[31][15]  ( .D(n9314), .CK(clk), .Q(\x_mult_f[31][15] ), 
        .QN(n3468) );
  DFF_X1 \adder_stage1_reg[0][0]  ( .D(n10169), .CK(clk), .Q(
        \adder_stage1[0][0] ) );
  DFF_X1 \adder_stage1_reg[0][1]  ( .D(n10168), .CK(clk), .Q(
        \adder_stage1[0][1] ) );
  DFF_X1 \adder_stage1_reg[0][2]  ( .D(n10167), .CK(clk), .Q(
        \adder_stage1[0][2] ) );
  DFF_X1 \adder_stage1_reg[0][3]  ( .D(n10166), .CK(clk), .Q(
        \adder_stage1[0][3] ) );
  DFF_X1 \adder_stage1_reg[0][4]  ( .D(n10165), .CK(clk), .Q(
        \adder_stage1[0][4] ) );
  DFF_X1 \adder_stage1_reg[0][5]  ( .D(n10164), .CK(clk), .Q(
        \adder_stage1[0][5] ) );
  DFF_X1 \adder_stage1_reg[0][6]  ( .D(n10163), .CK(clk), .Q(
        \adder_stage1[0][6] ) );
  DFF_X1 \adder_stage1_reg[0][7]  ( .D(n10162), .CK(clk), .Q(
        \adder_stage1[0][7] ) );
  DFF_X1 \adder_stage1_reg[0][8]  ( .D(n10161), .CK(clk), .Q(
        \adder_stage1[0][8] ) );
  DFF_X1 \adder_stage1_reg[0][9]  ( .D(n10160), .CK(clk), .Q(
        \adder_stage1[0][9] ) );
  DFF_X1 \adder_stage1_reg[0][10]  ( .D(n10159), .CK(clk), .Q(
        \adder_stage1[0][10] ) );
  DFF_X1 \adder_stage1_reg[0][11]  ( .D(n10158), .CK(clk), .Q(
        \adder_stage1[0][11] ) );
  DFF_X1 \adder_stage1_reg[0][12]  ( .D(n10157), .CK(clk), .Q(
        \adder_stage1[0][12] ) );
  DFF_X1 \adder_stage1_reg[0][13]  ( .D(n10156), .CK(clk), .Q(
        \adder_stage1[0][13] ) );
  DFF_X1 \adder_stage1_reg[0][14]  ( .D(n10155), .CK(clk), .Q(
        \adder_stage1[0][14] ) );
  DFF_X1 \adder_stage1_reg[0][15]  ( .D(n10154), .CK(clk), .Q(
        \adder_stage1[0][15] ) );
  DFF_X1 \adder_stage1_reg[0][20]  ( .D(n10153), .CK(clk), .Q(
        \adder_stage1[0][20] ), .QN(n8799) );
  DFF_X1 \adder_stage1_reg[1][0]  ( .D(n10152), .CK(clk), .Q(
        \adder_stage1[1][0] ) );
  DFF_X1 \adder_stage1_reg[1][1]  ( .D(n10151), .CK(clk), .Q(
        \adder_stage1[1][1] ) );
  DFF_X1 \adder_stage1_reg[1][2]  ( .D(n10150), .CK(clk), .Q(
        \adder_stage1[1][2] ) );
  DFF_X1 \adder_stage1_reg[1][3]  ( .D(n10149), .CK(clk), .Q(
        \adder_stage1[1][3] ) );
  DFF_X1 \adder_stage1_reg[1][4]  ( .D(n10148), .CK(clk), .Q(
        \adder_stage1[1][4] ) );
  DFF_X1 \adder_stage1_reg[1][5]  ( .D(n10147), .CK(clk), .Q(
        \adder_stage1[1][5] ) );
  DFF_X1 \adder_stage1_reg[1][6]  ( .D(n10146), .CK(clk), .Q(
        \adder_stage1[1][6] ) );
  DFF_X1 \adder_stage1_reg[1][7]  ( .D(n10145), .CK(clk), .Q(
        \adder_stage1[1][7] ) );
  DFF_X1 \adder_stage1_reg[1][8]  ( .D(n10144), .CK(clk), .Q(
        \adder_stage1[1][8] ) );
  DFF_X1 \adder_stage1_reg[1][9]  ( .D(n10143), .CK(clk), .Q(
        \adder_stage1[1][9] ) );
  DFF_X1 \adder_stage1_reg[1][10]  ( .D(n10142), .CK(clk), .Q(
        \adder_stage1[1][10] ) );
  DFF_X1 \adder_stage1_reg[1][11]  ( .D(n10141), .CK(clk), .Q(
        \adder_stage1[1][11] ) );
  DFF_X1 \adder_stage1_reg[1][12]  ( .D(n10140), .CK(clk), .Q(
        \adder_stage1[1][12] ) );
  DFF_X1 \adder_stage1_reg[1][13]  ( .D(n10139), .CK(clk), .Q(
        \adder_stage1[1][13] ) );
  DFF_X1 \adder_stage1_reg[1][14]  ( .D(n10138), .CK(clk), .Q(
        \adder_stage1[1][14] ) );
  DFF_X1 \adder_stage1_reg[1][15]  ( .D(n10137), .CK(clk), .Q(
        \adder_stage1[1][15] ) );
  DFF_X1 \adder_stage1_reg[1][20]  ( .D(n10136), .CK(clk), .Q(
        \adder_stage1[1][20] ), .QN(n3481) );
  DFF_X1 \adder_stage1_reg[2][0]  ( .D(n10135), .CK(clk), .Q(
        \adder_stage1[2][0] ), .QN(n3423) );
  DFF_X1 \adder_stage1_reg[2][1]  ( .D(n10134), .CK(clk), .Q(
        \adder_stage1[2][1] ) );
  DFF_X1 \adder_stage1_reg[2][2]  ( .D(n10133), .CK(clk), .Q(
        \adder_stage1[2][2] ) );
  DFF_X1 \adder_stage1_reg[2][3]  ( .D(n10132), .CK(clk), .Q(
        \adder_stage1[2][3] ) );
  DFF_X1 \adder_stage1_reg[2][4]  ( .D(n10131), .CK(clk), .Q(
        \adder_stage1[2][4] ) );
  DFF_X1 \adder_stage1_reg[2][5]  ( .D(n10130), .CK(clk), .Q(
        \adder_stage1[2][5] ) );
  DFF_X1 \adder_stage1_reg[2][6]  ( .D(n10129), .CK(clk), .Q(
        \adder_stage1[2][6] ) );
  DFF_X1 \adder_stage1_reg[2][7]  ( .D(n10128), .CK(clk), .Q(
        \adder_stage1[2][7] ) );
  DFF_X1 \adder_stage1_reg[2][8]  ( .D(n10127), .CK(clk), .Q(
        \adder_stage1[2][8] ), .QN(n3484) );
  DFF_X1 \adder_stage1_reg[2][9]  ( .D(n10126), .CK(clk), .Q(
        \adder_stage1[2][9] ) );
  DFF_X1 \adder_stage1_reg[2][10]  ( .D(n10125), .CK(clk), .Q(
        \adder_stage1[2][10] ) );
  DFF_X1 \adder_stage1_reg[2][11]  ( .D(n10124), .CK(clk), .Q(
        \adder_stage1[2][11] ) );
  DFF_X1 \adder_stage1_reg[2][12]  ( .D(n10123), .CK(clk), .Q(
        \adder_stage1[2][12] ) );
  DFF_X1 \adder_stage1_reg[2][14]  ( .D(n10122), .CK(clk), .Q(
        \adder_stage1[2][14] ) );
  DFF_X1 \adder_stage1_reg[2][15]  ( .D(n10121), .CK(clk), .Q(
        \adder_stage1[2][15] ), .QN(n3460) );
  DFF_X1 \adder_stage1_reg[3][0]  ( .D(n10120), .CK(clk), .Q(
        \adder_stage1[3][0] ), .QN(n3424) );
  DFF_X1 \adder_stage1_reg[3][1]  ( .D(n10119), .CK(clk), .Q(
        \adder_stage1[3][1] ) );
  DFF_X1 \adder_stage1_reg[3][2]  ( .D(n10118), .CK(clk), .Q(
        \adder_stage1[3][2] ) );
  DFF_X1 \adder_stage1_reg[3][3]  ( .D(n10117), .CK(clk), .Q(
        \adder_stage1[3][3] ) );
  DFF_X1 \adder_stage1_reg[3][4]  ( .D(n10116), .CK(clk), .Q(
        \adder_stage1[3][4] ) );
  DFF_X1 \adder_stage1_reg[3][5]  ( .D(n10115), .CK(clk), .Q(
        \adder_stage1[3][5] ) );
  DFF_X1 \adder_stage1_reg[3][6]  ( .D(n10114), .CK(clk), .Q(
        \adder_stage1[3][6] ) );
  DFF_X1 \adder_stage1_reg[3][7]  ( .D(n10113), .CK(clk), .Q(
        \adder_stage1[3][7] ) );
  DFF_X1 \adder_stage1_reg[3][8]  ( .D(n10112), .CK(clk), .Q(
        \adder_stage1[3][8] ), .QN(n3457) );
  DFF_X1 \adder_stage1_reg[3][9]  ( .D(n10111), .CK(clk), .Q(
        \adder_stage1[3][9] ) );
  DFF_X1 \adder_stage1_reg[3][10]  ( .D(n10110), .CK(clk), .Q(
        \adder_stage1[3][10] ) );
  DFF_X1 \adder_stage1_reg[3][11]  ( .D(n10109), .CK(clk), .Q(
        \adder_stage1[3][11] ) );
  DFF_X1 \adder_stage1_reg[3][12]  ( .D(n10108), .CK(clk), .Q(
        \adder_stage1[3][12] ) );
  DFF_X1 \adder_stage1_reg[3][13]  ( .D(n10107), .CK(clk), .Q(
        \adder_stage1[3][13] ) );
  DFF_X1 \adder_stage1_reg[3][14]  ( .D(n10106), .CK(clk), .Q(
        \adder_stage1[3][14] ) );
  DFF_X1 \adder_stage1_reg[3][15]  ( .D(n10105), .CK(clk), .Q(
        \adder_stage1[3][15] ) );
  DFF_X1 \adder_stage1_reg[3][20]  ( .D(n10104), .CK(clk), .Q(
        \adder_stage1[3][20] ), .QN(n3480) );
  DFF_X1 \adder_stage1_reg[4][0]  ( .D(n10103), .CK(clk), .Q(
        \adder_stage1[4][0] ) );
  DFF_X1 \adder_stage1_reg[4][1]  ( .D(n10102), .CK(clk), .Q(
        \adder_stage1[4][1] ) );
  DFF_X1 \adder_stage1_reg[4][2]  ( .D(n10101), .CK(clk), .Q(
        \adder_stage1[4][2] ) );
  DFF_X1 \adder_stage1_reg[4][3]  ( .D(n10100), .CK(clk), .Q(
        \adder_stage1[4][3] ) );
  DFF_X1 \adder_stage1_reg[4][4]  ( .D(n10099), .CK(clk), .Q(
        \adder_stage1[4][4] ) );
  DFF_X1 \adder_stage1_reg[4][5]  ( .D(n10098), .CK(clk), .Q(
        \adder_stage1[4][5] ) );
  DFF_X1 \adder_stage1_reg[4][6]  ( .D(n10097), .CK(clk), .Q(
        \adder_stage1[4][6] ) );
  DFF_X1 \adder_stage1_reg[4][7]  ( .D(n10096), .CK(clk), .Q(
        \adder_stage1[4][7] ) );
  DFF_X1 \adder_stage1_reg[4][8]  ( .D(n10095), .CK(clk), .Q(
        \adder_stage1[4][8] ) );
  DFF_X1 \adder_stage1_reg[4][9]  ( .D(n10094), .CK(clk), .Q(
        \adder_stage1[4][9] ) );
  DFF_X1 \adder_stage1_reg[4][10]  ( .D(n10093), .CK(clk), .Q(
        \adder_stage1[4][10] ) );
  DFF_X1 \adder_stage1_reg[4][11]  ( .D(n10092), .CK(clk), .Q(
        \adder_stage1[4][11] ) );
  DFF_X1 \adder_stage1_reg[4][12]  ( .D(n10091), .CK(clk), .Q(
        \adder_stage1[4][12] ) );
  DFF_X1 \adder_stage1_reg[4][13]  ( .D(n10090), .CK(clk), .Q(
        \adder_stage1[4][13] ) );
  DFF_X1 \adder_stage1_reg[4][14]  ( .D(n10089), .CK(clk), .Q(
        \adder_stage1[4][14] ) );
  DFF_X1 \adder_stage1_reg[4][15]  ( .D(n10088), .CK(clk), .Q(
        \adder_stage1[4][15] ) );
  DFF_X1 \adder_stage1_reg[4][20]  ( .D(n10087), .CK(clk), .Q(
        \adder_stage1[4][20] ), .QN(n8801) );
  DFF_X1 \adder_stage1_reg[5][0]  ( .D(n10086), .CK(clk), .Q(
        \adder_stage1[5][0] ) );
  DFF_X1 \adder_stage1_reg[5][1]  ( .D(n10085), .CK(clk), .Q(
        \adder_stage1[5][1] ) );
  DFF_X1 \adder_stage1_reg[5][2]  ( .D(n10084), .CK(clk), .Q(
        \adder_stage1[5][2] ) );
  DFF_X1 \adder_stage1_reg[5][3]  ( .D(n10083), .CK(clk), .Q(
        \adder_stage1[5][3] ) );
  DFF_X1 \adder_stage1_reg[5][4]  ( .D(n10082), .CK(clk), .Q(
        \adder_stage1[5][4] ) );
  DFF_X1 \adder_stage1_reg[5][5]  ( .D(n10081), .CK(clk), .Q(
        \adder_stage1[5][5] ) );
  DFF_X1 \adder_stage1_reg[5][6]  ( .D(n10080), .CK(clk), .Q(
        \adder_stage1[5][6] ) );
  DFF_X1 \adder_stage1_reg[5][7]  ( .D(n10079), .CK(clk), .Q(
        \adder_stage1[5][7] ) );
  DFF_X1 \adder_stage1_reg[5][8]  ( .D(n10078), .CK(clk), .Q(
        \adder_stage1[5][8] ) );
  DFF_X1 \adder_stage1_reg[5][9]  ( .D(n10077), .CK(clk), .Q(
        \adder_stage1[5][9] ) );
  DFF_X1 \adder_stage1_reg[5][10]  ( .D(n10076), .CK(clk), .Q(
        \adder_stage1[5][10] ) );
  DFF_X1 \adder_stage1_reg[5][11]  ( .D(n10075), .CK(clk), .Q(
        \adder_stage1[5][11] ) );
  DFF_X1 \adder_stage1_reg[5][12]  ( .D(n10074), .CK(clk), .Q(
        \adder_stage1[5][12] ) );
  DFF_X1 \adder_stage1_reg[5][13]  ( .D(n10073), .CK(clk), .Q(
        \adder_stage1[5][13] ) );
  DFF_X1 \adder_stage1_reg[5][14]  ( .D(n10072), .CK(clk), .Q(
        \adder_stage1[5][14] ) );
  DFF_X1 \adder_stage1_reg[5][20]  ( .D(n10071), .CK(clk), .Q(
        \adder_stage1[5][20] ), .QN(n8802) );
  DFF_X1 \adder_stage1_reg[6][0]  ( .D(n10070), .CK(clk), .Q(
        \adder_stage1[6][0] ) );
  DFF_X1 \adder_stage1_reg[6][1]  ( .D(n10069), .CK(clk), .Q(
        \adder_stage1[6][1] ) );
  DFF_X1 \adder_stage1_reg[6][2]  ( .D(n10068), .CK(clk), .Q(
        \adder_stage1[6][2] ) );
  DFF_X1 \adder_stage1_reg[6][3]  ( .D(n10067), .CK(clk), .Q(
        \adder_stage1[6][3] ) );
  DFF_X1 \adder_stage1_reg[6][4]  ( .D(n10066), .CK(clk), .Q(
        \adder_stage1[6][4] ) );
  DFF_X1 \adder_stage1_reg[6][5]  ( .D(n10065), .CK(clk), .Q(
        \adder_stage1[6][5] ) );
  DFF_X1 \adder_stage1_reg[6][6]  ( .D(n10064), .CK(clk), .Q(
        \adder_stage1[6][6] ) );
  DFF_X1 \adder_stage1_reg[6][7]  ( .D(n10063), .CK(clk), .Q(
        \adder_stage1[6][7] ) );
  DFF_X1 \adder_stage1_reg[6][8]  ( .D(n10062), .CK(clk), .Q(
        \adder_stage1[6][8] ) );
  DFF_X1 \adder_stage1_reg[6][9]  ( .D(n10061), .CK(clk), .Q(
        \adder_stage1[6][9] ), .QN(n3458) );
  DFF_X1 \adder_stage1_reg[6][10]  ( .D(n10060), .CK(clk), .Q(
        \adder_stage1[6][10] ) );
  DFF_X1 \adder_stage1_reg[6][11]  ( .D(n10059), .CK(clk), .Q(
        \adder_stage1[6][11] ) );
  DFF_X1 \adder_stage1_reg[6][12]  ( .D(n10058), .CK(clk), .Q(
        \adder_stage1[6][12] ) );
  DFF_X1 \adder_stage1_reg[6][13]  ( .D(n10057), .CK(clk), .Q(
        \adder_stage1[6][13] ) );
  DFF_X1 \adder_stage1_reg[6][14]  ( .D(n10056), .CK(clk), .Q(
        \adder_stage1[6][14] ) );
  DFF_X1 \adder_stage1_reg[6][15]  ( .D(n10055), .CK(clk), .Q(
        \adder_stage1[6][15] ) );
  DFF_X1 \adder_stage1_reg[6][20]  ( .D(n10054), .CK(clk), .Q(
        \adder_stage1[6][20] ), .QN(n3451) );
  DFF_X1 \adder_stage1_reg[7][0]  ( .D(n10053), .CK(clk), .Q(
        \adder_stage1[7][0] ) );
  DFF_X1 \adder_stage1_reg[7][1]  ( .D(n10052), .CK(clk), .Q(
        \adder_stage1[7][1] ) );
  DFF_X1 \adder_stage1_reg[7][2]  ( .D(n10051), .CK(clk), .Q(
        \adder_stage1[7][2] ) );
  DFF_X1 \adder_stage1_reg[7][3]  ( .D(n10050), .CK(clk), .Q(
        \adder_stage1[7][3] ) );
  DFF_X1 \adder_stage1_reg[7][4]  ( .D(n10049), .CK(clk), .Q(
        \adder_stage1[7][4] ) );
  DFF_X1 \adder_stage1_reg[7][5]  ( .D(n10048), .CK(clk), .Q(
        \adder_stage1[7][5] ) );
  DFF_X1 \adder_stage1_reg[7][6]  ( .D(n10047), .CK(clk), .Q(
        \adder_stage1[7][6] ) );
  DFF_X1 \adder_stage1_reg[7][7]  ( .D(n10046), .CK(clk), .Q(
        \adder_stage1[7][7] ) );
  DFF_X1 \adder_stage1_reg[7][8]  ( .D(n10045), .CK(clk), .Q(
        \adder_stage1[7][8] ) );
  DFF_X1 \adder_stage1_reg[7][9]  ( .D(n10044), .CK(clk), .Q(
        \adder_stage1[7][9] ), .QN(n3485) );
  DFF_X1 \adder_stage1_reg[7][10]  ( .D(n10043), .CK(clk), .Q(
        \adder_stage1[7][10] ) );
  DFF_X1 \adder_stage1_reg[7][11]  ( .D(n10042), .CK(clk), .Q(
        \adder_stage1[7][11] ) );
  DFF_X1 \adder_stage1_reg[7][12]  ( .D(n10041), .CK(clk), .Q(
        \adder_stage1[7][12] ) );
  DFF_X1 \adder_stage1_reg[7][13]  ( .D(n10040), .CK(clk), .Q(
        \adder_stage1[7][13] ) );
  DFF_X1 \adder_stage1_reg[7][14]  ( .D(n10039), .CK(clk), .Q(
        \adder_stage1[7][14] ) );
  DFF_X1 \adder_stage1_reg[7][15]  ( .D(n10038), .CK(clk), .Q(
        \adder_stage1[7][15] ) );
  DFF_X1 \adder_stage1_reg[7][20]  ( .D(n10037), .CK(clk), .Q(
        \adder_stage1[7][20] ), .QN(n3472) );
  DFF_X1 \adder_stage1_reg[8][0]  ( .D(n10036), .CK(clk), .Q(
        \adder_stage1[8][0] ) );
  DFF_X1 \adder_stage1_reg[8][1]  ( .D(n10035), .CK(clk), .Q(
        \adder_stage1[8][1] ) );
  DFF_X1 \adder_stage1_reg[8][2]  ( .D(n10034), .CK(clk), .Q(
        \adder_stage1[8][2] ) );
  DFF_X1 \adder_stage1_reg[8][3]  ( .D(n10033), .CK(clk), .Q(
        \adder_stage1[8][3] ) );
  DFF_X1 \adder_stage1_reg[8][4]  ( .D(n10032), .CK(clk), .Q(
        \adder_stage1[8][4] ) );
  DFF_X1 \adder_stage1_reg[8][5]  ( .D(n10031), .CK(clk), .Q(
        \adder_stage1[8][5] ) );
  DFF_X1 \adder_stage1_reg[8][6]  ( .D(n10030), .CK(clk), .Q(
        \adder_stage1[8][6] ) );
  DFF_X1 \adder_stage1_reg[8][7]  ( .D(n10029), .CK(clk), .Q(
        \adder_stage1[8][7] ) );
  DFF_X1 \adder_stage1_reg[8][8]  ( .D(n10028), .CK(clk), .Q(
        \adder_stage1[8][8] ) );
  DFF_X1 \adder_stage1_reg[8][9]  ( .D(n10027), .CK(clk), .Q(
        \adder_stage1[8][9] ) );
  DFF_X1 \adder_stage1_reg[8][10]  ( .D(n10026), .CK(clk), .Q(
        \adder_stage1[8][10] ) );
  DFF_X1 \adder_stage1_reg[8][11]  ( .D(n10025), .CK(clk), .Q(
        \adder_stage1[8][11] ) );
  DFF_X1 \adder_stage1_reg[8][12]  ( .D(n10024), .CK(clk), .Q(
        \adder_stage1[8][12] ) );
  DFF_X1 \adder_stage1_reg[8][13]  ( .D(n10023), .CK(clk), .Q(
        \adder_stage1[8][13] ) );
  DFF_X1 \adder_stage1_reg[8][14]  ( .D(n10022), .CK(clk), .Q(
        \adder_stage1[8][14] ) );
  DFF_X1 \adder_stage1_reg[8][15]  ( .D(n10021), .CK(clk), .Q(
        \adder_stage1[8][15] ) );
  DFF_X1 \adder_stage1_reg[8][20]  ( .D(n10020), .CK(clk), .Q(
        \adder_stage1[8][20] ), .QN(n3463) );
  DFF_X1 \adder_stage1_reg[9][0]  ( .D(n10019), .CK(clk), .Q(
        \adder_stage1[9][0] ) );
  DFF_X1 \adder_stage1_reg[9][1]  ( .D(n10018), .CK(clk), .Q(
        \adder_stage1[9][1] ) );
  DFF_X1 \adder_stage1_reg[9][2]  ( .D(n10017), .CK(clk), .Q(
        \adder_stage1[9][2] ) );
  DFF_X1 \adder_stage1_reg[9][3]  ( .D(n10016), .CK(clk), .Q(
        \adder_stage1[9][3] ) );
  DFF_X1 \adder_stage1_reg[9][4]  ( .D(n10015), .CK(clk), .Q(
        \adder_stage1[9][4] ) );
  DFF_X1 \adder_stage1_reg[9][5]  ( .D(n10014), .CK(clk), .Q(
        \adder_stage1[9][5] ) );
  DFF_X1 \adder_stage1_reg[9][6]  ( .D(n10013), .CK(clk), .Q(
        \adder_stage1[9][6] ) );
  DFF_X1 \adder_stage1_reg[9][7]  ( .D(n10012), .CK(clk), .Q(
        \adder_stage1[9][7] ) );
  DFF_X1 \adder_stage1_reg[9][8]  ( .D(n10011), .CK(clk), .Q(
        \adder_stage1[9][8] ) );
  DFF_X1 \adder_stage1_reg[9][9]  ( .D(n10010), .CK(clk), .Q(
        \adder_stage1[9][9] ) );
  DFF_X1 \adder_stage1_reg[9][10]  ( .D(n10009), .CK(clk), .Q(
        \adder_stage1[9][10] ) );
  DFF_X1 \adder_stage1_reg[9][11]  ( .D(n10008), .CK(clk), .Q(
        \adder_stage1[9][11] ) );
  DFF_X1 \adder_stage1_reg[9][12]  ( .D(n10007), .CK(clk), .Q(
        \adder_stage1[9][12] ) );
  DFF_X1 \adder_stage1_reg[9][13]  ( .D(n10006), .CK(clk), .Q(
        \adder_stage1[9][13] ) );
  DFF_X1 \adder_stage1_reg[9][14]  ( .D(n10005), .CK(clk), .Q(
        \adder_stage1[9][14] ) );
  DFF_X1 \adder_stage1_reg[9][15]  ( .D(n10004), .CK(clk), .Q(
        \adder_stage1[9][15] ) );
  DFF_X1 \adder_stage1_reg[9][20]  ( .D(n10003), .CK(clk), .Q(
        \adder_stage1[9][20] ), .QN(n8803) );
  DFF_X1 \adder_stage1_reg[10][0]  ( .D(n10002), .CK(clk), .Q(
        \adder_stage1[10][0] ) );
  DFF_X1 \adder_stage1_reg[10][1]  ( .D(n10001), .CK(clk), .Q(
        \adder_stage1[10][1] ) );
  DFF_X1 \adder_stage1_reg[10][2]  ( .D(n10000), .CK(clk), .Q(
        \adder_stage1[10][2] ) );
  DFF_X1 \adder_stage1_reg[10][4]  ( .D(n9999), .CK(clk), .Q(
        \adder_stage1[10][4] ) );
  DFF_X1 \adder_stage1_reg[10][5]  ( .D(n9998), .CK(clk), .Q(
        \adder_stage1[10][5] ) );
  DFF_X1 \adder_stage1_reg[10][6]  ( .D(n9997), .CK(clk), .Q(
        \adder_stage1[10][6] ) );
  DFF_X1 \adder_stage1_reg[10][7]  ( .D(n9996), .CK(clk), .Q(
        \adder_stage1[10][7] ) );
  DFF_X1 \adder_stage1_reg[10][8]  ( .D(n9995), .CK(clk), .Q(
        \adder_stage1[10][8] ) );
  DFF_X1 \adder_stage1_reg[10][9]  ( .D(n9994), .CK(clk), .Q(
        \adder_stage1[10][9] ) );
  DFF_X1 \adder_stage1_reg[10][10]  ( .D(n9993), .CK(clk), .Q(
        \adder_stage1[10][10] ) );
  DFF_X1 \adder_stage1_reg[10][11]  ( .D(n9992), .CK(clk), .Q(
        \adder_stage1[10][11] ) );
  DFF_X1 \adder_stage1_reg[10][12]  ( .D(n9991), .CK(clk), .Q(
        \adder_stage1[10][12] ) );
  DFF_X1 \adder_stage1_reg[10][13]  ( .D(n9990), .CK(clk), .Q(
        \adder_stage1[10][13] ) );
  DFF_X1 \adder_stage1_reg[10][14]  ( .D(n9989), .CK(clk), .Q(
        \adder_stage1[10][14] ) );
  DFF_X1 \adder_stage1_reg[10][15]  ( .D(n9988), .CK(clk), .Q(
        \adder_stage1[10][15] ) );
  DFF_X1 \adder_stage1_reg[10][20]  ( .D(n9987), .CK(clk), .Q(
        \adder_stage1[10][20] ), .QN(n3459) );
  DFF_X1 \adder_stage1_reg[11][0]  ( .D(n9986), .CK(clk), .Q(
        \adder_stage1[11][0] ) );
  DFF_X1 \adder_stage1_reg[11][1]  ( .D(n9985), .CK(clk), .Q(
        \adder_stage1[11][1] ) );
  DFF_X1 \adder_stage1_reg[11][2]  ( .D(n9984), .CK(clk), .Q(
        \adder_stage1[11][2] ) );
  DFF_X1 \adder_stage1_reg[11][3]  ( .D(n9983), .CK(clk), .Q(
        \adder_stage1[11][3] ) );
  DFF_X1 \adder_stage1_reg[11][4]  ( .D(n9982), .CK(clk), .Q(
        \adder_stage1[11][4] ) );
  DFF_X1 \adder_stage1_reg[11][5]  ( .D(n9981), .CK(clk), .Q(
        \adder_stage1[11][5] ) );
  DFF_X1 \adder_stage1_reg[11][6]  ( .D(n9980), .CK(clk), .Q(
        \adder_stage1[11][6] ) );
  DFF_X1 \adder_stage1_reg[11][7]  ( .D(n9979), .CK(clk), .Q(
        \adder_stage1[11][7] ) );
  DFF_X1 \adder_stage1_reg[11][8]  ( .D(n9978), .CK(clk), .Q(
        \adder_stage1[11][8] ) );
  DFF_X1 \adder_stage1_reg[11][10]  ( .D(n9976), .CK(clk), .Q(
        \adder_stage1[11][10] ) );
  DFF_X1 \adder_stage1_reg[11][11]  ( .D(n9975), .CK(clk), .Q(
        \adder_stage1[11][11] ) );
  DFF_X1 \adder_stage1_reg[11][12]  ( .D(n9974), .CK(clk), .Q(
        \adder_stage1[11][12] ) );
  DFF_X1 \adder_stage1_reg[11][13]  ( .D(n9973), .CK(clk), .Q(
        \adder_stage1[11][13] ) );
  DFF_X1 \adder_stage1_reg[11][14]  ( .D(n9972), .CK(clk), .Q(
        \adder_stage1[11][14] ) );
  DFF_X1 \adder_stage1_reg[11][15]  ( .D(n9971), .CK(clk), .Q(
        \adder_stage1[11][15] ) );
  DFF_X1 \adder_stage1_reg[11][20]  ( .D(n9970), .CK(clk), .Q(
        \adder_stage1[11][20] ), .QN(n3446) );
  DFF_X1 \adder_stage1_reg[12][0]  ( .D(n9969), .CK(clk), .Q(
        \adder_stage1[12][0] ) );
  DFF_X1 \adder_stage1_reg[12][1]  ( .D(n9968), .CK(clk), .Q(
        \adder_stage1[12][1] ) );
  DFF_X1 \adder_stage1_reg[12][2]  ( .D(n9967), .CK(clk), .Q(
        \adder_stage1[12][2] ) );
  DFF_X1 \adder_stage1_reg[12][3]  ( .D(n9966), .CK(clk), .Q(
        \adder_stage1[12][3] ) );
  DFF_X1 \adder_stage1_reg[12][4]  ( .D(n9965), .CK(clk), .Q(
        \adder_stage1[12][4] ) );
  DFF_X1 \adder_stage1_reg[12][5]  ( .D(n9964), .CK(clk), .Q(
        \adder_stage1[12][5] ) );
  DFF_X1 \adder_stage1_reg[12][6]  ( .D(n9963), .CK(clk), .Q(
        \adder_stage1[12][6] ) );
  DFF_X1 \adder_stage1_reg[12][8]  ( .D(n9961), .CK(clk), .Q(
        \adder_stage1[12][8] ) );
  DFF_X1 \adder_stage1_reg[12][9]  ( .D(n9960), .CK(clk), .Q(
        \adder_stage1[12][9] ) );
  DFF_X1 \adder_stage1_reg[12][10]  ( .D(n9959), .CK(clk), .Q(
        \adder_stage1[12][10] ) );
  DFF_X1 \adder_stage1_reg[12][11]  ( .D(n9958), .CK(clk), .Q(
        \adder_stage1[12][11] ) );
  DFF_X1 \adder_stage1_reg[12][12]  ( .D(n9957), .CK(clk), .Q(
        \adder_stage1[12][12] ) );
  DFF_X1 \adder_stage1_reg[12][13]  ( .D(n9956), .CK(clk), .Q(
        \adder_stage1[12][13] ) );
  DFF_X1 \adder_stage1_reg[12][14]  ( .D(n9955), .CK(clk), .Q(
        \adder_stage1[12][14] ) );
  DFF_X1 \adder_stage1_reg[12][15]  ( .D(n9954), .CK(clk), .Q(
        \adder_stage1[12][15] ) );
  DFF_X1 \adder_stage1_reg[12][20]  ( .D(n9953), .CK(clk), .Q(
        \adder_stage1[12][20] ), .QN(n3452) );
  DFF_X1 \adder_stage1_reg[13][0]  ( .D(n9952), .CK(clk), .Q(
        \adder_stage1[13][0] ) );
  DFF_X1 \adder_stage1_reg[13][1]  ( .D(n9951), .CK(clk), .Q(
        \adder_stage1[13][1] ) );
  DFF_X1 \adder_stage1_reg[13][2]  ( .D(n9950), .CK(clk), .Q(
        \adder_stage1[13][2] ) );
  DFF_X1 \adder_stage1_reg[13][3]  ( .D(n9949), .CK(clk), .Q(
        \adder_stage1[13][3] ) );
  DFF_X1 \adder_stage1_reg[13][4]  ( .D(n9948), .CK(clk), .Q(
        \adder_stage1[13][4] ) );
  DFF_X1 \adder_stage1_reg[13][5]  ( .D(n9947), .CK(clk), .Q(
        \adder_stage1[13][5] ) );
  DFF_X1 \adder_stage1_reg[13][6]  ( .D(n9946), .CK(clk), .Q(
        \adder_stage1[13][6] ) );
  DFF_X1 \adder_stage1_reg[13][7]  ( .D(n9945), .CK(clk), .Q(
        \adder_stage1[13][7] ) );
  DFF_X1 \adder_stage1_reg[13][8]  ( .D(n9944), .CK(clk), .Q(
        \adder_stage1[13][8] ) );
  DFF_X1 \adder_stage1_reg[13][9]  ( .D(n9943), .CK(clk), .Q(
        \adder_stage1[13][9] ) );
  DFF_X1 \adder_stage1_reg[13][10]  ( .D(n9942), .CK(clk), .Q(
        \adder_stage1[13][10] ) );
  DFF_X1 \adder_stage1_reg[13][11]  ( .D(n9941), .CK(clk), .Q(
        \adder_stage1[13][11] ) );
  DFF_X1 \adder_stage1_reg[13][12]  ( .D(n9940), .CK(clk), .Q(
        \adder_stage1[13][12] ) );
  DFF_X1 \adder_stage1_reg[13][13]  ( .D(n9939), .CK(clk), .Q(
        \adder_stage1[13][13] ) );
  DFF_X1 \adder_stage1_reg[13][14]  ( .D(n9938), .CK(clk), .Q(
        \adder_stage1[13][14] ) );
  DFF_X1 \adder_stage1_reg[13][15]  ( .D(n9937), .CK(clk), .Q(
        \adder_stage1[13][15] ) );
  DFF_X1 \adder_stage1_reg[13][20]  ( .D(n9936), .CK(clk), .Q(
        \adder_stage1[13][20] ), .QN(n3473) );
  DFF_X1 \adder_stage1_reg[14][0]  ( .D(n9935), .CK(clk), .Q(
        \adder_stage1[14][0] ) );
  DFF_X1 \adder_stage1_reg[14][1]  ( .D(n9934), .CK(clk), .Q(
        \adder_stage1[14][1] ) );
  DFF_X1 \adder_stage1_reg[14][2]  ( .D(n9933), .CK(clk), .Q(
        \adder_stage1[14][2] ) );
  DFF_X1 \adder_stage1_reg[14][3]  ( .D(n9932), .CK(clk), .Q(
        \adder_stage1[14][3] ) );
  DFF_X1 \adder_stage1_reg[14][4]  ( .D(n9931), .CK(clk), .Q(
        \adder_stage1[14][4] ) );
  DFF_X1 \adder_stage1_reg[14][5]  ( .D(n9930), .CK(clk), .Q(
        \adder_stage1[14][5] ) );
  DFF_X1 \adder_stage1_reg[14][6]  ( .D(n9929), .CK(clk), .Q(
        \adder_stage1[14][6] ) );
  DFF_X1 \adder_stage1_reg[14][7]  ( .D(n9928), .CK(clk), .Q(
        \adder_stage1[14][7] ) );
  DFF_X1 \adder_stage1_reg[14][8]  ( .D(n9927), .CK(clk), .Q(
        \adder_stage1[14][8] ) );
  DFF_X1 \adder_stage1_reg[14][9]  ( .D(n9926), .CK(clk), .Q(
        \adder_stage1[14][9] ) );
  DFF_X1 \adder_stage1_reg[14][10]  ( .D(n9925), .CK(clk), .Q(
        \adder_stage1[14][10] ) );
  DFF_X1 \adder_stage1_reg[14][11]  ( .D(n9924), .CK(clk), .Q(
        \adder_stage1[14][11] ) );
  DFF_X1 \adder_stage1_reg[14][12]  ( .D(n9923), .CK(clk), .Q(
        \adder_stage1[14][12] ) );
  DFF_X1 \adder_stage1_reg[14][13]  ( .D(n9922), .CK(clk), .Q(
        \adder_stage1[14][13] ) );
  DFF_X1 \adder_stage1_reg[14][14]  ( .D(n9921), .CK(clk), .Q(
        \adder_stage1[14][14] ) );
  DFF_X1 \adder_stage1_reg[14][15]  ( .D(n9920), .CK(clk), .Q(
        \adder_stage1[14][15] ) );
  DFF_X1 \adder_stage1_reg[14][20]  ( .D(n9919), .CK(clk), .Q(
        \adder_stage1[14][20] ), .QN(n3453) );
  DFF_X1 \adder_stage1_reg[15][0]  ( .D(n9918), .CK(clk), .Q(
        \adder_stage1[15][0] ) );
  DFF_X1 \adder_stage1_reg[15][1]  ( .D(n9917), .CK(clk), .Q(
        \adder_stage1[15][1] ) );
  DFF_X1 \adder_stage1_reg[15][2]  ( .D(n9916), .CK(clk), .Q(
        \adder_stage1[15][2] ) );
  DFF_X1 \adder_stage1_reg[15][3]  ( .D(n9915), .CK(clk), .Q(
        \adder_stage1[15][3] ) );
  DFF_X1 \adder_stage1_reg[15][4]  ( .D(n9914), .CK(clk), .Q(
        \adder_stage1[15][4] ) );
  DFF_X1 \adder_stage1_reg[15][5]  ( .D(n9913), .CK(clk), .Q(
        \adder_stage1[15][5] ) );
  DFF_X1 \adder_stage1_reg[15][6]  ( .D(n9912), .CK(clk), .Q(
        \adder_stage1[15][6] ) );
  DFF_X1 \adder_stage1_reg[15][7]  ( .D(n9911), .CK(clk), .Q(
        \adder_stage1[15][7] ) );
  DFF_X1 \adder_stage1_reg[15][8]  ( .D(n9910), .CK(clk), .Q(
        \adder_stage1[15][8] ) );
  DFF_X1 \adder_stage1_reg[15][9]  ( .D(n9909), .CK(clk), .Q(
        \adder_stage1[15][9] ) );
  DFF_X1 \adder_stage1_reg[15][10]  ( .D(n9908), .CK(clk), .Q(
        \adder_stage1[15][10] ) );
  DFF_X1 \adder_stage1_reg[15][11]  ( .D(n9907), .CK(clk), .Q(
        \adder_stage1[15][11] ) );
  DFF_X1 \adder_stage1_reg[15][12]  ( .D(n9906), .CK(clk), .Q(
        \adder_stage1[15][12] ) );
  DFF_X1 \adder_stage1_reg[15][20]  ( .D(n9905), .CK(clk), .Q(
        \adder_stage1[15][20] ), .QN(n3474) );
  DFF_X1 \adder_stage2_reg[0][0]  ( .D(n9904), .CK(clk), .Q(
        \adder_stage2[0][0] ) );
  DFF_X1 \adder_stage2_reg[0][1]  ( .D(n9903), .CK(clk), .Q(
        \adder_stage2[0][1] ) );
  DFF_X1 \adder_stage2_reg[0][2]  ( .D(n9902), .CK(clk), .Q(
        \adder_stage2[0][2] ) );
  DFF_X1 \adder_stage2_reg[0][3]  ( .D(n9901), .CK(clk), .Q(
        \adder_stage2[0][3] ) );
  DFF_X1 \adder_stage2_reg[0][4]  ( .D(n9900), .CK(clk), .Q(
        \adder_stage2[0][4] ) );
  DFF_X1 \adder_stage2_reg[0][5]  ( .D(n9899), .CK(clk), .Q(
        \adder_stage2[0][5] ) );
  DFF_X1 \adder_stage2_reg[0][6]  ( .D(n9898), .CK(clk), .Q(
        \adder_stage2[0][6] ) );
  DFF_X1 \adder_stage2_reg[0][7]  ( .D(n9897), .CK(clk), .Q(
        \adder_stage2[0][7] ) );
  DFF_X1 \adder_stage2_reg[0][8]  ( .D(n9896), .CK(clk), .Q(
        \adder_stage2[0][8] ) );
  DFF_X1 \adder_stage2_reg[0][9]  ( .D(n9895), .CK(clk), .Q(
        \adder_stage2[0][9] ) );
  DFF_X1 \adder_stage2_reg[0][10]  ( .D(n9894), .CK(clk), .Q(
        \adder_stage2[0][10] ) );
  DFF_X1 \adder_stage2_reg[0][11]  ( .D(n9893), .CK(clk), .Q(
        \adder_stage2[0][11] ) );
  DFF_X1 \adder_stage2_reg[0][12]  ( .D(n9892), .CK(clk), .Q(
        \adder_stage2[0][12] ) );
  DFF_X1 \adder_stage2_reg[0][13]  ( .D(n9891), .CK(clk), .Q(
        \adder_stage2[0][13] ) );
  DFF_X1 \adder_stage2_reg[0][14]  ( .D(n9890), .CK(clk), .Q(
        \adder_stage2[0][14] ) );
  DFF_X1 \adder_stage2_reg[0][15]  ( .D(n9889), .CK(clk), .Q(
        \adder_stage2[0][15] ) );
  DFF_X1 \adder_stage2_reg[0][16]  ( .D(n9888), .CK(clk), .Q(
        \adder_stage2[0][16] ) );
  DFF_X1 \adder_stage2_reg[0][17]  ( .D(n2059), .CK(clk), .Q(
        \adder_stage2[0][17] ), .QN(n8834) );
  DFF_X1 \adder_stage2_reg[0][18]  ( .D(n2058), .CK(clk), .Q(
        \adder_stage2[0][18] ), .QN(n8835) );
  DFF_X1 \adder_stage2_reg[0][19]  ( .D(n2057), .CK(clk), .Q(
        \adder_stage2[0][19] ), .QN(n8836) );
  DFF_X1 \adder_stage2_reg[0][20]  ( .D(n2056), .CK(clk), .Q(
        \adder_stage2[0][20] ), .QN(n8848) );
  DFF_X1 \adder_stage2_reg[1][0]  ( .D(n9887), .CK(clk), .Q(
        \adder_stage2[1][0] ) );
  DFF_X1 \adder_stage2_reg[1][1]  ( .D(n9886), .CK(clk), .Q(
        \adder_stage2[1][1] ) );
  DFF_X1 \adder_stage2_reg[1][2]  ( .D(n9885), .CK(clk), .Q(
        \adder_stage2[1][2] ) );
  DFF_X1 \adder_stage2_reg[1][3]  ( .D(n9884), .CK(clk), .Q(
        \adder_stage2[1][3] ) );
  DFF_X1 \adder_stage2_reg[1][4]  ( .D(n9883), .CK(clk), .Q(
        \adder_stage2[1][4] ) );
  DFF_X1 \adder_stage2_reg[1][5]  ( .D(n9882), .CK(clk), .Q(
        \adder_stage2[1][5] ) );
  DFF_X1 \adder_stage2_reg[1][6]  ( .D(n9881), .CK(clk), .Q(
        \adder_stage2[1][6] ) );
  DFF_X1 \adder_stage2_reg[1][7]  ( .D(n9880), .CK(clk), .Q(
        \adder_stage2[1][7] ) );
  DFF_X1 \adder_stage2_reg[1][8]  ( .D(n9879), .CK(clk), .Q(
        \adder_stage2[1][8] ) );
  DFF_X1 \adder_stage2_reg[1][9]  ( .D(n9878), .CK(clk), .Q(
        \adder_stage2[1][9] ) );
  DFF_X1 \adder_stage2_reg[1][10]  ( .D(n9877), .CK(clk), .Q(
        \adder_stage2[1][10] ) );
  DFF_X1 \adder_stage2_reg[1][11]  ( .D(n9876), .CK(clk), .Q(
        \adder_stage2[1][11] ) );
  DFF_X1 \adder_stage2_reg[1][12]  ( .D(n9875), .CK(clk), .Q(
        \adder_stage2[1][12] ) );
  DFF_X1 \adder_stage2_reg[1][13]  ( .D(n9874), .CK(clk), .Q(
        \adder_stage2[1][13] ) );
  DFF_X1 \adder_stage2_reg[1][14]  ( .D(n9873), .CK(clk), .Q(
        \adder_stage2[1][14] ) );
  DFF_X1 \adder_stage2_reg[1][15]  ( .D(n9872), .CK(clk), .Q(
        \adder_stage2[1][15] ) );
  DFF_X1 \adder_stage2_reg[1][16]  ( .D(n9871), .CK(clk), .Q(
        \adder_stage2[1][16] ) );
  DFF_X1 \adder_stage2_reg[1][17]  ( .D(n2038), .CK(clk), .Q(
        \adder_stage2[1][17] ), .QN(n8825) );
  DFF_X1 \adder_stage2_reg[1][18]  ( .D(n2037), .CK(clk), .Q(
        \adder_stage2[1][18] ), .QN(n8826) );
  DFF_X1 \adder_stage2_reg[1][19]  ( .D(n2036), .CK(clk), .Q(
        \adder_stage2[1][19] ), .QN(n8827) );
  DFF_X1 \adder_stage2_reg[1][20]  ( .D(n2035), .CK(clk), .Q(
        \adder_stage2[1][20] ), .QN(n8853) );
  DFF_X1 \adder_stage2_reg[2][0]  ( .D(n9870), .CK(clk), .Q(
        \adder_stage2[2][0] ) );
  DFF_X1 \adder_stage2_reg[2][1]  ( .D(n9869), .CK(clk), .Q(
        \adder_stage2[2][1] ) );
  DFF_X1 \adder_stage2_reg[2][2]  ( .D(n9868), .CK(clk), .Q(
        \adder_stage2[2][2] ) );
  DFF_X1 \adder_stage2_reg[2][3]  ( .D(n9867), .CK(clk), .Q(
        \adder_stage2[2][3] ) );
  DFF_X1 \adder_stage2_reg[2][4]  ( .D(n9866), .CK(clk), .Q(
        \adder_stage2[2][4] ) );
  DFF_X1 \adder_stage2_reg[2][5]  ( .D(n9865), .CK(clk), .Q(
        \adder_stage2[2][5] ) );
  DFF_X1 \adder_stage2_reg[2][6]  ( .D(n9864), .CK(clk), .Q(
        \adder_stage2[2][6] ) );
  DFF_X1 \adder_stage2_reg[2][7]  ( .D(n9863), .CK(clk), .Q(
        \adder_stage2[2][7] ) );
  DFF_X1 \adder_stage2_reg[2][8]  ( .D(n9862), .CK(clk), .Q(
        \adder_stage2[2][8] ) );
  DFF_X1 \adder_stage2_reg[2][9]  ( .D(n9861), .CK(clk), .Q(
        \adder_stage2[2][9] ) );
  DFF_X1 \adder_stage2_reg[2][10]  ( .D(n9860), .CK(clk), .Q(
        \adder_stage2[2][10] ) );
  DFF_X1 \adder_stage2_reg[2][11]  ( .D(n9859), .CK(clk), .Q(
        \adder_stage2[2][11] ) );
  DFF_X1 \adder_stage2_reg[2][12]  ( .D(n9858), .CK(clk), .Q(
        \adder_stage2[2][12] ) );
  DFF_X1 \adder_stage2_reg[2][13]  ( .D(n9857), .CK(clk), .Q(
        \adder_stage2[2][13] ) );
  DFF_X1 \adder_stage2_reg[2][14]  ( .D(n9856), .CK(clk), .Q(
        \adder_stage2[2][14] ) );
  DFF_X1 \adder_stage2_reg[2][15]  ( .D(n9855), .CK(clk), .Q(
        \adder_stage2[2][15] ) );
  DFF_X1 \adder_stage2_reg[2][16]  ( .D(n9854), .CK(clk), .Q(
        \adder_stage2[2][16] ) );
  DFF_X1 \adder_stage2_reg[2][17]  ( .D(n2017), .CK(clk), .Q(
        \adder_stage2[2][17] ), .QN(n8837) );
  DFF_X1 \adder_stage2_reg[2][18]  ( .D(n2016), .CK(clk), .Q(
        \adder_stage2[2][18] ), .QN(n8838) );
  DFF_X1 \adder_stage2_reg[2][19]  ( .D(n2015), .CK(clk), .Q(
        \adder_stage2[2][19] ), .QN(n8839) );
  DFF_X1 \adder_stage2_reg[2][20]  ( .D(n2014), .CK(clk), .Q(
        \adder_stage2[2][20] ), .QN(n8849) );
  DFF_X1 \adder_stage2_reg[3][0]  ( .D(n9853), .CK(clk), .Q(
        \adder_stage2[3][0] ) );
  DFF_X1 \adder_stage2_reg[3][1]  ( .D(n9852), .CK(clk), .Q(
        \adder_stage2[3][1] ) );
  DFF_X1 \adder_stage2_reg[3][2]  ( .D(n9851), .CK(clk), .Q(
        \adder_stage2[3][2] ) );
  DFF_X1 \adder_stage2_reg[3][3]  ( .D(n9850), .CK(clk), .Q(
        \adder_stage2[3][3] ) );
  DFF_X1 \adder_stage2_reg[3][4]  ( .D(n9849), .CK(clk), .Q(
        \adder_stage2[3][4] ) );
  DFF_X1 \adder_stage2_reg[3][5]  ( .D(n9848), .CK(clk), .Q(
        \adder_stage2[3][5] ) );
  DFF_X1 \adder_stage2_reg[3][6]  ( .D(n9847), .CK(clk), .Q(
        \adder_stage2[3][6] ) );
  DFF_X1 \adder_stage2_reg[3][7]  ( .D(n9846), .CK(clk), .Q(
        \adder_stage2[3][7] ) );
  DFF_X1 \adder_stage2_reg[3][8]  ( .D(n9845), .CK(clk), .Q(
        \adder_stage2[3][8] ) );
  DFF_X1 \adder_stage2_reg[3][9]  ( .D(n9844), .CK(clk), .Q(
        \adder_stage2[3][9] ) );
  DFF_X1 \adder_stage2_reg[3][10]  ( .D(n9843), .CK(clk), .Q(
        \adder_stage2[3][10] ) );
  DFF_X1 \adder_stage2_reg[3][12]  ( .D(n9841), .CK(clk), .Q(
        \adder_stage2[3][12] ) );
  DFF_X1 \adder_stage2_reg[3][13]  ( .D(n9840), .CK(clk), .Q(
        \adder_stage2[3][13] ) );
  DFF_X1 \adder_stage2_reg[3][14]  ( .D(n9839), .CK(clk), .Q(
        \adder_stage2[3][14] ) );
  DFF_X1 \adder_stage2_reg[3][15]  ( .D(n9838), .CK(clk), .Q(
        \adder_stage2[3][15] ) );
  DFF_X1 \adder_stage2_reg[3][16]  ( .D(n9837), .CK(clk), .Q(
        \adder_stage2[3][16] ) );
  DFF_X1 \adder_stage2_reg[3][17]  ( .D(n1996), .CK(clk), .Q(
        \adder_stage2[3][17] ), .QN(n8816) );
  DFF_X1 \adder_stage2_reg[3][18]  ( .D(n1995), .CK(clk), .Q(
        \adder_stage2[3][18] ), .QN(n8817) );
  DFF_X1 \adder_stage2_reg[3][19]  ( .D(n1994), .CK(clk), .Q(
        \adder_stage2[3][19] ), .QN(n8818) );
  DFF_X1 \adder_stage2_reg[3][20]  ( .D(n1993), .CK(clk), .Q(
        \adder_stage2[3][20] ), .QN(n8850) );
  DFF_X1 \adder_stage2_reg[4][0]  ( .D(n9836), .CK(clk), .Q(
        \adder_stage2[4][0] ) );
  DFF_X1 \adder_stage2_reg[4][1]  ( .D(n9835), .CK(clk), .Q(
        \adder_stage2[4][1] ) );
  DFF_X1 \adder_stage2_reg[4][2]  ( .D(n9834), .CK(clk), .Q(
        \adder_stage2[4][2] ) );
  DFF_X1 \adder_stage2_reg[4][3]  ( .D(n9833), .CK(clk), .Q(
        \adder_stage2[4][3] ) );
  DFF_X1 \adder_stage2_reg[4][4]  ( .D(n9832), .CK(clk), .Q(
        \adder_stage2[4][4] ) );
  DFF_X1 \adder_stage2_reg[4][5]  ( .D(n9831), .CK(clk), .Q(
        \adder_stage2[4][5] ) );
  DFF_X1 \adder_stage2_reg[4][6]  ( .D(n9830), .CK(clk), .Q(
        \adder_stage2[4][6] ) );
  DFF_X1 \adder_stage2_reg[4][7]  ( .D(n9829), .CK(clk), .Q(
        \adder_stage2[4][7] ) );
  DFF_X1 \adder_stage2_reg[4][8]  ( .D(n9828), .CK(clk), .Q(
        \adder_stage2[4][8] ) );
  DFF_X1 \adder_stage2_reg[4][9]  ( .D(n9827), .CK(clk), .Q(
        \adder_stage2[4][9] ) );
  DFF_X1 \adder_stage2_reg[4][10]  ( .D(n9826), .CK(clk), .Q(
        \adder_stage2[4][10] ) );
  DFF_X1 \adder_stage2_reg[4][11]  ( .D(n9825), .CK(clk), .Q(
        \adder_stage2[4][11] ) );
  DFF_X1 \adder_stage2_reg[4][12]  ( .D(n9824), .CK(clk), .Q(
        \adder_stage2[4][12] ) );
  DFF_X1 \adder_stage2_reg[4][13]  ( .D(n9823), .CK(clk), .Q(
        \adder_stage2[4][13] ) );
  DFF_X1 \adder_stage2_reg[4][14]  ( .D(n9822), .CK(clk), .Q(
        \adder_stage2[4][14] ) );
  DFF_X1 \adder_stage2_reg[4][15]  ( .D(n9821), .CK(clk), .Q(
        \adder_stage2[4][15] ) );
  DFF_X1 \adder_stage2_reg[4][16]  ( .D(n9820), .CK(clk), .Q(
        \adder_stage2[4][16] ) );
  DFF_X1 \adder_stage2_reg[4][17]  ( .D(n1975), .CK(clk), .Q(
        \adder_stage2[4][17] ), .QN(n8828) );
  DFF_X1 \adder_stage2_reg[4][18]  ( .D(n1974), .CK(clk), .Q(
        \adder_stage2[4][18] ), .QN(n8829) );
  DFF_X1 \adder_stage2_reg[4][19]  ( .D(n1973), .CK(clk), .Q(
        \adder_stage2[4][19] ), .QN(n8830) );
  DFF_X1 \adder_stage2_reg[4][20]  ( .D(n1972), .CK(clk), .Q(
        \adder_stage2[4][20] ), .QN(n8846) );
  DFF_X1 \adder_stage2_reg[5][0]  ( .D(n9819), .CK(clk), .Q(
        \adder_stage2[5][0] ) );
  DFF_X1 \adder_stage2_reg[5][1]  ( .D(n9818), .CK(clk), .Q(
        \adder_stage2[5][1] ) );
  DFF_X1 \adder_stage2_reg[5][2]  ( .D(n9817), .CK(clk), .Q(
        \adder_stage2[5][2] ) );
  DFF_X1 \adder_stage2_reg[5][4]  ( .D(n9815), .CK(clk), .Q(
        \adder_stage2[5][4] ) );
  DFF_X1 \adder_stage2_reg[5][5]  ( .D(n9814), .CK(clk), .Q(
        \adder_stage2[5][5] ) );
  DFF_X1 \adder_stage2_reg[5][6]  ( .D(n9813), .CK(clk), .Q(
        \adder_stage2[5][6] ) );
  DFF_X1 \adder_stage2_reg[5][7]  ( .D(n9812), .CK(clk), .Q(
        \adder_stage2[5][7] ) );
  DFF_X1 \adder_stage2_reg[5][8]  ( .D(n9811), .CK(clk), .Q(
        \adder_stage2[5][8] ) );
  DFF_X1 \adder_stage2_reg[5][9]  ( .D(n9810), .CK(clk), .Q(
        \adder_stage2[5][9] ) );
  DFF_X1 \adder_stage2_reg[5][10]  ( .D(n9809), .CK(clk), .Q(
        \adder_stage2[5][10] ) );
  DFF_X1 \adder_stage2_reg[5][11]  ( .D(n9808), .CK(clk), .Q(
        \adder_stage2[5][11] ) );
  DFF_X1 \adder_stage2_reg[5][12]  ( .D(n9807), .CK(clk), .Q(
        \adder_stage2[5][12] ) );
  DFF_X1 \adder_stage2_reg[5][13]  ( .D(n9806), .CK(clk), .Q(
        \adder_stage2[5][13] ) );
  DFF_X1 \adder_stage2_reg[5][14]  ( .D(n9805), .CK(clk), .Q(
        \adder_stage2[5][14] ) );
  DFF_X1 \adder_stage2_reg[5][15]  ( .D(n9804), .CK(clk), .Q(
        \adder_stage2[5][15] ) );
  DFF_X1 \adder_stage2_reg[5][17]  ( .D(n1954), .CK(clk), .Q(
        \adder_stage2[5][17] ), .QN(n8819) );
  DFF_X1 \adder_stage2_reg[5][18]  ( .D(n1953), .CK(clk), .Q(
        \adder_stage2[5][18] ), .QN(n8820) );
  DFF_X1 \adder_stage2_reg[5][19]  ( .D(n1952), .CK(clk), .Q(
        \adder_stage2[5][19] ), .QN(n8821) );
  DFF_X1 \adder_stage2_reg[5][20]  ( .D(n1951), .CK(clk), .Q(
        \adder_stage2[5][20] ), .QN(n8851) );
  DFF_X1 \adder_stage2_reg[6][0]  ( .D(n9803), .CK(clk), .Q(
        \adder_stage2[6][0] ) );
  DFF_X1 \adder_stage2_reg[6][1]  ( .D(n9802), .CK(clk), .Q(
        \adder_stage2[6][1] ) );
  DFF_X1 \adder_stage2_reg[6][2]  ( .D(n9801), .CK(clk), .Q(
        \adder_stage2[6][2] ) );
  DFF_X1 \adder_stage2_reg[6][3]  ( .D(n9800), .CK(clk), .Q(
        \adder_stage2[6][3] ) );
  DFF_X1 \adder_stage2_reg[6][4]  ( .D(n9799), .CK(clk), .Q(
        \adder_stage2[6][4] ) );
  DFF_X1 \adder_stage2_reg[6][5]  ( .D(n9798), .CK(clk), .Q(
        \adder_stage2[6][5] ) );
  DFF_X1 \adder_stage2_reg[6][6]  ( .D(n9797), .CK(clk), .Q(
        \adder_stage2[6][6] ) );
  DFF_X1 \adder_stage2_reg[6][7]  ( .D(n9796), .CK(clk), .Q(
        \adder_stage2[6][7] ) );
  DFF_X1 \adder_stage2_reg[6][8]  ( .D(n9795), .CK(clk), .Q(
        \adder_stage2[6][8] ) );
  DFF_X1 \adder_stage2_reg[6][9]  ( .D(n9794), .CK(clk), .Q(
        \adder_stage2[6][9] ) );
  DFF_X1 \adder_stage2_reg[6][10]  ( .D(n9793), .CK(clk), .Q(
        \adder_stage2[6][10] ) );
  DFF_X1 \adder_stage2_reg[6][11]  ( .D(n9792), .CK(clk), .Q(
        \adder_stage2[6][11] ) );
  DFF_X1 \adder_stage2_reg[6][12]  ( .D(n9791), .CK(clk), .Q(
        \adder_stage2[6][12] ) );
  DFF_X1 \adder_stage2_reg[6][13]  ( .D(n9790), .CK(clk), .Q(
        \adder_stage2[6][13] ) );
  DFF_X1 \adder_stage2_reg[6][14]  ( .D(n9789), .CK(clk), .Q(
        \adder_stage2[6][14] ) );
  DFF_X1 \adder_stage2_reg[6][15]  ( .D(n9788), .CK(clk), .Q(
        \adder_stage2[6][15] ) );
  DFF_X1 \adder_stage2_reg[6][16]  ( .D(n9787), .CK(clk), .Q(
        \adder_stage2[6][16] ) );
  DFF_X1 \adder_stage2_reg[6][17]  ( .D(n1933), .CK(clk), .Q(
        \adder_stage2[6][17] ), .QN(n8831) );
  DFF_X1 \adder_stage2_reg[6][18]  ( .D(n1932), .CK(clk), .Q(
        \adder_stage2[6][18] ), .QN(n8832) );
  DFF_X1 \adder_stage2_reg[6][19]  ( .D(n1931), .CK(clk), .Q(
        \adder_stage2[6][19] ), .QN(n8833) );
  DFF_X1 \adder_stage2_reg[6][20]  ( .D(n1930), .CK(clk), .Q(
        \adder_stage2[6][20] ), .QN(n8847) );
  DFF_X1 \adder_stage2_reg[7][1]  ( .D(n9785), .CK(clk), .Q(
        \adder_stage2[7][1] ) );
  DFF_X1 \adder_stage2_reg[7][2]  ( .D(n9784), .CK(clk), .Q(
        \adder_stage2[7][2] ) );
  DFF_X1 \adder_stage2_reg[7][3]  ( .D(n9783), .CK(clk), .Q(
        \adder_stage2[7][3] ) );
  DFF_X1 \adder_stage2_reg[7][4]  ( .D(n9782), .CK(clk), .Q(
        \adder_stage2[7][4] ) );
  DFF_X1 \adder_stage2_reg[7][5]  ( .D(n9781), .CK(clk), .Q(
        \adder_stage2[7][5] ) );
  DFF_X1 \adder_stage2_reg[7][6]  ( .D(n9780), .CK(clk), .Q(
        \adder_stage2[7][6] ) );
  DFF_X1 \adder_stage2_reg[7][7]  ( .D(n9779), .CK(clk), .Q(
        \adder_stage2[7][7] ) );
  DFF_X1 \adder_stage2_reg[7][8]  ( .D(n9778), .CK(clk), .Q(
        \adder_stage2[7][8] ) );
  DFF_X1 \adder_stage2_reg[7][9]  ( .D(n9777), .CK(clk), .Q(
        \adder_stage2[7][9] ) );
  DFF_X1 \adder_stage2_reg[7][10]  ( .D(n9776), .CK(clk), .Q(
        \adder_stage2[7][10] ) );
  DFF_X1 \adder_stage2_reg[7][11]  ( .D(n9775), .CK(clk), .Q(
        \adder_stage2[7][11] ) );
  DFF_X1 \adder_stage2_reg[7][12]  ( .D(n9774), .CK(clk), .Q(
        \adder_stage2[7][12] ) );
  DFF_X1 \adder_stage2_reg[7][13]  ( .D(n9773), .CK(clk), .Q(
        \adder_stage2[7][13] ) );
  DFF_X1 \adder_stage2_reg[7][14]  ( .D(n9772), .CK(clk), .Q(
        \adder_stage2[7][14] ) );
  DFF_X1 \adder_stage2_reg[7][15]  ( .D(n9771), .CK(clk), .Q(
        \adder_stage2[7][15] ) );
  DFF_X1 \adder_stage2_reg[7][16]  ( .D(n9770), .CK(clk), .Q(
        \adder_stage2[7][16] ) );
  DFF_X1 \adder_stage2_reg[7][17]  ( .D(n1912), .CK(clk), .Q(
        \adder_stage2[7][17] ), .QN(n8822) );
  DFF_X1 \adder_stage2_reg[7][18]  ( .D(n1911), .CK(clk), .Q(
        \adder_stage2[7][18] ), .QN(n8823) );
  DFF_X1 \adder_stage2_reg[7][19]  ( .D(n1910), .CK(clk), .Q(
        \adder_stage2[7][19] ), .QN(n8824) );
  DFF_X1 \adder_stage2_reg[7][20]  ( .D(n1909), .CK(clk), .Q(
        \adder_stage2[7][20] ), .QN(n8852) );
  DFF_X1 \adder_stage3_reg[0][0]  ( .D(n9769), .CK(clk), .Q(
        \adder_stage3[0][0] ) );
  DFF_X1 \adder_stage3_reg[0][1]  ( .D(n9768), .CK(clk), .Q(
        \adder_stage3[0][1] ) );
  DFF_X1 \adder_stage3_reg[0][2]  ( .D(n9767), .CK(clk), .Q(
        \adder_stage3[0][2] ) );
  DFF_X1 \adder_stage3_reg[0][3]  ( .D(n9766), .CK(clk), .Q(
        \adder_stage3[0][3] ) );
  DFF_X1 \adder_stage3_reg[0][4]  ( .D(n9765), .CK(clk), .Q(
        \adder_stage3[0][4] ) );
  DFF_X1 \adder_stage3_reg[0][5]  ( .D(n9764), .CK(clk), .Q(
        \adder_stage3[0][5] ) );
  DFF_X1 \adder_stage3_reg[0][6]  ( .D(n9763), .CK(clk), .Q(
        \adder_stage3[0][6] ) );
  DFF_X1 \adder_stage3_reg[0][7]  ( .D(n9762), .CK(clk), .Q(
        \adder_stage3[0][7] ) );
  DFF_X1 \adder_stage3_reg[0][8]  ( .D(n9761), .CK(clk), .Q(
        \adder_stage3[0][8] ) );
  DFF_X1 \adder_stage3_reg[0][9]  ( .D(n9760), .CK(clk), .Q(
        \adder_stage3[0][9] ) );
  DFF_X1 \adder_stage3_reg[0][10]  ( .D(n9759), .CK(clk), .Q(
        \adder_stage3[0][10] ) );
  DFF_X1 \adder_stage3_reg[0][11]  ( .D(n9758), .CK(clk), .Q(
        \adder_stage3[0][11] ) );
  DFF_X1 \adder_stage3_reg[0][12]  ( .D(n9757), .CK(clk), .Q(
        \adder_stage3[0][12] ) );
  DFF_X1 \adder_stage3_reg[0][13]  ( .D(n9756), .CK(clk), .Q(
        \adder_stage3[0][13] ) );
  DFF_X1 \adder_stage3_reg[0][14]  ( .D(n9755), .CK(clk), .Q(
        \adder_stage3[0][14] ) );
  DFF_X1 \adder_stage3_reg[0][15]  ( .D(n9754), .CK(clk), .Q(
        \adder_stage3[0][15] ) );
  DFF_X1 \adder_stage3_reg[0][16]  ( .D(n9753), .CK(clk), .Q(
        \adder_stage3[0][16] ) );
  DFF_X1 \adder_stage3_reg[0][17]  ( .D(n9752), .CK(clk), .Q(
        \adder_stage3[0][17] ) );
  DFF_X1 \adder_stage3_reg[0][18]  ( .D(n9751), .CK(clk), .Q(
        \adder_stage3[0][18] ) );
  DFF_X1 \adder_stage3_reg[0][19]  ( .D(n9750), .CK(clk), .Q(
        \adder_stage3[0][19] ) );
  DFF_X1 \adder_stage3_reg[0][20]  ( .D(n9749), .CK(clk), .Q(
        \adder_stage3[0][20] ) );
  DFF_X1 \adder_stage3_reg[1][0]  ( .D(n9748), .CK(clk), .Q(
        \adder_stage3[1][0] ) );
  DFF_X1 \adder_stage3_reg[1][1]  ( .D(n9747), .CK(clk), .Q(
        \adder_stage3[1][1] ) );
  DFF_X1 \adder_stage3_reg[1][2]  ( .D(n9746), .CK(clk), .Q(
        \adder_stage3[1][2] ) );
  DFF_X1 \adder_stage3_reg[1][3]  ( .D(n9745), .CK(clk), .Q(
        \adder_stage3[1][3] ) );
  DFF_X1 \adder_stage3_reg[1][4]  ( .D(n9744), .CK(clk), .Q(
        \adder_stage3[1][4] ) );
  DFF_X1 \adder_stage3_reg[1][5]  ( .D(n9743), .CK(clk), .Q(
        \adder_stage3[1][5] ) );
  DFF_X1 \adder_stage3_reg[1][6]  ( .D(n9742), .CK(clk), .Q(
        \adder_stage3[1][6] ) );
  DFF_X1 \adder_stage3_reg[1][7]  ( .D(n9741), .CK(clk), .Q(
        \adder_stage3[1][7] ) );
  DFF_X1 \adder_stage3_reg[1][8]  ( .D(n9740), .CK(clk), .Q(
        \adder_stage3[1][8] ) );
  DFF_X1 \adder_stage3_reg[1][9]  ( .D(n9739), .CK(clk), .Q(
        \adder_stage3[1][9] ) );
  DFF_X1 \adder_stage3_reg[1][10]  ( .D(n9738), .CK(clk), .Q(
        \adder_stage3[1][10] ) );
  DFF_X1 \adder_stage3_reg[1][11]  ( .D(n9737), .CK(clk), .Q(
        \adder_stage3[1][11] ) );
  DFF_X1 \adder_stage3_reg[1][12]  ( .D(n9736), .CK(clk), .Q(
        \adder_stage3[1][12] ) );
  DFF_X1 \adder_stage3_reg[1][13]  ( .D(n9735), .CK(clk), .Q(
        \adder_stage3[1][13] ) );
  DFF_X1 \adder_stage3_reg[1][14]  ( .D(n9734), .CK(clk), .Q(
        \adder_stage3[1][14] ) );
  DFF_X1 \adder_stage3_reg[1][15]  ( .D(n9733), .CK(clk), .Q(
        \adder_stage3[1][15] ) );
  DFF_X1 \adder_stage3_reg[1][16]  ( .D(n9732), .CK(clk), .Q(
        \adder_stage3[1][16] ) );
  DFF_X1 \adder_stage3_reg[1][17]  ( .D(n9731), .CK(clk), .Q(
        \adder_stage3[1][17] ) );
  DFF_X1 \adder_stage3_reg[1][20]  ( .D(n9730), .CK(clk), .Q(
        \adder_stage3[1][20] ) );
  DFF_X1 \adder_stage3_reg[2][0]  ( .D(n9729), .CK(clk), .Q(
        \adder_stage3[2][0] ) );
  DFF_X1 \adder_stage3_reg[2][1]  ( .D(n9728), .CK(clk), .Q(
        \adder_stage3[2][1] ) );
  DFF_X1 \adder_stage3_reg[2][2]  ( .D(n9727), .CK(clk), .Q(
        \adder_stage3[2][2] ) );
  DFF_X1 \adder_stage3_reg[2][3]  ( .D(n9726), .CK(clk), .Q(
        \adder_stage3[2][3] ) );
  DFF_X1 \adder_stage3_reg[2][4]  ( .D(n9725), .CK(clk), .Q(
        \adder_stage3[2][4] ) );
  DFF_X1 \adder_stage3_reg[2][5]  ( .D(n9724), .CK(clk), .Q(
        \adder_stage3[2][5] ) );
  DFF_X1 \adder_stage3_reg[2][6]  ( .D(n9723), .CK(clk), .Q(
        \adder_stage3[2][6] ) );
  DFF_X1 \adder_stage3_reg[2][7]  ( .D(n9722), .CK(clk), .Q(
        \adder_stage3[2][7] ) );
  DFF_X1 \adder_stage3_reg[2][8]  ( .D(n9721), .CK(clk), .Q(
        \adder_stage3[2][8] ) );
  DFF_X1 \adder_stage3_reg[2][9]  ( .D(n9720), .CK(clk), .Q(
        \adder_stage3[2][9] ) );
  DFF_X1 \adder_stage3_reg[2][10]  ( .D(n9719), .CK(clk), .Q(
        \adder_stage3[2][10] ) );
  DFF_X1 \adder_stage3_reg[2][11]  ( .D(n9718), .CK(clk), .Q(
        \adder_stage3[2][11] ) );
  DFF_X1 \adder_stage3_reg[2][12]  ( .D(n9717), .CK(clk), .Q(
        \adder_stage3[2][12] ) );
  DFF_X1 \adder_stage3_reg[2][13]  ( .D(n9716), .CK(clk), .Q(
        \adder_stage3[2][13] ) );
  DFF_X1 \adder_stage3_reg[2][14]  ( .D(n9715), .CK(clk), .Q(
        \adder_stage3[2][14] ) );
  DFF_X1 \adder_stage3_reg[2][15]  ( .D(n9714), .CK(clk), .Q(
        \adder_stage3[2][15] ) );
  DFF_X1 \adder_stage3_reg[2][16]  ( .D(n9713), .CK(clk), .Q(
        \adder_stage3[2][16] ) );
  DFF_X1 \adder_stage3_reg[2][17]  ( .D(n9712), .CK(clk), .Q(
        \adder_stage3[2][17] ) );
  DFF_X1 \adder_stage3_reg[2][18]  ( .D(n9711), .CK(clk), .Q(
        \adder_stage3[2][18] ) );
  DFF_X1 \adder_stage3_reg[2][19]  ( .D(n9710), .CK(clk), .Q(
        \adder_stage3[2][19] ) );
  DFF_X1 \adder_stage3_reg[3][0]  ( .D(n9708), .CK(clk), .Q(
        \adder_stage3[3][0] ) );
  DFF_X1 \adder_stage3_reg[3][1]  ( .D(n9707), .CK(clk), .Q(
        \adder_stage3[3][1] ) );
  DFF_X1 \adder_stage3_reg[3][2]  ( .D(n9706), .CK(clk), .Q(
        \adder_stage3[3][2] ) );
  DFF_X1 \adder_stage3_reg[3][4]  ( .D(n9704), .CK(clk), .Q(
        \adder_stage3[3][4] ) );
  DFF_X1 \adder_stage3_reg[3][5]  ( .D(n9703), .CK(clk), .Q(
        \adder_stage3[3][5] ) );
  DFF_X1 \adder_stage3_reg[3][6]  ( .D(n9702), .CK(clk), .Q(
        \adder_stage3[3][6] ) );
  DFF_X1 \adder_stage3_reg[3][7]  ( .D(n9701), .CK(clk), .Q(
        \adder_stage3[3][7] ) );
  DFF_X1 \adder_stage3_reg[3][8]  ( .D(n9700), .CK(clk), .Q(
        \adder_stage3[3][8] ) );
  DFF_X1 \adder_stage3_reg[3][9]  ( .D(n9699), .CK(clk), .Q(
        \adder_stage3[3][9] ) );
  DFF_X1 \adder_stage3_reg[3][10]  ( .D(n9698), .CK(clk), .Q(
        \adder_stage3[3][10] ) );
  DFF_X1 \adder_stage3_reg[3][12]  ( .D(n9696), .CK(clk), .Q(
        \adder_stage3[3][12] ) );
  DFF_X1 \adder_stage3_reg[3][13]  ( .D(n9695), .CK(clk), .Q(
        \adder_stage3[3][13] ) );
  DFF_X1 \adder_stage3_reg[3][14]  ( .D(n9694), .CK(clk), .Q(
        \adder_stage3[3][14] ) );
  DFF_X1 \adder_stage3_reg[3][15]  ( .D(n9693), .CK(clk), .Q(
        \adder_stage3[3][15] ) );
  DFF_X1 \adder_stage3_reg[3][16]  ( .D(n9692), .CK(clk), .Q(
        \adder_stage3[3][16] ) );
  DFF_X1 \adder_stage3_reg[3][17]  ( .D(n9691), .CK(clk), .Q(
        \adder_stage3[3][17] ) );
  DFF_X1 \adder_stage3_reg[3][18]  ( .D(n9690), .CK(clk), .Q(
        \adder_stage3[3][18] ) );
  DFF_X1 \adder_stage3_reg[3][19]  ( .D(n9689), .CK(clk), .Q(
        \adder_stage3[3][19] ) );
  DFF_X1 \adder_stage3_reg[3][20]  ( .D(n9688), .CK(clk), .Q(
        \adder_stage3[3][20] ) );
  DFF_X1 \adder_stage4_reg[0][0]  ( .D(n9687), .CK(clk), .Q(
        \adder_stage4[0][0] ) );
  DFF_X1 \adder_stage4_reg[0][1]  ( .D(n9686), .CK(clk), .Q(
        \adder_stage4[0][1] ) );
  DFF_X1 \adder_stage4_reg[0][2]  ( .D(n9685), .CK(clk), .Q(
        \adder_stage4[0][2] ) );
  DFF_X1 \adder_stage4_reg[0][3]  ( .D(n9684), .CK(clk), .Q(
        \adder_stage4[0][3] ), .QN(n3417) );
  DFF_X1 \adder_stage4_reg[0][4]  ( .D(n9683), .CK(clk), .Q(
        \adder_stage4[0][4] ) );
  DFF_X1 \adder_stage4_reg[0][5]  ( .D(n9682), .CK(clk), .Q(
        \adder_stage4[0][5] ) );
  DFF_X1 \adder_stage4_reg[0][6]  ( .D(n9681), .CK(clk), .Q(
        \adder_stage4[0][6] ) );
  DFF_X1 \adder_stage4_reg[0][7]  ( .D(n9680), .CK(clk), .Q(
        \adder_stage4[0][7] ) );
  DFF_X1 \adder_stage4_reg[0][8]  ( .D(n9679), .CK(clk), .Q(
        \adder_stage4[0][8] ) );
  DFF_X1 \adder_stage4_reg[0][9]  ( .D(n9678), .CK(clk), .Q(
        \adder_stage4[0][9] ) );
  DFF_X1 \adder_stage4_reg[0][10]  ( .D(n9677), .CK(clk), .Q(
        \adder_stage4[0][10] ) );
  DFF_X1 \adder_stage4_reg[0][11]  ( .D(n9676), .CK(clk), .Q(
        \adder_stage4[0][11] ) );
  DFF_X1 \adder_stage4_reg[0][12]  ( .D(n9675), .CK(clk), .Q(
        \adder_stage4[0][12] ) );
  DFF_X1 \adder_stage4_reg[0][13]  ( .D(n9674), .CK(clk), .Q(
        \adder_stage4[0][13] ) );
  DFF_X1 \adder_stage4_reg[0][14]  ( .D(n9673), .CK(clk), .Q(
        \adder_stage4[0][14] ) );
  DFF_X1 \adder_stage4_reg[0][15]  ( .D(n9672), .CK(clk), .Q(
        \adder_stage4[0][15] ) );
  DFF_X1 \adder_stage4_reg[0][16]  ( .D(n9671), .CK(clk), .Q(
        \adder_stage4[0][16] ) );
  DFF_X1 \adder_stage4_reg[0][17]  ( .D(n9670), .CK(clk), .Q(
        \adder_stage4[0][17] ) );
  DFF_X1 \adder_stage4_reg[0][18]  ( .D(n9669), .CK(clk), .Q(
        \adder_stage4[0][18] ) );
  DFF_X1 \adder_stage4_reg[0][19]  ( .D(n9668), .CK(clk), .Q(
        \adder_stage4[0][19] ) );
  DFF_X1 \adder_stage4_reg[0][20]  ( .D(n9667), .CK(clk), .Q(
        \adder_stage4[0][20] ) );
  DFF_X1 \adder_stage4_reg[1][0]  ( .D(n9666), .CK(clk), .Q(
        \adder_stage4[1][0] ) );
  DFF_X1 \adder_stage4_reg[1][1]  ( .D(n9665), .CK(clk), .Q(
        \adder_stage4[1][1] ) );
  DFF_X1 \adder_stage4_reg[1][2]  ( .D(n9664), .CK(clk), .Q(
        \adder_stage4[1][2] ) );
  DFF_X1 \adder_stage4_reg[1][3]  ( .D(n9663), .CK(clk), .Q(
        \adder_stage4[1][3] ), .QN(n3418) );
  DFF_X1 \adder_stage4_reg[1][4]  ( .D(n9662), .CK(clk), .Q(
        \adder_stage4[1][4] ) );
  DFF_X1 \adder_stage4_reg[1][5]  ( .D(n9661), .CK(clk), .Q(
        \adder_stage4[1][5] ) );
  DFF_X1 \adder_stage4_reg[1][6]  ( .D(n9660), .CK(clk), .Q(
        \adder_stage4[1][6] ) );
  DFF_X1 \adder_stage4_reg[1][7]  ( .D(n9659), .CK(clk), .Q(
        \adder_stage4[1][7] ) );
  DFF_X1 \adder_stage4_reg[1][8]  ( .D(n9658), .CK(clk), .Q(
        \adder_stage4[1][8] ) );
  DFF_X1 \adder_stage4_reg[1][9]  ( .D(n9657), .CK(clk), .Q(
        \adder_stage4[1][9] ) );
  DFF_X1 \adder_stage4_reg[1][10]  ( .D(n9656), .CK(clk), .Q(
        \adder_stage4[1][10] ) );
  DFF_X1 \adder_stage4_reg[1][11]  ( .D(n9655), .CK(clk), .Q(
        \adder_stage4[1][11] ) );
  DFF_X1 \adder_stage4_reg[1][12]  ( .D(n9654), .CK(clk), .Q(
        \adder_stage4[1][12] ) );
  DFF_X1 \adder_stage4_reg[1][13]  ( .D(n9653), .CK(clk), .Q(
        \adder_stage4[1][13] ) );
  DFF_X1 \adder_stage4_reg[1][14]  ( .D(n9652), .CK(clk), .Q(
        \adder_stage4[1][14] ) );
  DFF_X1 \adder_stage4_reg[1][15]  ( .D(n9651), .CK(clk), .Q(
        \adder_stage4[1][15] ) );
  DFF_X1 \adder_stage4_reg[1][16]  ( .D(n9650), .CK(clk), .Q(
        \adder_stage4[1][16] ) );
  DFF_X1 \adder_stage4_reg[1][17]  ( .D(n9649), .CK(clk), .Q(
        \adder_stage4[1][17] ) );
  DFF_X1 \adder_stage4_reg[1][18]  ( .D(n9648), .CK(clk), .Q(
        \adder_stage4[1][18] ) );
  DFF_X1 \adder_stage4_reg[1][19]  ( .D(n9647), .CK(clk), .Q(
        \adder_stage4[1][19] ) );
  DFF_X1 \adder_stage4_reg[1][20]  ( .D(n9646), .CK(clk), .Q(
        \adder_stage4[1][20] ) );
  conv_128_32_opt_DW_mult_pipe_J1_0 \multiplier[31].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8903), .tc(1'b1), .a({\xmem_data[31][7] , 
        \xmem_data[31][6] , \xmem_data[31][5] , \xmem_data[31][4] , 
        \xmem_data[31][3] , \xmem_data[31][2] , \xmem_data[31][1] , 
        \xmem_data[31][0] }), .b({\fmem_data[31][7] , \fmem_data[31][6] , 
        \fmem_data[31][5] , \fmem_data[31][4] , \fmem_data[31][3] , 
        \fmem_data[31][2] , \fmem_data[31][1] , \fmem_data[31][0] }), 
        .product({\x_mult_f_int[31][15] , \x_mult_f_int[31][14] , 
        \x_mult_f_int[31][13] , \x_mult_f_int[31][12] , \x_mult_f_int[31][11] , 
        \x_mult_f_int[31][10] , \x_mult_f_int[31][9] , \x_mult_f_int[31][8] , 
        \x_mult_f_int[31][7] , \x_mult_f_int[31][6] , \x_mult_f_int[31][5] , 
        \x_mult_f_int[31][4] , \x_mult_f_int[31][3] , \x_mult_f_int[31][2] , 
        \x_mult_f_int[31][1] , \x_mult_f_int[31][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_1 \multiplier[30].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8901), .tc(1'b1), .a({\xmem_data[30][7] , 
        \xmem_data[30][6] , \xmem_data[30][5] , \xmem_data[30][4] , 
        \xmem_data[30][3] , \xmem_data[30][2] , \xmem_data[30][1] , 
        \xmem_data[30][0] }), .b({\fmem_data[30][7] , \fmem_data[30][6] , 
        \fmem_data[30][5] , \fmem_data[30][4] , \fmem_data[30][3] , 
        \fmem_data[30][2] , \fmem_data[30][1] , \fmem_data[30][0] }), 
        .product({\x_mult_f_int[30][15] , \x_mult_f_int[30][14] , 
        \x_mult_f_int[30][13] , \x_mult_f_int[30][12] , \x_mult_f_int[30][11] , 
        \x_mult_f_int[30][10] , \x_mult_f_int[30][9] , \x_mult_f_int[30][8] , 
        \x_mult_f_int[30][7] , \x_mult_f_int[30][6] , \x_mult_f_int[30][5] , 
        \x_mult_f_int[30][4] , \x_mult_f_int[30][3] , \x_mult_f_int[30][2] , 
        \x_mult_f_int[30][1] , \x_mult_f_int[30][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_2 \multiplier[29].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8901), .tc(1'b1), .a({\xmem_data[29][7] , 
        \xmem_data[29][6] , \xmem_data[29][5] , \xmem_data[29][4] , 
        \xmem_data[29][3] , \xmem_data[29][2] , \xmem_data[29][1] , 
        \xmem_data[29][0] }), .b({\fmem_data[29][7] , \fmem_data[29][6] , 
        \fmem_data[29][5] , \fmem_data[29][4] , \fmem_data[29][3] , 
        \fmem_data[29][2] , \fmem_data[29][1] , \fmem_data[29][0] }), 
        .product({\x_mult_f_int[29][15] , \x_mult_f_int[29][14] , 
        \x_mult_f_int[29][13] , \x_mult_f_int[29][12] , \x_mult_f_int[29][11] , 
        \x_mult_f_int[29][10] , \x_mult_f_int[29][9] , \x_mult_f_int[29][8] , 
        \x_mult_f_int[29][7] , \x_mult_f_int[29][6] , \x_mult_f_int[29][5] , 
        \x_mult_f_int[29][4] , \x_mult_f_int[29][3] , \x_mult_f_int[29][2] , 
        \x_mult_f_int[29][1] , \x_mult_f_int[29][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_3 \multiplier[28].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8911), .tc(1'b1), .a({\xmem_data[28][7] , 
        \xmem_data[28][6] , \xmem_data[28][5] , \xmem_data[28][4] , 
        \xmem_data[28][3] , \xmem_data[28][2] , \xmem_data[28][1] , 
        \xmem_data[28][0] }), .b({\fmem_data[28][7] , \fmem_data[28][6] , 
        \fmem_data[28][5] , \fmem_data[28][4] , \fmem_data[28][3] , 
        \fmem_data[28][2] , \fmem_data[28][1] , \fmem_data[28][0] }), 
        .product({\x_mult_f_int[28][15] , \x_mult_f_int[28][14] , 
        \x_mult_f_int[28][13] , \x_mult_f_int[28][12] , \x_mult_f_int[28][11] , 
        \x_mult_f_int[28][10] , \x_mult_f_int[28][9] , \x_mult_f_int[28][8] , 
        \x_mult_f_int[28][7] , \x_mult_f_int[28][6] , \x_mult_f_int[28][5] , 
        \x_mult_f_int[28][4] , \x_mult_f_int[28][3] , \x_mult_f_int[28][2] , 
        \x_mult_f_int[28][1] , \x_mult_f_int[28][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_4 \multiplier[27].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8909), .tc(1'b1), .a({\xmem_data[27][7] , 
        \xmem_data[27][6] , \xmem_data[27][5] , \xmem_data[27][4] , 
        \xmem_data[27][3] , \xmem_data[27][2] , \xmem_data[27][1] , 
        \xmem_data[27][0] }), .b({\fmem_data[27][7] , \fmem_data[27][6] , 
        \fmem_data[27][5] , \fmem_data[27][4] , \fmem_data[27][3] , 
        \fmem_data[27][2] , \fmem_data[27][1] , \fmem_data[27][0] }), 
        .product({\x_mult_f_int[27][15] , \x_mult_f_int[27][14] , 
        \x_mult_f_int[27][13] , \x_mult_f_int[27][12] , \x_mult_f_int[27][11] , 
        \x_mult_f_int[27][10] , \x_mult_f_int[27][9] , \x_mult_f_int[27][8] , 
        \x_mult_f_int[27][7] , \x_mult_f_int[27][6] , \x_mult_f_int[27][5] , 
        \x_mult_f_int[27][4] , \x_mult_f_int[27][3] , \x_mult_f_int[27][2] , 
        \x_mult_f_int[27][1] , \x_mult_f_int[27][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_5 \multiplier[26].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8901), .tc(1'b1), .a({\xmem_data[26][7] , 
        \xmem_data[26][6] , \xmem_data[26][5] , \xmem_data[26][4] , 
        \xmem_data[26][3] , \xmem_data[26][2] , \xmem_data[26][1] , 
        \xmem_data[26][0] }), .b({\fmem_data[26][7] , \fmem_data[26][6] , 
        \fmem_data[26][5] , \fmem_data[26][4] , \fmem_data[26][3] , 
        \fmem_data[26][2] , \fmem_data[26][1] , \fmem_data[26][0] }), 
        .product({\x_mult_f_int[26][15] , \x_mult_f_int[26][14] , 
        \x_mult_f_int[26][13] , \x_mult_f_int[26][12] , \x_mult_f_int[26][11] , 
        \x_mult_f_int[26][10] , \x_mult_f_int[26][9] , \x_mult_f_int[26][8] , 
        \x_mult_f_int[26][7] , \x_mult_f_int[26][6] , \x_mult_f_int[26][5] , 
        \x_mult_f_int[26][4] , \x_mult_f_int[26][3] , \x_mult_f_int[26][2] , 
        \x_mult_f_int[26][1] , \x_mult_f_int[26][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_6 \multiplier[25].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8911), .tc(1'b1), .a({\xmem_data[25][7] , 
        \xmem_data[25][6] , \xmem_data[25][5] , \xmem_data[25][4] , 
        \xmem_data[25][3] , \xmem_data[25][2] , \xmem_data[25][1] , 
        \xmem_data[25][0] }), .b({\fmem_data[25][7] , \fmem_data[25][6] , 
        \fmem_data[25][5] , \fmem_data[25][4] , \fmem_data[25][3] , 
        \fmem_data[25][2] , \fmem_data[25][1] , \fmem_data[25][0] }), 
        .product({\x_mult_f_int[25][15] , \x_mult_f_int[25][14] , 
        \x_mult_f_int[25][13] , \x_mult_f_int[25][12] , \x_mult_f_int[25][11] , 
        \x_mult_f_int[25][10] , \x_mult_f_int[25][9] , \x_mult_f_int[25][8] , 
        \x_mult_f_int[25][7] , \x_mult_f_int[25][6] , \x_mult_f_int[25][5] , 
        \x_mult_f_int[25][4] , \x_mult_f_int[25][3] , \x_mult_f_int[25][2] , 
        \x_mult_f_int[25][1] , \x_mult_f_int[25][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_7 \multiplier[24].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8903), .tc(1'b1), .a({\xmem_data[24][7] , 
        \xmem_data[24][6] , \xmem_data[24][5] , \xmem_data[24][4] , 
        \xmem_data[24][3] , \xmem_data[24][2] , \xmem_data[24][1] , 
        \xmem_data[24][0] }), .b({\fmem_data[24][7] , \fmem_data[24][6] , 
        \fmem_data[24][5] , \fmem_data[24][4] , \fmem_data[24][3] , 
        \fmem_data[24][2] , \fmem_data[24][1] , \fmem_data[24][0] }), 
        .product({\x_mult_f_int[24][15] , \x_mult_f_int[24][14] , 
        \x_mult_f_int[24][13] , \x_mult_f_int[24][12] , \x_mult_f_int[24][11] , 
        \x_mult_f_int[24][10] , \x_mult_f_int[24][9] , \x_mult_f_int[24][8] , 
        \x_mult_f_int[24][7] , \x_mult_f_int[24][6] , \x_mult_f_int[24][5] , 
        \x_mult_f_int[24][4] , \x_mult_f_int[24][3] , \x_mult_f_int[24][2] , 
        \x_mult_f_int[24][1] , \x_mult_f_int[24][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_8 \multiplier[23].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n3650), .tc(1'b1), .a({\xmem_data[23][7] , 
        \xmem_data[23][6] , \xmem_data[23][5] , \xmem_data[23][4] , 
        \xmem_data[23][3] , \xmem_data[23][2] , \xmem_data[23][1] , 
        \xmem_data[23][0] }), .b({\fmem_data[23][7] , \fmem_data[23][6] , 
        \fmem_data[23][5] , \fmem_data[23][4] , \fmem_data[23][3] , 
        \fmem_data[23][2] , \fmem_data[23][1] , \fmem_data[23][0] }), 
        .product({\x_mult_f_int[23][15] , \x_mult_f_int[23][14] , 
        \x_mult_f_int[23][13] , \x_mult_f_int[23][12] , \x_mult_f_int[23][11] , 
        \x_mult_f_int[23][10] , \x_mult_f_int[23][9] , \x_mult_f_int[23][8] , 
        \x_mult_f_int[23][7] , \x_mult_f_int[23][6] , \x_mult_f_int[23][5] , 
        \x_mult_f_int[23][4] , \x_mult_f_int[23][3] , \x_mult_f_int[23][2] , 
        \x_mult_f_int[23][1] , \x_mult_f_int[23][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_9 \multiplier[22].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8903), .tc(1'b1), .a({\xmem_data[22][7] , 
        \xmem_data[22][6] , \xmem_data[22][5] , \xmem_data[22][4] , 
        \xmem_data[22][3] , \xmem_data[22][2] , \xmem_data[22][1] , 
        \xmem_data[22][0] }), .b({\fmem_data[22][7] , \fmem_data[22][6] , 
        \fmem_data[22][5] , \fmem_data[22][4] , \fmem_data[22][3] , 
        \fmem_data[22][2] , \fmem_data[22][1] , \fmem_data[22][0] }), 
        .product({\x_mult_f_int[22][15] , \x_mult_f_int[22][14] , 
        \x_mult_f_int[22][13] , \x_mult_f_int[22][12] , \x_mult_f_int[22][11] , 
        \x_mult_f_int[22][10] , \x_mult_f_int[22][9] , \x_mult_f_int[22][8] , 
        \x_mult_f_int[22][7] , \x_mult_f_int[22][6] , \x_mult_f_int[22][5] , 
        \x_mult_f_int[22][4] , \x_mult_f_int[22][3] , \x_mult_f_int[22][2] , 
        \x_mult_f_int[22][1] , \x_mult_f_int[22][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_10 \multiplier[21].x_f_mult_inst  ( .clk(clk), .rst_n(n8905), .en(n8910), .tc(1'b1), .a({\xmem_data[21][7] , 
        \xmem_data[21][6] , \xmem_data[21][5] , \xmem_data[21][4] , 
        \xmem_data[21][3] , \xmem_data[21][2] , \xmem_data[21][1] , 
        \xmem_data[21][0] }), .b({\fmem_data[21][7] , \fmem_data[21][6] , 
        \fmem_data[21][5] , \fmem_data[21][4] , \fmem_data[21][3] , 
        \fmem_data[21][2] , \fmem_data[21][1] , \fmem_data[21][0] }), 
        .product({\x_mult_f_int[21][15] , \x_mult_f_int[21][14] , 
        \x_mult_f_int[21][13] , \x_mult_f_int[21][12] , \x_mult_f_int[21][11] , 
        \x_mult_f_int[21][10] , \x_mult_f_int[21][9] , \x_mult_f_int[21][8] , 
        \x_mult_f_int[21][7] , \x_mult_f_int[21][6] , \x_mult_f_int[21][5] , 
        \x_mult_f_int[21][4] , \x_mult_f_int[21][3] , \x_mult_f_int[21][2] , 
        \x_mult_f_int[21][1] , \x_mult_f_int[21][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_11 \multiplier[20].x_f_mult_inst  ( .clk(clk), .rst_n(n8905), .en(n8909), .tc(1'b1), .a({\xmem_data[20][7] , 
        \xmem_data[20][6] , \xmem_data[20][5] , \xmem_data[20][4] , 
        \xmem_data[20][3] , \xmem_data[20][2] , \xmem_data[20][1] , 
        \xmem_data[20][0] }), .b({\fmem_data[20][7] , \fmem_data[20][6] , 
        \fmem_data[20][5] , \fmem_data[20][4] , \fmem_data[20][3] , 
        \fmem_data[20][2] , \fmem_data[20][1] , \fmem_data[20][0] }), 
        .product({\x_mult_f_int[20][15] , \x_mult_f_int[20][14] , 
        \x_mult_f_int[20][13] , \x_mult_f_int[20][12] , \x_mult_f_int[20][11] , 
        \x_mult_f_int[20][10] , \x_mult_f_int[20][9] , \x_mult_f_int[20][8] , 
        \x_mult_f_int[20][7] , \x_mult_f_int[20][6] , \x_mult_f_int[20][5] , 
        \x_mult_f_int[20][4] , \x_mult_f_int[20][3] , \x_mult_f_int[20][2] , 
        \x_mult_f_int[20][1] , \x_mult_f_int[20][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_12 \multiplier[19].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8908), .tc(1'b1), .a({\xmem_data[19][7] , 
        \xmem_data[19][6] , \xmem_data[19][5] , \xmem_data[19][4] , 
        \xmem_data[19][3] , \xmem_data[19][2] , \xmem_data[19][1] , 
        \xmem_data[19][0] }), .b({\fmem_data[19][7] , \fmem_data[19][6] , 
        \fmem_data[19][5] , \fmem_data[19][4] , \fmem_data[19][3] , 
        \fmem_data[19][2] , \fmem_data[19][1] , \fmem_data[19][0] }), 
        .product({\x_mult_f_int[19][15] , \x_mult_f_int[19][14] , 
        \x_mult_f_int[19][13] , \x_mult_f_int[19][12] , \x_mult_f_int[19][11] , 
        \x_mult_f_int[19][10] , \x_mult_f_int[19][9] , \x_mult_f_int[19][8] , 
        \x_mult_f_int[19][7] , \x_mult_f_int[19][6] , \x_mult_f_int[19][5] , 
        \x_mult_f_int[19][4] , \x_mult_f_int[19][3] , \x_mult_f_int[19][2] , 
        \x_mult_f_int[19][1] , \x_mult_f_int[19][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_13 \multiplier[18].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8908), .tc(1'b1), .a({\xmem_data[18][7] , 
        \xmem_data[18][6] , \xmem_data[18][5] , \xmem_data[18][4] , 
        \xmem_data[18][3] , \xmem_data[18][2] , \xmem_data[18][1] , 
        \xmem_data[18][0] }), .b({\fmem_data[18][7] , \fmem_data[18][6] , 
        \fmem_data[18][5] , \fmem_data[18][4] , \fmem_data[18][3] , 
        \fmem_data[18][2] , \fmem_data[18][1] , \fmem_data[18][0] }), 
        .product({\x_mult_f_int[18][15] , \x_mult_f_int[18][14] , 
        \x_mult_f_int[18][13] , \x_mult_f_int[18][12] , \x_mult_f_int[18][11] , 
        \x_mult_f_int[18][10] , \x_mult_f_int[18][9] , \x_mult_f_int[18][8] , 
        \x_mult_f_int[18][7] , \x_mult_f_int[18][6] , \x_mult_f_int[18][5] , 
        \x_mult_f_int[18][4] , \x_mult_f_int[18][3] , \x_mult_f_int[18][2] , 
        \x_mult_f_int[18][1] , \x_mult_f_int[18][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_14 \multiplier[17].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8903), .tc(1'b1), .a({\xmem_data[17][7] , 
        \xmem_data[17][6] , \xmem_data[17][5] , \xmem_data[17][4] , 
        \xmem_data[17][3] , \xmem_data[17][2] , \xmem_data[17][1] , 
        \xmem_data[17][0] }), .b({\fmem_data[17][7] , \fmem_data[17][6] , 
        \fmem_data[17][5] , \fmem_data[17][4] , \fmem_data[17][3] , 
        \fmem_data[17][2] , \fmem_data[17][1] , \fmem_data[17][0] }), 
        .product({\x_mult_f_int[17][15] , \x_mult_f_int[17][14] , 
        \x_mult_f_int[17][13] , \x_mult_f_int[17][12] , \x_mult_f_int[17][11] , 
        \x_mult_f_int[17][10] , \x_mult_f_int[17][9] , \x_mult_f_int[17][8] , 
        \x_mult_f_int[17][7] , \x_mult_f_int[17][6] , \x_mult_f_int[17][5] , 
        \x_mult_f_int[17][4] , \x_mult_f_int[17][3] , \x_mult_f_int[17][2] , 
        \x_mult_f_int[17][1] , \x_mult_f_int[17][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_15 \multiplier[16].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n3650), .tc(1'b1), .a({\xmem_data[16][7] , 
        \xmem_data[16][6] , \xmem_data[16][5] , \xmem_data[16][4] , 
        \xmem_data[16][3] , \xmem_data[16][2] , \xmem_data[16][1] , 
        \xmem_data[16][0] }), .b({\fmem_data[16][7] , \fmem_data[16][6] , 
        \fmem_data[16][5] , \fmem_data[16][4] , \fmem_data[16][3] , 
        \fmem_data[16][2] , \fmem_data[16][1] , \fmem_data[16][0] }), 
        .product({\x_mult_f_int[16][15] , \x_mult_f_int[16][14] , 
        \x_mult_f_int[16][13] , \x_mult_f_int[16][12] , \x_mult_f_int[16][11] , 
        \x_mult_f_int[16][10] , \x_mult_f_int[16][9] , \x_mult_f_int[16][8] , 
        \x_mult_f_int[16][7] , \x_mult_f_int[16][6] , \x_mult_f_int[16][5] , 
        \x_mult_f_int[16][4] , \x_mult_f_int[16][3] , \x_mult_f_int[16][2] , 
        \x_mult_f_int[16][1] , \x_mult_f_int[16][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_16 \multiplier[15].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8901), .tc(1'b1), .a({\xmem_data[15][7] , 
        \xmem_data[15][6] , \xmem_data[15][5] , \xmem_data[15][4] , 
        \xmem_data[15][3] , \xmem_data[15][2] , \xmem_data[15][1] , 
        \xmem_data[15][0] }), .b({\fmem_data[15][7] , \fmem_data[15][6] , 
        \fmem_data[15][5] , \fmem_data[15][4] , \fmem_data[15][3] , 
        \fmem_data[15][2] , \fmem_data[15][1] , \fmem_data[15][0] }), 
        .product({\x_mult_f_int[15][15] , \x_mult_f_int[15][14] , 
        \x_mult_f_int[15][13] , \x_mult_f_int[15][12] , \x_mult_f_int[15][11] , 
        \x_mult_f_int[15][10] , \x_mult_f_int[15][9] , \x_mult_f_int[15][8] , 
        \x_mult_f_int[15][7] , \x_mult_f_int[15][6] , \x_mult_f_int[15][5] , 
        \x_mult_f_int[15][4] , \x_mult_f_int[15][3] , \x_mult_f_int[15][2] , 
        \x_mult_f_int[15][1] , \x_mult_f_int[15][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_17 \multiplier[14].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8903), .tc(1'b1), .a({\xmem_data[14][7] , 
        \xmem_data[14][6] , \xmem_data[14][5] , \xmem_data[14][4] , 
        \xmem_data[14][3] , \xmem_data[14][2] , \xmem_data[14][1] , 
        \xmem_data[14][0] }), .b({\fmem_data[14][7] , \fmem_data[14][6] , 
        \fmem_data[14][5] , \fmem_data[14][4] , \fmem_data[14][3] , 
        \fmem_data[14][2] , \fmem_data[14][1] , \fmem_data[14][0] }), 
        .product({\x_mult_f_int[14][15] , \x_mult_f_int[14][14] , 
        \x_mult_f_int[14][13] , \x_mult_f_int[14][12] , \x_mult_f_int[14][11] , 
        \x_mult_f_int[14][10] , \x_mult_f_int[14][9] , \x_mult_f_int[14][8] , 
        \x_mult_f_int[14][7] , \x_mult_f_int[14][6] , \x_mult_f_int[14][5] , 
        \x_mult_f_int[14][4] , \x_mult_f_int[14][3] , \x_mult_f_int[14][2] , 
        \x_mult_f_int[14][1] , \x_mult_f_int[14][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_18 \multiplier[13].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8902), .tc(1'b1), .a({\xmem_data[13][7] , 
        \xmem_data[13][6] , \xmem_data[13][5] , \xmem_data[13][4] , 
        \xmem_data[13][3] , \xmem_data[13][2] , \xmem_data[13][1] , 
        \xmem_data[13][0] }), .b({\fmem_data[13][7] , \fmem_data[13][6] , 
        \fmem_data[13][5] , \fmem_data[13][4] , \fmem_data[13][3] , 
        \fmem_data[13][2] , \fmem_data[13][1] , \fmem_data[13][0] }), 
        .product({\x_mult_f_int[13][15] , \x_mult_f_int[13][14] , 
        \x_mult_f_int[13][13] , \x_mult_f_int[13][12] , \x_mult_f_int[13][11] , 
        \x_mult_f_int[13][10] , \x_mult_f_int[13][9] , \x_mult_f_int[13][8] , 
        \x_mult_f_int[13][7] , \x_mult_f_int[13][6] , \x_mult_f_int[13][5] , 
        \x_mult_f_int[13][4] , \x_mult_f_int[13][3] , \x_mult_f_int[13][2] , 
        \x_mult_f_int[13][1] , \x_mult_f_int[13][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_19 \multiplier[12].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8902), .tc(1'b1), .a({\xmem_data[12][7] , 
        \xmem_data[12][6] , \xmem_data[12][5] , \xmem_data[12][4] , 
        \xmem_data[12][3] , \xmem_data[12][2] , \xmem_data[12][1] , 
        \xmem_data[12][0] }), .b({\fmem_data[12][7] , \fmem_data[12][6] , 
        \fmem_data[12][5] , \fmem_data[12][4] , \fmem_data[12][3] , 
        \fmem_data[12][2] , \fmem_data[12][1] , \fmem_data[12][0] }), 
        .product({\x_mult_f_int[12][15] , \x_mult_f_int[12][14] , 
        \x_mult_f_int[12][13] , \x_mult_f_int[12][12] , \x_mult_f_int[12][11] , 
        \x_mult_f_int[12][10] , \x_mult_f_int[12][9] , \x_mult_f_int[12][8] , 
        \x_mult_f_int[12][7] , \x_mult_f_int[12][6] , \x_mult_f_int[12][5] , 
        \x_mult_f_int[12][4] , \x_mult_f_int[12][3] , \x_mult_f_int[12][2] , 
        \x_mult_f_int[12][1] , \x_mult_f_int[12][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_20 \multiplier[11].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n8901), .tc(1'b1), .a({\xmem_data[11][7] , 
        \xmem_data[11][6] , \xmem_data[11][5] , \xmem_data[11][4] , 
        \xmem_data[11][3] , \xmem_data[11][2] , \xmem_data[11][1] , 
        \xmem_data[11][0] }), .b({\fmem_data[11][7] , \fmem_data[11][6] , 
        \fmem_data[11][5] , \fmem_data[11][4] , \fmem_data[11][3] , 
        \fmem_data[11][2] , \fmem_data[11][1] , \fmem_data[11][0] }), 
        .product({\x_mult_f_int[11][15] , \x_mult_f_int[11][14] , 
        \x_mult_f_int[11][13] , \x_mult_f_int[11][12] , \x_mult_f_int[11][11] , 
        \x_mult_f_int[11][10] , \x_mult_f_int[11][9] , \x_mult_f_int[11][8] , 
        \x_mult_f_int[11][7] , \x_mult_f_int[11][6] , \x_mult_f_int[11][5] , 
        \x_mult_f_int[11][4] , \x_mult_f_int[11][3] , \x_mult_f_int[11][2] , 
        \x_mult_f_int[11][1] , \x_mult_f_int[11][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_21 \multiplier[10].x_f_mult_inst  ( .clk(clk), .rst_n(n8906), .en(n3650), .tc(1'b1), .a({\xmem_data[10][7] , 
        \xmem_data[10][6] , \xmem_data[10][5] , \xmem_data[10][4] , 
        \xmem_data[10][3] , \xmem_data[10][2] , \xmem_data[10][1] , 
        \xmem_data[10][0] }), .b({\fmem_data[10][7] , \fmem_data[10][6] , 
        \fmem_data[10][5] , \fmem_data[10][4] , \fmem_data[10][3] , 
        \fmem_data[10][2] , \fmem_data[10][1] , \fmem_data[10][0] }), 
        .product({\x_mult_f_int[10][15] , \x_mult_f_int[10][14] , 
        \x_mult_f_int[10][13] , \x_mult_f_int[10][12] , \x_mult_f_int[10][11] , 
        \x_mult_f_int[10][10] , \x_mult_f_int[10][9] , \x_mult_f_int[10][8] , 
        \x_mult_f_int[10][7] , \x_mult_f_int[10][6] , \x_mult_f_int[10][5] , 
        \x_mult_f_int[10][4] , \x_mult_f_int[10][3] , \x_mult_f_int[10][2] , 
        \x_mult_f_int[10][1] , \x_mult_f_int[10][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_22 \multiplier[9].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8906), .en(n8902), .tc(1'b1), .a({\xmem_data[9][7] , 
        \xmem_data[9][6] , \xmem_data[9][5] , \xmem_data[9][4] , 
        \xmem_data[9][3] , \xmem_data[9][2] , \xmem_data[9][1] , 
        \xmem_data[9][0] }), .b({\fmem_data[9][7] , \fmem_data[9][6] , 
        \fmem_data[9][5] , \fmem_data[9][4] , \fmem_data[9][3] , 
        \fmem_data[9][2] , \fmem_data[9][1] , \fmem_data[9][0] }), .product({
        \x_mult_f_int[9][15] , \x_mult_f_int[9][14] , \x_mult_f_int[9][13] , 
        \x_mult_f_int[9][12] , \x_mult_f_int[9][11] , \x_mult_f_int[9][10] , 
        \x_mult_f_int[9][9] , \x_mult_f_int[9][8] , \x_mult_f_int[9][7] , 
        \x_mult_f_int[9][6] , \x_mult_f_int[9][5] , \x_mult_f_int[9][4] , 
        \x_mult_f_int[9][3] , \x_mult_f_int[9][2] , \x_mult_f_int[9][1] , 
        \x_mult_f_int[9][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_23 \multiplier[8].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8906), .en(n8902), .tc(1'b1), .a({\xmem_data[8][7] , 
        \xmem_data[8][6] , \xmem_data[8][5] , \xmem_data[8][4] , 
        \xmem_data[8][3] , \xmem_data[8][2] , \xmem_data[8][1] , 
        \xmem_data[8][0] }), .b({\fmem_data[8][7] , \fmem_data[8][6] , 
        \fmem_data[8][5] , \fmem_data[8][4] , \fmem_data[8][3] , 
        \fmem_data[8][2] , \fmem_data[8][1] , \fmem_data[8][0] }), .product({
        \x_mult_f_int[8][15] , \x_mult_f_int[8][14] , \x_mult_f_int[8][13] , 
        \x_mult_f_int[8][12] , \x_mult_f_int[8][11] , \x_mult_f_int[8][10] , 
        \x_mult_f_int[8][9] , \x_mult_f_int[8][8] , \x_mult_f_int[8][7] , 
        \x_mult_f_int[8][6] , \x_mult_f_int[8][5] , \x_mult_f_int[8][4] , 
        \x_mult_f_int[8][3] , \x_mult_f_int[8][2] , \x_mult_f_int[8][1] , 
        \x_mult_f_int[8][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_24 \multiplier[7].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n8902), .tc(1'b1), .a({\xmem_data[7][7] , 
        \xmem_data[7][6] , \xmem_data[7][5] , \xmem_data[7][4] , 
        \xmem_data[7][3] , \xmem_data[7][2] , \xmem_data[7][1] , 
        \xmem_data[7][0] }), .b({\fmem_data[7][7] , \fmem_data[7][6] , 
        \fmem_data[7][5] , \fmem_data[7][4] , \fmem_data[7][3] , 
        \fmem_data[7][2] , \fmem_data[7][1] , \fmem_data[7][0] }), .product({
        \x_mult_f_int[7][15] , \x_mult_f_int[7][14] , \x_mult_f_int[7][13] , 
        \x_mult_f_int[7][12] , \x_mult_f_int[7][11] , \x_mult_f_int[7][10] , 
        \x_mult_f_int[7][9] , \x_mult_f_int[7][8] , \x_mult_f_int[7][7] , 
        \x_mult_f_int[7][6] , \x_mult_f_int[7][5] , \x_mult_f_int[7][4] , 
        \x_mult_f_int[7][3] , \x_mult_f_int[7][2] , \x_mult_f_int[7][1] , 
        \x_mult_f_int[7][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_25 \multiplier[6].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n8903), .tc(1'b1), .a({\xmem_data[6][7] , 
        \xmem_data[6][6] , \xmem_data[6][5] , \xmem_data[6][4] , 
        \xmem_data[6][3] , \xmem_data[6][2] , \xmem_data[6][1] , 
        \xmem_data[6][0] }), .b({\fmem_data[6][7] , \fmem_data[6][6] , 
        \fmem_data[6][5] , \fmem_data[6][4] , \fmem_data[6][3] , 
        \fmem_data[6][2] , \fmem_data[6][1] , \fmem_data[6][0] }), .product({
        \x_mult_f_int[6][15] , \x_mult_f_int[6][14] , \x_mult_f_int[6][13] , 
        \x_mult_f_int[6][12] , \x_mult_f_int[6][11] , \x_mult_f_int[6][10] , 
        \x_mult_f_int[6][9] , \x_mult_f_int[6][8] , \x_mult_f_int[6][7] , 
        \x_mult_f_int[6][6] , \x_mult_f_int[6][5] , \x_mult_f_int[6][4] , 
        \x_mult_f_int[6][3] , \x_mult_f_int[6][2] , \x_mult_f_int[6][1] , 
        \x_mult_f_int[6][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_26 \multiplier[5].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n3650), .tc(1'b1), .a({\xmem_data[5][7] , 
        \xmem_data[5][6] , \xmem_data[5][5] , \xmem_data[5][4] , 
        \xmem_data[5][3] , \xmem_data[5][2] , \xmem_data[5][1] , 
        \xmem_data[5][0] }), .b({\fmem_data[5][7] , \fmem_data[5][6] , 
        \fmem_data[5][5] , \fmem_data[5][4] , \fmem_data[5][3] , 
        \fmem_data[5][2] , \fmem_data[5][1] , \fmem_data[5][0] }), .product({
        \x_mult_f_int[5][15] , \x_mult_f_int[5][14] , \x_mult_f_int[5][13] , 
        \x_mult_f_int[5][12] , \x_mult_f_int[5][11] , \x_mult_f_int[5][10] , 
        \x_mult_f_int[5][9] , \x_mult_f_int[5][8] , \x_mult_f_int[5][7] , 
        \x_mult_f_int[5][6] , \x_mult_f_int[5][5] , \x_mult_f_int[5][4] , 
        \x_mult_f_int[5][3] , \x_mult_f_int[5][2] , \x_mult_f_int[5][1] , 
        \x_mult_f_int[5][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_27 \multiplier[4].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n8901), .tc(1'b1), .a({\xmem_data[4][7] , 
        \xmem_data[4][6] , \xmem_data[4][5] , \xmem_data[4][4] , 
        \xmem_data[4][3] , \xmem_data[4][2] , \xmem_data[4][1] , 
        \xmem_data[4][0] }), .b({\fmem_data[4][7] , \fmem_data[4][6] , 
        \fmem_data[4][5] , \fmem_data[4][4] , \fmem_data[4][3] , 
        \fmem_data[4][2] , \fmem_data[4][1] , \fmem_data[4][0] }), .product({
        \x_mult_f_int[4][15] , \x_mult_f_int[4][14] , \x_mult_f_int[4][13] , 
        \x_mult_f_int[4][12] , \x_mult_f_int[4][11] , \x_mult_f_int[4][10] , 
        \x_mult_f_int[4][9] , \x_mult_f_int[4][8] , \x_mult_f_int[4][7] , 
        \x_mult_f_int[4][6] , \x_mult_f_int[4][5] , \x_mult_f_int[4][4] , 
        \x_mult_f_int[4][3] , \x_mult_f_int[4][2] , \x_mult_f_int[4][1] , 
        \x_mult_f_int[4][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_28 \multiplier[3].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n8902), .tc(1'b1), .a({\xmem_data[3][7] , 
        \xmem_data[3][6] , \xmem_data[3][5] , \xmem_data[3][4] , 
        \xmem_data[3][3] , \xmem_data[3][2] , \xmem_data[3][1] , 
        \xmem_data[3][0] }), .b({\fmem_data[3][7] , \fmem_data[3][6] , 
        \fmem_data[3][5] , \fmem_data[3][4] , \fmem_data[3][3] , 
        \fmem_data[3][2] , \fmem_data[3][1] , \fmem_data[3][0] }), .product({
        \x_mult_f_int[3][15] , \x_mult_f_int[3][14] , \x_mult_f_int[3][13] , 
        \x_mult_f_int[3][12] , \x_mult_f_int[3][11] , \x_mult_f_int[3][10] , 
        \x_mult_f_int[3][9] , \x_mult_f_int[3][8] , \x_mult_f_int[3][7] , 
        \x_mult_f_int[3][6] , \x_mult_f_int[3][5] , \x_mult_f_int[3][4] , 
        \x_mult_f_int[3][3] , \x_mult_f_int[3][2] , \x_mult_f_int[3][1] , 
        \x_mult_f_int[3][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_29 \multiplier[2].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8905), .en(n8902), .tc(1'b1), .a({\xmem_data[2][7] , 
        \xmem_data[2][6] , \xmem_data[2][5] , \xmem_data[2][4] , 
        \xmem_data[2][3] , \xmem_data[2][2] , \xmem_data[2][1] , 
        \xmem_data[2][0] }), .b({\fmem_data[2][7] , \fmem_data[2][6] , 
        \fmem_data[2][5] , \fmem_data[2][4] , \fmem_data[2][3] , 
        \fmem_data[2][2] , \fmem_data[2][1] , \fmem_data[2][0] }), .product({
        \x_mult_f_int[2][15] , \x_mult_f_int[2][14] , \x_mult_f_int[2][13] , 
        \x_mult_f_int[2][12] , \x_mult_f_int[2][11] , \x_mult_f_int[2][10] , 
        \x_mult_f_int[2][9] , \x_mult_f_int[2][8] , \x_mult_f_int[2][7] , 
        \x_mult_f_int[2][6] , \x_mult_f_int[2][5] , \x_mult_f_int[2][4] , 
        \x_mult_f_int[2][3] , \x_mult_f_int[2][2] , \x_mult_f_int[2][1] , 
        \x_mult_f_int[2][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_30 \multiplier[1].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n3650), .tc(1'b1), .a({\xmem_data[1][7] , 
        \xmem_data[1][6] , \xmem_data[1][5] , \xmem_data[1][4] , 
        \xmem_data[1][3] , \xmem_data[1][2] , \xmem_data[1][1] , 
        \xmem_data[1][0] }), .b({\fmem_data[1][7] , \fmem_data[1][6] , 
        \fmem_data[1][5] , \fmem_data[1][4] , \fmem_data[1][3] , 
        \fmem_data[1][2] , \fmem_data[1][1] , \fmem_data[1][0] }), .product({
        \x_mult_f_int[1][15] , \x_mult_f_int[1][14] , \x_mult_f_int[1][13] , 
        \x_mult_f_int[1][12] , \x_mult_f_int[1][11] , \x_mult_f_int[1][10] , 
        \x_mult_f_int[1][9] , \x_mult_f_int[1][8] , \x_mult_f_int[1][7] , 
        \x_mult_f_int[1][6] , \x_mult_f_int[1][5] , \x_mult_f_int[1][4] , 
        \x_mult_f_int[1][3] , \x_mult_f_int[1][2] , \x_mult_f_int[1][1] , 
        \x_mult_f_int[1][0] }) );
  conv_128_32_opt_DW_mult_pipe_J1_31 \multiplier[0].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8907), .en(n3650), .tc(1'b1), .a({\xmem_data[0][7] , 
        \xmem_data[0][6] , \xmem_data[0][5] , \xmem_data[0][4] , 
        \xmem_data[0][3] , \xmem_data[0][2] , \xmem_data[0][1] , 
        \xmem_data[0][0] }), .b({\fmem_data[0][7] , \fmem_data[0][6] , 
        \fmem_data[0][5] , \fmem_data[0][4] , \fmem_data[0][3] , 
        \fmem_data[0][2] , \fmem_data[0][1] , \fmem_data[0][0] }), .product({
        \x_mult_f_int[0][15] , \x_mult_f_int[0][14] , \x_mult_f_int[0][13] , 
        \x_mult_f_int[0][12] , \x_mult_f_int[0][11] , \x_mult_f_int[0][10] , 
        \x_mult_f_int[0][9] , \x_mult_f_int[0][8] , \x_mult_f_int[0][7] , 
        \x_mult_f_int[0][6] , \x_mult_f_int[0][5] , \x_mult_f_int[0][4] , 
        \x_mult_f_int[0][3] , \x_mult_f_int[0][2] , \x_mult_f_int[0][1] , 
        \x_mult_f_int[0][0] }) );
  DFF_X1 \adder_stage3_reg[3][3]  ( .D(n9705), .CK(clk), .Q(
        \adder_stage3[3][3] ) );
  DFF_X1 \x_mult_f_reg[3][0]  ( .D(n9333), .CK(clk), .Q(\x_mult_f[3][0] ) );
  DFF_X1 \x_mult_f_reg[28][0]  ( .D(n9383), .CK(clk), .Q(\x_mult_f[28][0] ) );
  DFF_X1 \x_mult_f_reg[3][1]  ( .D(n9332), .CK(clk), .Q(\x_mult_f[3][1] ) );
  DFF_X1 \adder_stage2_reg[7][0]  ( .D(n9786), .CK(clk), .Q(
        \adder_stage2[7][0] ) );
  DFF_X1 \x_mult_f_reg[14][7]  ( .D(n9103), .CK(clk), .Q(\x_mult_f[14][7] ) );
  DFF_X1 \adder_stage1_reg[12][7]  ( .D(n9962), .CK(clk), .Q(
        \adder_stage1[12][7] ) );
  DFF_X1 \x_mult_f_reg[25][5]  ( .D(n9240), .CK(clk), .Q(\x_mult_f[25][5] ) );
  DFF_X1 \adder_stage1_reg[11][9]  ( .D(n9977), .CK(clk), .Q(
        \adder_stage1[11][9] ) );
  DFF_X1 \adder_stage3_reg[3][11]  ( .D(n9697), .CK(clk), .Q(
        \adder_stage3[3][11] ) );
  DFF_X1 \adder_stage2_reg[3][11]  ( .D(n9842), .CK(clk), .Q(
        \adder_stage2[3][11] ) );
  DFF_X1 \adder_stage2_reg[5][3]  ( .D(n9816), .CK(clk), .Q(
        \adder_stage2[5][3] ) );
  DFF_X1 \x_mult_f_reg[23][3]  ( .D(n9222), .CK(clk), .Q(\x_mult_f[23][3] ) );
  DFF_X1 \x_mult_f_reg[17][5]  ( .D(n9136), .CK(clk), .Q(\x_mult_f[17][5] ) );
  DFF_X1 \x_mult_f_reg[11][15]  ( .D(n8867), .CK(clk), .Q(n8793), .QN(
        \x_mult_f[11][15] ) );
  DFFS_X1 \ctrl_inst/state_reg[1]  ( .D(n3387), .CK(clk), .SN(1'b1), .Q(
        \ctrl_inst/state [1]), .QN(n8815) );
  DFF_X1 \adder_stage1_reg[10][3]  ( .D(n8892), .CK(clk), .QN(
        \adder_stage1[10][3] ) );
  DFF_X1 \x_mult_f_reg[31][7]  ( .D(n8898), .CK(clk), .QN(\x_mult_f[31][7] )
         );
  DFF_X1 \x_mult_f_reg[17][15]  ( .D(n8868), .CK(clk), .Q(n8794), .QN(
        \x_mult_f[17][15] ) );
  DFF_X1 \x_mult_f_reg[17][14]  ( .D(n8861), .CK(clk), .QN(\x_mult_f[17][14] )
         );
  DFF_X1 \x_mult_f_reg[17][13]  ( .D(n8859), .CK(clk), .QN(\x_mult_f[17][13] )
         );
  DFF_X1 \x_mult_f_reg[17][12]  ( .D(n8860), .CK(clk), .QN(\x_mult_f[17][12] )
         );
  DFF_X1 \x_mult_f_reg[16][9]  ( .D(n8888), .CK(clk), .QN(\x_mult_f[16][9] )
         );
  DFF_X1 \x_mult_f_reg[16][8]  ( .D(n8889), .CK(clk), .QN(\x_mult_f[16][8] )
         );
  DFF_X1 \x_mult_f_reg[16][7]  ( .D(n8890), .CK(clk), .QN(\x_mult_f[16][7] )
         );
  DFF_X1 \x_mult_f_reg[16][6]  ( .D(n8891), .CK(clk), .QN(\x_mult_f[16][6] )
         );
  DFF_X1 \x_mult_f_reg[5][15]  ( .D(n8866), .CK(clk), .Q(n8790), .QN(
        \x_mult_f[5][15] ) );
  DFF_X1 \adder_stage1_reg[15][14]  ( .D(n8864), .CK(clk), .QN(
        \adder_stage1[15][14] ) );
  DFF_X1 \adder_stage1_reg[15][13]  ( .D(n8900), .CK(clk), .QN(
        \adder_stage1[15][13] ) );
  DFF_X1 \x_mult_f_reg[4][9]  ( .D(n8872), .CK(clk), .QN(\x_mult_f[4][9] ) );
  DFF_X1 \x_mult_f_reg[4][8]  ( .D(n8873), .CK(clk), .QN(\x_mult_f[4][8] ) );
  DFF_X1 \x_mult_f_reg[4][7]  ( .D(n8874), .CK(clk), .QN(\x_mult_f[4][7] ) );
  DFF_X1 \x_mult_f_reg[4][6]  ( .D(n8875), .CK(clk), .QN(\x_mult_f[4][6] ) );
  DFF_X1 \x_mult_f_reg[24][8]  ( .D(n8896), .CK(clk), .QN(\x_mult_f[24][8] )
         );
  DFF_X1 \x_mult_f_reg[24][7]  ( .D(n8897), .CK(clk), .QN(\x_mult_f[24][7] )
         );
  DFF_X1 \x_mult_f_reg[5][14]  ( .D(n8856), .CK(clk), .QN(\x_mult_f[5][14] )
         );
  DFF_X1 \x_mult_f_reg[5][9]  ( .D(n8878), .CK(clk), .QN(\x_mult_f[5][9] ) );
  DFF_X1 \adder_stage1_reg[2][13]  ( .D(n8883), .CK(clk), .QN(
        \adder_stage1[2][13] ) );
  DFF_X1 \x_mult_f_reg[24][15]  ( .D(n8869), .CK(clk), .Q(n8797), .QN(
        \x_mult_f[24][15] ) );
  DFF_X1 \x_mult_f_reg[24][14]  ( .D(n8862), .CK(clk), .QN(\x_mult_f[24][14] )
         );
  DFF_X1 \x_mult_f_reg[24][13]  ( .D(n8855), .CK(clk), .QN(\x_mult_f[24][13] )
         );
  DFF_X1 \x_mult_f_reg[24][11]  ( .D(n8893), .CK(clk), .QN(\x_mult_f[24][11] )
         );
  DFF_X1 \x_mult_f_reg[24][10]  ( .D(n8894), .CK(clk), .QN(\x_mult_f[24][10] )
         );
  DFF_X1 \x_mult_f_reg[24][9]  ( .D(n8895), .CK(clk), .QN(\x_mult_f[24][9] )
         );
  DFF_X1 \adder_stage1_reg[5][15]  ( .D(n8863), .CK(clk), .QN(
        \adder_stage1[5][15] ) );
  DFF_X1 \x_mult_f_reg[31][6]  ( .D(n8899), .CK(clk), .QN(\x_mult_f[31][6] )
         );
  DFF_X1 \adder_stage1_reg[15][15]  ( .D(n8854), .CK(clk), .QN(
        \adder_stage1[15][15] ) );
  DFF_X1 \adder_stage3_reg[1][19]  ( .D(n8884), .CK(clk), .QN(
        \adder_stage3[1][19] ) );
  DFF_X1 \adder_stage3_reg[1][18]  ( .D(n8885), .CK(clk), .QN(
        \adder_stage3[1][18] ) );
  DFF_X1 \x_mult_f_reg[5][12]  ( .D(n8858), .CK(clk), .QN(\x_mult_f[5][12] )
         );
  DFF_X1 \x_mult_f_reg[5][11]  ( .D(n8876), .CK(clk), .QN(\x_mult_f[5][11] )
         );
  DFF_X1 \x_mult_f_reg[5][10]  ( .D(n8877), .CK(clk), .QN(\x_mult_f[5][10] )
         );
  DFF_X1 \x_mult_f_reg[5][7]  ( .D(n8880), .CK(clk), .QN(\x_mult_f[5][7] ) );
  DFF_X1 \adder_stage1_reg[2][20]  ( .D(n8882), .CK(clk), .Q(n8800), .QN(
        \adder_stage1[2][20] ) );
  DFF_X1 \x_mult_f_reg[5][8]  ( .D(n8879), .CK(clk), .QN(\x_mult_f[5][8] ) );
  DFF_X1 \x_mult_f_reg[5][6]  ( .D(n8881), .CK(clk), .QN(\x_mult_f[5][6] ) );
  DFF_X1 \x_mult_f_reg[16][12]  ( .D(n8857), .CK(clk), .QN(\x_mult_f[16][12] )
         );
  DFF_X1 \x_mult_f_reg[16][11]  ( .D(n8886), .CK(clk), .QN(\x_mult_f[16][11] )
         );
  DFF_X1 \x_mult_f_reg[16][10]  ( .D(n8887), .CK(clk), .QN(\x_mult_f[16][10] )
         );
  DFF_X1 \adder_stage2_reg[5][16]  ( .D(n8865), .CK(clk), .QN(
        \adder_stage2[5][16] ) );
  DFF_X1 \ctrl_inst/m_valid_reg  ( .D(n8870), .CK(clk), .Q(n8787), .QN(
        m_valid_y) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[1]  ( .D(n3394), .CK(clk), .Q(
        fmem_addr[1]), .QN(n8808) );
  DFF_X1 \ctrl_fmem_write_inst/s_ready_reg  ( .D(n3392), .CK(clk), .Q(
        s_ready_f), .QN(n8811) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[0]  ( .D(n3121), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [0]), .QN(n8810) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[1]  ( .D(n3120), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [1]), .QN(n8840) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[4]  ( .D(n3397), .CK(clk), .Q(
        fmem_addr[4]), .QN(n8845) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[0]  ( .D(n3395), .CK(clk), .Q(
        fmem_addr[0]), .QN(n8805) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[6]  ( .D(n8871), .CK(clk), .Q(n8842), 
        .QN(\ctrl_inst/xmem_tracker [6]) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[2]  ( .D(n3119), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [2]), .QN(n8814) );
  DFF_X1 \adder_stage3_reg[2][20]  ( .D(n9709), .CK(clk), .Q(
        \adder_stage3[2][20] ) );
  BUF_X1 U3404 ( .A(n5384), .Z(n5175) );
  BUF_X1 U3405 ( .A(n5384), .Z(n6307) );
  BUF_X2 U3406 ( .A(n5181), .Z(n8298) );
  CLKBUF_X1 U3407 ( .A(n3445), .Z(n3409) );
  INV_X1 U3408 ( .A(n8778), .ZN(n8770) );
  BUF_X1 U3409 ( .A(n4097), .Z(n4671) );
  OR2_X2 U3410 ( .A1(n3650), .A2(n3649), .ZN(n3445) );
  INV_X1 U3411 ( .A(n3682), .ZN(n3400) );
  NAND2_X2 U3412 ( .A1(n8778), .A2(n3400), .ZN(n3649) );
  NOR2_X2 U3413 ( .A1(conv_done), .A2(reset), .ZN(n8778) );
  NAND2_X1 U3414 ( .A1(n3402), .A2(n3401), .ZN(n9226) );
  NAND2_X1 U3415 ( .A1(n8088), .A2(\x_mult_f[24][5] ), .ZN(n3401) );
  NAND2_X1 U3416 ( .A1(n4257), .A2(\x_mult_f_int[24][5] ), .ZN(n3402) );
  NAND2_X1 U3417 ( .A1(n3404), .A2(n3403), .ZN(n10051) );
  NAND2_X1 U3418 ( .A1(n8088), .A2(\adder_stage1[7][2] ), .ZN(n3403) );
  NAND2_X1 U3419 ( .A1(n8281), .A2(n5832), .ZN(n3404) );
  NAND2_X1 U3420 ( .A1(n3406), .A2(n3405), .ZN(n9356) );
  NAND2_X1 U3421 ( .A1(n8088), .A2(\x_mult_f[15][1] ), .ZN(n3405) );
  NAND2_X1 U3422 ( .A1(n8153), .A2(\x_mult_f_int[15][1] ), .ZN(n3406) );
  NOR2_X1 U3423 ( .A1(\adder_stage1[12][3] ), .A2(\adder_stage1[13][3] ), .ZN(
        n6987) );
  NOR2_X1 U3424 ( .A1(\adder_stage1[8][3] ), .A2(\adder_stage1[9][3] ), .ZN(
        n4800) );
  NOR2_X1 U3425 ( .A1(\x_mult_f[0][3] ), .A2(\x_mult_f[1][3] ), .ZN(n5657) );
  OR2_X1 U3426 ( .A1(m_ready_y), .A2(\ctrl_inst/s_ready_fsm ), .ZN(n3494) );
  INV_X2 U3427 ( .A(n5247), .ZN(n7614) );
  INV_X1 U3428 ( .A(n8045), .ZN(n8306) );
  INV_X1 U3429 ( .A(n8045), .ZN(n8338) );
  INV_X2 U3430 ( .A(n8045), .ZN(n7855) );
  BUF_X2 U3431 ( .A(n7163), .Z(n8189) );
  NOR2_X1 U3432 ( .A1(n3685), .A2(n3684), .ZN(n3983) );
  INV_X4 U3433 ( .A(n5247), .ZN(n7920) );
  BUF_X1 U3434 ( .A(n6093), .Z(n4314) );
  INV_X4 U3435 ( .A(n7989), .ZN(n8273) );
  BUF_X2 U3436 ( .A(n5449), .Z(n7862) );
  BUF_X2 U3437 ( .A(n5181), .Z(n6279) );
  CLKBUF_X2 U3438 ( .A(n4671), .Z(n4444) );
  CLKBUF_X2 U3439 ( .A(n4671), .Z(n6352) );
  BUF_X1 U3440 ( .A(n4771), .Z(n4990) );
  BUF_X1 U3441 ( .A(n5406), .Z(n7979) );
  BUF_X1 U3442 ( .A(n3445), .Z(n6720) );
  CLKBUF_X2 U3443 ( .A(n4671), .Z(n4645) );
  BUF_X1 U3444 ( .A(n5124), .Z(n5449) );
  BUF_X2 U3445 ( .A(n5332), .Z(n3407) );
  BUF_X2 U3446 ( .A(n5406), .Z(n3408) );
  BUF_X1 U3447 ( .A(n4097), .Z(n5124) );
  BUF_X2 U3448 ( .A(n3445), .Z(n4771) );
  INV_X1 U3449 ( .A(n3666), .ZN(n8388) );
  NOR2_X1 U3450 ( .A1(n8504), .A2(n8754), .ZN(n8512) );
  NOR2_X1 U3451 ( .A1(n8504), .A2(n8688), .ZN(n8451) );
  NOR2_X1 U3452 ( .A1(n8504), .A2(n8699), .ZN(n8461) );
  NOR2_X1 U3453 ( .A1(n8504), .A2(n8710), .ZN(n8471) );
  NOR2_X1 U3454 ( .A1(n8504), .A2(n8742), .ZN(n8501) );
  NOR2_X1 U3455 ( .A1(n8504), .A2(n8775), .ZN(n8481) );
  NOR2_X1 U3456 ( .A1(n8504), .A2(n8731), .ZN(n8491) );
  NOR2_X1 U3457 ( .A1(n8731), .A2(n8586), .ZN(n8573) );
  NOR2_X1 U3458 ( .A1(n8775), .A2(n8586), .ZN(n8563) );
  NOR2_X1 U3459 ( .A1(n8710), .A2(n8586), .ZN(n8553) );
  NOR2_X1 U3460 ( .A1(n8699), .A2(n8586), .ZN(n8543) );
  NOR2_X1 U3461 ( .A1(n8688), .A2(n8586), .ZN(n8533) );
  NOR2_X1 U3462 ( .A1(n8766), .A2(n8586), .ZN(n8523) );
  NOR2_X1 U3463 ( .A1(n8754), .A2(n8586), .ZN(n8594) );
  NOR2_X1 U3464 ( .A1(n8742), .A2(n8586), .ZN(n8583) );
  OR2_X1 U3465 ( .A1(n8809), .A2(n8515), .ZN(n8504) );
  OR2_X1 U3466 ( .A1(n3681), .A2(n3486), .ZN(n3496) );
  OR2_X1 U3467 ( .A1(fmem_addr[3]), .A2(n8515), .ZN(n8586) );
  NOR2_X1 U3468 ( .A1(\x_mult_f[30][5] ), .A2(\x_mult_f[31][5] ), .ZN(n7444)
         );
  NOR2_X1 U3469 ( .A1(\x_mult_f[12][3] ), .A2(\x_mult_f[13][3] ), .ZN(n5881)
         );
  CLKBUF_X1 U3470 ( .A(n6631), .Z(n3410) );
  CLKBUF_X1 U3471 ( .A(n7957), .Z(n3411) );
  CLKBUF_X1 U3472 ( .A(n7320), .Z(n3412) );
  AOI21_X1 U3473 ( .B1(n5735), .B2(n5734), .A(n5733), .ZN(n3413) );
  INV_X1 U3474 ( .A(n5735), .ZN(n3414) );
  AOI21_X1 U3475 ( .B1(n5557), .B2(n5555), .A(n5534), .ZN(n5727) );
  AND2_X1 U3476 ( .A1(n3415), .A2(n3416), .ZN(n5853) );
  AND2_X1 U3477 ( .A1(n3417), .A2(n3418), .ZN(n3638) );
  AOI21_X1 U3478 ( .B1(n6704), .B2(n6844), .A(n6703), .ZN(n6783) );
  AOI21_X1 U3479 ( .B1(n5285), .B2(n5792), .A(n5284), .ZN(n5782) );
  CLKBUF_X1 U3480 ( .A(n7938), .Z(n3419) );
  OAI21_X1 U3481 ( .B1(n3799), .B2(n3798), .A(n3797), .ZN(n7938) );
  AOI21_X1 U3482 ( .B1(n3527), .B2(n3578), .A(n3526), .ZN(n3420) );
  NOR2_X2 U3483 ( .A1(\x_mult_f[30][3] ), .A2(\x_mult_f[31][3] ), .ZN(n4430)
         );
  CLKBUF_X1 U3484 ( .A(n7032), .Z(n3421) );
  NOR2_X2 U3485 ( .A1(\adder_stage4[0][9] ), .A2(\adder_stage4[1][9] ), .ZN(
        n3616) );
  CLKBUF_X1 U3486 ( .A(n6063), .Z(n3422) );
  NAND2_X1 U3487 ( .A1(\ctrl_inst/xmem_tracker [4]), .A2(
        \ctrl_inst/xmem_tracker [2]), .ZN(n3651) );
  INV_X1 U3488 ( .A(n4344), .ZN(n3508) );
  OAI21_X1 U3489 ( .B1(n5084), .B2(n3507), .A(n5086), .ZN(n4343) );
  INV_X1 U3490 ( .A(n5087), .ZN(n3507) );
  AOI21_X1 U3491 ( .B1(n3506), .B2(n5096), .A(n3505), .ZN(n5084) );
  INV_X1 U3492 ( .A(n5100), .ZN(n3505) );
  NAND2_X1 U3493 ( .A1(\adder_stage1[2][15] ), .A2(\adder_stage1[3][15] ), 
        .ZN(n8006) );
  NOR2_X1 U3494 ( .A1(\adder_stage1[3][15] ), .A2(\adder_stage1[2][15] ), .ZN(
        n8007) );
  INV_X1 U3495 ( .A(n3680), .ZN(n3495) );
  AOI21_X1 U3496 ( .B1(n6956), .B2(n6986), .A(n6955), .ZN(n6976) );
  INV_X1 U3497 ( .A(n8133), .ZN(n7997) );
  NOR2_X1 U3498 ( .A1(n3446), .A2(n3459), .ZN(n7998) );
  NAND2_X1 U3499 ( .A1(n3459), .A2(n3446), .ZN(n7996) );
  AOI21_X1 U3500 ( .B1(n4779), .B2(n4799), .A(n4778), .ZN(n4794) );
  CLKBUF_X1 U3501 ( .A(n4324), .Z(n4334) );
  AOI21_X1 U3502 ( .B1(n4154), .B2(n5602), .A(n4153), .ZN(n4184) );
  NOR2_X1 U3503 ( .A1(n5099), .A2(n3504), .ZN(n5083) );
  INV_X1 U3504 ( .A(n5097), .ZN(n3504) );
  CLKBUF_X1 U3505 ( .A(n6778), .Z(n6721) );
  CLKBUF_X1 U3506 ( .A(n4476), .Z(n4455) );
  AOI21_X1 U3507 ( .B1(n4446), .B2(n5656), .A(n4445), .ZN(n4493) );
  CLKBUF_X1 U3508 ( .A(n4771), .Z(n7989) );
  CLKBUF_X1 U3509 ( .A(n6093), .Z(n7343) );
  NAND2_X1 U3510 ( .A1(fmem_addr[3]), .A2(n8677), .ZN(n8666) );
  NAND2_X1 U3511 ( .A1(n8677), .A2(n8809), .ZN(n8753) );
  NOR2_X1 U3512 ( .A1(n3651), .A2(n3483), .ZN(n3652) );
  AND2_X1 U3513 ( .A1(\ctrl_inst/xmem_tracker [1]), .A2(
        \ctrl_inst/xmem_tracker [0]), .ZN(n3658) );
  NAND2_X1 U3514 ( .A1(n3490), .A2(n3489), .ZN(n3648) );
  AND2_X1 U3515 ( .A1(\ctrl_inst/xmem_tracker [5]), .A2(
        \ctrl_inst/xmem_tracker [6]), .ZN(n3490) );
  NOR2_X1 U3516 ( .A1(n3488), .A2(n3651), .ZN(n3489) );
  NAND2_X1 U3517 ( .A1(xmem_full), .A2(n8811), .ZN(n3682) );
  AOI21_X1 U3518 ( .B1(n3534), .B2(n3533), .A(n3532), .ZN(n3539) );
  INV_X2 U3519 ( .A(n3649), .ZN(n8907) );
  NAND2_X1 U3520 ( .A1(s_ready_f), .A2(s_valid_f), .ZN(n8772) );
  INV_X1 U3521 ( .A(n8772), .ZN(n8771) );
  NAND2_X1 U3522 ( .A1(m_ready_y), .A2(m_valid_y), .ZN(n3681) );
  NAND2_X1 U3523 ( .A1(\adder_stage1[15][15] ), .A2(\adder_stage1[14][15] ), 
        .ZN(n7812) );
  NOR2_X1 U3524 ( .A1(\adder_stage1[15][15] ), .A2(\adder_stage1[14][15] ), 
        .ZN(n7813) );
  CLKBUF_X1 U3525 ( .A(n7814), .Z(n3430) );
  CLKBUF_X1 U3526 ( .A(n8218), .Z(n8222) );
  CLKBUF_X1 U3527 ( .A(n6589), .Z(n3429) );
  CLKBUF_X1 U3528 ( .A(n7159), .Z(n3436) );
  CLKBUF_X1 U3529 ( .A(n6156), .Z(n3437) );
  CLKBUF_X1 U3530 ( .A(n7925), .Z(n3425) );
  CLKBUF_X1 U3531 ( .A(n7452), .Z(n3435) );
  CLKBUF_X1 U3532 ( .A(n6918), .Z(n3433) );
  CLKBUF_X1 U3533 ( .A(n5352), .Z(n8018) );
  AOI21_X1 U3534 ( .B1(n4343), .B2(n3482), .A(n3508), .ZN(n3509) );
  AOI21_X1 U3535 ( .B1(n5098), .B2(n3456), .A(n4343), .ZN(n4346) );
  NAND2_X1 U3536 ( .A1(n5085), .A2(n5084), .ZN(n5089) );
  NAND2_X1 U3537 ( .A1(n5098), .A2(n5083), .ZN(n5085) );
  AOI21_X1 U3538 ( .B1(n5098), .B2(n5097), .A(n5096), .ZN(n5102) );
  CLKBUF_X1 U3539 ( .A(n6744), .Z(n3441) );
  NAND2_X1 U3540 ( .A1(\x_mult_f[5][2] ), .A2(\x_mult_f[4][2] ), .ZN(n6866) );
  INV_X2 U3541 ( .A(n8045), .ZN(n8336) );
  INV_X1 U3542 ( .A(n3444), .ZN(n8779) );
  INV_X1 U3543 ( .A(n8451), .ZN(n8452) );
  INV_X1 U3544 ( .A(n8461), .ZN(n8462) );
  INV_X1 U3545 ( .A(n8471), .ZN(n8472) );
  INV_X1 U3546 ( .A(n8481), .ZN(n8482) );
  INV_X1 U3547 ( .A(n8491), .ZN(n8492) );
  INV_X1 U3548 ( .A(n8501), .ZN(n8502) );
  INV_X1 U3549 ( .A(n8512), .ZN(n8513) );
  INV_X1 U3550 ( .A(n8523), .ZN(n8524) );
  INV_X1 U3551 ( .A(n8533), .ZN(n8534) );
  INV_X1 U3552 ( .A(n8543), .ZN(n8544) );
  INV_X1 U3553 ( .A(n8553), .ZN(n8554) );
  INV_X1 U3554 ( .A(n8563), .ZN(n8564) );
  INV_X1 U3555 ( .A(n8573), .ZN(n8574) );
  INV_X1 U3556 ( .A(n8583), .ZN(n8584) );
  INV_X1 U3557 ( .A(n8594), .ZN(n8595) );
  NOR2_X1 U3558 ( .A1(n8766), .A2(n8666), .ZN(n8604) );
  NOR2_X1 U3559 ( .A1(n8666), .A2(n8688), .ZN(n8613) );
  INV_X1 U3560 ( .A(n8613), .ZN(n8614) );
  NOR2_X1 U3561 ( .A1(n8666), .A2(n8699), .ZN(n8623) );
  INV_X1 U3562 ( .A(n8623), .ZN(n8624) );
  NOR2_X1 U3563 ( .A1(n8666), .A2(n8710), .ZN(n8633) );
  INV_X1 U3564 ( .A(n8633), .ZN(n8634) );
  NOR2_X1 U3565 ( .A1(n8666), .A2(n8775), .ZN(n8643) );
  INV_X1 U3566 ( .A(n8643), .ZN(n8644) );
  NOR2_X1 U3567 ( .A1(n8666), .A2(n8731), .ZN(n8653) );
  INV_X1 U3568 ( .A(n8653), .ZN(n8654) );
  NOR2_X1 U3569 ( .A1(n8666), .A2(n8742), .ZN(n8663) );
  INV_X1 U3570 ( .A(n8663), .ZN(n8664) );
  NOR2_X1 U3571 ( .A1(n8666), .A2(n8754), .ZN(n8674) );
  INV_X1 U3572 ( .A(n8674), .ZN(n8675) );
  NOR2_X1 U3573 ( .A1(n8766), .A2(n8753), .ZN(n8685) );
  INV_X1 U3574 ( .A(n8685), .ZN(n8686) );
  NOR2_X1 U3575 ( .A1(n8688), .A2(n8753), .ZN(n8696) );
  INV_X1 U3576 ( .A(n8696), .ZN(n8697) );
  NOR2_X1 U3577 ( .A1(n8699), .A2(n8753), .ZN(n8707) );
  INV_X1 U3578 ( .A(n8707), .ZN(n8708) );
  NOR2_X1 U3579 ( .A1(n8710), .A2(n8753), .ZN(n8718) );
  INV_X1 U3580 ( .A(n8718), .ZN(n8719) );
  NOR2_X1 U3581 ( .A1(n8775), .A2(n8753), .ZN(n8728) );
  INV_X1 U3582 ( .A(n8728), .ZN(n8729) );
  NOR2_X1 U3583 ( .A1(n8731), .A2(n8753), .ZN(n8739) );
  INV_X1 U3584 ( .A(n8739), .ZN(n8740) );
  NOR2_X1 U3585 ( .A1(n8742), .A2(n8753), .ZN(n8750) );
  INV_X1 U3586 ( .A(n8750), .ZN(n8751) );
  NOR2_X1 U3587 ( .A1(n8754), .A2(n8753), .ZN(n8762) );
  INV_X1 U3588 ( .A(n8762), .ZN(n8763) );
  INV_X1 U3589 ( .A(n8604), .ZN(n8768) );
  INV_X1 U3590 ( .A(n3648), .ZN(n3979) );
  CLKBUF_X1 U3591 ( .A(n8353), .Z(n8367) );
  XNOR2_X1 U3592 ( .A(n8133), .B(n8132), .ZN(n8134) );
  XNOR2_X1 U3593 ( .A(n3459), .B(n3446), .ZN(n8132) );
  CLKBUF_X1 U3594 ( .A(n8403), .Z(n8408) );
  NOR2_X1 U3595 ( .A1(n8045), .A2(n3460), .ZN(n8046) );
  INV_X8 U3596 ( .A(n3649), .ZN(n8905) );
  NOR2_X2 U3597 ( .A1(\adder_stage4[0][11] ), .A2(\adder_stage4[1][11] ), .ZN(
        n3583) );
  NOR2_X1 U3598 ( .A1(\x_mult_f[4][3] ), .A2(\x_mult_f[5][3] ), .ZN(n6869) );
  AOI21_X2 U3599 ( .B1(n5374), .B2(n5373), .A(n5372), .ZN(n8202) );
  AOI21_X2 U3600 ( .B1(n5916), .B2(n5426), .A(n5425), .ZN(n8193) );
  AOI21_X2 U3601 ( .B1(n6994), .B2(n6964), .A(n6963), .ZN(n7663) );
  OR2_X1 U3602 ( .A1(n3423), .A2(n3424), .ZN(n7238) );
  AOI21_X1 U3603 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n7349) );
  AOI21_X1 U3604 ( .B1(n7925), .B2(n7923), .A(n6278), .ZN(n3426) );
  AOI21_X1 U3605 ( .B1(n5352), .B2(n5227), .A(n5226), .ZN(n3427) );
  AOI21_X1 U3606 ( .B1(n6504), .B2(n6537), .A(n6503), .ZN(n3428) );
  AOI21_X1 U3607 ( .B1(n6063), .B2(n6062), .A(n6061), .ZN(n3431) );
  AOI21_X1 U3608 ( .B1(n5140), .B2(n6918), .A(n5139), .ZN(n3432) );
  NOR2_X2 U3609 ( .A1(\x_mult_f[28][3] ), .A2(\x_mult_f[29][3] ), .ZN(n5611)
         );
  AOI21_X1 U3610 ( .B1(n7452), .B2(n5644), .A(n5643), .ZN(n3434) );
  NAND2_X1 U3611 ( .A1(n8349), .A2(n3496), .ZN(n3438) );
  NAND2_X1 U3612 ( .A1(n8349), .A2(n3496), .ZN(n3439) );
  NAND2_X1 U3613 ( .A1(n8349), .A2(n3496), .ZN(n3650) );
  AOI21_X1 U3614 ( .B1(n5467), .B2(n6744), .A(n5466), .ZN(n3440) );
  AND2_X1 U3615 ( .A1(n3650), .A2(n8907), .ZN(n4097) );
  INV_X2 U3616 ( .A(n8372), .ZN(n8911) );
  NAND2_X1 U3617 ( .A1(n8010), .A2(n6279), .ZN(n3442) );
  AOI21_X1 U3618 ( .B1(n3421), .B2(n7030), .A(n6286), .ZN(n3443) );
  AOI21_X2 U3619 ( .B1(n5934), .B2(n5932), .A(n5290), .ZN(n7912) );
  XNOR2_X1 U3620 ( .A(n3430), .B(n7567), .ZN(n7568) );
  OAI21_X1 U3621 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n8001) );
  AOI21_X1 U3622 ( .B1(n8218), .B2(n8220), .A(n7566), .ZN(n7814) );
  NOR2_X1 U3623 ( .A1(\adder_stage1[14][3] ), .A2(\adder_stage1[15][3] ), .ZN(
        n6615) );
  OR2_X1 U3624 ( .A1(n8766), .A2(n8504), .ZN(n3444) );
  XNOR2_X1 U3625 ( .A(n3443), .B(n6287), .ZN(n6288) );
  OAI21_X1 U3626 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n8129) );
  AOI21_X1 U3627 ( .B1(n7032), .B2(n7030), .A(n6286), .ZN(n8008) );
  INV_X1 U3628 ( .A(n3439), .ZN(n8372) );
  BUF_X1 U3629 ( .A(n6093), .Z(n7163) );
  BUF_X1 U3630 ( .A(n5332), .Z(n8004) );
  BUF_X2 U3631 ( .A(n7979), .Z(n8000) );
  BUF_X2 U3632 ( .A(n8045), .Z(n7978) );
  INV_X1 U3633 ( .A(n3407), .ZN(n8323) );
  INV_X1 U3634 ( .A(n3407), .ZN(n8097) );
  INV_X1 U3635 ( .A(n3407), .ZN(n7556) );
  INV_X1 U3636 ( .A(n7979), .ZN(n7952) );
  INV_X1 U3637 ( .A(n4771), .ZN(n8088) );
  BUF_X1 U3638 ( .A(n5124), .Z(n5181) );
  BUF_X1 U3639 ( .A(n4671), .Z(n5767) );
  AND2_X1 U3640 ( .A1(n5083), .A2(n5087), .ZN(n3456) );
  BUF_X2 U3641 ( .A(n5384), .Z(n6636) );
  INV_X1 U3642 ( .A(n8045), .ZN(n8427) );
  INV_X1 U3643 ( .A(n8045), .ZN(n8409) );
  INV_X1 U3644 ( .A(n8045), .ZN(n7864) );
  INV_X4 U3645 ( .A(n8388), .ZN(n8391) );
  INV_X1 U3646 ( .A(n5099), .ZN(n3506) );
  INV_X1 U3647 ( .A(n3445), .ZN(n8340) );
  BUF_X1 U3648 ( .A(n3445), .Z(n5406) );
  BUF_X1 U3649 ( .A(n5124), .Z(n6093) );
  BUF_X1 U3650 ( .A(n5124), .Z(n6238) );
  OR2_X1 U3651 ( .A1(\x_mult_f[12][13] ), .A2(\x_mult_f[13][13] ), .ZN(n3482)
         );
  AND2_X1 U3652 ( .A1(n3495), .A2(n8806), .ZN(n3486) );
  AND2_X1 U3653 ( .A1(n3456), .A2(n3482), .ZN(n3487) );
  NAND3_X1 U3655 ( .A1(\ctrl_inst/xmem_tracker [1]), .A2(
        \ctrl_inst/xmem_tracker [0]), .A3(\ctrl_inst/xmem_tracker [3]), .ZN(
        n3488) );
  NAND2_X1 U3656 ( .A1(n8812), .A2(n8787), .ZN(n3491) );
  NAND2_X1 U3657 ( .A1(n3491), .A2(n8806), .ZN(n3492) );
  NAND2_X1 U3658 ( .A1(\ctrl_inst/state [0]), .A2(n8815), .ZN(n3680) );
  NOR2_X1 U3659 ( .A1(n3492), .A2(n3680), .ZN(n3493) );
  NAND4_X2 U3660 ( .A1(n3494), .A2(n3648), .A3(s_valid_x), .A4(n3493), .ZN(
        n8349) );
  BUF_X4 U3661 ( .A(n3439), .Z(n8901) );
  INV_X2 U3662 ( .A(n8372), .ZN(n8908) );
  INV_X1 U3663 ( .A(n8372), .ZN(n8910) );
  INV_X1 U3664 ( .A(n8372), .ZN(n8909) );
  NOR2_X1 U3665 ( .A1(\x_mult_f[12][1] ), .A2(\x_mult_f[13][1] ), .ZN(n5937)
         );
  NAND2_X1 U3666 ( .A1(\x_mult_f[12][0] ), .A2(\x_mult_f[13][0] ), .ZN(n5978)
         );
  NAND2_X1 U3667 ( .A1(\x_mult_f[12][1] ), .A2(\x_mult_f[13][1] ), .ZN(n5938)
         );
  OAI21_X1 U3668 ( .B1(n5937), .B2(n5978), .A(n5938), .ZN(n5880) );
  NOR2_X1 U3669 ( .A1(\x_mult_f[12][2] ), .A2(\x_mult_f[13][2] ), .ZN(n5892)
         );
  NOR2_X1 U3670 ( .A1(n5892), .A2(n5881), .ZN(n3498) );
  NAND2_X1 U3671 ( .A1(\x_mult_f[12][2] ), .A2(\x_mult_f[13][2] ), .ZN(n5893)
         );
  NAND2_X1 U3672 ( .A1(\x_mult_f[12][3] ), .A2(\x_mult_f[13][3] ), .ZN(n5882)
         );
  OAI21_X1 U3673 ( .B1(n5881), .B2(n5893), .A(n5882), .ZN(n3497) );
  AOI21_X1 U3674 ( .B1(n5880), .B2(n3498), .A(n3497), .ZN(n5757) );
  NOR2_X1 U3675 ( .A1(\x_mult_f[12][4] ), .A2(\x_mult_f[13][4] ), .ZN(n5888)
         );
  NOR2_X1 U3676 ( .A1(\x_mult_f[12][5] ), .A2(\x_mult_f[13][5] ), .ZN(n5947)
         );
  NOR2_X1 U3677 ( .A1(n5888), .A2(n5947), .ZN(n5759) );
  NOR2_X1 U3678 ( .A1(\x_mult_f[12][6] ), .A2(\x_mult_f[13][6] ), .ZN(n5924)
         );
  NOR2_X1 U3679 ( .A1(\x_mult_f[12][7] ), .A2(\x_mult_f[13][7] ), .ZN(n5760)
         );
  NOR2_X1 U3680 ( .A1(n5924), .A2(n5760), .ZN(n3500) );
  NAND2_X1 U3681 ( .A1(n5759), .A2(n3500), .ZN(n3502) );
  NAND2_X1 U3682 ( .A1(\x_mult_f[12][4] ), .A2(\x_mult_f[13][4] ), .ZN(n5943)
         );
  NAND2_X1 U3683 ( .A1(\x_mult_f[12][5] ), .A2(\x_mult_f[13][5] ), .ZN(n5948)
         );
  OAI21_X1 U3684 ( .B1(n5947), .B2(n5943), .A(n5948), .ZN(n5758) );
  NAND2_X1 U3685 ( .A1(\x_mult_f[12][6] ), .A2(\x_mult_f[13][6] ), .ZN(n5925)
         );
  NAND2_X1 U3686 ( .A1(\x_mult_f[12][7] ), .A2(\x_mult_f[13][7] ), .ZN(n5761)
         );
  OAI21_X1 U3687 ( .B1(n5760), .B2(n5925), .A(n5761), .ZN(n3499) );
  AOI21_X1 U3688 ( .B1(n3500), .B2(n5758), .A(n3499), .ZN(n3501) );
  OAI21_X1 U3689 ( .B1(n5757), .B2(n3502), .A(n3501), .ZN(n5837) );
  OR2_X1 U3690 ( .A1(\x_mult_f[12][8] ), .A2(\x_mult_f[13][8] ), .ZN(n5835) );
  NAND2_X1 U3691 ( .A1(\x_mult_f[12][8] ), .A2(\x_mult_f[13][8] ), .ZN(n5834)
         );
  INV_X1 U3692 ( .A(n5834), .ZN(n3503) );
  AOI21_X1 U3693 ( .B1(n5837), .B2(n5835), .A(n3503), .ZN(n5877) );
  NOR2_X1 U3694 ( .A1(\x_mult_f[12][9] ), .A2(\x_mult_f[13][9] ), .ZN(n5873)
         );
  NAND2_X1 U3695 ( .A1(\x_mult_f[12][9] ), .A2(\x_mult_f[13][9] ), .ZN(n5874)
         );
  OAI21_X1 U3696 ( .B1(n5877), .B2(n5873), .A(n5874), .ZN(n5098) );
  NOR2_X1 U3697 ( .A1(\x_mult_f[12][11] ), .A2(\x_mult_f[13][11] ), .ZN(n5099)
         );
  OR2_X1 U3698 ( .A1(\x_mult_f[12][10] ), .A2(\x_mult_f[13][10] ), .ZN(n5097)
         );
  OR2_X1 U3699 ( .A1(\x_mult_f[12][12] ), .A2(\x_mult_f[13][12] ), .ZN(n5087)
         );
  NAND2_X1 U3700 ( .A1(n5098), .A2(n3487), .ZN(n3510) );
  NAND2_X1 U3701 ( .A1(\x_mult_f[12][10] ), .A2(\x_mult_f[13][10] ), .ZN(n5092) );
  INV_X1 U3702 ( .A(n5092), .ZN(n5096) );
  NAND2_X1 U3703 ( .A1(\x_mult_f[12][11] ), .A2(\x_mult_f[13][11] ), .ZN(n5100) );
  NAND2_X1 U3704 ( .A1(\x_mult_f[12][12] ), .A2(\x_mult_f[13][12] ), .ZN(n5086) );
  NAND2_X1 U3705 ( .A1(\x_mult_f[12][13] ), .A2(\x_mult_f[13][13] ), .ZN(n4344) );
  NAND2_X1 U3706 ( .A1(n3510), .A2(n3509), .ZN(n7905) );
  BUF_X4 U3707 ( .A(n3438), .Z(n8903) );
  BUF_X2 U3708 ( .A(n4894), .Z(n8334) );
  NAND2_X1 U3709 ( .A1(n3511), .A2(n8334), .ZN(n3513) );
  NAND2_X1 U3710 ( .A1(n7525), .A2(\adder_stage1[6][15] ), .ZN(n3512) );
  NAND2_X1 U3711 ( .A1(n3513), .A2(n3512), .ZN(n10055) );
  NOR2_X1 U3712 ( .A1(\adder_stage4[0][1] ), .A2(\adder_stage4[1][1] ), .ZN(
        n3517) );
  INV_X1 U3713 ( .A(n3517), .ZN(n3514) );
  NAND2_X1 U3714 ( .A1(\adder_stage4[0][1] ), .A2(\adder_stage4[1][1] ), .ZN(
        n3516) );
  NAND2_X1 U3715 ( .A1(n3514), .A2(n3516), .ZN(n3515) );
  NAND2_X1 U3716 ( .A1(\adder_stage4[0][0] ), .A2(\adder_stage4[1][0] ), .ZN(
        n3566) );
  XOR2_X1 U3717 ( .A(n3515), .B(n3566), .Z(m_data_out_y[1]) );
  NOR2_X1 U3718 ( .A1(\adder_stage4[0][2] ), .A2(\adder_stage4[1][2] ), .ZN(
        n3643) );
  NOR2_X1 U3719 ( .A1(n3643), .A2(n3638), .ZN(n3519) );
  OAI21_X1 U3720 ( .B1(n3517), .B2(n3566), .A(n3516), .ZN(n3637) );
  NAND2_X1 U3721 ( .A1(\adder_stage4[0][2] ), .A2(\adder_stage4[1][2] ), .ZN(
        n3644) );
  NAND2_X1 U3722 ( .A1(\adder_stage4[0][3] ), .A2(\adder_stage4[1][3] ), .ZN(
        n3639) );
  OAI21_X1 U3723 ( .B1(n3638), .B2(n3644), .A(n3639), .ZN(n3518) );
  AOI21_X1 U3724 ( .B1(n3519), .B2(n3637), .A(n3518), .ZN(n3601) );
  NOR2_X1 U3725 ( .A1(\adder_stage4[0][4] ), .A2(\adder_stage4[1][4] ), .ZN(
        n3626) );
  NOR2_X1 U3726 ( .A1(\adder_stage4[0][5] ), .A2(\adder_stage4[1][5] ), .ZN(
        n3628) );
  NOR2_X1 U3727 ( .A1(n3626), .A2(n3628), .ZN(n3603) );
  NOR2_X1 U3728 ( .A1(\adder_stage4[0][6] ), .A2(\adder_stage4[1][6] ), .ZN(
        n3621) );
  NOR2_X1 U3729 ( .A1(\adder_stage4[0][7] ), .A2(\adder_stage4[1][7] ), .ZN(
        n3604) );
  NOR2_X1 U3730 ( .A1(n3621), .A2(n3604), .ZN(n3521) );
  NAND2_X1 U3731 ( .A1(n3603), .A2(n3521), .ZN(n3523) );
  NAND2_X1 U3732 ( .A1(\adder_stage4[0][4] ), .A2(\adder_stage4[1][4] ), .ZN(
        n3633) );
  NAND2_X1 U3733 ( .A1(\adder_stage4[0][5] ), .A2(\adder_stage4[1][5] ), .ZN(
        n3629) );
  OAI21_X1 U3734 ( .B1(n3628), .B2(n3633), .A(n3629), .ZN(n3602) );
  NAND2_X1 U3735 ( .A1(\adder_stage4[0][6] ), .A2(\adder_stage4[1][6] ), .ZN(
        n3622) );
  NAND2_X1 U3736 ( .A1(\adder_stage4[0][7] ), .A2(\adder_stage4[1][7] ), .ZN(
        n3605) );
  OAI21_X1 U3737 ( .B1(n3604), .B2(n3622), .A(n3605), .ZN(n3520) );
  AOI21_X1 U3738 ( .B1(n3521), .B2(n3602), .A(n3520), .ZN(n3522) );
  OAI21_X1 U3739 ( .B1(n3601), .B2(n3523), .A(n3522), .ZN(n3534) );
  INV_X1 U3740 ( .A(n3534), .ZN(n3615) );
  NOR2_X1 U3741 ( .A1(\adder_stage4[0][8] ), .A2(\adder_stage4[1][8] ), .ZN(
        n3614) );
  INV_X1 U3742 ( .A(n3614), .ZN(n3524) );
  NAND2_X1 U3743 ( .A1(\adder_stage4[0][8] ), .A2(\adder_stage4[1][8] ), .ZN(
        n3613) );
  NAND2_X1 U3744 ( .A1(n3524), .A2(n3613), .ZN(n3525) );
  XOR2_X1 U3745 ( .A(n3615), .B(n3525), .Z(m_data_out_y[8]) );
  NOR2_X1 U3746 ( .A1(n3614), .A2(n3616), .ZN(n3577) );
  NOR2_X1 U3747 ( .A1(\adder_stage4[0][10] ), .A2(\adder_stage4[1][10] ), .ZN(
        n3581) );
  NOR2_X1 U3748 ( .A1(n3581), .A2(n3583), .ZN(n3527) );
  NAND2_X1 U3749 ( .A1(n3577), .A2(n3527), .ZN(n3556) );
  NOR2_X1 U3750 ( .A1(\adder_stage4[0][12] ), .A2(\adder_stage4[1][12] ), .ZN(
        n3557) );
  NOR2_X1 U3751 ( .A1(\adder_stage4[0][13] ), .A2(\adder_stage4[1][13] ), .ZN(
        n3592) );
  NOR2_X1 U3752 ( .A1(n3557), .A2(n3592), .ZN(n3559) );
  NOR2_X1 U3753 ( .A1(\adder_stage4[0][14] ), .A2(\adder_stage4[1][14] ), .ZN(
        n3564) );
  NOR2_X1 U3754 ( .A1(\adder_stage4[0][15] ), .A2(\adder_stage4[1][15] ), .ZN(
        n3572) );
  NOR2_X1 U3755 ( .A1(n3564), .A2(n3572), .ZN(n3529) );
  NAND2_X1 U3756 ( .A1(n3559), .A2(n3529), .ZN(n3531) );
  NOR2_X1 U3757 ( .A1(n3556), .A2(n3531), .ZN(n3533) );
  NAND2_X1 U3758 ( .A1(\adder_stage4[0][9] ), .A2(\adder_stage4[1][9] ), .ZN(
        n3617) );
  OAI21_X1 U3759 ( .B1(n3616), .B2(n3613), .A(n3617), .ZN(n3578) );
  NAND2_X1 U3760 ( .A1(\adder_stage4[0][10] ), .A2(\adder_stage4[1][10] ), 
        .ZN(n3597) );
  NAND2_X1 U3761 ( .A1(\adder_stage4[0][11] ), .A2(\adder_stage4[1][11] ), 
        .ZN(n3584) );
  OAI21_X1 U3762 ( .B1(n3583), .B2(n3597), .A(n3584), .ZN(n3526) );
  AOI21_X1 U3763 ( .B1(n3527), .B2(n3578), .A(n3526), .ZN(n3555) );
  NAND2_X1 U3764 ( .A1(\adder_stage4[0][12] ), .A2(\adder_stage4[1][12] ), 
        .ZN(n3588) );
  NAND2_X1 U3765 ( .A1(\adder_stage4[0][13] ), .A2(\adder_stage4[1][13] ), 
        .ZN(n3593) );
  OAI21_X1 U3766 ( .B1(n3592), .B2(n3588), .A(n3593), .ZN(n3560) );
  NAND2_X1 U3767 ( .A1(\adder_stage4[0][14] ), .A2(\adder_stage4[1][14] ), 
        .ZN(n3568) );
  NAND2_X1 U3768 ( .A1(\adder_stage4[0][15] ), .A2(\adder_stage4[1][15] ), 
        .ZN(n3573) );
  OAI21_X1 U3769 ( .B1(n3572), .B2(n3568), .A(n3573), .ZN(n3528) );
  AOI21_X1 U3770 ( .B1(n3529), .B2(n3560), .A(n3528), .ZN(n3530) );
  OAI21_X1 U3771 ( .B1(n3555), .B2(n3531), .A(n3530), .ZN(n3532) );
  NOR2_X1 U3772 ( .A1(\adder_stage4[0][16] ), .A2(\adder_stage4[1][16] ), .ZN(
        n3538) );
  INV_X1 U3773 ( .A(n3538), .ZN(n3535) );
  NAND2_X1 U3774 ( .A1(\adder_stage4[0][16] ), .A2(\adder_stage4[1][16] ), 
        .ZN(n3537) );
  NAND2_X1 U3775 ( .A1(n3535), .A2(n3537), .ZN(n3536) );
  XOR2_X1 U3776 ( .A(n3539), .B(n3536), .Z(m_data_out_y[16]) );
  OAI21_X1 U3777 ( .B1(n3539), .B2(n3538), .A(n3537), .ZN(n3612) );
  OR2_X1 U3778 ( .A1(\adder_stage4[0][17] ), .A2(\adder_stage4[1][17] ), .ZN(
        n3610) );
  NAND2_X1 U3779 ( .A1(\adder_stage4[0][17] ), .A2(\adder_stage4[1][17] ), 
        .ZN(n3609) );
  INV_X1 U3780 ( .A(n3609), .ZN(n3540) );
  AOI21_X1 U3781 ( .B1(n3612), .B2(n3610), .A(n3540), .ZN(n3545) );
  NOR2_X1 U3782 ( .A1(\adder_stage4[0][18] ), .A2(\adder_stage4[1][18] ), .ZN(
        n3544) );
  INV_X1 U3783 ( .A(n3544), .ZN(n3541) );
  NAND2_X1 U3784 ( .A1(\adder_stage4[0][18] ), .A2(\adder_stage4[1][18] ), 
        .ZN(n3543) );
  NAND2_X1 U3785 ( .A1(n3541), .A2(n3543), .ZN(n3542) );
  XOR2_X1 U3786 ( .A(n3545), .B(n3542), .Z(m_data_out_y[18]) );
  OAI21_X1 U3787 ( .B1(n3545), .B2(n3544), .A(n3543), .ZN(n3550) );
  OR2_X1 U3788 ( .A1(\adder_stage4[0][19] ), .A2(\adder_stage4[1][19] ), .ZN(
        n3549) );
  NAND2_X1 U3789 ( .A1(\adder_stage4[0][19] ), .A2(\adder_stage4[1][19] ), 
        .ZN(n3547) );
  NAND2_X1 U3790 ( .A1(n3549), .A2(n3547), .ZN(n3546) );
  XNOR2_X1 U3791 ( .A(n3550), .B(n3546), .ZN(m_data_out_y[19]) );
  INV_X1 U3792 ( .A(n3547), .ZN(n3548) );
  AOI21_X1 U3793 ( .B1(n3550), .B2(n3549), .A(n3548), .ZN(n3554) );
  OR2_X1 U3794 ( .A1(\adder_stage4[0][20] ), .A2(\adder_stage4[1][20] ), .ZN(
        n3552) );
  NAND2_X1 U3795 ( .A1(\adder_stage4[0][20] ), .A2(\adder_stage4[1][20] ), 
        .ZN(n3551) );
  NAND2_X1 U3796 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  XOR2_X1 U3797 ( .A(n3554), .B(n3553), .Z(m_data_out_y[20]) );
  OAI21_X1 U3798 ( .B1(n3615), .B2(n3556), .A(n3420), .ZN(n3591) );
  INV_X1 U3799 ( .A(n3591), .ZN(n3563) );
  INV_X1 U3800 ( .A(n3557), .ZN(n3590) );
  NAND2_X1 U3801 ( .A1(n3590), .A2(n3588), .ZN(n3558) );
  XOR2_X1 U3802 ( .A(n3563), .B(n3558), .Z(m_data_out_y[12]) );
  INV_X1 U3803 ( .A(n3559), .ZN(n3562) );
  INV_X1 U3804 ( .A(n3560), .ZN(n3561) );
  OAI21_X1 U3805 ( .B1(n3563), .B2(n3562), .A(n3561), .ZN(n3571) );
  INV_X1 U3806 ( .A(n3564), .ZN(n3570) );
  NAND2_X1 U3807 ( .A1(n3570), .A2(n3568), .ZN(n3565) );
  XNOR2_X1 U3808 ( .A(n3571), .B(n3565), .ZN(m_data_out_y[14]) );
  OR2_X1 U3809 ( .A1(\adder_stage4[0][0] ), .A2(\adder_stage4[1][0] ), .ZN(
        n3567) );
  AND2_X1 U3810 ( .A1(n3567), .A2(n3566), .ZN(m_data_out_y[0]) );
  INV_X1 U3811 ( .A(n3568), .ZN(n3569) );
  AOI21_X1 U3812 ( .B1(n3571), .B2(n3570), .A(n3569), .ZN(n3576) );
  INV_X1 U3813 ( .A(n3572), .ZN(n3574) );
  NAND2_X1 U3814 ( .A1(n3574), .A2(n3573), .ZN(n3575) );
  XOR2_X1 U3815 ( .A(n3576), .B(n3575), .Z(m_data_out_y[15]) );
  INV_X1 U3816 ( .A(n3577), .ZN(n3580) );
  INV_X1 U3817 ( .A(n3578), .ZN(n3579) );
  OAI21_X1 U3818 ( .B1(n3615), .B2(n3580), .A(n3579), .ZN(n3600) );
  INV_X1 U3819 ( .A(n3581), .ZN(n3598) );
  INV_X1 U3820 ( .A(n3597), .ZN(n3582) );
  AOI21_X1 U3821 ( .B1(n3600), .B2(n3598), .A(n3582), .ZN(n3587) );
  INV_X1 U3822 ( .A(n3583), .ZN(n3585) );
  NAND2_X1 U3823 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  XOR2_X1 U3824 ( .A(n3587), .B(n3586), .Z(m_data_out_y[11]) );
  INV_X1 U3825 ( .A(n3588), .ZN(n3589) );
  AOI21_X1 U3826 ( .B1(n3591), .B2(n3590), .A(n3589), .ZN(n3596) );
  INV_X1 U3827 ( .A(n3592), .ZN(n3594) );
  NAND2_X1 U3828 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  XOR2_X1 U3829 ( .A(n3596), .B(n3595), .Z(m_data_out_y[13]) );
  NAND2_X1 U3830 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  XNOR2_X1 U3831 ( .A(n3600), .B(n3599), .ZN(m_data_out_y[10]) );
  INV_X1 U3832 ( .A(n3601), .ZN(n3636) );
  AOI21_X1 U3833 ( .B1(n3636), .B2(n3603), .A(n3602), .ZN(n3625) );
  OAI21_X1 U3834 ( .B1(n3625), .B2(n3621), .A(n3622), .ZN(n3608) );
  INV_X1 U3835 ( .A(n3604), .ZN(n3606) );
  NAND2_X1 U3836 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U3837 ( .A(n3608), .B(n3607), .ZN(m_data_out_y[7]) );
  NAND2_X1 U3838 ( .A1(n3610), .A2(n3609), .ZN(n3611) );
  XNOR2_X1 U3839 ( .A(n3612), .B(n3611), .ZN(m_data_out_y[17]) );
  OAI21_X1 U3840 ( .B1(n3615), .B2(n3614), .A(n3613), .ZN(n3620) );
  INV_X1 U3841 ( .A(n3616), .ZN(n3618) );
  NAND2_X1 U3842 ( .A1(n3618), .A2(n3617), .ZN(n3619) );
  XNOR2_X1 U3843 ( .A(n3620), .B(n3619), .ZN(m_data_out_y[9]) );
  INV_X1 U3844 ( .A(n3621), .ZN(n3623) );
  NAND2_X1 U3845 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  XOR2_X1 U3846 ( .A(n3625), .B(n3624), .Z(m_data_out_y[6]) );
  INV_X1 U3847 ( .A(n3626), .ZN(n3634) );
  INV_X1 U3848 ( .A(n3633), .ZN(n3627) );
  AOI21_X1 U3849 ( .B1(n3636), .B2(n3634), .A(n3627), .ZN(n3632) );
  INV_X1 U3850 ( .A(n3628), .ZN(n3630) );
  NAND2_X1 U3851 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  XOR2_X1 U3852 ( .A(n3632), .B(n3631), .Z(m_data_out_y[5]) );
  NAND2_X1 U3853 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  XNOR2_X1 U3854 ( .A(n3636), .B(n3635), .ZN(m_data_out_y[4]) );
  INV_X1 U3855 ( .A(n3637), .ZN(n3647) );
  OAI21_X1 U3856 ( .B1(n3647), .B2(n3643), .A(n3644), .ZN(n3642) );
  INV_X1 U3857 ( .A(n3638), .ZN(n3640) );
  NAND2_X1 U3858 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  XNOR2_X1 U3859 ( .A(n3642), .B(n3641), .ZN(m_data_out_y[3]) );
  INV_X1 U3860 ( .A(n3643), .ZN(n3645) );
  NAND2_X1 U3861 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  XOR2_X1 U3862 ( .A(n3647), .B(n3646), .Z(m_data_out_y[2]) );
  AOI21_X1 U3863 ( .B1(n8812), .B2(n3681), .A(n3979), .ZN(s_ready_x) );
  INV_X4 U3864 ( .A(n3649), .ZN(n8906) );
  BUF_X4 U3865 ( .A(n3438), .Z(n8902) );
  NAND2_X1 U3866 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n3666) );
  NOR2_X1 U3867 ( .A1(\ctrl_inst/state [1]), .A2(\ctrl_inst/state [0]), .ZN(
        n3984) );
  NAND2_X1 U3868 ( .A1(n3984), .A2(n8806), .ZN(n8392) );
  NAND2_X1 U3869 ( .A1(n8807), .A2(n8842), .ZN(n8347) );
  NOR2_X1 U3870 ( .A1(n8392), .A2(n8347), .ZN(n3654) );
  NAND2_X1 U3871 ( .A1(n3652), .A2(n3658), .ZN(n8348) );
  INV_X1 U3872 ( .A(n8348), .ZN(n3653) );
  NAND2_X1 U3873 ( .A1(n3654), .A2(n3653), .ZN(n8383) );
  AOI21_X1 U3874 ( .B1(n8388), .B2(n8383), .A(n8770), .ZN(n8374) );
  NAND2_X1 U3875 ( .A1(n8383), .A2(n8778), .ZN(n3655) );
  NOR2_X1 U3876 ( .A1(n3666), .A2(n3655), .ZN(n8375) );
  XOR2_X1 U3877 ( .A(\ctrl_inst/xmem_tracker [1]), .B(
        \ctrl_inst/xmem_tracker [0]), .Z(n3656) );
  AOI22_X1 U3878 ( .A1(n8374), .A2(\ctrl_inst/xmem_tracker [1]), .B1(n8375), 
        .B2(n3656), .ZN(n3657) );
  INV_X1 U3879 ( .A(n3657), .ZN(n10421) );
  NAND2_X1 U3880 ( .A1(n8375), .A2(n3658), .ZN(n3671) );
  NAND3_X1 U3881 ( .A1(n3671), .A2(n8778), .A3(\ctrl_inst/xmem_tracker [2]), 
        .ZN(n3659) );
  OAI21_X1 U3882 ( .B1(\ctrl_inst/xmem_tracker [2]), .B2(n3671), .A(n3659), 
        .ZN(n10420) );
  INV_X1 U3883 ( .A(n3681), .ZN(n3668) );
  NAND3_X1 U3884 ( .A1(n8806), .A2(n8813), .A3(\ctrl_inst/state [1]), .ZN(
        n3977) );
  NOR3_X1 U3885 ( .A1(n8388), .A2(n3979), .A3(n3977), .ZN(n8379) );
  NOR2_X1 U3886 ( .A1(\ctrl_inst/pline_cntr [0]), .A2(
        \ctrl_inst/pline_cntr [1]), .ZN(n3662) );
  NOR2_X1 U3887 ( .A1(\ctrl_inst/pline_cntr [2]), .A2(
        \ctrl_inst/pline_cntr [3]), .ZN(n3660) );
  NAND2_X1 U3888 ( .A1(n3662), .A2(n3660), .ZN(n8371) );
  NAND2_X1 U3889 ( .A1(n3984), .A2(\ctrl_inst/state [2]), .ZN(n8345) );
  NOR2_X1 U3890 ( .A1(n8371), .A2(n8345), .ZN(n3661) );
  NAND2_X1 U3891 ( .A1(n8911), .A2(n3661), .ZN(n8395) );
  NAND2_X1 U3892 ( .A1(n8814), .A2(\ctrl_inst/pline_cntr [3]), .ZN(n3664) );
  INV_X1 U3893 ( .A(n3662), .ZN(n3663) );
  NOR2_X1 U3894 ( .A1(n3664), .A2(n3663), .ZN(n8352) );
  OAI211_X1 U3895 ( .C1(n8352), .C2(\ctrl_inst/state [1]), .A(
        \ctrl_inst/state [0]), .B(n8806), .ZN(n3665) );
  NOR2_X1 U3896 ( .A1(n3666), .A2(n3665), .ZN(n8382) );
  NOR2_X1 U3897 ( .A1(n8382), .A2(reset), .ZN(n3667) );
  NAND2_X1 U3898 ( .A1(n8395), .A2(n3667), .ZN(n3685) );
  AOI21_X1 U3899 ( .B1(n3668), .B2(n8379), .A(n3685), .ZN(n3670) );
  INV_X1 U3900 ( .A(reset), .ZN(n8394) );
  NAND2_X1 U3901 ( .A1(\ctrl_inst/state [0]), .A2(n8394), .ZN(n3669) );
  NOR2_X1 U3902 ( .A1(n3669), .A2(\ctrl_inst/state [2]), .ZN(n8355) );
  OAI22_X1 U3903 ( .A1(n3670), .A2(n8355), .B1(m_valid_y), .B2(n3685), .ZN(
        n8870) );
  NOR2_X1 U3904 ( .A1(n3671), .A2(n8843), .ZN(n3674) );
  AOI22_X1 U3905 ( .A1(n3674), .A2(\ctrl_inst/xmem_tracker [3]), .B1(
        \ctrl_inst/xmem_tracker [4]), .B2(n8778), .ZN(n3673) );
  INV_X1 U3906 ( .A(n8375), .ZN(n3672) );
  NOR2_X1 U3907 ( .A1(n3672), .A2(n8348), .ZN(n3677) );
  NOR2_X1 U3908 ( .A1(n3673), .A2(n3677), .ZN(n10418) );
  AOI22_X1 U3909 ( .A1(n3677), .A2(\ctrl_inst/xmem_tracker [5]), .B1(
        \ctrl_inst/xmem_tracker [6]), .B2(n8778), .ZN(n8871) );
  INV_X1 U3910 ( .A(n3674), .ZN(n3676) );
  NAND3_X1 U3911 ( .A1(n3676), .A2(n8778), .A3(\ctrl_inst/xmem_tracker [3]), 
        .ZN(n3675) );
  OAI21_X1 U3912 ( .B1(\ctrl_inst/xmem_tracker [3]), .B2(n3676), .A(n3675), 
        .ZN(n10419) );
  INV_X1 U3913 ( .A(n3677), .ZN(n3679) );
  NAND3_X1 U3914 ( .A1(n3679), .A2(n8778), .A3(\ctrl_inst/xmem_tracker [5]), 
        .ZN(n3678) );
  OAI21_X1 U3915 ( .B1(\ctrl_inst/xmem_tracker [5]), .B2(n3679), .A(n3678), 
        .ZN(n3378) );
  OR2_X1 U3916 ( .A1(n3680), .A2(n8806), .ZN(n8369) );
  NOR2_X1 U3917 ( .A1(n3681), .A2(n3977), .ZN(n3683) );
  NOR2_X1 U3918 ( .A1(n8383), .A2(n3682), .ZN(n8378) );
  AOI21_X1 U3919 ( .B1(n3666), .B2(n3683), .A(n8378), .ZN(n8384) );
  OAI21_X1 U3920 ( .B1(conv_done), .B2(n8369), .A(n8384), .ZN(n3684) );
  NOR2_X1 U3921 ( .A1(n3983), .A2(reset), .ZN(n3985) );
  NAND2_X1 U3922 ( .A1(n3985), .A2(n8379), .ZN(n3986) );
  INV_X1 U3923 ( .A(n8355), .ZN(n8781) );
  MUX2_X1 U3924 ( .A(n8781), .B(n8815), .S(n3983), .Z(n3686) );
  NAND2_X1 U3925 ( .A1(n3986), .A2(n3686), .ZN(n3387) );
  BUF_X2 U3926 ( .A(n4444), .Z(n8251) );
  NOR2_X1 U3927 ( .A1(\adder_stage1[6][2] ), .A2(\adder_stage1[7][2] ), .ZN(
        n3761) );
  NOR2_X1 U3928 ( .A1(\adder_stage1[6][3] ), .A2(\adder_stage1[7][3] ), .ZN(
        n3763) );
  NOR2_X1 U3929 ( .A1(n3761), .A2(n3763), .ZN(n3688) );
  NOR2_X1 U3930 ( .A1(\adder_stage1[6][1] ), .A2(\adder_stage1[7][1] ), .ZN(
        n3937) );
  NAND2_X1 U3931 ( .A1(\adder_stage1[6][0] ), .A2(\adder_stage1[7][0] ), .ZN(
        n3940) );
  NAND2_X1 U3932 ( .A1(\adder_stage1[6][1] ), .A2(\adder_stage1[7][1] ), .ZN(
        n3938) );
  OAI21_X1 U3933 ( .B1(n3937), .B2(n3940), .A(n3938), .ZN(n3727) );
  NAND2_X1 U3934 ( .A1(\adder_stage1[6][2] ), .A2(\adder_stage1[7][2] ), .ZN(
        n3760) );
  NAND2_X1 U3935 ( .A1(\adder_stage1[6][3] ), .A2(\adder_stage1[7][3] ), .ZN(
        n3764) );
  OAI21_X1 U3936 ( .B1(n3763), .B2(n3760), .A(n3764), .ZN(n3687) );
  AOI21_X1 U3937 ( .B1(n3688), .B2(n3727), .A(n3687), .ZN(n5422) );
  INV_X1 U3938 ( .A(n5422), .ZN(n3813) );
  NOR2_X1 U3939 ( .A1(\adder_stage1[6][4] ), .A2(\adder_stage1[7][4] ), .ZN(
        n3742) );
  NOR2_X1 U3940 ( .A1(\adder_stage1[6][5] ), .A2(\adder_stage1[7][5] ), .ZN(
        n3814) );
  NOR2_X1 U3941 ( .A1(n3742), .A2(n3814), .ZN(n5413) );
  NAND2_X1 U3942 ( .A1(\adder_stage1[6][4] ), .A2(\adder_stage1[7][4] ), .ZN(
        n3810) );
  NAND2_X1 U3943 ( .A1(\adder_stage1[6][5] ), .A2(\adder_stage1[7][5] ), .ZN(
        n3815) );
  OAI21_X1 U3944 ( .B1(n3814), .B2(n3810), .A(n3815), .ZN(n5418) );
  AOI21_X1 U3945 ( .B1(n3813), .B2(n5413), .A(n5418), .ZN(n3757) );
  NOR2_X1 U3946 ( .A1(\adder_stage1[6][6] ), .A2(\adder_stage1[7][6] ), .ZN(
        n5412) );
  NAND2_X1 U3947 ( .A1(\adder_stage1[6][6] ), .A2(\adder_stage1[7][6] ), .ZN(
        n5415) );
  OAI21_X1 U3948 ( .B1(n3757), .B2(n5412), .A(n5415), .ZN(n3691) );
  NOR2_X1 U3949 ( .A1(\adder_stage1[6][7] ), .A2(\adder_stage1[7][7] ), .ZN(
        n5416) );
  INV_X1 U3950 ( .A(n5416), .ZN(n3689) );
  NAND2_X1 U3951 ( .A1(\adder_stage1[6][7] ), .A2(\adder_stage1[7][7] ), .ZN(
        n5414) );
  NAND2_X1 U3952 ( .A1(n3689), .A2(n5414), .ZN(n3690) );
  XNOR2_X1 U3953 ( .A(n3691), .B(n3690), .ZN(n3692) );
  AOI22_X1 U3954 ( .A1(n8336), .A2(\adder_stage2[3][7] ), .B1(n8251), .B2(
        n3692), .ZN(n3693) );
  INV_X1 U3955 ( .A(n3693), .ZN(n9846) );
  NOR2_X1 U3956 ( .A1(\adder_stage2[2][2] ), .A2(\adder_stage2[3][2] ), .ZN(
        n3860) );
  NOR2_X1 U3957 ( .A1(\adder_stage2[2][3] ), .A2(\adder_stage2[3][3] ), .ZN(
        n3826) );
  NOR2_X1 U3958 ( .A1(n3860), .A2(n3826), .ZN(n3695) );
  NOR2_X1 U3959 ( .A1(\adder_stage2[2][1] ), .A2(\adder_stage2[3][1] ), .ZN(
        n3846) );
  NAND2_X1 U3960 ( .A1(\adder_stage2[2][0] ), .A2(\adder_stage2[3][0] ), .ZN(
        n3849) );
  NAND2_X1 U3961 ( .A1(\adder_stage2[2][1] ), .A2(\adder_stage2[3][1] ), .ZN(
        n3847) );
  OAI21_X1 U3962 ( .B1(n3846), .B2(n3849), .A(n3847), .ZN(n3825) );
  NAND2_X1 U3963 ( .A1(\adder_stage2[2][2] ), .A2(\adder_stage2[3][2] ), .ZN(
        n3861) );
  NAND2_X1 U3964 ( .A1(\adder_stage2[2][3] ), .A2(\adder_stage2[3][3] ), .ZN(
        n3827) );
  OAI21_X1 U3965 ( .B1(n3826), .B2(n3861), .A(n3827), .ZN(n3694) );
  AOI21_X1 U3966 ( .B1(n3695), .B2(n3825), .A(n3694), .ZN(n3853) );
  NOR2_X1 U3967 ( .A1(\adder_stage2[2][4] ), .A2(\adder_stage2[3][4] ), .ZN(
        n3910) );
  NOR2_X1 U3968 ( .A1(\adder_stage2[2][5] ), .A2(\adder_stage2[3][5] ), .ZN(
        n3912) );
  NOR2_X1 U3969 ( .A1(n3910), .A2(n3912), .ZN(n3855) );
  NOR2_X1 U3970 ( .A1(\adder_stage2[2][6] ), .A2(\adder_stage2[3][6] ), .ZN(
        n3968) );
  NOR2_X1 U3971 ( .A1(\adder_stage2[2][7] ), .A2(\adder_stage2[3][7] ), .ZN(
        n3970) );
  NOR2_X1 U3972 ( .A1(n3968), .A2(n3970), .ZN(n3697) );
  NAND2_X1 U3973 ( .A1(n3855), .A2(n3697), .ZN(n3699) );
  NAND2_X1 U3974 ( .A1(\adder_stage2[2][4] ), .A2(\adder_stage2[3][4] ), .ZN(
        n3961) );
  NAND2_X1 U3975 ( .A1(\adder_stage2[2][5] ), .A2(\adder_stage2[3][5] ), .ZN(
        n3913) );
  OAI21_X1 U3976 ( .B1(n3912), .B2(n3961), .A(n3913), .ZN(n3854) );
  NAND2_X1 U3977 ( .A1(\adder_stage2[2][6] ), .A2(\adder_stage2[3][6] ), .ZN(
        n3967) );
  NAND2_X1 U3978 ( .A1(\adder_stage2[2][7] ), .A2(\adder_stage2[3][7] ), .ZN(
        n3971) );
  OAI21_X1 U3979 ( .B1(n3970), .B2(n3967), .A(n3971), .ZN(n3696) );
  AOI21_X1 U3980 ( .B1(n3697), .B2(n3854), .A(n3696), .ZN(n3698) );
  OAI21_X1 U3981 ( .B1(n3853), .B2(n3699), .A(n3698), .ZN(n3732) );
  NOR2_X1 U3982 ( .A1(\adder_stage2[2][10] ), .A2(\adder_stage2[3][10] ), .ZN(
        n3837) );
  NOR2_X1 U3983 ( .A1(\adder_stage2[3][11] ), .A2(\adder_stage2[2][11] ), .ZN(
        n3839) );
  NOR2_X1 U3984 ( .A1(n3837), .A2(n3839), .ZN(n3701) );
  NOR2_X1 U3985 ( .A1(\adder_stage2[2][8] ), .A2(\adder_stage2[3][8] ), .ZN(
        n3747) );
  NOR2_X1 U3986 ( .A1(\adder_stage2[2][9] ), .A2(\adder_stage2[3][9] ), .ZN(
        n3748) );
  NOR2_X1 U3987 ( .A1(n3747), .A2(n3748), .ZN(n3833) );
  NAND2_X1 U3988 ( .A1(n3701), .A2(n3833), .ZN(n3928) );
  NOR2_X1 U3989 ( .A1(\adder_stage2[2][12] ), .A2(\adder_stage2[3][12] ), .ZN(
        n3930) );
  NOR2_X1 U3990 ( .A1(n3928), .A2(n3930), .ZN(n3703) );
  NAND2_X1 U3991 ( .A1(\adder_stage2[2][8] ), .A2(\adder_stage2[3][8] ), .ZN(
        n3746) );
  NAND2_X1 U3992 ( .A1(\adder_stage2[2][9] ), .A2(\adder_stage2[3][9] ), .ZN(
        n3749) );
  OAI21_X1 U3993 ( .B1(n3748), .B2(n3746), .A(n3749), .ZN(n3834) );
  NAND2_X1 U3994 ( .A1(\adder_stage2[2][10] ), .A2(\adder_stage2[3][10] ), 
        .ZN(n3955) );
  NAND2_X1 U3995 ( .A1(\adder_stage2[2][11] ), .A2(\adder_stage2[3][11] ), 
        .ZN(n3840) );
  OAI21_X1 U3996 ( .B1(n3839), .B2(n3955), .A(n3840), .ZN(n3700) );
  AOI21_X1 U3997 ( .B1(n3701), .B2(n3834), .A(n3700), .ZN(n3927) );
  NAND2_X1 U3998 ( .A1(\adder_stage2[2][12] ), .A2(\adder_stage2[3][12] ), 
        .ZN(n3931) );
  OAI21_X1 U3999 ( .B1(n3927), .B2(n3930), .A(n3931), .ZN(n3702) );
  AOI21_X1 U4000 ( .B1(n3732), .B2(n3703), .A(n3702), .ZN(n3869) );
  NOR2_X1 U4001 ( .A1(\adder_stage2[2][13] ), .A2(\adder_stage2[3][13] ), .ZN(
        n3868) );
  INV_X1 U4002 ( .A(n3868), .ZN(n3704) );
  NAND2_X1 U4003 ( .A1(\adder_stage2[2][13] ), .A2(\adder_stage2[3][13] ), 
        .ZN(n3867) );
  NAND2_X1 U4004 ( .A1(n3704), .A2(n3867), .ZN(n3705) );
  XOR2_X1 U4005 ( .A(n3869), .B(n3705), .Z(n3706) );
  AOI22_X1 U4006 ( .A1(n8273), .A2(\adder_stage3[1][13] ), .B1(n8251), .B2(
        n3706), .ZN(n3707) );
  INV_X1 U4007 ( .A(n3707), .ZN(n9735) );
  BUF_X2 U4008 ( .A(n6352), .Z(n8272) );
  NOR2_X1 U4009 ( .A1(\adder_stage3[0][9] ), .A2(\adder_stage3[1][9] ), .ZN(
        n3988) );
  NAND2_X1 U4010 ( .A1(\adder_stage3[0][8] ), .A2(\adder_stage3[1][8] ), .ZN(
        n4019) );
  NAND2_X1 U4011 ( .A1(\adder_stage3[0][9] ), .A2(\adder_stage3[1][9] ), .ZN(
        n3989) );
  OAI21_X1 U4012 ( .B1(n3988), .B2(n4019), .A(n3989), .ZN(n4006) );
  NOR2_X1 U4013 ( .A1(\adder_stage3[0][11] ), .A2(\adder_stage3[1][11] ), .ZN(
        n4011) );
  NAND2_X1 U4014 ( .A1(\adder_stage3[0][10] ), .A2(\adder_stage3[1][10] ), 
        .ZN(n4025) );
  NAND2_X1 U4015 ( .A1(\adder_stage3[0][11] ), .A2(\adder_stage3[1][11] ), 
        .ZN(n4012) );
  OAI21_X1 U4016 ( .B1(n4011), .B2(n4025), .A(n4012), .ZN(n3995) );
  OR2_X1 U4017 ( .A1(n4006), .A2(n3995), .ZN(n3712) );
  NAND2_X1 U4018 ( .A1(\adder_stage3[0][12] ), .A2(\adder_stage3[1][12] ), 
        .ZN(n3999) );
  INV_X1 U4019 ( .A(n3999), .ZN(n3711) );
  NOR2_X1 U4020 ( .A1(\adder_stage3[0][10] ), .A2(\adder_stage3[1][10] ), .ZN(
        n4009) );
  NOR2_X1 U4021 ( .A1(n4009), .A2(n4011), .ZN(n3996) );
  NOR2_X1 U4022 ( .A1(n3996), .A2(n3711), .ZN(n3709) );
  INV_X1 U4023 ( .A(n3995), .ZN(n3708) );
  NOR2_X1 U4024 ( .A1(\adder_stage3[0][12] ), .A2(\adder_stage3[1][12] ), .ZN(
        n3713) );
  INV_X1 U4025 ( .A(n3713), .ZN(n4000) );
  AOI21_X1 U4026 ( .B1(n3709), .B2(n3708), .A(n3713), .ZN(n3710) );
  OAI21_X1 U4027 ( .B1(n3712), .B2(n3711), .A(n3710), .ZN(n4040) );
  NOR2_X1 U4028 ( .A1(\adder_stage3[0][13] ), .A2(\adder_stage3[1][13] ), .ZN(
        n3721) );
  NAND2_X1 U4029 ( .A1(\adder_stage3[0][13] ), .A2(\adder_stage3[1][13] ), 
        .ZN(n4041) );
  NOR2_X1 U4030 ( .A1(\adder_stage3[0][8] ), .A2(\adder_stage3[1][8] ), .ZN(
        n4018) );
  NOR2_X1 U4031 ( .A1(n4018), .A2(n3988), .ZN(n4005) );
  NAND2_X1 U4032 ( .A1(n4005), .A2(n3996), .ZN(n3998) );
  NOR2_X1 U4033 ( .A1(n3998), .A2(n3713), .ZN(n4038) );
  NOR2_X1 U4034 ( .A1(\adder_stage3[0][1] ), .A2(\adder_stage3[1][1] ), .ZN(
        n4878) );
  NAND2_X1 U4035 ( .A1(\adder_stage3[0][0] ), .A2(\adder_stage3[1][0] ), .ZN(
        n6089) );
  NAND2_X1 U4036 ( .A1(\adder_stage3[0][1] ), .A2(\adder_stage3[1][1] ), .ZN(
        n4879) );
  OAI21_X1 U4037 ( .B1(n4878), .B2(n6089), .A(n4879), .ZN(n4089) );
  NOR2_X1 U4038 ( .A1(\adder_stage3[0][2] ), .A2(\adder_stage3[1][2] ), .ZN(
        n4871) );
  NOR2_X1 U4039 ( .A1(\adder_stage3[0][3] ), .A2(\adder_stage3[1][3] ), .ZN(
        n4090) );
  NOR2_X1 U4040 ( .A1(n4871), .A2(n4090), .ZN(n3715) );
  NAND2_X1 U4041 ( .A1(\adder_stage3[0][2] ), .A2(\adder_stage3[1][2] ), .ZN(
        n4872) );
  NAND2_X1 U4042 ( .A1(\adder_stage3[0][3] ), .A2(\adder_stage3[1][3] ), .ZN(
        n4091) );
  OAI21_X1 U4043 ( .B1(n4090), .B2(n4872), .A(n4091), .ZN(n3714) );
  AOI21_X1 U4044 ( .B1(n4089), .B2(n3715), .A(n3714), .ZN(n4057) );
  NOR2_X1 U4045 ( .A1(\adder_stage3[0][4] ), .A2(\adder_stage3[1][4] ), .ZN(
        n4058) );
  NOR2_X1 U4046 ( .A1(\adder_stage3[0][5] ), .A2(\adder_stage3[1][5] ), .ZN(
        n4060) );
  NOR2_X1 U4047 ( .A1(n4058), .A2(n4060), .ZN(n4068) );
  NOR2_X1 U4048 ( .A1(\adder_stage3[0][6] ), .A2(\adder_stage3[1][6] ), .ZN(
        n4076) );
  NOR2_X1 U4049 ( .A1(\adder_stage3[0][7] ), .A2(\adder_stage3[1][7] ), .ZN(
        n4069) );
  NOR2_X1 U4050 ( .A1(n4076), .A2(n4069), .ZN(n3717) );
  NAND2_X1 U4051 ( .A1(n4068), .A2(n3717), .ZN(n3719) );
  NAND2_X1 U4052 ( .A1(\adder_stage3[0][4] ), .A2(\adder_stage3[1][4] ), .ZN(
        n4083) );
  NAND2_X1 U4053 ( .A1(\adder_stage3[0][5] ), .A2(\adder_stage3[1][5] ), .ZN(
        n4061) );
  OAI21_X1 U4054 ( .B1(n4060), .B2(n4083), .A(n4061), .ZN(n4067) );
  NAND2_X1 U4055 ( .A1(\adder_stage3[0][6] ), .A2(\adder_stage3[1][6] ), .ZN(
        n4077) );
  NAND2_X1 U4056 ( .A1(\adder_stage3[0][7] ), .A2(\adder_stage3[1][7] ), .ZN(
        n4070) );
  OAI21_X1 U4057 ( .B1(n4069), .B2(n4077), .A(n4070), .ZN(n3716) );
  AOI21_X1 U4058 ( .B1(n4067), .B2(n3717), .A(n3716), .ZN(n3718) );
  OAI21_X1 U4059 ( .B1(n4057), .B2(n3719), .A(n3718), .ZN(n4037) );
  INV_X1 U4060 ( .A(n3721), .ZN(n4042) );
  NAND3_X1 U4061 ( .A1(n4038), .A2(n4037), .A3(n4042), .ZN(n3720) );
  OAI211_X1 U4062 ( .C1(n4040), .C2(n3721), .A(n4041), .B(n3720), .ZN(n4034)
         );
  OR2_X1 U4063 ( .A1(\adder_stage3[0][14] ), .A2(\adder_stage3[1][14] ), .ZN(
        n4032) );
  NAND2_X1 U4064 ( .A1(\adder_stage3[0][14] ), .A2(\adder_stage3[1][14] ), 
        .ZN(n4031) );
  INV_X1 U4065 ( .A(n4031), .ZN(n3722) );
  AOI21_X1 U4066 ( .B1(n4034), .B2(n4032), .A(n3722), .ZN(n7472) );
  NOR2_X1 U4067 ( .A1(\adder_stage3[0][15] ), .A2(\adder_stage3[1][15] ), .ZN(
        n7471) );
  INV_X1 U4068 ( .A(n7471), .ZN(n3723) );
  NAND2_X1 U4069 ( .A1(\adder_stage3[0][15] ), .A2(\adder_stage3[1][15] ), 
        .ZN(n7470) );
  NAND2_X1 U4070 ( .A1(n3723), .A2(n7470), .ZN(n3724) );
  XOR2_X1 U4071 ( .A(n7472), .B(n3724), .Z(n3725) );
  AOI22_X1 U4072 ( .A1(n8273), .A2(\adder_stage4[0][15] ), .B1(n8272), .B2(
        n3725), .ZN(n3726) );
  INV_X1 U4073 ( .A(n3726), .ZN(n9672) );
  INV_X1 U4074 ( .A(n3727), .ZN(n3762) );
  INV_X1 U4075 ( .A(n3761), .ZN(n3728) );
  NAND2_X1 U4076 ( .A1(n3728), .A2(n3760), .ZN(n3729) );
  XOR2_X1 U4077 ( .A(n3762), .B(n3729), .Z(n3730) );
  AOI22_X1 U4078 ( .A1(n7855), .A2(\adder_stage2[3][2] ), .B1(n8251), .B2(
        n3730), .ZN(n3731) );
  INV_X1 U4079 ( .A(n3731), .ZN(n9851) );
  INV_X1 U4080 ( .A(n3732), .ZN(n3929) );
  INV_X1 U4081 ( .A(n3747), .ZN(n3733) );
  NAND2_X1 U4082 ( .A1(n3733), .A2(n3746), .ZN(n3734) );
  XOR2_X1 U4083 ( .A(n3929), .B(n3734), .Z(n3735) );
  AOI22_X1 U4084 ( .A1(n8273), .A2(\adder_stage3[1][8] ), .B1(n8272), .B2(
        n3735), .ZN(n3736) );
  INV_X1 U4085 ( .A(n3736), .ZN(n9740) );
  BUF_X2 U4086 ( .A(n4444), .Z(n4311) );
  NOR2_X1 U4087 ( .A1(\x_mult_f[2][2] ), .A2(\x_mult_f[3][2] ), .ZN(n3944) );
  NOR2_X1 U4088 ( .A1(\x_mult_f[2][3] ), .A2(\x_mult_f[3][3] ), .ZN(n3920) );
  NOR2_X1 U4089 ( .A1(n3944), .A2(n3920), .ZN(n3738) );
  NOR2_X1 U4090 ( .A1(\x_mult_f[2][1] ), .A2(\x_mult_f[3][1] ), .ZN(n4305) );
  NAND2_X1 U4091 ( .A1(\x_mult_f[2][0] ), .A2(\x_mult_f[3][0] ), .ZN(n4308) );
  NAND2_X1 U4092 ( .A1(\x_mult_f[2][1] ), .A2(\x_mult_f[3][1] ), .ZN(n4306) );
  OAI21_X1 U4093 ( .B1(n4305), .B2(n4308), .A(n4306), .ZN(n3919) );
  NAND2_X1 U4094 ( .A1(\x_mult_f[2][2] ), .A2(\x_mult_f[3][2] ), .ZN(n3945) );
  NAND2_X1 U4095 ( .A1(\x_mult_f[2][3] ), .A2(\x_mult_f[3][3] ), .ZN(n3921) );
  OAI21_X1 U4096 ( .B1(n3920), .B2(n3945), .A(n3921), .ZN(n3737) );
  AOI21_X1 U4097 ( .B1(n3738), .B2(n3919), .A(n3737), .ZN(n3799) );
  INV_X1 U4098 ( .A(n3799), .ZN(n3902) );
  NOR2_X1 U4099 ( .A1(\x_mult_f[2][4] ), .A2(\x_mult_f[3][4] ), .ZN(n3794) );
  INV_X1 U4100 ( .A(n3794), .ZN(n3901) );
  NAND2_X1 U4101 ( .A1(\x_mult_f[2][4] ), .A2(\x_mult_f[3][4] ), .ZN(n3899) );
  NAND2_X1 U4102 ( .A1(n3901), .A2(n3899), .ZN(n3739) );
  XNOR2_X1 U4103 ( .A(n3902), .B(n3739), .ZN(n3740) );
  AOI22_X1 U4104 ( .A1(n8088), .A2(\adder_stage1[1][4] ), .B1(n4311), .B2(
        n3740), .ZN(n3741) );
  INV_X1 U4105 ( .A(n3741), .ZN(n10148) );
  INV_X1 U4106 ( .A(n3742), .ZN(n3812) );
  NAND2_X1 U4107 ( .A1(n3812), .A2(n3810), .ZN(n3743) );
  XNOR2_X1 U4108 ( .A(n3813), .B(n3743), .ZN(n3744) );
  AOI22_X1 U4109 ( .A1(n8336), .A2(\adder_stage2[3][4] ), .B1(n8251), .B2(
        n3744), .ZN(n3745) );
  INV_X1 U4110 ( .A(n3745), .ZN(n9849) );
  OAI21_X1 U4111 ( .B1(n3929), .B2(n3747), .A(n3746), .ZN(n3752) );
  INV_X1 U4112 ( .A(n3748), .ZN(n3750) );
  NAND2_X1 U4113 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  XNOR2_X1 U4114 ( .A(n3752), .B(n3751), .ZN(n3753) );
  AOI22_X1 U4115 ( .A1(n8306), .A2(\adder_stage3[1][9] ), .B1(n8272), .B2(
        n3753), .ZN(n3754) );
  INV_X1 U4116 ( .A(n3754), .ZN(n9739) );
  INV_X1 U4117 ( .A(n5412), .ZN(n3755) );
  NAND2_X1 U4118 ( .A1(n3755), .A2(n5415), .ZN(n3756) );
  XOR2_X1 U4119 ( .A(n3757), .B(n3756), .Z(n3758) );
  AOI22_X1 U4120 ( .A1(n7855), .A2(\adder_stage2[3][6] ), .B1(n8251), .B2(
        n3758), .ZN(n3759) );
  INV_X1 U4121 ( .A(n3759), .ZN(n9847) );
  OAI21_X1 U4122 ( .B1(n3762), .B2(n3761), .A(n3760), .ZN(n3767) );
  INV_X1 U4123 ( .A(n3763), .ZN(n3765) );
  NAND2_X1 U4124 ( .A1(n3765), .A2(n3764), .ZN(n3766) );
  XNOR2_X1 U4125 ( .A(n3767), .B(n3766), .ZN(n3768) );
  AOI22_X1 U4126 ( .A1(n8336), .A2(\adder_stage2[3][3] ), .B1(n8251), .B2(
        n3768), .ZN(n3769) );
  INV_X1 U4127 ( .A(n3769), .ZN(n9850) );
  OR2_X1 U4128 ( .A1(\adder_stage2[2][0] ), .A2(\adder_stage2[3][0] ), .ZN(
        n3770) );
  AND2_X1 U4129 ( .A1(n3770), .A2(n3849), .ZN(n3771) );
  AOI22_X1 U4130 ( .A1(n8273), .A2(\adder_stage3[1][0] ), .B1(n8272), .B2(
        n3771), .ZN(n3772) );
  INV_X1 U4131 ( .A(n3772), .ZN(n9748) );
  NOR2_X1 U4132 ( .A1(\adder_stage1[0][2] ), .A2(\adder_stage1[1][2] ), .ZN(
        n4757) );
  NOR2_X1 U4133 ( .A1(\adder_stage1[0][3] ), .A2(\adder_stage1[1][3] ), .ZN(
        n4750) );
  NOR2_X1 U4134 ( .A1(n4757), .A2(n4750), .ZN(n3774) );
  NOR2_X1 U4135 ( .A1(\adder_stage1[0][1] ), .A2(\adder_stage1[1][1] ), .ZN(
        n4742) );
  NAND2_X1 U4136 ( .A1(\adder_stage1[0][0] ), .A2(\adder_stage1[1][0] ), .ZN(
        n4745) );
  NAND2_X1 U4137 ( .A1(\adder_stage1[0][1] ), .A2(\adder_stage1[1][1] ), .ZN(
        n4743) );
  OAI21_X1 U4138 ( .B1(n4742), .B2(n4745), .A(n4743), .ZN(n4749) );
  NAND2_X1 U4139 ( .A1(\adder_stage1[0][2] ), .A2(\adder_stage1[1][2] ), .ZN(
        n4758) );
  NAND2_X1 U4140 ( .A1(\adder_stage1[0][3] ), .A2(\adder_stage1[1][3] ), .ZN(
        n4751) );
  OAI21_X1 U4141 ( .B1(n4750), .B2(n4758), .A(n4751), .ZN(n3773) );
  AOI21_X1 U4142 ( .B1(n3774), .B2(n4749), .A(n3773), .ZN(n4672) );
  NOR2_X1 U4143 ( .A1(\adder_stage1[0][4] ), .A2(\adder_stage1[1][4] ), .ZN(
        n4673) );
  NOR2_X1 U4144 ( .A1(\adder_stage1[0][5] ), .A2(\adder_stage1[1][5] ), .ZN(
        n4675) );
  NOR2_X1 U4145 ( .A1(n4673), .A2(n4675), .ZN(n4683) );
  NOR2_X1 U4146 ( .A1(\adder_stage1[0][6] ), .A2(\adder_stage1[1][6] ), .ZN(
        n4712) );
  NOR2_X1 U4147 ( .A1(\adder_stage1[0][7] ), .A2(\adder_stage1[1][7] ), .ZN(
        n4714) );
  NOR2_X1 U4148 ( .A1(n4712), .A2(n4714), .ZN(n3776) );
  NAND2_X1 U4149 ( .A1(n4683), .A2(n3776), .ZN(n3778) );
  NAND2_X1 U4150 ( .A1(\adder_stage1[0][4] ), .A2(\adder_stage1[1][4] ), .ZN(
        n4764) );
  NAND2_X1 U4151 ( .A1(\adder_stage1[0][5] ), .A2(\adder_stage1[1][5] ), .ZN(
        n4676) );
  OAI21_X1 U4152 ( .B1(n4675), .B2(n4764), .A(n4676), .ZN(n4682) );
  NAND2_X1 U4153 ( .A1(\adder_stage1[0][6] ), .A2(\adder_stage1[1][6] ), .ZN(
        n4711) );
  NAND2_X1 U4154 ( .A1(\adder_stage1[0][7] ), .A2(\adder_stage1[1][7] ), .ZN(
        n4715) );
  OAI21_X1 U4155 ( .B1(n4714), .B2(n4711), .A(n4715), .ZN(n3775) );
  AOI21_X1 U4156 ( .B1(n3776), .B2(n4682), .A(n3775), .ZN(n3777) );
  OAI21_X1 U4157 ( .B1(n4672), .B2(n3778), .A(n3777), .ZN(n4688) );
  NOR2_X1 U4158 ( .A1(\adder_stage1[0][8] ), .A2(\adder_stage1[1][8] ), .ZN(
        n4689) );
  INV_X1 U4159 ( .A(n4689), .ZN(n4706) );
  OR2_X1 U4160 ( .A1(\adder_stage1[0][9] ), .A2(\adder_stage1[1][9] ), .ZN(
        n4691) );
  NAND2_X1 U4161 ( .A1(n4706), .A2(n4691), .ZN(n4697) );
  NOR2_X1 U4162 ( .A1(\adder_stage1[0][10] ), .A2(\adder_stage1[1][10] ), .ZN(
        n4698) );
  NOR2_X1 U4163 ( .A1(n4697), .A2(n4698), .ZN(n3782) );
  NAND2_X1 U4164 ( .A1(\adder_stage1[0][8] ), .A2(\adder_stage1[1][8] ), .ZN(
        n4705) );
  INV_X1 U4165 ( .A(n4705), .ZN(n3780) );
  NAND2_X1 U4166 ( .A1(\adder_stage1[0][9] ), .A2(\adder_stage1[1][9] ), .ZN(
        n4690) );
  INV_X1 U4167 ( .A(n4690), .ZN(n3779) );
  AOI21_X1 U4168 ( .B1(n4691), .B2(n3780), .A(n3779), .ZN(n4696) );
  NAND2_X1 U4169 ( .A1(\adder_stage1[0][10] ), .A2(\adder_stage1[1][10] ), 
        .ZN(n4699) );
  OAI21_X1 U4170 ( .B1(n4696), .B2(n4698), .A(n4699), .ZN(n3781) );
  AOI21_X1 U4171 ( .B1(n4688), .B2(n3782), .A(n3781), .ZN(n7310) );
  NOR2_X1 U4172 ( .A1(\adder_stage1[0][12] ), .A2(\adder_stage1[1][12] ), .ZN(
        n3783) );
  NOR2_X1 U4173 ( .A1(\adder_stage1[0][11] ), .A2(\adder_stage1[1][11] ), .ZN(
        n3892) );
  NOR3_X1 U4174 ( .A1(n7310), .A2(n3783), .A3(n3892), .ZN(n3786) );
  NAND2_X1 U4175 ( .A1(\adder_stage1[0][12] ), .A2(\adder_stage1[1][12] ), 
        .ZN(n3893) );
  INV_X1 U4176 ( .A(n3783), .ZN(n3894) );
  NAND2_X1 U4177 ( .A1(\adder_stage1[0][11] ), .A2(\adder_stage1[1][11] ), 
        .ZN(n3891) );
  INV_X1 U4178 ( .A(n3891), .ZN(n3784) );
  NAND2_X1 U4179 ( .A1(n3894), .A2(n3784), .ZN(n3785) );
  NAND2_X1 U4180 ( .A1(n3893), .A2(n3785), .ZN(n3880) );
  NOR2_X1 U4181 ( .A1(n3786), .A2(n3880), .ZN(n3788) );
  NOR2_X1 U4182 ( .A1(\adder_stage1[0][13] ), .A2(\adder_stage1[1][13] ), .ZN(
        n3875) );
  INV_X1 U4183 ( .A(n3875), .ZN(n3879) );
  NAND2_X1 U4184 ( .A1(\adder_stage1[0][13] ), .A2(\adder_stage1[1][13] ), 
        .ZN(n3877) );
  NAND2_X1 U4185 ( .A1(n3879), .A2(n3877), .ZN(n3787) );
  XOR2_X1 U4186 ( .A(n3788), .B(n3787), .Z(n3789) );
  AOI22_X1 U4187 ( .A1(n8398), .A2(\adder_stage2[0][13] ), .B1(n4311), .B2(
        n3789), .ZN(n3790) );
  INV_X1 U4188 ( .A(n3790), .ZN(n9891) );
  OR2_X1 U4189 ( .A1(\adder_stage1[6][0] ), .A2(\adder_stage1[7][0] ), .ZN(
        n3791) );
  AND2_X1 U4190 ( .A1(n3791), .A2(n3940), .ZN(n3792) );
  AOI22_X1 U4191 ( .A1(n8088), .A2(\adder_stage2[3][0] ), .B1(n8251), .B2(
        n3792), .ZN(n3793) );
  INV_X1 U4192 ( .A(n3793), .ZN(n9853) );
  NOR2_X1 U4193 ( .A1(\x_mult_f[2][5] ), .A2(\x_mult_f[3][5] ), .ZN(n3903) );
  NOR2_X1 U4194 ( .A1(n3794), .A2(n3903), .ZN(n3805) );
  NOR2_X1 U4195 ( .A1(\x_mult_f[2][6] ), .A2(\x_mult_f[3][6] ), .ZN(n4048) );
  NOR2_X1 U4196 ( .A1(\x_mult_f[2][7] ), .A2(\x_mult_f[3][7] ), .ZN(n4050) );
  NOR2_X1 U4197 ( .A1(n4048), .A2(n4050), .ZN(n3796) );
  NAND2_X1 U4198 ( .A1(n3805), .A2(n3796), .ZN(n3798) );
  NAND2_X1 U4199 ( .A1(\x_mult_f[2][5] ), .A2(\x_mult_f[3][5] ), .ZN(n3904) );
  OAI21_X1 U4200 ( .B1(n3903), .B2(n3899), .A(n3904), .ZN(n3804) );
  NAND2_X1 U4201 ( .A1(\x_mult_f[2][6] ), .A2(\x_mult_f[3][6] ), .ZN(n4047) );
  NAND2_X1 U4202 ( .A1(\x_mult_f[2][7] ), .A2(\x_mult_f[3][7] ), .ZN(n4051) );
  OAI21_X1 U4203 ( .B1(n4050), .B2(n4047), .A(n4051), .ZN(n3795) );
  AOI21_X1 U4204 ( .B1(n3796), .B2(n3804), .A(n3795), .ZN(n3797) );
  OR2_X1 U4205 ( .A1(\x_mult_f[2][8] ), .A2(\x_mult_f[3][8] ), .ZN(n4266) );
  NAND2_X1 U4206 ( .A1(\x_mult_f[2][8] ), .A2(\x_mult_f[3][8] ), .ZN(n3951) );
  INV_X1 U4207 ( .A(n3951), .ZN(n4270) );
  AOI21_X1 U4208 ( .B1(n7938), .B2(n4266), .A(n4270), .ZN(n3801) );
  OR2_X1 U4209 ( .A1(\x_mult_f[2][9] ), .A2(\x_mult_f[3][9] ), .ZN(n4269) );
  NAND2_X1 U4210 ( .A1(\x_mult_f[2][9] ), .A2(\x_mult_f[3][9] ), .ZN(n4267) );
  NAND2_X1 U4211 ( .A1(n4269), .A2(n4267), .ZN(n3800) );
  XOR2_X1 U4212 ( .A(n3801), .B(n3800), .Z(n3802) );
  AOI22_X1 U4213 ( .A1(n8088), .A2(\adder_stage1[1][9] ), .B1(n4311), .B2(
        n3802), .ZN(n3803) );
  INV_X1 U4214 ( .A(n3803), .ZN(n10143) );
  AOI21_X1 U4215 ( .B1(n3902), .B2(n3805), .A(n3804), .ZN(n4049) );
  INV_X1 U4216 ( .A(n4048), .ZN(n3806) );
  NAND2_X1 U4217 ( .A1(n3806), .A2(n4047), .ZN(n3807) );
  XOR2_X1 U4218 ( .A(n4049), .B(n3807), .Z(n3808) );
  AOI22_X1 U4219 ( .A1(n8088), .A2(\adder_stage1[1][6] ), .B1(n4311), .B2(
        n3808), .ZN(n3809) );
  INV_X1 U4220 ( .A(n3809), .ZN(n10146) );
  INV_X1 U4221 ( .A(n3810), .ZN(n3811) );
  AOI21_X1 U4222 ( .B1(n3813), .B2(n3812), .A(n3811), .ZN(n3818) );
  INV_X1 U4223 ( .A(n3814), .ZN(n3816) );
  NAND2_X1 U4224 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  XOR2_X1 U4225 ( .A(n3818), .B(n3817), .Z(n3819) );
  AOI22_X1 U4226 ( .A1(n8057), .A2(\adder_stage2[3][5] ), .B1(n8251), .B2(
        n3819), .ZN(n3820) );
  INV_X1 U4227 ( .A(n3820), .ZN(n9848) );
  INV_X1 U4228 ( .A(n3892), .ZN(n3821) );
  NAND2_X1 U4229 ( .A1(n3821), .A2(n3891), .ZN(n3822) );
  XOR2_X1 U4230 ( .A(n7310), .B(n3822), .Z(n3823) );
  AOI22_X1 U4231 ( .A1(n7972), .A2(\adder_stage2[0][11] ), .B1(n4311), .B2(
        n3823), .ZN(n3824) );
  INV_X1 U4232 ( .A(n3824), .ZN(n9893) );
  INV_X1 U4233 ( .A(n3825), .ZN(n3864) );
  OAI21_X1 U4234 ( .B1(n3864), .B2(n3860), .A(n3861), .ZN(n3830) );
  INV_X1 U4235 ( .A(n3826), .ZN(n3828) );
  NAND2_X1 U4236 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  XNOR2_X1 U4237 ( .A(n3830), .B(n3829), .ZN(n3831) );
  AOI22_X1 U4238 ( .A1(n8273), .A2(\adder_stage3[1][3] ), .B1(n8272), .B2(
        n3831), .ZN(n3832) );
  INV_X1 U4239 ( .A(n3832), .ZN(n9745) );
  INV_X1 U4240 ( .A(n3833), .ZN(n3836) );
  INV_X1 U4241 ( .A(n3834), .ZN(n3835) );
  OAI21_X1 U4242 ( .B1(n3929), .B2(n3836), .A(n3835), .ZN(n3958) );
  INV_X1 U4243 ( .A(n3837), .ZN(n3956) );
  INV_X1 U4244 ( .A(n3955), .ZN(n3838) );
  AOI21_X1 U4245 ( .B1(n3958), .B2(n3956), .A(n3838), .ZN(n3843) );
  INV_X1 U4246 ( .A(n3839), .ZN(n3841) );
  NAND2_X1 U4247 ( .A1(n3841), .A2(n3840), .ZN(n3842) );
  XOR2_X1 U4248 ( .A(n3843), .B(n3842), .Z(n3844) );
  AOI22_X1 U4249 ( .A1(n8319), .A2(\adder_stage3[1][11] ), .B1(n8251), .B2(
        n3844), .ZN(n3845) );
  INV_X1 U4250 ( .A(n3845), .ZN(n9737) );
  INV_X1 U4251 ( .A(n3846), .ZN(n3848) );
  NAND2_X1 U4252 ( .A1(n3848), .A2(n3847), .ZN(n3850) );
  XOR2_X1 U4253 ( .A(n3850), .B(n3849), .Z(n3851) );
  AOI22_X1 U4254 ( .A1(n8273), .A2(\adder_stage3[1][1] ), .B1(n8272), .B2(
        n3851), .ZN(n3852) );
  INV_X1 U4255 ( .A(n3852), .ZN(n9747) );
  INV_X1 U4256 ( .A(n3853), .ZN(n3964) );
  AOI21_X1 U4257 ( .B1(n3964), .B2(n3855), .A(n3854), .ZN(n3969) );
  INV_X1 U4258 ( .A(n3968), .ZN(n3856) );
  NAND2_X1 U4259 ( .A1(n3856), .A2(n3967), .ZN(n3857) );
  XOR2_X1 U4260 ( .A(n3969), .B(n3857), .Z(n3858) );
  AOI22_X1 U4261 ( .A1(n7640), .A2(\adder_stage3[1][6] ), .B1(n8272), .B2(
        n3858), .ZN(n3859) );
  INV_X1 U4262 ( .A(n3859), .ZN(n9742) );
  INV_X1 U4263 ( .A(n3860), .ZN(n3862) );
  NAND2_X1 U4264 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  XOR2_X1 U4265 ( .A(n3864), .B(n3863), .Z(n3865) );
  AOI22_X1 U4266 ( .A1(n8273), .A2(\adder_stage3[1][2] ), .B1(n8272), .B2(
        n3865), .ZN(n3866) );
  INV_X1 U4267 ( .A(n3866), .ZN(n9746) );
  OAI21_X1 U4268 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n3888) );
  OR2_X1 U4269 ( .A1(\adder_stage2[2][14] ), .A2(\adder_stage2[3][14] ), .ZN(
        n3886) );
  NAND2_X1 U4270 ( .A1(\adder_stage2[2][14] ), .A2(\adder_stage2[3][14] ), 
        .ZN(n3885) );
  INV_X1 U4271 ( .A(n3885), .ZN(n3870) );
  AOI21_X1 U4272 ( .B1(n3888), .B2(n3886), .A(n3870), .ZN(n5584) );
  NOR2_X1 U4273 ( .A1(\adder_stage2[2][15] ), .A2(\adder_stage2[3][15] ), .ZN(
        n5583) );
  INV_X1 U4274 ( .A(n5583), .ZN(n3871) );
  NAND2_X1 U4275 ( .A1(\adder_stage2[2][15] ), .A2(\adder_stage2[3][15] ), 
        .ZN(n5582) );
  NAND2_X1 U4276 ( .A1(n3871), .A2(n5582), .ZN(n3872) );
  XOR2_X1 U4277 ( .A(n5584), .B(n3872), .Z(n3873) );
  AOI22_X1 U4278 ( .A1(n8309), .A2(\adder_stage3[1][15] ), .B1(n8251), .B2(
        n3873), .ZN(n3874) );
  INV_X1 U4279 ( .A(n3874), .ZN(n9733) );
  NOR2_X1 U4280 ( .A1(n3875), .A2(n3892), .ZN(n3876) );
  NAND2_X1 U4281 ( .A1(n3894), .A2(n3876), .ZN(n7309) );
  INV_X1 U4282 ( .A(n3877), .ZN(n3878) );
  AOI21_X1 U4283 ( .B1(n3880), .B2(n3879), .A(n3878), .ZN(n7313) );
  OAI21_X1 U4284 ( .B1(n7310), .B2(n7309), .A(n7313), .ZN(n3882) );
  OR2_X1 U4285 ( .A1(\adder_stage1[0][14] ), .A2(\adder_stage1[1][14] ), .ZN(
        n7308) );
  NAND2_X1 U4286 ( .A1(\adder_stage1[0][14] ), .A2(\adder_stage1[1][14] ), 
        .ZN(n7311) );
  NAND2_X1 U4287 ( .A1(n7308), .A2(n7311), .ZN(n3881) );
  XNOR2_X1 U4288 ( .A(n3882), .B(n3881), .ZN(n3883) );
  AOI22_X1 U4289 ( .A1(n7640), .A2(\adder_stage2[0][14] ), .B1(n4311), .B2(
        n3883), .ZN(n3884) );
  INV_X1 U4290 ( .A(n3884), .ZN(n9890) );
  NAND2_X1 U4291 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  XNOR2_X1 U4292 ( .A(n3888), .B(n3887), .ZN(n3889) );
  AOI22_X1 U4293 ( .A1(n7177), .A2(\adder_stage3[1][14] ), .B1(n8251), .B2(
        n3889), .ZN(n3890) );
  INV_X1 U4294 ( .A(n3890), .ZN(n9734) );
  OAI21_X1 U4295 ( .B1(n7310), .B2(n3892), .A(n3891), .ZN(n3896) );
  NAND2_X1 U4296 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  XNOR2_X1 U4297 ( .A(n3896), .B(n3895), .ZN(n3897) );
  AOI22_X1 U4298 ( .A1(n7622), .A2(\adder_stage2[0][12] ), .B1(n4311), .B2(
        n3897), .ZN(n3898) );
  INV_X1 U4299 ( .A(n3898), .ZN(n9892) );
  INV_X1 U4300 ( .A(n3899), .ZN(n3900) );
  AOI21_X1 U4301 ( .B1(n3902), .B2(n3901), .A(n3900), .ZN(n3907) );
  INV_X1 U4302 ( .A(n3903), .ZN(n3905) );
  NAND2_X1 U4303 ( .A1(n3905), .A2(n3904), .ZN(n3906) );
  XOR2_X1 U4304 ( .A(n3907), .B(n3906), .Z(n3908) );
  AOI22_X1 U4305 ( .A1(n8088), .A2(\adder_stage1[1][5] ), .B1(n4311), .B2(
        n3908), .ZN(n3909) );
  INV_X1 U4306 ( .A(n3909), .ZN(n10147) );
  INV_X1 U4307 ( .A(n3910), .ZN(n3962) );
  INV_X1 U4308 ( .A(n3961), .ZN(n3911) );
  AOI21_X1 U4309 ( .B1(n3964), .B2(n3962), .A(n3911), .ZN(n3916) );
  INV_X1 U4310 ( .A(n3912), .ZN(n3914) );
  NAND2_X1 U4311 ( .A1(n3914), .A2(n3913), .ZN(n3915) );
  XOR2_X1 U4312 ( .A(n3916), .B(n3915), .Z(n3917) );
  AOI22_X1 U4313 ( .A1(n7074), .A2(\adder_stage3[1][5] ), .B1(n8272), .B2(
        n3917), .ZN(n3918) );
  INV_X1 U4314 ( .A(n3918), .ZN(n9743) );
  INV_X1 U4315 ( .A(n3919), .ZN(n3948) );
  OAI21_X1 U4316 ( .B1(n3948), .B2(n3944), .A(n3945), .ZN(n3924) );
  INV_X1 U4317 ( .A(n3920), .ZN(n3922) );
  NAND2_X1 U4318 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  XNOR2_X1 U4319 ( .A(n3924), .B(n3923), .ZN(n3925) );
  AOI22_X1 U4320 ( .A1(n8088), .A2(\adder_stage1[1][3] ), .B1(n4311), .B2(
        n3925), .ZN(n3926) );
  INV_X1 U4321 ( .A(n3926), .ZN(n10149) );
  OAI21_X1 U4322 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3934) );
  INV_X1 U4323 ( .A(n3930), .ZN(n3932) );
  NAND2_X1 U4324 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  XNOR2_X1 U4325 ( .A(n3934), .B(n3933), .ZN(n3935) );
  AOI22_X1 U4326 ( .A1(n6854), .A2(\adder_stage3[1][12] ), .B1(n8251), .B2(
        n3935), .ZN(n3936) );
  INV_X1 U4327 ( .A(n3936), .ZN(n9736) );
  INV_X1 U4328 ( .A(n3937), .ZN(n3939) );
  NAND2_X1 U4329 ( .A1(n3939), .A2(n3938), .ZN(n3941) );
  XOR2_X1 U4330 ( .A(n3941), .B(n3940), .Z(n3942) );
  AOI22_X1 U4331 ( .A1(n7855), .A2(\adder_stage2[3][1] ), .B1(n8251), .B2(
        n3942), .ZN(n3943) );
  INV_X1 U4332 ( .A(n3943), .ZN(n9852) );
  INV_X1 U4333 ( .A(n3944), .ZN(n3946) );
  NAND2_X1 U4334 ( .A1(n3946), .A2(n3945), .ZN(n3947) );
  XOR2_X1 U4335 ( .A(n3948), .B(n3947), .Z(n3949) );
  AOI22_X1 U4336 ( .A1(n8088), .A2(\adder_stage1[1][2] ), .B1(n4311), .B2(
        n3949), .ZN(n3950) );
  INV_X1 U4337 ( .A(n3950), .ZN(n10150) );
  NAND2_X1 U4338 ( .A1(n4266), .A2(n3951), .ZN(n3952) );
  XNOR2_X1 U4339 ( .A(n3419), .B(n3952), .ZN(n3953) );
  AOI22_X1 U4340 ( .A1(n8088), .A2(\adder_stage1[1][8] ), .B1(n4311), .B2(
        n3953), .ZN(n3954) );
  INV_X1 U4341 ( .A(n3954), .ZN(n10144) );
  NAND2_X1 U4342 ( .A1(n3956), .A2(n3955), .ZN(n3957) );
  XNOR2_X1 U4343 ( .A(n3958), .B(n3957), .ZN(n3959) );
  AOI22_X1 U4344 ( .A1(n8273), .A2(\adder_stage3[1][10] ), .B1(n8272), .B2(
        n3959), .ZN(n3960) );
  INV_X1 U4345 ( .A(n3960), .ZN(n9738) );
  NAND2_X1 U4346 ( .A1(n3962), .A2(n3961), .ZN(n3963) );
  XNOR2_X1 U4347 ( .A(n3964), .B(n3963), .ZN(n3965) );
  AOI22_X1 U4348 ( .A1(n8398), .A2(\adder_stage3[1][4] ), .B1(n8272), .B2(
        n3965), .ZN(n3966) );
  INV_X1 U4349 ( .A(n3966), .ZN(n9744) );
  OAI21_X1 U4350 ( .B1(n3969), .B2(n3968), .A(n3967), .ZN(n3974) );
  INV_X1 U4351 ( .A(n3970), .ZN(n3972) );
  NAND2_X1 U4352 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  XNOR2_X1 U4353 ( .A(n3974), .B(n3973), .ZN(n3975) );
  AOI22_X1 U4354 ( .A1(n8401), .A2(\adder_stage3[1][7] ), .B1(n8272), .B2(
        n3975), .ZN(n3976) );
  INV_X1 U4355 ( .A(n3976), .ZN(n9741) );
  INV_X1 U4356 ( .A(n3983), .ZN(n3981) );
  INV_X1 U4357 ( .A(n3977), .ZN(n3978) );
  NAND3_X1 U4358 ( .A1(n3985), .A2(n3979), .A3(n3978), .ZN(n3980) );
  NOR2_X1 U4359 ( .A1(n8345), .A2(reset), .ZN(n8365) );
  INV_X1 U4360 ( .A(n8365), .ZN(n8373) );
  OAI211_X1 U4361 ( .C1(n3981), .C2(n8806), .A(n3980), .B(n8373), .ZN(n3386)
         );
  BUF_X1 U4362 ( .A(n3445), .Z(n5332) );
  BUF_X2 U4363 ( .A(n5332), .Z(n5247) );
  INV_X2 U4364 ( .A(n5247), .ZN(n6273) );
  AOI22_X1 U4365 ( .A1(n6273), .A2(\x_mult_f[21][4] ), .B1(n8272), .B2(
        \x_mult_f_int[21][4] ), .ZN(n3982) );
  INV_X1 U4366 ( .A(n3982), .ZN(n9193) );
  AOI22_X1 U4367 ( .A1(n3985), .A2(n3984), .B1(\ctrl_inst/state [0]), .B2(
        n3983), .ZN(n3987) );
  NAND2_X1 U4368 ( .A1(n3987), .A2(n3986), .ZN(n3388) );
  INV_X1 U4369 ( .A(n4037), .ZN(n4022) );
  OAI21_X1 U4370 ( .B1(n4022), .B2(n4018), .A(n4019), .ZN(n3992) );
  INV_X1 U4371 ( .A(n3988), .ZN(n3990) );
  NAND2_X1 U4372 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  XNOR2_X1 U4373 ( .A(n3992), .B(n3991), .ZN(n3993) );
  AOI22_X1 U4374 ( .A1(n8273), .A2(\adder_stage4[0][9] ), .B1(n7507), .B2(
        n3993), .ZN(n3994) );
  INV_X1 U4375 ( .A(n3994), .ZN(n9678) );
  AOI21_X1 U4376 ( .B1(n4006), .B2(n3996), .A(n3995), .ZN(n3997) );
  OAI21_X1 U4377 ( .B1(n4022), .B2(n3998), .A(n3997), .ZN(n4002) );
  NAND2_X1 U4378 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  XNOR2_X1 U4379 ( .A(n4002), .B(n4001), .ZN(n4003) );
  AOI22_X1 U4380 ( .A1(n8273), .A2(\adder_stage4[0][12] ), .B1(n7507), .B2(
        n4003), .ZN(n4004) );
  INV_X1 U4381 ( .A(n4004), .ZN(n9675) );
  INV_X1 U4382 ( .A(n4005), .ZN(n4008) );
  INV_X1 U4383 ( .A(n4006), .ZN(n4007) );
  OAI21_X1 U4384 ( .B1(n4022), .B2(n4008), .A(n4007), .ZN(n4028) );
  INV_X1 U4385 ( .A(n4009), .ZN(n4026) );
  INV_X1 U4386 ( .A(n4025), .ZN(n4010) );
  AOI21_X1 U4387 ( .B1(n4028), .B2(n4026), .A(n4010), .ZN(n4015) );
  INV_X1 U4388 ( .A(n4011), .ZN(n4013) );
  NAND2_X1 U4389 ( .A1(n4013), .A2(n4012), .ZN(n4014) );
  XOR2_X1 U4390 ( .A(n4015), .B(n4014), .Z(n4016) );
  AOI22_X1 U4391 ( .A1(n8273), .A2(\adder_stage4[0][11] ), .B1(n7507), .B2(
        n4016), .ZN(n4017) );
  INV_X1 U4392 ( .A(n4017), .ZN(n9676) );
  INV_X1 U4393 ( .A(n4018), .ZN(n4020) );
  NAND2_X1 U4394 ( .A1(n4020), .A2(n4019), .ZN(n4021) );
  XOR2_X1 U4395 ( .A(n4022), .B(n4021), .Z(n4023) );
  AOI22_X1 U4396 ( .A1(n8273), .A2(\adder_stage4[0][8] ), .B1(n7507), .B2(
        n4023), .ZN(n4024) );
  INV_X1 U4397 ( .A(n4024), .ZN(n9679) );
  NAND2_X1 U4398 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  XNOR2_X1 U4399 ( .A(n4028), .B(n4027), .ZN(n4029) );
  AOI22_X1 U4400 ( .A1(n8273), .A2(\adder_stage4[0][10] ), .B1(n7507), .B2(
        n4029), .ZN(n4030) );
  INV_X1 U4401 ( .A(n4030), .ZN(n9677) );
  NAND2_X1 U4402 ( .A1(n4032), .A2(n4031), .ZN(n4033) );
  XNOR2_X1 U4403 ( .A(n4034), .B(n4033), .ZN(n4035) );
  AOI22_X1 U4404 ( .A1(n8273), .A2(\adder_stage4[0][14] ), .B1(n8209), .B2(
        n4035), .ZN(n4036) );
  INV_X1 U4405 ( .A(n4036), .ZN(n9673) );
  NAND2_X1 U4406 ( .A1(n4038), .A2(n4037), .ZN(n4039) );
  AND2_X1 U4407 ( .A1(n4040), .A2(n4039), .ZN(n4044) );
  NAND2_X1 U4408 ( .A1(n4042), .A2(n4041), .ZN(n4043) );
  XOR2_X1 U4409 ( .A(n4044), .B(n4043), .Z(n4045) );
  AOI22_X1 U4410 ( .A1(n8273), .A2(\adder_stage4[0][13] ), .B1(n6272), .B2(
        n4045), .ZN(n4046) );
  INV_X1 U4411 ( .A(n4046), .ZN(n9674) );
  INV_X2 U4412 ( .A(n5247), .ZN(n7525) );
  OAI21_X1 U4413 ( .B1(n4049), .B2(n4048), .A(n4047), .ZN(n4054) );
  INV_X1 U4414 ( .A(n4050), .ZN(n4052) );
  NAND2_X1 U4415 ( .A1(n4052), .A2(n4051), .ZN(n4053) );
  XNOR2_X1 U4416 ( .A(n4054), .B(n4053), .ZN(n4055) );
  AOI22_X1 U4417 ( .A1(n7525), .A2(\adder_stage1[1][7] ), .B1(n4311), .B2(
        n4055), .ZN(n4056) );
  INV_X1 U4418 ( .A(n4056), .ZN(n10145) );
  INV_X1 U4419 ( .A(n4057), .ZN(n4086) );
  INV_X1 U4420 ( .A(n4058), .ZN(n4084) );
  INV_X1 U4421 ( .A(n4083), .ZN(n4059) );
  AOI21_X1 U4422 ( .B1(n4086), .B2(n4084), .A(n4059), .ZN(n4064) );
  INV_X1 U4423 ( .A(n4060), .ZN(n4062) );
  NAND2_X1 U4424 ( .A1(n4062), .A2(n4061), .ZN(n4063) );
  XOR2_X1 U4425 ( .A(n4064), .B(n4063), .Z(n4065) );
  AOI22_X1 U4426 ( .A1(n8118), .A2(\adder_stage4[0][5] ), .B1(n6036), .B2(
        n4065), .ZN(n4066) );
  INV_X1 U4427 ( .A(n4066), .ZN(n9682) );
  AOI21_X1 U4428 ( .B1(n4086), .B2(n4068), .A(n4067), .ZN(n4080) );
  OAI21_X1 U4429 ( .B1(n4080), .B2(n4076), .A(n4077), .ZN(n4073) );
  INV_X1 U4430 ( .A(n4069), .ZN(n4071) );
  NAND2_X1 U4431 ( .A1(n4071), .A2(n4070), .ZN(n4072) );
  XNOR2_X1 U4432 ( .A(n4073), .B(n4072), .ZN(n4074) );
  AOI22_X1 U4433 ( .A1(n7640), .A2(\adder_stage4[0][7] ), .B1(n8024), .B2(
        n4074), .ZN(n4075) );
  INV_X1 U4434 ( .A(n4075), .ZN(n9680) );
  INV_X1 U4435 ( .A(n4076), .ZN(n4078) );
  NAND2_X1 U4436 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  XOR2_X1 U4437 ( .A(n4080), .B(n4079), .Z(n4081) );
  AOI22_X1 U4438 ( .A1(n8309), .A2(\adder_stage4[0][6] ), .B1(n7507), .B2(
        n4081), .ZN(n4082) );
  INV_X1 U4439 ( .A(n4082), .ZN(n9681) );
  NAND2_X1 U4440 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  XNOR2_X1 U4441 ( .A(n4086), .B(n4085), .ZN(n4087) );
  AOI22_X1 U4442 ( .A1(n7698), .A2(\adder_stage4[0][4] ), .B1(n7507), .B2(
        n4087), .ZN(n4088) );
  INV_X1 U4443 ( .A(n4088), .ZN(n9683) );
  INV_X1 U4444 ( .A(n4089), .ZN(n4875) );
  OAI21_X1 U4445 ( .B1(n4875), .B2(n4871), .A(n4872), .ZN(n4094) );
  INV_X1 U4446 ( .A(n4090), .ZN(n4092) );
  NAND2_X1 U4447 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  XNOR2_X1 U4448 ( .A(n4094), .B(n4093), .ZN(n4095) );
  AOI22_X1 U4449 ( .A1(n7640), .A2(\adder_stage4[0][3] ), .B1(n8209), .B2(
        n4095), .ZN(n4096) );
  INV_X1 U4450 ( .A(n4096), .ZN(n9684) );
  BUF_X2 U4451 ( .A(n4314), .Z(n8258) );
  NOR2_X1 U4452 ( .A1(\adder_stage2[4][2] ), .A2(\adder_stage2[5][2] ), .ZN(
        n5480) );
  NOR2_X1 U4453 ( .A1(\adder_stage2[5][3] ), .A2(\adder_stage2[4][3] ), .ZN(
        n5482) );
  NOR2_X1 U4454 ( .A1(n5480), .A2(n5482), .ZN(n4099) );
  NOR2_X1 U4455 ( .A1(\adder_stage2[4][1] ), .A2(\adder_stage2[5][1] ), .ZN(
        n4358) );
  NAND2_X1 U4456 ( .A1(\adder_stage2[4][0] ), .A2(\adder_stage2[5][0] ), .ZN(
        n4361) );
  NAND2_X1 U4457 ( .A1(\adder_stage2[4][1] ), .A2(\adder_stage2[5][1] ), .ZN(
        n4359) );
  OAI21_X1 U4458 ( .B1(n4358), .B2(n4361), .A(n4359), .ZN(n4353) );
  NAND2_X1 U4459 ( .A1(\adder_stage2[4][2] ), .A2(\adder_stage2[5][2] ), .ZN(
        n5479) );
  NAND2_X1 U4460 ( .A1(\adder_stage2[4][3] ), .A2(\adder_stage2[5][3] ), .ZN(
        n5483) );
  OAI21_X1 U4461 ( .B1(n5482), .B2(n5479), .A(n5483), .ZN(n4098) );
  AOI21_X1 U4462 ( .B1(n4099), .B2(n4353), .A(n4098), .ZN(n4208) );
  NOR2_X1 U4463 ( .A1(\adder_stage2[4][4] ), .A2(\adder_stage2[5][4] ), .ZN(
        n4209) );
  NOR2_X1 U4464 ( .A1(\adder_stage2[4][5] ), .A2(\adder_stage2[5][5] ), .ZN(
        n4211) );
  NOR2_X1 U4465 ( .A1(n4209), .A2(n4211), .ZN(n4219) );
  NOR2_X1 U4466 ( .A1(\adder_stage2[4][6] ), .A2(\adder_stage2[5][6] ), .ZN(
        n4243) );
  NOR2_X1 U4467 ( .A1(\adder_stage2[4][7] ), .A2(\adder_stage2[5][7] ), .ZN(
        n4220) );
  NOR2_X1 U4468 ( .A1(n4243), .A2(n4220), .ZN(n4101) );
  NAND2_X1 U4469 ( .A1(n4219), .A2(n4101), .ZN(n4123) );
  NAND2_X1 U4470 ( .A1(\adder_stage2[4][4] ), .A2(\adder_stage2[5][4] ), .ZN(
        n5473) );
  NAND2_X1 U4471 ( .A1(\adder_stage2[4][5] ), .A2(\adder_stage2[5][5] ), .ZN(
        n4212) );
  OAI21_X1 U4472 ( .B1(n4211), .B2(n5473), .A(n4212), .ZN(n4218) );
  NAND2_X1 U4473 ( .A1(\adder_stage2[4][6] ), .A2(\adder_stage2[5][6] ), .ZN(
        n4244) );
  NAND2_X1 U4474 ( .A1(\adder_stage2[4][7] ), .A2(\adder_stage2[5][7] ), .ZN(
        n4221) );
  OAI21_X1 U4475 ( .B1(n4220), .B2(n4244), .A(n4221), .ZN(n4100) );
  AOI21_X1 U4476 ( .B1(n4101), .B2(n4218), .A(n4100), .ZN(n4126) );
  OAI21_X1 U4477 ( .B1(n4208), .B2(n4123), .A(n4126), .ZN(n4118) );
  INV_X1 U4478 ( .A(n4118), .ZN(n4263) );
  NOR2_X1 U4479 ( .A1(\adder_stage2[4][8] ), .A2(\adder_stage2[5][8] ), .ZN(
        n4259) );
  NOR2_X1 U4480 ( .A1(\adder_stage2[4][9] ), .A2(\adder_stage2[5][9] ), .ZN(
        n4159) );
  NOR2_X1 U4481 ( .A1(n4259), .A2(n4159), .ZN(n4111) );
  INV_X1 U4482 ( .A(n4111), .ZN(n4103) );
  NAND2_X1 U4483 ( .A1(\adder_stage2[4][8] ), .A2(\adder_stage2[5][8] ), .ZN(
        n4260) );
  NAND2_X1 U4484 ( .A1(\adder_stage2[4][9] ), .A2(\adder_stage2[5][9] ), .ZN(
        n4160) );
  OAI21_X1 U4485 ( .B1(n4159), .B2(n4260), .A(n4160), .ZN(n4115) );
  INV_X1 U4486 ( .A(n4115), .ZN(n4102) );
  OAI21_X1 U4487 ( .B1(n4263), .B2(n4103), .A(n4102), .ZN(n4175) );
  NOR2_X1 U4488 ( .A1(\adder_stage2[4][10] ), .A2(\adder_stage2[5][10] ), .ZN(
        n4110) );
  INV_X1 U4489 ( .A(n4110), .ZN(n4173) );
  NAND2_X1 U4490 ( .A1(\adder_stage2[4][10] ), .A2(\adder_stage2[5][10] ), 
        .ZN(n4172) );
  INV_X1 U4491 ( .A(n4172), .ZN(n4104) );
  AOI21_X1 U4492 ( .B1(n4175), .B2(n4173), .A(n4104), .ZN(n4107) );
  NOR2_X1 U4493 ( .A1(\adder_stage2[4][11] ), .A2(\adder_stage2[5][11] ), .ZN(
        n4113) );
  INV_X1 U4494 ( .A(n4113), .ZN(n4105) );
  NAND2_X1 U4495 ( .A1(\adder_stage2[4][11] ), .A2(\adder_stage2[5][11] ), 
        .ZN(n4112) );
  NAND2_X1 U4496 ( .A1(n4105), .A2(n4112), .ZN(n4106) );
  XOR2_X1 U4497 ( .A(n4107), .B(n4106), .Z(n4108) );
  AOI22_X1 U4498 ( .A1(n7669), .A2(\adder_stage3[2][11] ), .B1(n8258), .B2(
        n4108), .ZN(n4109) );
  INV_X1 U4499 ( .A(n4109), .ZN(n9718) );
  NOR2_X1 U4500 ( .A1(n4110), .A2(n4113), .ZN(n4116) );
  NAND2_X1 U4501 ( .A1(n4111), .A2(n4116), .ZN(n4146) );
  NOR2_X1 U4502 ( .A1(\adder_stage2[4][12] ), .A2(\adder_stage2[5][12] ), .ZN(
        n4130) );
  NOR2_X1 U4503 ( .A1(n4146), .A2(n4130), .ZN(n4128) );
  OAI21_X1 U4504 ( .B1(n4113), .B2(n4172), .A(n4112), .ZN(n4114) );
  AOI21_X1 U4505 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4145) );
  NAND2_X1 U4506 ( .A1(\adder_stage2[4][12] ), .A2(\adder_stage2[5][12] ), 
        .ZN(n4147) );
  OAI21_X1 U4507 ( .B1(n4145), .B2(n4130), .A(n4147), .ZN(n4117) );
  AOI21_X1 U4508 ( .B1(n4128), .B2(n4118), .A(n4117), .ZN(n4120) );
  OR2_X1 U4509 ( .A1(\adder_stage2[4][13] ), .A2(\adder_stage2[5][13] ), .ZN(
        n4134) );
  NAND2_X1 U4510 ( .A1(\adder_stage2[4][13] ), .A2(\adder_stage2[5][13] ), 
        .ZN(n4131) );
  NAND2_X1 U4511 ( .A1(n4134), .A2(n4131), .ZN(n4119) );
  XOR2_X1 U4512 ( .A(n4120), .B(n4119), .Z(n4121) );
  AOI22_X1 U4513 ( .A1(n8176), .A2(\adder_stage3[2][13] ), .B1(n8258), .B2(
        n4121), .ZN(n4122) );
  INV_X1 U4514 ( .A(n4122), .ZN(n9716) );
  INV_X1 U4515 ( .A(n4123), .ZN(n4124) );
  NAND2_X1 U4516 ( .A1(n4134), .A2(n4124), .ZN(n4127) );
  INV_X1 U4517 ( .A(n4134), .ZN(n4125) );
  OAI22_X1 U4518 ( .A1(n4208), .A2(n4127), .B1(n4126), .B2(n4125), .ZN(n4129)
         );
  NAND2_X1 U4519 ( .A1(n4129), .A2(n4128), .ZN(n4139) );
  INV_X1 U4520 ( .A(n4130), .ZN(n4148) );
  NAND2_X1 U4521 ( .A1(n4134), .A2(n4148), .ZN(n4136) );
  INV_X1 U4522 ( .A(n4147), .ZN(n4133) );
  INV_X1 U4523 ( .A(n4131), .ZN(n4132) );
  AOI21_X1 U4524 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4135) );
  OAI21_X1 U4525 ( .B1(n4145), .B2(n4136), .A(n4135), .ZN(n4137) );
  INV_X1 U4526 ( .A(n4137), .ZN(n4138) );
  NAND2_X1 U4527 ( .A1(n4139), .A2(n4138), .ZN(n4169) );
  OR2_X1 U4528 ( .A1(\adder_stage2[4][14] ), .A2(\adder_stage2[5][14] ), .ZN(
        n4167) );
  NAND2_X1 U4529 ( .A1(\adder_stage2[4][14] ), .A2(\adder_stage2[5][14] ), 
        .ZN(n4166) );
  INV_X1 U4530 ( .A(n4166), .ZN(n4140) );
  AOI21_X1 U4531 ( .B1(n4169), .B2(n4167), .A(n4140), .ZN(n4889) );
  NOR2_X1 U4532 ( .A1(\adder_stage2[4][15] ), .A2(\adder_stage2[5][15] ), .ZN(
        n4888) );
  INV_X1 U4533 ( .A(n4888), .ZN(n4141) );
  NAND2_X1 U4534 ( .A1(\adder_stage2[4][15] ), .A2(\adder_stage2[5][15] ), 
        .ZN(n4887) );
  NAND2_X1 U4535 ( .A1(n4141), .A2(n4887), .ZN(n4142) );
  XOR2_X1 U4536 ( .A(n4889), .B(n4142), .Z(n4143) );
  AOI22_X1 U4537 ( .A1(n8319), .A2(\adder_stage3[2][15] ), .B1(n8258), .B2(
        n4143), .ZN(n4144) );
  INV_X1 U4538 ( .A(n4144), .ZN(n9714) );
  OAI21_X1 U4539 ( .B1(n4263), .B2(n4146), .A(n4145), .ZN(n4150) );
  NAND2_X1 U4540 ( .A1(n4148), .A2(n4147), .ZN(n4149) );
  XNOR2_X1 U4541 ( .A(n4150), .B(n4149), .ZN(n4151) );
  AOI22_X1 U4542 ( .A1(n7959), .A2(\adder_stage3[2][12] ), .B1(n8258), .B2(
        n4151), .ZN(n4152) );
  INV_X1 U4543 ( .A(n4152), .ZN(n9717) );
  INV_X2 U4544 ( .A(n3408), .ZN(n7928) );
  BUF_X2 U4545 ( .A(n4314), .Z(n4257) );
  NOR2_X1 U4546 ( .A1(\x_mult_f[28][2] ), .A2(\x_mult_f[29][2] ), .ZN(n5609)
         );
  NOR2_X1 U4547 ( .A1(n5609), .A2(n5611), .ZN(n4154) );
  NOR2_X1 U4548 ( .A1(\x_mult_f[28][1] ), .A2(\x_mult_f[29][1] ), .ZN(n5593)
         );
  NAND2_X1 U4549 ( .A1(\x_mult_f[28][0] ), .A2(\x_mult_f[29][0] ), .ZN(n5631)
         );
  NAND2_X1 U4550 ( .A1(\x_mult_f[28][1] ), .A2(\x_mult_f[29][1] ), .ZN(n5594)
         );
  OAI21_X1 U4551 ( .B1(n5593), .B2(n5631), .A(n5594), .ZN(n5602) );
  NAND2_X1 U4552 ( .A1(\x_mult_f[28][2] ), .A2(\x_mult_f[29][2] ), .ZN(n5608)
         );
  NAND2_X1 U4553 ( .A1(\x_mult_f[28][3] ), .A2(\x_mult_f[29][3] ), .ZN(n5612)
         );
  OAI21_X1 U4554 ( .B1(n5611), .B2(n5608), .A(n5612), .ZN(n4153) );
  INV_X1 U4555 ( .A(n4184), .ZN(n7950) );
  NOR2_X1 U4556 ( .A1(\x_mult_f[28][4] ), .A2(\x_mult_f[29][4] ), .ZN(n7404)
         );
  NOR2_X1 U4557 ( .A1(\x_mult_f[28][5] ), .A2(\x_mult_f[29][5] ), .ZN(n7406)
         );
  NOR2_X1 U4558 ( .A1(n7404), .A2(n7406), .ZN(n4178) );
  NAND2_X1 U4559 ( .A1(\x_mult_f[28][4] ), .A2(\x_mult_f[29][4] ), .ZN(n7947)
         );
  NAND2_X1 U4560 ( .A1(\x_mult_f[28][5] ), .A2(\x_mult_f[29][5] ), .ZN(n7407)
         );
  OAI21_X1 U4561 ( .B1(n7406), .B2(n7947), .A(n7407), .ZN(n4180) );
  AOI21_X1 U4562 ( .B1(n7950), .B2(n4178), .A(n4180), .ZN(n4190) );
  NOR2_X1 U4563 ( .A1(\x_mult_f[28][6] ), .A2(\x_mult_f[29][6] ), .ZN(n4189)
         );
  INV_X1 U4564 ( .A(n4189), .ZN(n4155) );
  NAND2_X1 U4565 ( .A1(\x_mult_f[28][6] ), .A2(\x_mult_f[29][6] ), .ZN(n4188)
         );
  NAND2_X1 U4566 ( .A1(n4155), .A2(n4188), .ZN(n4156) );
  XOR2_X1 U4567 ( .A(n4190), .B(n4156), .Z(n4157) );
  AOI22_X1 U4568 ( .A1(n7928), .A2(\adder_stage1[14][6] ), .B1(n4257), .B2(
        n4157), .ZN(n4158) );
  INV_X1 U4569 ( .A(n4158), .ZN(n9929) );
  OAI21_X1 U4570 ( .B1(n4263), .B2(n4259), .A(n4260), .ZN(n4163) );
  INV_X1 U4571 ( .A(n4159), .ZN(n4161) );
  NAND2_X1 U4572 ( .A1(n4161), .A2(n4160), .ZN(n4162) );
  XNOR2_X1 U4573 ( .A(n4163), .B(n4162), .ZN(n4164) );
  AOI22_X1 U4574 ( .A1(n7928), .A2(\adder_stage3[2][9] ), .B1(n8258), .B2(
        n4164), .ZN(n4165) );
  INV_X1 U4575 ( .A(n4165), .ZN(n9720) );
  NAND2_X1 U4576 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  XNOR2_X1 U4577 ( .A(n4169), .B(n4168), .ZN(n4170) );
  AOI22_X1 U4578 ( .A1(n7074), .A2(\adder_stage3[2][14] ), .B1(n8258), .B2(
        n4170), .ZN(n4171) );
  INV_X1 U4579 ( .A(n4171), .ZN(n9715) );
  NAND2_X1 U4580 ( .A1(n4173), .A2(n4172), .ZN(n4174) );
  XNOR2_X1 U4581 ( .A(n4175), .B(n4174), .ZN(n4176) );
  AOI22_X1 U4582 ( .A1(n8434), .A2(\adder_stage3[2][10] ), .B1(n8258), .B2(
        n4176), .ZN(n4177) );
  INV_X1 U4583 ( .A(n4177), .ZN(n9719) );
  NOR2_X1 U4584 ( .A1(\x_mult_f[28][7] ), .A2(\x_mult_f[29][7] ), .ZN(n4191)
         );
  NOR2_X1 U4585 ( .A1(n4189), .A2(n4191), .ZN(n4181) );
  NAND2_X1 U4586 ( .A1(n4178), .A2(n4181), .ZN(n4183) );
  NAND2_X1 U4587 ( .A1(\x_mult_f[28][7] ), .A2(\x_mult_f[29][7] ), .ZN(n4192)
         );
  OAI21_X1 U4588 ( .B1(n4191), .B2(n4188), .A(n4192), .ZN(n4179) );
  AOI21_X1 U4589 ( .B1(n4181), .B2(n4180), .A(n4179), .ZN(n4182) );
  OAI21_X1 U4590 ( .B1(n4184), .B2(n4183), .A(n4182), .ZN(n4324) );
  OR2_X1 U4591 ( .A1(\x_mult_f[28][8] ), .A2(\x_mult_f[29][8] ), .ZN(n4326) );
  NAND2_X1 U4592 ( .A1(\x_mult_f[28][8] ), .A2(\x_mult_f[29][8] ), .ZN(n4315)
         );
  NAND2_X1 U4593 ( .A1(n4326), .A2(n4315), .ZN(n4185) );
  XNOR2_X1 U4594 ( .A(n4324), .B(n4185), .ZN(n4186) );
  AOI22_X1 U4595 ( .A1(n7928), .A2(\adder_stage1[14][8] ), .B1(n4257), .B2(
        n4186), .ZN(n4187) );
  INV_X1 U4596 ( .A(n4187), .ZN(n9927) );
  OAI21_X1 U4597 ( .B1(n4190), .B2(n4189), .A(n4188), .ZN(n4195) );
  INV_X1 U4598 ( .A(n4191), .ZN(n4193) );
  NAND2_X1 U4599 ( .A1(n4193), .A2(n4192), .ZN(n4194) );
  XNOR2_X1 U4600 ( .A(n4195), .B(n4194), .ZN(n4196) );
  AOI22_X1 U4601 ( .A1(n7928), .A2(\adder_stage1[14][7] ), .B1(n4257), .B2(
        n4196), .ZN(n4197) );
  INV_X1 U4602 ( .A(n4197), .ZN(n9928) );
  INV_X2 U4603 ( .A(n3409), .ZN(n8176) );
  AOI22_X1 U4604 ( .A1(n8176), .A2(\x_mult_f[24][0] ), .B1(n4257), .B2(
        \x_mult_f_int[24][0] ), .ZN(n4198) );
  INV_X1 U4605 ( .A(n4198), .ZN(n9375) );
  AOI22_X1 U4606 ( .A1(n8176), .A2(\x_mult_f[24][1] ), .B1(n4257), .B2(
        \x_mult_f_int[24][1] ), .ZN(n4199) );
  INV_X1 U4607 ( .A(n4199), .ZN(n9374) );
  AOI22_X1 U4608 ( .A1(n8176), .A2(\x_mult_f[24][2] ), .B1(n4257), .B2(
        \x_mult_f_int[24][2] ), .ZN(n4200) );
  INV_X1 U4609 ( .A(n4200), .ZN(n9229) );
  AOI22_X1 U4610 ( .A1(n6854), .A2(\x_mult_f[26][4] ), .B1(n4257), .B2(
        \x_mult_f_int[26][4] ), .ZN(n4201) );
  INV_X1 U4611 ( .A(n4201), .ZN(n9255) );
  NOR2_X1 U4612 ( .A1(\x_mult_f[26][2] ), .A2(\x_mult_f[27][2] ), .ZN(n4251)
         );
  NOR2_X1 U4613 ( .A1(\x_mult_f[26][3] ), .A2(\x_mult_f[27][3] ), .ZN(n4236)
         );
  NOR2_X1 U4614 ( .A1(n4251), .A2(n4236), .ZN(n4204) );
  NOR2_X1 U4615 ( .A1(\x_mult_f[26][1] ), .A2(\x_mult_f[27][1] ), .ZN(n6300)
         );
  NAND2_X1 U4616 ( .A1(\x_mult_f[26][0] ), .A2(\x_mult_f[27][0] ), .ZN(n6303)
         );
  NAND2_X1 U4617 ( .A1(\x_mult_f[26][1] ), .A2(\x_mult_f[27][1] ), .ZN(n6301)
         );
  OAI21_X1 U4618 ( .B1(n6300), .B2(n6303), .A(n6301), .ZN(n4235) );
  NAND2_X1 U4619 ( .A1(\x_mult_f[26][2] ), .A2(\x_mult_f[27][2] ), .ZN(n4252)
         );
  NAND2_X1 U4620 ( .A1(\x_mult_f[26][3] ), .A2(\x_mult_f[27][3] ), .ZN(n4237)
         );
  OAI21_X1 U4621 ( .B1(n4236), .B2(n4252), .A(n4237), .ZN(n4203) );
  AOI21_X1 U4622 ( .B1(n4204), .B2(n4235), .A(n4203), .ZN(n4851) );
  INV_X1 U4623 ( .A(n4851), .ZN(n7379) );
  NOR2_X1 U4624 ( .A1(\x_mult_f[26][4] ), .A2(\x_mult_f[27][4] ), .ZN(n4843)
         );
  INV_X1 U4625 ( .A(n4843), .ZN(n4228) );
  NAND2_X1 U4626 ( .A1(\x_mult_f[26][4] ), .A2(\x_mult_f[27][4] ), .ZN(n4845)
         );
  NAND2_X1 U4627 ( .A1(n4228), .A2(n4845), .ZN(n4205) );
  XNOR2_X1 U4628 ( .A(n7379), .B(n4205), .ZN(n4206) );
  AOI22_X1 U4629 ( .A1(n8057), .A2(\adder_stage1[13][4] ), .B1(n4257), .B2(
        n4206), .ZN(n4207) );
  INV_X1 U4630 ( .A(n4207), .ZN(n9948) );
  INV_X1 U4631 ( .A(n4208), .ZN(n5476) );
  INV_X1 U4632 ( .A(n4209), .ZN(n5474) );
  INV_X1 U4633 ( .A(n5473), .ZN(n4210) );
  AOI21_X1 U4634 ( .B1(n5476), .B2(n5474), .A(n4210), .ZN(n4215) );
  INV_X1 U4635 ( .A(n4211), .ZN(n4213) );
  NAND2_X1 U4636 ( .A1(n4213), .A2(n4212), .ZN(n4214) );
  XOR2_X1 U4637 ( .A(n4215), .B(n4214), .Z(n4216) );
  AOI22_X1 U4638 ( .A1(n8296), .A2(\adder_stage3[2][5] ), .B1(n8258), .B2(
        n4216), .ZN(n4217) );
  INV_X1 U4639 ( .A(n4217), .ZN(n9724) );
  AOI21_X1 U4640 ( .B1(n5476), .B2(n4219), .A(n4218), .ZN(n4247) );
  OAI21_X1 U4641 ( .B1(n4247), .B2(n4243), .A(n4244), .ZN(n4224) );
  INV_X1 U4642 ( .A(n4220), .ZN(n4222) );
  NAND2_X1 U4643 ( .A1(n4222), .A2(n4221), .ZN(n4223) );
  XNOR2_X1 U4644 ( .A(n4224), .B(n4223), .ZN(n4225) );
  AOI22_X1 U4645 ( .A1(n8325), .A2(\adder_stage3[2][7] ), .B1(n8258), .B2(
        n4225), .ZN(n4226) );
  INV_X1 U4646 ( .A(n4226), .ZN(n9722) );
  INV_X1 U4647 ( .A(n4845), .ZN(n4227) );
  AOI21_X1 U4648 ( .B1(n7379), .B2(n4228), .A(n4227), .ZN(n4231) );
  NOR2_X1 U4649 ( .A1(\x_mult_f[26][5] ), .A2(\x_mult_f[27][5] ), .ZN(n4846)
         );
  INV_X1 U4650 ( .A(n4846), .ZN(n4229) );
  NAND2_X1 U4651 ( .A1(\x_mult_f[26][5] ), .A2(\x_mult_f[27][5] ), .ZN(n4844)
         );
  NAND2_X1 U4652 ( .A1(n4229), .A2(n4844), .ZN(n4230) );
  XOR2_X1 U4653 ( .A(n4231), .B(n4230), .Z(n4232) );
  AOI22_X1 U4654 ( .A1(n7855), .A2(\adder_stage1[13][5] ), .B1(n4257), .B2(
        n4232), .ZN(n4233) );
  INV_X1 U4655 ( .A(n4233), .ZN(n9947) );
  AOI22_X1 U4656 ( .A1(n8330), .A2(\x_mult_f[24][3] ), .B1(n4257), .B2(
        \x_mult_f_int[24][3] ), .ZN(n4234) );
  INV_X1 U4657 ( .A(n4234), .ZN(n9228) );
  INV_X1 U4658 ( .A(n4235), .ZN(n4255) );
  OAI21_X1 U4659 ( .B1(n4255), .B2(n4251), .A(n4252), .ZN(n4240) );
  INV_X1 U4660 ( .A(n4236), .ZN(n4238) );
  NAND2_X1 U4661 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  XNOR2_X1 U4662 ( .A(n4240), .B(n4239), .ZN(n4241) );
  AOI22_X1 U4663 ( .A1(n8057), .A2(\adder_stage1[13][3] ), .B1(n4257), .B2(
        n4241), .ZN(n4242) );
  INV_X1 U4664 ( .A(n4242), .ZN(n9949) );
  INV_X1 U4665 ( .A(n4243), .ZN(n4245) );
  NAND2_X1 U4666 ( .A1(n4245), .A2(n4244), .ZN(n4246) );
  XOR2_X1 U4667 ( .A(n4247), .B(n4246), .Z(n4248) );
  AOI22_X1 U4668 ( .A1(n8328), .A2(\adder_stage3[2][6] ), .B1(n8258), .B2(
        n4248), .ZN(n4249) );
  INV_X1 U4669 ( .A(n4249), .ZN(n9723) );
  AOI22_X1 U4670 ( .A1(n7640), .A2(\x_mult_f[24][4] ), .B1(n4257), .B2(
        \x_mult_f_int[24][4] ), .ZN(n4250) );
  INV_X1 U4671 ( .A(n4250), .ZN(n9227) );
  INV_X1 U4672 ( .A(n4251), .ZN(n4253) );
  NAND2_X1 U4673 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  XOR2_X1 U4674 ( .A(n4255), .B(n4254), .Z(n4256) );
  AOI22_X1 U4675 ( .A1(n7972), .A2(\adder_stage1[13][2] ), .B1(n4257), .B2(
        n4256), .ZN(n4258) );
  INV_X1 U4676 ( .A(n4258), .ZN(n9950) );
  INV_X1 U4677 ( .A(n4259), .ZN(n4261) );
  NAND2_X1 U4678 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  XOR2_X1 U4679 ( .A(n4263), .B(n4262), .Z(n4264) );
  AOI22_X1 U4680 ( .A1(n8434), .A2(\adder_stage3[2][8] ), .B1(n8258), .B2(
        n4264), .ZN(n4265) );
  INV_X1 U4681 ( .A(n4265), .ZN(n9721) );
  BUF_X2 U4682 ( .A(n4444), .Z(n8054) );
  AND2_X1 U4683 ( .A1(n4266), .A2(n4269), .ZN(n5107) );
  NAND2_X1 U4684 ( .A1(n7938), .A2(n5107), .ZN(n4271) );
  INV_X1 U4685 ( .A(n4267), .ZN(n4268) );
  AOI21_X1 U4686 ( .B1(n4270), .B2(n4269), .A(n4268), .ZN(n7936) );
  NAND2_X1 U4687 ( .A1(n4271), .A2(n7936), .ZN(n4273) );
  OR2_X1 U4688 ( .A1(\x_mult_f[2][10] ), .A2(\x_mult_f[3][10] ), .ZN(n5108) );
  NAND2_X1 U4689 ( .A1(\x_mult_f[2][10] ), .A2(\x_mult_f[3][10] ), .ZN(n7934)
         );
  NAND2_X1 U4690 ( .A1(n5108), .A2(n7934), .ZN(n4272) );
  XNOR2_X1 U4691 ( .A(n4273), .B(n4272), .ZN(n4274) );
  AOI22_X1 U4692 ( .A1(n8088), .A2(\adder_stage1[1][10] ), .B1(n8054), .B2(
        n4274), .ZN(n4275) );
  INV_X1 U4693 ( .A(n4275), .ZN(n10142) );
  AOI22_X1 U4694 ( .A1(n6273), .A2(\x_mult_f[21][3] ), .B1(n8258), .B2(
        \x_mult_f_int[21][3] ), .ZN(n4276) );
  INV_X1 U4695 ( .A(n4276), .ZN(n9194) );
  INV_X2 U4696 ( .A(n4771), .ZN(n8057) );
  AOI22_X1 U4697 ( .A1(n8057), .A2(\x_mult_f[3][4] ), .B1(n8054), .B2(
        \x_mult_f_int[3][4] ), .ZN(n4277) );
  INV_X1 U4698 ( .A(n4277), .ZN(n8966) );
  AOI22_X1 U4699 ( .A1(n8057), .A2(\x_mult_f[3][1] ), .B1(n8054), .B2(
        \x_mult_f_int[3][1] ), .ZN(n4278) );
  INV_X1 U4700 ( .A(n4278), .ZN(n9332) );
  AOI22_X1 U4701 ( .A1(n8057), .A2(\x_mult_f[3][0] ), .B1(n8054), .B2(
        \x_mult_f_int[3][0] ), .ZN(n4279) );
  INV_X1 U4702 ( .A(n4279), .ZN(n9333) );
  AOI22_X1 U4703 ( .A1(n8057), .A2(\x_mult_f[3][2] ), .B1(n8054), .B2(
        \x_mult_f_int[3][2] ), .ZN(n4280) );
  INV_X1 U4704 ( .A(n4280), .ZN(n8968) );
  AOI22_X1 U4705 ( .A1(n8057), .A2(\x_mult_f[3][5] ), .B1(n8054), .B2(
        \x_mult_f_int[3][5] ), .ZN(n4281) );
  INV_X1 U4706 ( .A(n4281), .ZN(n8965) );
  AOI22_X1 U4707 ( .A1(n8057), .A2(\x_mult_f[3][3] ), .B1(n8054), .B2(
        \x_mult_f_int[3][3] ), .ZN(n4282) );
  INV_X1 U4708 ( .A(n4282), .ZN(n8967) );
  BUF_X2 U4709 ( .A(n6238), .Z(n8281) );
  AOI22_X1 U4710 ( .A1(n7952), .A2(\x_mult_f[30][1] ), .B1(n8281), .B2(
        \x_mult_f_int[30][1] ), .ZN(n4283) );
  INV_X1 U4711 ( .A(n4283), .ZN(n9386) );
  AOI22_X1 U4712 ( .A1(n7952), .A2(\x_mult_f[30][3] ), .B1(n8281), .B2(
        \x_mult_f_int[30][3] ), .ZN(n4284) );
  INV_X1 U4713 ( .A(n4284), .ZN(n9312) );
  AOI22_X1 U4714 ( .A1(n7952), .A2(\x_mult_f[30][2] ), .B1(n8281), .B2(
        \x_mult_f_int[30][2] ), .ZN(n4285) );
  INV_X1 U4715 ( .A(n4285), .ZN(n9313) );
  AOI22_X1 U4716 ( .A1(n7952), .A2(\x_mult_f[30][4] ), .B1(n8281), .B2(
        \x_mult_f_int[30][4] ), .ZN(n4286) );
  INV_X1 U4717 ( .A(n4286), .ZN(n9311) );
  AOI22_X1 U4718 ( .A1(n7952), .A2(\x_mult_f[30][5] ), .B1(n8281), .B2(
        \x_mult_f_int[30][5] ), .ZN(n4287) );
  INV_X1 U4719 ( .A(n4287), .ZN(n9310) );
  NOR2_X1 U4720 ( .A1(\adder_stage3[2][1] ), .A2(\adder_stage3[3][1] ), .ZN(
        n8275) );
  NAND2_X1 U4721 ( .A1(\adder_stage3[2][0] ), .A2(\adder_stage3[3][0] ), .ZN(
        n8278) );
  NAND2_X1 U4722 ( .A1(\adder_stage3[2][1] ), .A2(\adder_stage3[3][1] ), .ZN(
        n8276) );
  OAI21_X1 U4723 ( .B1(n8275), .B2(n8278), .A(n8276), .ZN(n4543) );
  INV_X1 U4724 ( .A(n4543), .ZN(n4295) );
  NOR2_X1 U4725 ( .A1(\adder_stage3[2][2] ), .A2(\adder_stage3[3][2] ), .ZN(
        n4538) );
  NAND2_X1 U4726 ( .A1(\adder_stage3[2][2] ), .A2(\adder_stage3[3][2] ), .ZN(
        n4540) );
  OAI21_X1 U4727 ( .B1(n4295), .B2(n4538), .A(n4540), .ZN(n4290) );
  NOR2_X1 U4728 ( .A1(\adder_stage3[2][3] ), .A2(\adder_stage3[3][3] ), .ZN(
        n4541) );
  INV_X1 U4729 ( .A(n4541), .ZN(n4288) );
  NAND2_X1 U4730 ( .A1(\adder_stage3[2][3] ), .A2(\adder_stage3[3][3] ), .ZN(
        n4539) );
  NAND2_X1 U4731 ( .A1(n4288), .A2(n4539), .ZN(n4289) );
  XNOR2_X1 U4732 ( .A(n4290), .B(n4289), .ZN(n4291) );
  AOI22_X1 U4733 ( .A1(n8057), .A2(\adder_stage4[1][3] ), .B1(n8281), .B2(
        n4291), .ZN(n4292) );
  INV_X1 U4734 ( .A(n4292), .ZN(n9663) );
  INV_X1 U4735 ( .A(n4538), .ZN(n4293) );
  NAND2_X1 U4736 ( .A1(n4293), .A2(n4540), .ZN(n4294) );
  XOR2_X1 U4737 ( .A(n4295), .B(n4294), .Z(n4296) );
  AOI22_X1 U4738 ( .A1(n6273), .A2(\adder_stage4[1][2] ), .B1(n8281), .B2(
        n4296), .ZN(n4297) );
  INV_X1 U4739 ( .A(n4297), .ZN(n9664) );
  AOI22_X1 U4740 ( .A1(n8168), .A2(\x_mult_f[28][5] ), .B1(n8281), .B2(
        \x_mult_f_int[28][5] ), .ZN(n4298) );
  INV_X1 U4741 ( .A(n4298), .ZN(n9282) );
  AOI22_X1 U4742 ( .A1(n6273), .A2(\x_mult_f[21][2] ), .B1(n8281), .B2(
        \x_mult_f_int[21][2] ), .ZN(n4299) );
  INV_X1 U4743 ( .A(n4299), .ZN(n9195) );
  AOI22_X1 U4744 ( .A1(n7614), .A2(\x_mult_f[21][0] ), .B1(n8281), .B2(
        \x_mult_f_int[21][0] ), .ZN(n4300) );
  INV_X1 U4745 ( .A(n4300), .ZN(n9369) );
  AOI22_X1 U4746 ( .A1(n7614), .A2(\x_mult_f[21][1] ), .B1(n8281), .B2(
        \x_mult_f_int[21][1] ), .ZN(n4301) );
  INV_X1 U4747 ( .A(n4301), .ZN(n9368) );
  OR2_X1 U4748 ( .A1(\x_mult_f[2][0] ), .A2(\x_mult_f[3][0] ), .ZN(n4302) );
  AND2_X1 U4749 ( .A1(n4302), .A2(n4308), .ZN(n4303) );
  AOI22_X1 U4750 ( .A1(n8057), .A2(\adder_stage1[1][0] ), .B1(n4311), .B2(
        n4303), .ZN(n4304) );
  INV_X1 U4751 ( .A(n4304), .ZN(n10152) );
  INV_X1 U4752 ( .A(n4305), .ZN(n4307) );
  NAND2_X1 U4753 ( .A1(n4307), .A2(n4306), .ZN(n4309) );
  XOR2_X1 U4754 ( .A(n4309), .B(n4308), .Z(n4310) );
  AOI22_X1 U4755 ( .A1(n7640), .A2(\adder_stage1[1][1] ), .B1(n4311), .B2(
        n4310), .ZN(n4312) );
  INV_X1 U4756 ( .A(n4312), .ZN(n10151) );
  AOI22_X1 U4757 ( .A1(n6877), .A2(\x_mult_f[26][5] ), .B1(n8281), .B2(
        \x_mult_f_int[26][5] ), .ZN(n4313) );
  INV_X1 U4758 ( .A(n4313), .ZN(n9254) );
  BUF_X2 U4759 ( .A(n4314), .Z(n7927) );
  OR2_X1 U4760 ( .A1(\x_mult_f[28][9] ), .A2(\x_mult_f[29][9] ), .ZN(n4328) );
  AND2_X1 U4761 ( .A1(n4326), .A2(n4328), .ZN(n4333) );
  OR2_X1 U4762 ( .A1(\x_mult_f[28][10] ), .A2(\x_mult_f[29][10] ), .ZN(n4338)
         );
  AND2_X1 U4763 ( .A1(n4333), .A2(n4338), .ZN(n4319) );
  INV_X1 U4764 ( .A(n4315), .ZN(n4325) );
  NAND2_X1 U4765 ( .A1(\x_mult_f[28][9] ), .A2(\x_mult_f[29][9] ), .ZN(n4327)
         );
  INV_X1 U4766 ( .A(n4327), .ZN(n4316) );
  AOI21_X1 U4767 ( .B1(n4325), .B2(n4328), .A(n4316), .ZN(n4335) );
  INV_X1 U4768 ( .A(n4338), .ZN(n4317) );
  NAND2_X1 U4769 ( .A1(\x_mult_f[28][10] ), .A2(\x_mult_f[29][10] ), .ZN(n4337) );
  OAI21_X1 U4770 ( .B1(n4335), .B2(n4317), .A(n4337), .ZN(n4318) );
  AOI21_X1 U4771 ( .B1(n4319), .B2(n4324), .A(n4318), .ZN(n6277) );
  NOR2_X1 U4772 ( .A1(\x_mult_f[28][11] ), .A2(\x_mult_f[29][11] ), .ZN(n6276)
         );
  INV_X1 U4773 ( .A(n6276), .ZN(n4320) );
  NAND2_X1 U4774 ( .A1(\x_mult_f[28][11] ), .A2(\x_mult_f[29][11] ), .ZN(n6275) );
  NAND2_X1 U4775 ( .A1(n4320), .A2(n6275), .ZN(n4321) );
  XOR2_X1 U4776 ( .A(n6277), .B(n4321), .Z(n4322) );
  AOI22_X1 U4777 ( .A1(n7928), .A2(\adder_stage1[14][11] ), .B1(n7927), .B2(
        n4322), .ZN(n4323) );
  INV_X1 U4778 ( .A(n4323), .ZN(n9924) );
  AOI21_X1 U4779 ( .B1(n4334), .B2(n4326), .A(n4325), .ZN(n4330) );
  NAND2_X1 U4780 ( .A1(n4328), .A2(n4327), .ZN(n4329) );
  XOR2_X1 U4781 ( .A(n4330), .B(n4329), .Z(n4331) );
  AOI22_X1 U4782 ( .A1(n7928), .A2(\adder_stage1[14][9] ), .B1(n7927), .B2(
        n4331), .ZN(n4332) );
  INV_X1 U4783 ( .A(n4332), .ZN(n9926) );
  NAND2_X1 U4784 ( .A1(n4334), .A2(n4333), .ZN(n4336) );
  NAND2_X1 U4785 ( .A1(n4336), .A2(n4335), .ZN(n4340) );
  NAND2_X1 U4786 ( .A1(n4338), .A2(n4337), .ZN(n4339) );
  XNOR2_X1 U4787 ( .A(n4340), .B(n4339), .ZN(n4341) );
  AOI22_X1 U4788 ( .A1(n7928), .A2(\adder_stage1[14][10] ), .B1(n7927), .B2(
        n4341), .ZN(n4342) );
  INV_X1 U4789 ( .A(n4342), .ZN(n9925) );
  NAND2_X1 U4790 ( .A1(n3482), .A2(n4344), .ZN(n4345) );
  XOR2_X1 U4791 ( .A(n4346), .B(n4345), .Z(n4347) );
  AOI22_X1 U4792 ( .A1(n4347), .A2(n8334), .B1(n7622), .B2(
        \adder_stage1[6][13] ), .ZN(n4348) );
  INV_X1 U4793 ( .A(n4348), .ZN(n10057) );
  BUF_X1 U4794 ( .A(n5449), .Z(n4894) );
  BUF_X2 U4795 ( .A(n4894), .Z(n8332) );
  AOI22_X1 U4796 ( .A1(\x_mult_f_int[24][6] ), .A2(n8332), .B1(n8428), .B2(
        \x_mult_f[24][6] ), .ZN(n4349) );
  INV_X1 U4797 ( .A(n4349), .ZN(n9225) );
  OR2_X1 U4798 ( .A1(\adder_stage2[4][0] ), .A2(\adder_stage2[5][0] ), .ZN(
        n4350) );
  AND2_X1 U4799 ( .A1(n4350), .A2(n4361), .ZN(n4351) );
  AOI22_X1 U4800 ( .A1(n7959), .A2(\adder_stage3[2][0] ), .B1(n7927), .B2(
        n4351), .ZN(n4352) );
  INV_X1 U4801 ( .A(n4352), .ZN(n9729) );
  INV_X1 U4802 ( .A(n4353), .ZN(n5481) );
  INV_X1 U4803 ( .A(n5480), .ZN(n4354) );
  NAND2_X1 U4804 ( .A1(n4354), .A2(n5479), .ZN(n4355) );
  XOR2_X1 U4805 ( .A(n5481), .B(n4355), .Z(n4356) );
  AOI22_X1 U4806 ( .A1(n8057), .A2(\adder_stage3[2][2] ), .B1(n7927), .B2(
        n4356), .ZN(n4357) );
  INV_X1 U4807 ( .A(n4357), .ZN(n9727) );
  INV_X1 U4808 ( .A(n4358), .ZN(n4360) );
  NAND2_X1 U4809 ( .A1(n4360), .A2(n4359), .ZN(n4362) );
  XOR2_X1 U4810 ( .A(n4362), .B(n4361), .Z(n4363) );
  AOI22_X1 U4811 ( .A1(n7074), .A2(\adder_stage3[2][1] ), .B1(n7927), .B2(
        n4363), .ZN(n4364) );
  INV_X1 U4812 ( .A(n4364), .ZN(n9728) );
  BUF_X2 U4813 ( .A(n6238), .Z(n8153) );
  AOI22_X1 U4814 ( .A1(n8057), .A2(\x_mult_f[15][2] ), .B1(n8153), .B2(
        \x_mult_f_int[15][2] ), .ZN(n4365) );
  INV_X1 U4815 ( .A(n4365), .ZN(n9122) );
  AOI22_X1 U4816 ( .A1(n7669), .A2(\x_mult_f[15][3] ), .B1(n8153), .B2(
        \x_mult_f_int[15][3] ), .ZN(n4366) );
  INV_X1 U4817 ( .A(n4366), .ZN(n9121) );
  NOR2_X1 U4818 ( .A1(\x_mult_f[14][2] ), .A2(\x_mult_f[15][2] ), .ZN(n5827)
         );
  NOR2_X1 U4819 ( .A1(\x_mult_f[14][3] ), .A2(\x_mult_f[15][3] ), .ZN(n5820)
         );
  NOR2_X1 U4820 ( .A1(n5827), .A2(n5820), .ZN(n4368) );
  NOR2_X1 U4821 ( .A1(\x_mult_f[14][1] ), .A2(\x_mult_f[15][1] ), .ZN(n5840)
         );
  NAND2_X1 U4822 ( .A1(\x_mult_f[14][0] ), .A2(\x_mult_f[15][0] ), .ZN(n5846)
         );
  NAND2_X1 U4823 ( .A1(\x_mult_f[14][1] ), .A2(\x_mult_f[15][1] ), .ZN(n5841)
         );
  OAI21_X1 U4824 ( .B1(n5840), .B2(n5846), .A(n5841), .ZN(n5819) );
  NAND2_X1 U4825 ( .A1(\x_mult_f[14][2] ), .A2(\x_mult_f[15][2] ), .ZN(n5828)
         );
  NAND2_X1 U4826 ( .A1(\x_mult_f[14][3] ), .A2(\x_mult_f[15][3] ), .ZN(n5821)
         );
  OAI21_X1 U4827 ( .B1(n5820), .B2(n5828), .A(n5821), .ZN(n4367) );
  AOI21_X1 U4828 ( .B1(n4368), .B2(n5819), .A(n4367), .ZN(n4396) );
  NOR2_X1 U4829 ( .A1(\x_mult_f[14][4] ), .A2(\x_mult_f[15][4] ), .ZN(n5804)
         );
  NOR2_X1 U4830 ( .A1(\x_mult_f[14][5] ), .A2(\x_mult_f[15][5] ), .ZN(n5806)
         );
  NOR2_X1 U4831 ( .A1(n5804), .A2(n5806), .ZN(n4398) );
  NOR2_X1 U4832 ( .A1(\x_mult_f[14][6] ), .A2(\x_mult_f[15][6] ), .ZN(n5797)
         );
  NOR2_X1 U4833 ( .A1(\x_mult_f[14][7] ), .A2(\x_mult_f[15][7] ), .ZN(n4399)
         );
  NOR2_X1 U4834 ( .A1(n5797), .A2(n4399), .ZN(n4370) );
  NAND2_X1 U4835 ( .A1(n4398), .A2(n4370), .ZN(n4372) );
  NAND2_X1 U4836 ( .A1(\x_mult_f[15][4] ), .A2(\x_mult_f[14][4] ), .ZN(n5813)
         );
  NAND2_X1 U4837 ( .A1(\x_mult_f[14][5] ), .A2(\x_mult_f[15][5] ), .ZN(n5807)
         );
  OAI21_X1 U4838 ( .B1(n5806), .B2(n5813), .A(n5807), .ZN(n4397) );
  NAND2_X1 U4839 ( .A1(\x_mult_f[14][6] ), .A2(\x_mult_f[15][6] ), .ZN(n5798)
         );
  NAND2_X1 U4840 ( .A1(\x_mult_f[14][7] ), .A2(\x_mult_f[15][7] ), .ZN(n4400)
         );
  OAI21_X1 U4841 ( .B1(n4399), .B2(n5798), .A(n4400), .ZN(n4369) );
  AOI21_X1 U4842 ( .B1(n4370), .B2(n4397), .A(n4369), .ZN(n4371) );
  OAI21_X1 U4843 ( .B1(n4396), .B2(n4372), .A(n4371), .ZN(n4380) );
  OR2_X1 U4844 ( .A1(\x_mult_f[14][8] ), .A2(\x_mult_f[15][8] ), .ZN(n4379) );
  NAND2_X1 U4845 ( .A1(\x_mult_f[14][8] ), .A2(\x_mult_f[15][8] ), .ZN(n4377)
         );
  NAND2_X1 U4846 ( .A1(n4379), .A2(n4377), .ZN(n4373) );
  XNOR2_X1 U4847 ( .A(n4380), .B(n4373), .ZN(n4374) );
  AOI22_X1 U4848 ( .A1(n8057), .A2(\adder_stage1[7][8] ), .B1(n8153), .B2(
        n4374), .ZN(n4375) );
  INV_X1 U4849 ( .A(n4375), .ZN(n10045) );
  AOI22_X1 U4850 ( .A1(n8336), .A2(\x_mult_f[15][5] ), .B1(n8153), .B2(
        \x_mult_f_int[15][5] ), .ZN(n4376) );
  INV_X1 U4851 ( .A(n4376), .ZN(n9119) );
  INV_X1 U4852 ( .A(n4377), .ZN(n4378) );
  AOI21_X1 U4853 ( .B1(n4380), .B2(n4379), .A(n4378), .ZN(n4389) );
  NOR2_X1 U4854 ( .A1(\x_mult_f[14][9] ), .A2(\x_mult_f[15][9] ), .ZN(n4388)
         );
  INV_X1 U4855 ( .A(n4388), .ZN(n4381) );
  NAND2_X1 U4856 ( .A1(\x_mult_f[14][9] ), .A2(\x_mult_f[15][9] ), .ZN(n4387)
         );
  NAND2_X1 U4857 ( .A1(n4381), .A2(n4387), .ZN(n4382) );
  XOR2_X1 U4858 ( .A(n4389), .B(n4382), .Z(n4383) );
  AOI22_X1 U4859 ( .A1(n8176), .A2(\adder_stage1[7][9] ), .B1(n8153), .B2(
        n4383), .ZN(n4384) );
  INV_X1 U4860 ( .A(n4384), .ZN(n10044) );
  AOI22_X1 U4861 ( .A1(n7525), .A2(\x_mult_f[14][1] ), .B1(n8153), .B2(
        \x_mult_f_int[14][1] ), .ZN(n4386) );
  INV_X1 U4862 ( .A(n4386), .ZN(n9354) );
  OAI21_X1 U4863 ( .B1(n4389), .B2(n4388), .A(n4387), .ZN(n8145) );
  OR2_X1 U4864 ( .A1(\x_mult_f[14][10] ), .A2(\x_mult_f[15][10] ), .ZN(n6879)
         );
  NAND2_X1 U4865 ( .A1(\x_mult_f[14][10] ), .A2(\x_mult_f[15][10] ), .ZN(n4406) );
  NAND2_X1 U4866 ( .A1(n6879), .A2(n4406), .ZN(n4390) );
  XNOR2_X1 U4867 ( .A(n8145), .B(n4390), .ZN(n4391) );
  AOI22_X1 U4868 ( .A1(n7855), .A2(\adder_stage1[7][10] ), .B1(n8153), .B2(
        n4391), .ZN(n4392) );
  INV_X1 U4869 ( .A(n4392), .ZN(n10043) );
  AOI22_X1 U4870 ( .A1(n8057), .A2(\x_mult_f[15][4] ), .B1(n8153), .B2(
        \x_mult_f_int[15][4] ), .ZN(n4393) );
  INV_X1 U4871 ( .A(n4393), .ZN(n9120) );
  AOI22_X1 U4872 ( .A1(n7855), .A2(\x_mult_f[15][0] ), .B1(n8153), .B2(
        \x_mult_f_int[15][0] ), .ZN(n4394) );
  INV_X1 U4873 ( .A(n4394), .ZN(n9357) );
  AOI22_X1 U4874 ( .A1(n6273), .A2(\x_mult_f[14][0] ), .B1(n8153), .B2(
        \x_mult_f_int[14][0] ), .ZN(n4395) );
  INV_X1 U4875 ( .A(n4395), .ZN(n9355) );
  INV_X1 U4876 ( .A(n4396), .ZN(n5816) );
  AOI21_X1 U4877 ( .B1(n5816), .B2(n4398), .A(n4397), .ZN(n5801) );
  OAI21_X1 U4878 ( .B1(n5801), .B2(n5797), .A(n5798), .ZN(n4403) );
  INV_X1 U4879 ( .A(n4399), .ZN(n4401) );
  NAND2_X1 U4880 ( .A1(n4401), .A2(n4400), .ZN(n4402) );
  XNOR2_X1 U4881 ( .A(n4403), .B(n4402), .ZN(n4404) );
  AOI22_X1 U4882 ( .A1(n8401), .A2(\adder_stage1[7][7] ), .B1(n8153), .B2(
        n4404), .ZN(n4405) );
  INV_X1 U4883 ( .A(n4405), .ZN(n10046) );
  INV_X1 U4884 ( .A(n4406), .ZN(n6884) );
  AOI21_X1 U4885 ( .B1(n8145), .B2(n6879), .A(n6884), .ZN(n4408) );
  OR2_X1 U4886 ( .A1(\x_mult_f[14][11] ), .A2(\x_mult_f[15][11] ), .ZN(n6883)
         );
  NAND2_X1 U4887 ( .A1(\x_mult_f[14][11] ), .A2(\x_mult_f[15][11] ), .ZN(n6881) );
  NAND2_X1 U4888 ( .A1(n6883), .A2(n6881), .ZN(n4407) );
  XOR2_X1 U4889 ( .A(n4408), .B(n4407), .Z(n4409) );
  AOI22_X1 U4890 ( .A1(n8057), .A2(\adder_stage1[7][11] ), .B1(n8153), .B2(
        n4409), .ZN(n4410) );
  INV_X1 U4891 ( .A(n4410), .ZN(n10042) );
  BUF_X2 U4892 ( .A(n3445), .Z(n8045) );
  AOI22_X1 U4893 ( .A1(\x_mult_f_int[25][11] ), .A2(n8332), .B1(n7864), .B2(
        \x_mult_f[25][11] ), .ZN(n4411) );
  INV_X1 U4894 ( .A(n4411), .ZN(n9234) );
  AOI22_X1 U4895 ( .A1(\x_mult_f_int[25][10] ), .A2(n8332), .B1(n7864), .B2(
        \x_mult_f[25][10] ), .ZN(n4412) );
  INV_X1 U4896 ( .A(n4412), .ZN(n9235) );
  AOI22_X1 U4897 ( .A1(\x_mult_f_int[25][9] ), .A2(n8332), .B1(n7864), .B2(
        \x_mult_f[25][9] ), .ZN(n4413) );
  INV_X1 U4898 ( .A(n4413), .ZN(n9236) );
  NOR2_X1 U4899 ( .A1(\x_mult_f[30][1] ), .A2(\x_mult_f[31][1] ), .ZN(n4437)
         );
  NAND2_X1 U4900 ( .A1(\x_mult_f[30][0] ), .A2(\x_mult_f[31][0] ), .ZN(n4440)
         );
  NAND2_X1 U4901 ( .A1(\x_mult_f[30][1] ), .A2(\x_mult_f[31][1] ), .ZN(n4438)
         );
  OAI21_X1 U4902 ( .B1(n4437), .B2(n4440), .A(n4438), .ZN(n4432) );
  INV_X1 U4903 ( .A(n4432), .ZN(n4421) );
  NOR2_X1 U4904 ( .A1(\x_mult_f[30][2] ), .A2(\x_mult_f[31][2] ), .ZN(n4427)
         );
  NAND2_X1 U4905 ( .A1(\x_mult_f[31][2] ), .A2(\x_mult_f[30][2] ), .ZN(n4429)
         );
  OAI21_X1 U4906 ( .B1(n4421), .B2(n4427), .A(n4429), .ZN(n4416) );
  INV_X1 U4907 ( .A(n4430), .ZN(n4414) );
  NAND2_X1 U4908 ( .A1(\x_mult_f[30][3] ), .A2(\x_mult_f[31][3] ), .ZN(n4428)
         );
  NAND2_X1 U4909 ( .A1(n4414), .A2(n4428), .ZN(n4415) );
  XNOR2_X1 U4910 ( .A(n4416), .B(n4415), .ZN(n4417) );
  AOI22_X1 U4911 ( .A1(n8118), .A2(\adder_stage1[15][3] ), .B1(n7927), .B2(
        n4417), .ZN(n4418) );
  INV_X1 U4912 ( .A(n4418), .ZN(n9915) );
  INV_X1 U4913 ( .A(n4427), .ZN(n4419) );
  NAND2_X1 U4914 ( .A1(n4419), .A2(n4429), .ZN(n4420) );
  XOR2_X1 U4915 ( .A(n4421), .B(n4420), .Z(n4422) );
  AOI22_X1 U4916 ( .A1(n8434), .A2(\adder_stage1[15][2] ), .B1(n7927), .B2(
        n4422), .ZN(n4423) );
  INV_X1 U4917 ( .A(n4423), .ZN(n9916) );
  OR2_X1 U4918 ( .A1(\x_mult_f[30][0] ), .A2(\x_mult_f[31][0] ), .ZN(n4424) );
  AND2_X1 U4919 ( .A1(n4424), .A2(n4440), .ZN(n4425) );
  AOI22_X1 U4920 ( .A1(n6877), .A2(\adder_stage1[15][0] ), .B1(n7927), .B2(
        n4425), .ZN(n4426) );
  INV_X1 U4921 ( .A(n4426), .ZN(n9918) );
  NOR2_X1 U4922 ( .A1(n4427), .A2(n4430), .ZN(n4433) );
  OAI21_X1 U4923 ( .B1(n4430), .B2(n4429), .A(n4428), .ZN(n4431) );
  INV_X1 U4924 ( .A(n7349), .ZN(n7443) );
  NOR2_X1 U4925 ( .A1(\x_mult_f[30][4] ), .A2(\x_mult_f[31][4] ), .ZN(n5618)
         );
  INV_X1 U4926 ( .A(n5618), .ZN(n7442) );
  NAND2_X1 U4927 ( .A1(\x_mult_f[30][4] ), .A2(\x_mult_f[31][4] ), .ZN(n7440)
         );
  NAND2_X1 U4928 ( .A1(n7442), .A2(n7440), .ZN(n4434) );
  XNOR2_X1 U4929 ( .A(n7443), .B(n4434), .ZN(n4435) );
  AOI22_X1 U4930 ( .A1(n7614), .A2(\adder_stage1[15][4] ), .B1(n7927), .B2(
        n4435), .ZN(n4436) );
  INV_X1 U4931 ( .A(n4436), .ZN(n9914) );
  INV_X1 U4932 ( .A(n4437), .ZN(n4439) );
  NAND2_X1 U4933 ( .A1(n4439), .A2(n4438), .ZN(n4441) );
  XOR2_X1 U4934 ( .A(n4441), .B(n4440), .Z(n4442) );
  AOI22_X1 U4935 ( .A1(n7640), .A2(\adder_stage1[15][1] ), .B1(n7927), .B2(
        n4442), .ZN(n4443) );
  INV_X1 U4936 ( .A(n4443), .ZN(n9917) );
  INV_X2 U4937 ( .A(n7979), .ZN(n8118) );
  BUF_X2 U4938 ( .A(n4444), .Z(n5707) );
  NOR2_X1 U4939 ( .A1(\x_mult_f[0][4] ), .A2(\x_mult_f[1][4] ), .ZN(n4494) );
  NOR2_X1 U4940 ( .A1(\x_mult_f[0][5] ), .A2(\x_mult_f[1][5] ), .ZN(n4496) );
  NOR2_X1 U4941 ( .A1(n4494), .A2(n4496), .ZN(n5692) );
  NOR2_X1 U4942 ( .A1(\x_mult_f[1][6] ), .A2(\x_mult_f[0][6] ), .ZN(n5699) );
  NOR2_X1 U4943 ( .A1(\x_mult_f[0][7] ), .A2(\x_mult_f[1][7] ), .ZN(n5701) );
  NOR2_X1 U4944 ( .A1(n5699), .A2(n5701), .ZN(n4448) );
  NAND2_X1 U4945 ( .A1(n5692), .A2(n4448), .ZN(n4450) );
  NOR2_X1 U4946 ( .A1(\x_mult_f[0][2] ), .A2(\x_mult_f[1][2] ), .ZN(n5676) );
  NOR2_X1 U4947 ( .A1(n5676), .A2(n5657), .ZN(n4446) );
  NOR2_X1 U4948 ( .A1(\x_mult_f[0][1] ), .A2(\x_mult_f[1][1] ), .ZN(n5664) );
  NAND2_X1 U4949 ( .A1(\x_mult_f[0][0] ), .A2(\x_mult_f[1][0] ), .ZN(n5667) );
  NAND2_X1 U4950 ( .A1(\x_mult_f[0][1] ), .A2(\x_mult_f[1][1] ), .ZN(n5665) );
  OAI21_X1 U4951 ( .B1(n5664), .B2(n5667), .A(n5665), .ZN(n5656) );
  NAND2_X1 U4952 ( .A1(\x_mult_f[0][2] ), .A2(\x_mult_f[1][2] ), .ZN(n5677) );
  NAND2_X1 U4953 ( .A1(\x_mult_f[0][3] ), .A2(\x_mult_f[1][3] ), .ZN(n5658) );
  OAI21_X1 U4954 ( .B1(n5657), .B2(n5677), .A(n5658), .ZN(n4445) );
  NAND2_X1 U4955 ( .A1(\x_mult_f[0][4] ), .A2(\x_mult_f[1][4] ), .ZN(n5671) );
  NAND2_X1 U4956 ( .A1(\x_mult_f[0][5] ), .A2(\x_mult_f[1][5] ), .ZN(n4497) );
  OAI21_X1 U4957 ( .B1(n4496), .B2(n5671), .A(n4497), .ZN(n5691) );
  NAND2_X1 U4958 ( .A1(\x_mult_f[0][6] ), .A2(\x_mult_f[1][6] ), .ZN(n5698) );
  NAND2_X1 U4959 ( .A1(\x_mult_f[0][7] ), .A2(\x_mult_f[1][7] ), .ZN(n5702) );
  OAI21_X1 U4960 ( .B1(n5701), .B2(n5698), .A(n5702), .ZN(n4447) );
  AOI21_X1 U4961 ( .B1(n4448), .B2(n5691), .A(n4447), .ZN(n4449) );
  OAI21_X1 U4962 ( .B1(n4450), .B2(n4493), .A(n4449), .ZN(n4476) );
  OR2_X1 U4963 ( .A1(\x_mult_f[0][8] ), .A2(\x_mult_f[1][8] ), .ZN(n4466) );
  NAND2_X1 U4964 ( .A1(\x_mult_f[0][8] ), .A2(\x_mult_f[1][8] ), .ZN(n4465) );
  INV_X1 U4965 ( .A(n4465), .ZN(n4459) );
  AOI21_X1 U4966 ( .B1(n4455), .B2(n4466), .A(n4459), .ZN(n4452) );
  OR2_X1 U4967 ( .A1(\x_mult_f[0][9] ), .A2(\x_mult_f[1][9] ), .ZN(n4458) );
  NAND2_X1 U4968 ( .A1(\x_mult_f[0][9] ), .A2(\x_mult_f[1][9] ), .ZN(n4456) );
  NAND2_X1 U4969 ( .A1(n4458), .A2(n4456), .ZN(n4451) );
  XOR2_X1 U4970 ( .A(n4452), .B(n4451), .Z(n4453) );
  AOI22_X1 U4971 ( .A1(n8118), .A2(\adder_stage1[0][9] ), .B1(n5707), .B2(
        n4453), .ZN(n4454) );
  INV_X1 U4972 ( .A(n4454), .ZN(n10160) );
  AND2_X1 U4973 ( .A1(n4466), .A2(n4458), .ZN(n4470) );
  NAND2_X1 U4974 ( .A1(n4455), .A2(n4470), .ZN(n4460) );
  INV_X1 U4975 ( .A(n4456), .ZN(n4457) );
  AOI21_X1 U4976 ( .B1(n4459), .B2(n4458), .A(n4457), .ZN(n4474) );
  NAND2_X1 U4977 ( .A1(n4460), .A2(n4474), .ZN(n4462) );
  OR2_X1 U4978 ( .A1(\x_mult_f[0][10] ), .A2(\x_mult_f[1][10] ), .ZN(n4471) );
  NAND2_X1 U4979 ( .A1(\x_mult_f[0][10] ), .A2(\x_mult_f[1][10] ), .ZN(n4472)
         );
  NAND2_X1 U4980 ( .A1(n4471), .A2(n4472), .ZN(n4461) );
  XNOR2_X1 U4981 ( .A(n4462), .B(n4461), .ZN(n4463) );
  AOI22_X1 U4982 ( .A1(n8118), .A2(\adder_stage1[0][10] ), .B1(n5707), .B2(
        n4463), .ZN(n4464) );
  INV_X1 U4983 ( .A(n4464), .ZN(n10159) );
  NAND2_X1 U4984 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  XNOR2_X1 U4985 ( .A(n4476), .B(n4467), .ZN(n4468) );
  AOI22_X1 U4986 ( .A1(n8118), .A2(\adder_stage1[0][8] ), .B1(n5707), .B2(
        n4468), .ZN(n4469) );
  INV_X1 U4987 ( .A(n4469), .ZN(n10161) );
  AND2_X1 U4988 ( .A1(n4470), .A2(n4471), .ZN(n4477) );
  INV_X1 U4989 ( .A(n4471), .ZN(n4473) );
  OAI21_X1 U4990 ( .B1(n4474), .B2(n4473), .A(n4472), .ZN(n4475) );
  AOI21_X1 U4991 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4484) );
  NOR2_X1 U4992 ( .A1(\x_mult_f[0][11] ), .A2(\x_mult_f[1][11] ), .ZN(n4483)
         );
  INV_X1 U4993 ( .A(n4483), .ZN(n4478) );
  NAND2_X1 U4994 ( .A1(\x_mult_f[0][11] ), .A2(\x_mult_f[1][11] ), .ZN(n4482)
         );
  NAND2_X1 U4995 ( .A1(n4478), .A2(n4482), .ZN(n4479) );
  XOR2_X1 U4996 ( .A(n4484), .B(n4479), .Z(n4480) );
  AOI22_X1 U4997 ( .A1(n8118), .A2(\adder_stage1[0][11] ), .B1(n5707), .B2(
        n4480), .ZN(n4481) );
  INV_X1 U4998 ( .A(n4481), .ZN(n10158) );
  OAI21_X1 U4999 ( .B1(n4484), .B2(n4483), .A(n4482), .ZN(n6063) );
  OR2_X1 U5000 ( .A1(\x_mult_f[0][12] ), .A2(\x_mult_f[1][12] ), .ZN(n6062) );
  NAND2_X1 U5001 ( .A1(\x_mult_f[0][12] ), .A2(\x_mult_f[1][12] ), .ZN(n6060)
         );
  NAND2_X1 U5002 ( .A1(n6062), .A2(n6060), .ZN(n4485) );
  XNOR2_X1 U5003 ( .A(n3422), .B(n4485), .ZN(n4486) );
  AOI22_X1 U5004 ( .A1(n8118), .A2(\adder_stage1[0][12] ), .B1(n5707), .B2(
        n4486), .ZN(n4487) );
  INV_X1 U5005 ( .A(n4487), .ZN(n10157) );
  AOI22_X1 U5006 ( .A1(n7952), .A2(\x_mult_f[30][0] ), .B1(n4645), .B2(
        \x_mult_f_int[30][0] ), .ZN(n4488) );
  INV_X1 U5007 ( .A(n4488), .ZN(n9387) );
  AOI22_X1 U5008 ( .A1(n7864), .A2(\x_mult_f[26][2] ), .B1(n8216), .B2(
        \x_mult_f_int[26][2] ), .ZN(n4489) );
  INV_X1 U5009 ( .A(n4489), .ZN(n9257) );
  AOI22_X1 U5010 ( .A1(n8273), .A2(\x_mult_f[27][5] ), .B1(n8265), .B2(
        \x_mult_f_int[27][5] ), .ZN(n4490) );
  INV_X1 U5011 ( .A(n4490), .ZN(n9268) );
  AOI22_X1 U5012 ( .A1(n8328), .A2(\x_mult_f[26][1] ), .B1(n8105), .B2(
        \x_mult_f_int[26][1] ), .ZN(n4491) );
  INV_X1 U5013 ( .A(n4491), .ZN(n9378) );
  AOI22_X1 U5014 ( .A1(n8296), .A2(\x_mult_f[26][0] ), .B1(n8167), .B2(
        \x_mult_f_int[26][0] ), .ZN(n4492) );
  INV_X1 U5015 ( .A(n4492), .ZN(n9379) );
  INV_X2 U5016 ( .A(n7979), .ZN(n7074) );
  INV_X1 U5017 ( .A(n4493), .ZN(n5693) );
  INV_X1 U5018 ( .A(n4494), .ZN(n5672) );
  INV_X1 U5019 ( .A(n5671), .ZN(n4495) );
  AOI21_X1 U5020 ( .B1(n5693), .B2(n5672), .A(n4495), .ZN(n4500) );
  INV_X1 U5021 ( .A(n4496), .ZN(n4498) );
  NAND2_X1 U5022 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  XOR2_X1 U5023 ( .A(n4500), .B(n4499), .Z(n4501) );
  AOI22_X1 U5024 ( .A1(n7074), .A2(\adder_stage1[0][5] ), .B1(n5707), .B2(
        n4501), .ZN(n4502) );
  INV_X1 U5025 ( .A(n4502), .ZN(n10164) );
  NOR2_X1 U5026 ( .A1(\x_mult_f[24][1] ), .A2(\x_mult_f[25][1] ), .ZN(n4523)
         );
  NAND2_X1 U5027 ( .A1(\x_mult_f[24][0] ), .A2(\x_mult_f[25][0] ), .ZN(n4529)
         );
  NAND2_X1 U5028 ( .A1(\x_mult_f[24][1] ), .A2(\x_mult_f[25][1] ), .ZN(n4524)
         );
  OAI21_X1 U5029 ( .B1(n4523), .B2(n4529), .A(n4524), .ZN(n4511) );
  INV_X1 U5030 ( .A(n4511), .ZN(n4520) );
  NOR2_X1 U5031 ( .A1(\x_mult_f[24][2] ), .A2(\x_mult_f[25][2] ), .ZN(n4516)
         );
  NAND2_X1 U5032 ( .A1(\x_mult_f[24][2] ), .A2(\x_mult_f[25][2] ), .ZN(n4517)
         );
  OAI21_X1 U5033 ( .B1(n4520), .B2(n4516), .A(n4517), .ZN(n4505) );
  NOR2_X1 U5034 ( .A1(\x_mult_f[24][3] ), .A2(\x_mult_f[25][3] ), .ZN(n4509)
         );
  INV_X1 U5035 ( .A(n4509), .ZN(n4503) );
  NAND2_X1 U5036 ( .A1(\x_mult_f[24][3] ), .A2(\x_mult_f[25][3] ), .ZN(n4508)
         );
  NAND2_X1 U5037 ( .A1(n4503), .A2(n4508), .ZN(n4504) );
  XNOR2_X1 U5038 ( .A(n4505), .B(n4504), .ZN(n4506) );
  AOI22_X1 U5039 ( .A1(n7177), .A2(\adder_stage1[12][3] ), .B1(n7507), .B2(
        n4506), .ZN(n4507) );
  INV_X1 U5040 ( .A(n4507), .ZN(n9966) );
  NOR2_X1 U5041 ( .A1(n4516), .A2(n4509), .ZN(n4512) );
  OAI21_X1 U5042 ( .B1(n4509), .B2(n4517), .A(n4508), .ZN(n4510) );
  AOI21_X1 U5043 ( .B1(n4512), .B2(n4511), .A(n4510), .ZN(n5640) );
  INV_X1 U5044 ( .A(n5640), .ZN(n6021) );
  NOR2_X1 U5045 ( .A1(\x_mult_f[24][4] ), .A2(\x_mult_f[25][4] ), .ZN(n5635)
         );
  INV_X1 U5046 ( .A(n5635), .ZN(n6020) );
  NAND2_X1 U5047 ( .A1(\x_mult_f[24][4] ), .A2(\x_mult_f[25][4] ), .ZN(n6018)
         );
  NAND2_X1 U5048 ( .A1(n6020), .A2(n6018), .ZN(n4513) );
  XNOR2_X1 U5049 ( .A(n6021), .B(n4513), .ZN(n4514) );
  AOI22_X1 U5050 ( .A1(n8245), .A2(\adder_stage1[12][4] ), .B1(n8024), .B2(
        n4514), .ZN(n4515) );
  INV_X1 U5051 ( .A(n4515), .ZN(n9965) );
  INV_X1 U5052 ( .A(n4516), .ZN(n4518) );
  NAND2_X1 U5053 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  XOR2_X1 U5054 ( .A(n4520), .B(n4519), .Z(n4521) );
  AOI22_X1 U5055 ( .A1(n8273), .A2(\adder_stage1[12][2] ), .B1(n6279), .B2(
        n4521), .ZN(n4522) );
  INV_X1 U5056 ( .A(n4522), .ZN(n9967) );
  INV_X1 U5057 ( .A(n4523), .ZN(n4525) );
  NAND2_X1 U5058 ( .A1(n4525), .A2(n4524), .ZN(n4526) );
  XOR2_X1 U5059 ( .A(n4526), .B(n4529), .Z(n4527) );
  AOI22_X1 U5060 ( .A1(n7920), .A2(\adder_stage1[12][1] ), .B1(n8216), .B2(
        n4527), .ZN(n4528) );
  INV_X1 U5061 ( .A(n4528), .ZN(n9968) );
  OR2_X1 U5062 ( .A1(\x_mult_f[24][0] ), .A2(\x_mult_f[25][0] ), .ZN(n4530) );
  AND2_X1 U5063 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  AOI22_X1 U5064 ( .A1(n7855), .A2(\adder_stage1[12][0] ), .B1(n8265), .B2(
        n4531), .ZN(n4532) );
  INV_X1 U5065 ( .A(n4532), .ZN(n9969) );
  AOI22_X1 U5066 ( .A1(\x_mult_f_int[13][6] ), .A2(n4257), .B1(n7972), .B2(
        \x_mult_f[13][6] ), .ZN(n4533) );
  INV_X1 U5067 ( .A(n4533), .ZN(n9090) );
  AOI22_X1 U5068 ( .A1(\x_mult_f_int[13][7] ), .A2(n8281), .B1(n8296), .B2(
        \x_mult_f[13][7] ), .ZN(n4534) );
  INV_X1 U5069 ( .A(n4534), .ZN(n9089) );
  AOI22_X1 U5070 ( .A1(\x_mult_f_int[13][8] ), .A2(n5981), .B1(n8176), .B2(
        \x_mult_f[13][8] ), .ZN(n4535) );
  INV_X1 U5071 ( .A(n4535), .ZN(n9088) );
  AOI22_X1 U5072 ( .A1(\x_mult_f_int[13][10] ), .A2(n6875), .B1(n8340), .B2(
        \x_mult_f[13][10] ), .ZN(n4536) );
  INV_X1 U5073 ( .A(n4536), .ZN(n9086) );
  AOI22_X1 U5074 ( .A1(\x_mult_f_int[13][9] ), .A2(n8292), .B1(n7972), .B2(
        \x_mult_f[13][9] ), .ZN(n4537) );
  INV_X1 U5075 ( .A(n4537), .ZN(n9087) );
  NOR2_X1 U5076 ( .A1(n4538), .A2(n4541), .ZN(n4544) );
  OAI21_X1 U5077 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4542) );
  AOI21_X1 U5078 ( .B1(n4544), .B2(n4543), .A(n4542), .ZN(n6190) );
  INV_X1 U5079 ( .A(n6190), .ZN(n6685) );
  NOR2_X1 U5080 ( .A1(\adder_stage3[2][4] ), .A2(\adder_stage3[3][4] ), .ZN(
        n6182) );
  INV_X1 U5081 ( .A(n6182), .ZN(n4549) );
  NAND2_X1 U5082 ( .A1(\adder_stage3[2][4] ), .A2(\adder_stage3[3][4] ), .ZN(
        n6184) );
  NAND2_X1 U5083 ( .A1(n4549), .A2(n6184), .ZN(n4545) );
  XNOR2_X1 U5084 ( .A(n6685), .B(n4545), .ZN(n4546) );
  AOI22_X1 U5085 ( .A1(n8336), .A2(\adder_stage4[1][4] ), .B1(n5707), .B2(
        n4546), .ZN(n4547) );
  INV_X1 U5086 ( .A(n4547), .ZN(n9662) );
  INV_X1 U5087 ( .A(n6184), .ZN(n4548) );
  AOI21_X1 U5088 ( .B1(n6685), .B2(n4549), .A(n4548), .ZN(n4552) );
  NOR2_X1 U5089 ( .A1(\adder_stage3[2][5] ), .A2(\adder_stage3[3][5] ), .ZN(
        n6185) );
  INV_X1 U5090 ( .A(n6185), .ZN(n4550) );
  NAND2_X1 U5091 ( .A1(\adder_stage3[2][5] ), .A2(\adder_stage3[3][5] ), .ZN(
        n6183) );
  NAND2_X1 U5092 ( .A1(n4550), .A2(n6183), .ZN(n4551) );
  XOR2_X1 U5093 ( .A(n4552), .B(n4551), .Z(n4553) );
  AOI22_X1 U5094 ( .A1(n8088), .A2(\adder_stage4[1][5] ), .B1(n4311), .B2(
        n4553), .ZN(n4554) );
  INV_X1 U5095 ( .A(n4554), .ZN(n9661) );
  INV_X2 U5096 ( .A(n7979), .ZN(n6854) );
  NOR2_X1 U5097 ( .A1(\x_mult_f[10][1] ), .A2(\x_mult_f[11][1] ), .ZN(n4568)
         );
  NAND2_X1 U5098 ( .A1(\x_mult_f[10][0] ), .A2(\x_mult_f[11][0] ), .ZN(n4571)
         );
  NAND2_X1 U5099 ( .A1(\x_mult_f[10][1] ), .A2(\x_mult_f[11][1] ), .ZN(n4569)
         );
  OAI21_X1 U5100 ( .B1(n4568), .B2(n4571), .A(n4569), .ZN(n4652) );
  INV_X1 U5101 ( .A(n4652), .ZN(n4565) );
  NOR2_X1 U5102 ( .A1(\x_mult_f[10][2] ), .A2(\x_mult_f[11][2] ), .ZN(n4647)
         );
  NAND2_X1 U5103 ( .A1(\x_mult_f[10][2] ), .A2(\x_mult_f[11][2] ), .ZN(n4649)
         );
  OAI21_X1 U5104 ( .B1(n4565), .B2(n4647), .A(n4649), .ZN(n4557) );
  NOR2_X1 U5105 ( .A1(\x_mult_f[10][3] ), .A2(\x_mult_f[11][3] ), .ZN(n4650)
         );
  INV_X1 U5106 ( .A(n4650), .ZN(n4555) );
  NAND2_X1 U5107 ( .A1(\x_mult_f[10][3] ), .A2(\x_mult_f[11][3] ), .ZN(n4648)
         );
  NAND2_X1 U5108 ( .A1(n4555), .A2(n4648), .ZN(n4556) );
  XNOR2_X1 U5109 ( .A(n4557), .B(n4556), .ZN(n4558) );
  AOI22_X1 U5110 ( .A1(n6854), .A2(\adder_stage1[5][3] ), .B1(n6036), .B2(
        n4558), .ZN(n4559) );
  INV_X1 U5111 ( .A(n4559), .ZN(n10083) );
  OR2_X1 U5112 ( .A1(\x_mult_f[10][0] ), .A2(\x_mult_f[11][0] ), .ZN(n4560) );
  AND2_X1 U5113 ( .A1(n4560), .A2(n4571), .ZN(n4561) );
  AOI22_X1 U5114 ( .A1(n6854), .A2(\adder_stage1[5][0] ), .B1(n8209), .B2(
        n4561), .ZN(n4562) );
  INV_X1 U5115 ( .A(n4562), .ZN(n10086) );
  INV_X1 U5116 ( .A(n4647), .ZN(n4563) );
  NAND2_X1 U5117 ( .A1(n4563), .A2(n4649), .ZN(n4564) );
  XOR2_X1 U5118 ( .A(n4565), .B(n4564), .Z(n4566) );
  AOI22_X1 U5119 ( .A1(n6854), .A2(\adder_stage1[5][2] ), .B1(n6272), .B2(
        n4566), .ZN(n4567) );
  INV_X1 U5120 ( .A(n4567), .ZN(n10084) );
  INV_X1 U5121 ( .A(n4568), .ZN(n4570) );
  NAND2_X1 U5122 ( .A1(n4570), .A2(n4569), .ZN(n4572) );
  XOR2_X1 U5123 ( .A(n4572), .B(n4571), .Z(n4573) );
  AOI22_X1 U5124 ( .A1(n6854), .A2(\adder_stage1[5][1] ), .B1(n8024), .B2(
        n4573), .ZN(n4574) );
  INV_X1 U5125 ( .A(n4574), .ZN(n10085) );
  AOI22_X1 U5126 ( .A1(n7920), .A2(\x_mult_f[28][4] ), .B1(n8054), .B2(
        \x_mult_f_int[28][4] ), .ZN(n4575) );
  INV_X1 U5127 ( .A(n4575), .ZN(n9283) );
  AOI22_X1 U5128 ( .A1(n8168), .A2(\x_mult_f[28][0] ), .B1(n8251), .B2(
        \x_mult_f_int[28][0] ), .ZN(n4576) );
  INV_X1 U5129 ( .A(n4576), .ZN(n9383) );
  NOR2_X1 U5130 ( .A1(\adder_stage1[4][2] ), .A2(\adder_stage1[5][2] ), .ZN(
        n4911) );
  NOR2_X1 U5131 ( .A1(\adder_stage1[4][3] ), .A2(\adder_stage1[5][3] ), .ZN(
        n4913) );
  NOR2_X1 U5132 ( .A1(n4911), .A2(n4913), .ZN(n4578) );
  NOR2_X1 U5133 ( .A1(\adder_stage1[4][1] ), .A2(\adder_stage1[5][1] ), .ZN(
        n4920) );
  NAND2_X1 U5134 ( .A1(\adder_stage1[4][0] ), .A2(\adder_stage1[5][0] ), .ZN(
        n4923) );
  NAND2_X1 U5135 ( .A1(\adder_stage1[4][1] ), .A2(\adder_stage1[5][1] ), .ZN(
        n4921) );
  OAI21_X1 U5136 ( .B1(n4920), .B2(n4923), .A(n4921), .ZN(n4905) );
  NAND2_X1 U5137 ( .A1(\adder_stage1[4][2] ), .A2(\adder_stage1[5][2] ), .ZN(
        n4910) );
  NAND2_X1 U5138 ( .A1(\adder_stage1[4][3] ), .A2(\adder_stage1[5][3] ), .ZN(
        n4914) );
  OAI21_X1 U5139 ( .B1(n4913), .B2(n4910), .A(n4914), .ZN(n4577) );
  AOI21_X1 U5140 ( .B1(n4578), .B2(n4905), .A(n4577), .ZN(n4927) );
  NOR2_X1 U5141 ( .A1(\adder_stage1[4][4] ), .A2(\adder_stage1[5][4] ), .ZN(
        n4928) );
  NOR2_X1 U5142 ( .A1(\adder_stage1[4][5] ), .A2(\adder_stage1[5][5] ), .ZN(
        n8111) );
  NOR2_X1 U5143 ( .A1(n4928), .A2(n8111), .ZN(n5044) );
  NOR2_X1 U5144 ( .A1(\adder_stage1[4][7] ), .A2(\adder_stage1[5][7] ), .ZN(
        n5052) );
  NOR2_X1 U5145 ( .A1(\adder_stage1[4][6] ), .A2(\adder_stage1[5][6] ), .ZN(
        n5050) );
  NOR2_X1 U5146 ( .A1(n5052), .A2(n5050), .ZN(n4580) );
  NAND2_X1 U5147 ( .A1(n5044), .A2(n4580), .ZN(n4582) );
  NAND2_X1 U5148 ( .A1(\adder_stage1[4][4] ), .A2(\adder_stage1[5][4] ), .ZN(
        n8107) );
  NAND2_X1 U5149 ( .A1(\adder_stage1[4][5] ), .A2(\adder_stage1[5][5] ), .ZN(
        n8112) );
  OAI21_X1 U5150 ( .B1(n8111), .B2(n8107), .A(n8112), .ZN(n5043) );
  NAND2_X1 U5151 ( .A1(\adder_stage1[4][6] ), .A2(\adder_stage1[5][6] ), .ZN(
        n5049) );
  NAND2_X1 U5152 ( .A1(\adder_stage1[4][7] ), .A2(\adder_stage1[5][7] ), .ZN(
        n5053) );
  OAI21_X1 U5153 ( .B1(n5052), .B2(n5049), .A(n5053), .ZN(n4579) );
  AOI21_X1 U5154 ( .B1(n4580), .B2(n5043), .A(n4579), .ZN(n4581) );
  OAI21_X1 U5155 ( .B1(n4927), .B2(n4582), .A(n4581), .ZN(n7052) );
  NOR2_X1 U5156 ( .A1(\adder_stage1[4][8] ), .A2(\adder_stage1[5][8] ), .ZN(
        n7053) );
  INV_X1 U5157 ( .A(n7053), .ZN(n7070) );
  OR2_X1 U5158 ( .A1(\adder_stage1[4][9] ), .A2(\adder_stage1[5][9] ), .ZN(
        n7055) );
  NAND2_X1 U5159 ( .A1(n7070), .A2(n7055), .ZN(n7061) );
  NOR2_X1 U5160 ( .A1(\adder_stage1[4][10] ), .A2(\adder_stage1[5][10] ), .ZN(
        n7062) );
  NOR2_X1 U5161 ( .A1(n7061), .A2(n7062), .ZN(n4586) );
  NAND2_X1 U5162 ( .A1(\adder_stage1[4][8] ), .A2(\adder_stage1[5][8] ), .ZN(
        n7069) );
  INV_X1 U5163 ( .A(n7069), .ZN(n4584) );
  NAND2_X1 U5164 ( .A1(\adder_stage1[4][9] ), .A2(\adder_stage1[5][9] ), .ZN(
        n7054) );
  INV_X1 U5165 ( .A(n7054), .ZN(n4583) );
  AOI21_X1 U5166 ( .B1(n7055), .B2(n4584), .A(n4583), .ZN(n7060) );
  NAND2_X1 U5167 ( .A1(\adder_stage1[4][10] ), .A2(\adder_stage1[5][10] ), 
        .ZN(n7063) );
  OAI21_X1 U5168 ( .B1(n7060), .B2(n7062), .A(n7063), .ZN(n4585) );
  AOI21_X1 U5169 ( .B1(n7052), .B2(n4586), .A(n4585), .ZN(n7049) );
  OR2_X1 U5170 ( .A1(\adder_stage1[4][12] ), .A2(\adder_stage1[5][12] ), .ZN(
        n5061) );
  NOR2_X1 U5171 ( .A1(\adder_stage1[4][11] ), .A2(\adder_stage1[5][11] ), .ZN(
        n5059) );
  INV_X1 U5172 ( .A(n5059), .ZN(n7047) );
  NAND2_X1 U5173 ( .A1(n5061), .A2(n7047), .ZN(n4596) );
  INV_X1 U5174 ( .A(n4596), .ZN(n4587) );
  NOR2_X1 U5175 ( .A1(\adder_stage1[4][13] ), .A2(\adder_stage1[5][13] ), .ZN(
        n4590) );
  INV_X1 U5176 ( .A(n4590), .ZN(n4601) );
  NAND2_X1 U5177 ( .A1(n4587), .A2(n4601), .ZN(n5400) );
  NAND2_X1 U5178 ( .A1(\adder_stage1[4][11] ), .A2(\adder_stage1[5][11] ), 
        .ZN(n7046) );
  INV_X1 U5179 ( .A(n7046), .ZN(n4589) );
  NAND2_X1 U5180 ( .A1(\adder_stage1[4][12] ), .A2(\adder_stage1[5][12] ), 
        .ZN(n5060) );
  INV_X1 U5181 ( .A(n5060), .ZN(n4588) );
  AOI21_X1 U5182 ( .B1(n5061), .B2(n4589), .A(n4588), .ZN(n4597) );
  NAND2_X1 U5183 ( .A1(\adder_stage1[4][13] ), .A2(\adder_stage1[5][13] ), 
        .ZN(n4600) );
  OAI21_X1 U5184 ( .B1(n4597), .B2(n4590), .A(n4600), .ZN(n4591) );
  INV_X1 U5185 ( .A(n4591), .ZN(n5403) );
  OAI21_X1 U5186 ( .B1(n7049), .B2(n5400), .A(n5403), .ZN(n4593) );
  OR2_X1 U5187 ( .A1(\adder_stage1[4][14] ), .A2(\adder_stage1[5][14] ), .ZN(
        n5399) );
  NAND2_X1 U5188 ( .A1(\adder_stage1[4][14] ), .A2(\adder_stage1[5][14] ), 
        .ZN(n5401) );
  NAND2_X1 U5189 ( .A1(n5399), .A2(n5401), .ZN(n4592) );
  XNOR2_X1 U5190 ( .A(n4593), .B(n4592), .ZN(n4594) );
  AOI22_X1 U5191 ( .A1(n7074), .A2(\adder_stage2[2][14] ), .B1(n5767), .B2(
        n4594), .ZN(n4595) );
  INV_X1 U5192 ( .A(n4595), .ZN(n9856) );
  NOR2_X1 U5193 ( .A1(n7049), .A2(n4596), .ZN(n4599) );
  INV_X1 U5194 ( .A(n4597), .ZN(n4598) );
  NOR2_X1 U5195 ( .A1(n4599), .A2(n4598), .ZN(n4603) );
  NAND2_X1 U5196 ( .A1(n4601), .A2(n4600), .ZN(n4602) );
  XOR2_X1 U5197 ( .A(n4603), .B(n4602), .Z(n4604) );
  AOI22_X1 U5198 ( .A1(n7074), .A2(\adder_stage2[2][13] ), .B1(n7507), .B2(
        n4604), .ZN(n4605) );
  INV_X1 U5199 ( .A(n4605), .ZN(n9857) );
  NOR2_X1 U5200 ( .A1(\x_mult_f[20][2] ), .A2(\x_mult_f[21][2] ), .ZN(n8155)
         );
  NOR2_X1 U5201 ( .A1(\x_mult_f[20][3] ), .A2(\x_mult_f[21][3] ), .ZN(n7598)
         );
  NOR2_X1 U5202 ( .A1(n8155), .A2(n7598), .ZN(n4607) );
  NOR2_X1 U5203 ( .A1(\x_mult_f[20][1] ), .A2(\x_mult_f[21][1] ), .ZN(n7089)
         );
  NAND2_X1 U5204 ( .A1(\x_mult_f[20][0] ), .A2(\x_mult_f[21][0] ), .ZN(n7092)
         );
  NAND2_X1 U5205 ( .A1(\x_mult_f[20][1] ), .A2(\x_mult_f[21][1] ), .ZN(n7090)
         );
  OAI21_X1 U5206 ( .B1(n7089), .B2(n7092), .A(n7090), .ZN(n7597) );
  NAND2_X1 U5207 ( .A1(\x_mult_f[21][2] ), .A2(\x_mult_f[20][2] ), .ZN(n8156)
         );
  NAND2_X1 U5208 ( .A1(\x_mult_f[20][3] ), .A2(\x_mult_f[21][3] ), .ZN(n7599)
         );
  OAI21_X1 U5209 ( .B1(n7598), .B2(n8156), .A(n7599), .ZN(n4606) );
  AOI21_X1 U5210 ( .B1(n4607), .B2(n7597), .A(n4606), .ZN(n4638) );
  NOR2_X1 U5211 ( .A1(\x_mult_f[20][4] ), .A2(\x_mult_f[21][4] ), .ZN(n6946)
         );
  NOR2_X1 U5212 ( .A1(\x_mult_f[20][5] ), .A2(\x_mult_f[21][5] ), .ZN(n7608)
         );
  NOR2_X1 U5213 ( .A1(n6946), .A2(n7608), .ZN(n4640) );
  NOR2_X1 U5214 ( .A1(\x_mult_f[20][6] ), .A2(\x_mult_f[21][6] ), .ZN(n6074)
         );
  NOR2_X1 U5215 ( .A1(\x_mult_f[20][7] ), .A2(\x_mult_f[21][7] ), .ZN(n6076)
         );
  NOR2_X1 U5216 ( .A1(n6074), .A2(n6076), .ZN(n4609) );
  NAND2_X1 U5217 ( .A1(n4640), .A2(n4609), .ZN(n4611) );
  NAND2_X1 U5218 ( .A1(\x_mult_f[20][4] ), .A2(\x_mult_f[21][4] ), .ZN(n7604)
         );
  NAND2_X1 U5219 ( .A1(\x_mult_f[20][5] ), .A2(\x_mult_f[21][5] ), .ZN(n7609)
         );
  OAI21_X1 U5220 ( .B1(n7608), .B2(n7604), .A(n7609), .ZN(n4639) );
  NAND2_X1 U5221 ( .A1(\x_mult_f[20][6] ), .A2(\x_mult_f[21][6] ), .ZN(n6073)
         );
  NAND2_X1 U5222 ( .A1(\x_mult_f[20][7] ), .A2(\x_mult_f[21][7] ), .ZN(n6077)
         );
  OAI21_X1 U5223 ( .B1(n6076), .B2(n6073), .A(n6077), .ZN(n4608) );
  AOI21_X1 U5224 ( .B1(n4609), .B2(n4639), .A(n4608), .ZN(n4610) );
  OAI21_X1 U5225 ( .B1(n4638), .B2(n4611), .A(n4610), .ZN(n6086) );
  OR2_X1 U5226 ( .A1(\x_mult_f[20][8] ), .A2(\x_mult_f[21][8] ), .ZN(n6084) );
  NAND2_X1 U5227 ( .A1(\x_mult_f[20][8] ), .A2(\x_mult_f[21][8] ), .ZN(n6083)
         );
  INV_X1 U5228 ( .A(n6083), .ZN(n4612) );
  AOI21_X1 U5229 ( .B1(n6086), .B2(n6084), .A(n4612), .ZN(n4620) );
  NOR2_X1 U5230 ( .A1(\x_mult_f[20][9] ), .A2(\x_mult_f[21][9] ), .ZN(n4616)
         );
  NAND2_X1 U5231 ( .A1(\x_mult_f[20][9] ), .A2(\x_mult_f[21][9] ), .ZN(n4617)
         );
  OAI21_X1 U5232 ( .B1(n4620), .B2(n4616), .A(n4617), .ZN(n6631) );
  OR2_X1 U5233 ( .A1(\x_mult_f[20][10] ), .A2(\x_mult_f[21][10] ), .ZN(n4628)
         );
  NAND2_X1 U5234 ( .A1(\x_mult_f[20][10] ), .A2(\x_mult_f[21][10] ), .ZN(n4623) );
  NAND2_X1 U5235 ( .A1(n4628), .A2(n4623), .ZN(n4613) );
  XNOR2_X1 U5236 ( .A(n3410), .B(n4613), .ZN(n4614) );
  AOI22_X1 U5237 ( .A1(n7614), .A2(\adder_stage1[10][10] ), .B1(n7919), .B2(
        n4614), .ZN(n4615) );
  INV_X1 U5238 ( .A(n4615), .ZN(n9993) );
  INV_X1 U5239 ( .A(n4616), .ZN(n4618) );
  NAND2_X1 U5240 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  XOR2_X1 U5241 ( .A(n4620), .B(n4619), .Z(n4621) );
  AOI22_X1 U5242 ( .A1(n7614), .A2(\adder_stage1[10][9] ), .B1(n6609), .B2(
        n4621), .ZN(n4622) );
  INV_X1 U5243 ( .A(n4622), .ZN(n9994) );
  INV_X1 U5244 ( .A(n4623), .ZN(n4632) );
  AOI21_X1 U5245 ( .B1(n6631), .B2(n4628), .A(n4632), .ZN(n4625) );
  OR2_X1 U5246 ( .A1(\x_mult_f[20][11] ), .A2(\x_mult_f[21][11] ), .ZN(n4631)
         );
  NAND2_X1 U5247 ( .A1(\x_mult_f[20][11] ), .A2(\x_mult_f[21][11] ), .ZN(n4629) );
  NAND2_X1 U5248 ( .A1(n4631), .A2(n4629), .ZN(n4624) );
  XOR2_X1 U5249 ( .A(n4625), .B(n4624), .Z(n4626) );
  AOI22_X1 U5250 ( .A1(n7614), .A2(\adder_stage1[10][11] ), .B1(n7919), .B2(
        n4626), .ZN(n4627) );
  INV_X1 U5251 ( .A(n4627), .ZN(n9992) );
  AND2_X1 U5252 ( .A1(n4628), .A2(n4631), .ZN(n5147) );
  NAND2_X1 U5253 ( .A1(n6631), .A2(n5147), .ZN(n4633) );
  INV_X1 U5254 ( .A(n4629), .ZN(n4630) );
  AOI21_X1 U5255 ( .B1(n4632), .B2(n4631), .A(n4630), .ZN(n5151) );
  NAND2_X1 U5256 ( .A1(n4633), .A2(n5151), .ZN(n4635) );
  NOR2_X1 U5257 ( .A1(\x_mult_f[20][12] ), .A2(\x_mult_f[21][12] ), .ZN(n5150)
         );
  INV_X1 U5258 ( .A(n5150), .ZN(n5146) );
  NAND2_X1 U5259 ( .A1(\x_mult_f[20][12] ), .A2(\x_mult_f[21][12] ), .ZN(n5149) );
  NAND2_X1 U5260 ( .A1(n5146), .A2(n5149), .ZN(n4634) );
  XNOR2_X1 U5261 ( .A(n4635), .B(n4634), .ZN(n4636) );
  AOI22_X1 U5262 ( .A1(n7614), .A2(\adder_stage1[10][12] ), .B1(n4311), .B2(
        n4636), .ZN(n4637) );
  INV_X1 U5263 ( .A(n4637), .ZN(n9991) );
  INV_X1 U5264 ( .A(n4638), .ZN(n7607) );
  AOI21_X1 U5265 ( .B1(n7607), .B2(n4640), .A(n4639), .ZN(n6075) );
  INV_X1 U5266 ( .A(n6074), .ZN(n4641) );
  NAND2_X1 U5267 ( .A1(n4641), .A2(n6073), .ZN(n4642) );
  XOR2_X1 U5268 ( .A(n6075), .B(n4642), .Z(n4643) );
  AOI22_X1 U5269 ( .A1(n7614), .A2(\adder_stage1[10][6] ), .B1(n8054), .B2(
        n4643), .ZN(n4644) );
  INV_X1 U5270 ( .A(n4644), .ZN(n9997) );
  BUF_X2 U5271 ( .A(n4645), .Z(n8314) );
  INV_X2 U5272 ( .A(n8045), .ZN(n8313) );
  AOI22_X1 U5273 ( .A1(\x_mult_f_int[11][8] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][8] ), .ZN(n4646) );
  INV_X1 U5274 ( .A(n4646), .ZN(n9060) );
  OR2_X1 U5275 ( .A1(\x_mult_f[10][10] ), .A2(\x_mult_f[11][10] ), .ZN(n6325)
         );
  OR2_X1 U5276 ( .A1(\x_mult_f[10][11] ), .A2(\x_mult_f[11][11] ), .ZN(n6327)
         );
  AND2_X1 U5277 ( .A1(n6325), .A2(n6327), .ZN(n8069) );
  NOR2_X1 U5278 ( .A1(\x_mult_f[10][12] ), .A2(\x_mult_f[11][12] ), .ZN(n4661)
         );
  INV_X1 U5279 ( .A(n4661), .ZN(n8074) );
  AND2_X1 U5280 ( .A1(n8069), .A2(n8074), .ZN(n5439) );
  OR2_X1 U5281 ( .A1(\x_mult_f[10][13] ), .A2(\x_mult_f[11][13] ), .ZN(n5441)
         );
  AND2_X1 U5282 ( .A1(n5439), .A2(n5441), .ZN(n4659) );
  NOR2_X1 U5283 ( .A1(n4647), .A2(n4650), .ZN(n4653) );
  OAI21_X1 U5284 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(n4651) );
  AOI21_X1 U5285 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n6379) );
  NOR2_X1 U5286 ( .A1(\x_mult_f[10][4] ), .A2(\x_mult_f[11][4] ), .ZN(n6387)
         );
  NOR2_X1 U5287 ( .A1(\x_mult_f[10][5] ), .A2(\x_mult_f[11][5] ), .ZN(n6389)
         );
  NOR2_X1 U5288 ( .A1(n6387), .A2(n6389), .ZN(n6381) );
  NOR2_X1 U5289 ( .A1(\x_mult_f[10][7] ), .A2(\x_mult_f[11][7] ), .ZN(n6401)
         );
  NOR2_X1 U5290 ( .A1(\x_mult_f[10][6] ), .A2(\x_mult_f[11][6] ), .ZN(n6399)
         );
  NOR2_X1 U5291 ( .A1(n6401), .A2(n6399), .ZN(n4655) );
  NAND2_X1 U5292 ( .A1(n6381), .A2(n4655), .ZN(n4657) );
  NAND2_X1 U5293 ( .A1(\x_mult_f[10][4] ), .A2(\x_mult_f[11][4] ), .ZN(n6849)
         );
  NAND2_X1 U5294 ( .A1(\x_mult_f[10][5] ), .A2(\x_mult_f[11][5] ), .ZN(n6390)
         );
  OAI21_X1 U5295 ( .B1(n6389), .B2(n6849), .A(n6390), .ZN(n6380) );
  NAND2_X1 U5296 ( .A1(\x_mult_f[10][6] ), .A2(\x_mult_f[11][6] ), .ZN(n6398)
         );
  NAND2_X1 U5297 ( .A1(\x_mult_f[10][7] ), .A2(\x_mult_f[11][7] ), .ZN(n6402)
         );
  OAI21_X1 U5298 ( .B1(n6401), .B2(n6398), .A(n6402), .ZN(n4654) );
  AOI21_X1 U5299 ( .B1(n4655), .B2(n6380), .A(n4654), .ZN(n4656) );
  OAI21_X1 U5300 ( .B1(n6379), .B2(n4657), .A(n4656), .ZN(n6341) );
  OR2_X1 U5301 ( .A1(\x_mult_f[10][8] ), .A2(\x_mult_f[11][8] ), .ZN(n6339) );
  NAND2_X1 U5302 ( .A1(\x_mult_f[10][8] ), .A2(\x_mult_f[11][8] ), .ZN(n6338)
         );
  INV_X1 U5303 ( .A(n6338), .ZN(n4658) );
  AOI21_X1 U5304 ( .B1(n6341), .B2(n6339), .A(n4658), .ZN(n6313) );
  NOR2_X1 U5305 ( .A1(\x_mult_f[10][9] ), .A2(\x_mult_f[11][9] ), .ZN(n6309)
         );
  NAND2_X1 U5306 ( .A1(\x_mult_f[10][9] ), .A2(\x_mult_f[11][9] ), .ZN(n6310)
         );
  OAI21_X1 U5307 ( .B1(n6313), .B2(n6309), .A(n6310), .ZN(n8070) );
  NAND2_X1 U5308 ( .A1(n4659), .A2(n8070), .ZN(n4664) );
  NAND2_X1 U5309 ( .A1(\x_mult_f[10][10] ), .A2(\x_mult_f[11][10] ), .ZN(n6320) );
  INV_X1 U5310 ( .A(n6320), .ZN(n6324) );
  NAND2_X1 U5311 ( .A1(\x_mult_f[10][11] ), .A2(\x_mult_f[11][11] ), .ZN(n6326) );
  INV_X1 U5312 ( .A(n6326), .ZN(n4660) );
  AOI21_X1 U5313 ( .B1(n6324), .B2(n6327), .A(n4660), .ZN(n8071) );
  NAND2_X1 U5314 ( .A1(\x_mult_f[10][12] ), .A2(\x_mult_f[11][12] ), .ZN(n8073) );
  OAI21_X1 U5315 ( .B1(n8071), .B2(n4661), .A(n8073), .ZN(n5438) );
  NAND2_X1 U5316 ( .A1(\x_mult_f[10][13] ), .A2(\x_mult_f[11][13] ), .ZN(n5440) );
  INV_X1 U5317 ( .A(n5440), .ZN(n4662) );
  AOI21_X1 U5318 ( .B1(n5438), .B2(n5441), .A(n4662), .ZN(n4663) );
  NAND2_X1 U5319 ( .A1(n4664), .A2(n4663), .ZN(n4884) );
  INV_X1 U5320 ( .A(n4665), .ZN(n4666) );
  AOI22_X1 U5321 ( .A1(n4666), .A2(n8314), .B1(n8313), .B2(
        \adder_stage1[5][20] ), .ZN(n4667) );
  INV_X1 U5322 ( .A(n4667), .ZN(n10071) );
  AOI22_X1 U5323 ( .A1(\x_mult_f_int[11][7] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][7] ), .ZN(n4668) );
  INV_X1 U5324 ( .A(n4668), .ZN(n9061) );
  AOI22_X1 U5325 ( .A1(\x_mult_f_int[11][9] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][9] ), .ZN(n4669) );
  INV_X1 U5326 ( .A(n4669), .ZN(n9059) );
  AOI22_X1 U5327 ( .A1(\x_mult_f_int[11][6] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][6] ), .ZN(n4670) );
  INV_X1 U5328 ( .A(n4670), .ZN(n9062) );
  BUF_X2 U5329 ( .A(n7163), .Z(n4840) );
  INV_X1 U5330 ( .A(n4672), .ZN(n4767) );
  INV_X1 U5331 ( .A(n4673), .ZN(n4765) );
  INV_X1 U5332 ( .A(n4764), .ZN(n4674) );
  AOI21_X1 U5333 ( .B1(n4767), .B2(n4765), .A(n4674), .ZN(n4679) );
  INV_X1 U5334 ( .A(n4675), .ZN(n4677) );
  NAND2_X1 U5335 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  XOR2_X1 U5336 ( .A(n4679), .B(n4678), .Z(n4680) );
  AOI22_X1 U5337 ( .A1(n7669), .A2(\adder_stage2[0][5] ), .B1(n4840), .B2(
        n4680), .ZN(n4681) );
  INV_X1 U5338 ( .A(n4681), .ZN(n9899) );
  AOI21_X1 U5339 ( .B1(n4767), .B2(n4683), .A(n4682), .ZN(n4713) );
  INV_X1 U5340 ( .A(n4712), .ZN(n4684) );
  NAND2_X1 U5341 ( .A1(n4684), .A2(n4711), .ZN(n4685) );
  XOR2_X1 U5342 ( .A(n4713), .B(n4685), .Z(n4686) );
  AOI22_X1 U5343 ( .A1(n8176), .A2(\adder_stage2[0][6] ), .B1(n4840), .B2(
        n4686), .ZN(n4687) );
  INV_X1 U5344 ( .A(n4687), .ZN(n9898) );
  INV_X1 U5345 ( .A(n4688), .ZN(n4708) );
  OAI21_X1 U5346 ( .B1(n4708), .B2(n4689), .A(n4705), .ZN(n4693) );
  NAND2_X1 U5347 ( .A1(n4691), .A2(n4690), .ZN(n4692) );
  XNOR2_X1 U5348 ( .A(n4693), .B(n4692), .ZN(n4694) );
  AOI22_X1 U5349 ( .A1(n7622), .A2(\adder_stage2[0][9] ), .B1(n4840), .B2(
        n4694), .ZN(n4695) );
  INV_X1 U5350 ( .A(n4695), .ZN(n9895) );
  OAI21_X1 U5351 ( .B1(n4708), .B2(n4697), .A(n4696), .ZN(n4702) );
  INV_X1 U5352 ( .A(n4698), .ZN(n4700) );
  NAND2_X1 U5353 ( .A1(n4700), .A2(n4699), .ZN(n4701) );
  XNOR2_X1 U5354 ( .A(n4702), .B(n4701), .ZN(n4703) );
  AOI22_X1 U5355 ( .A1(n8273), .A2(\adder_stage2[0][10] ), .B1(n4840), .B2(
        n4703), .ZN(n4704) );
  INV_X1 U5356 ( .A(n4704), .ZN(n9894) );
  NAND2_X1 U5357 ( .A1(n4706), .A2(n4705), .ZN(n4707) );
  XOR2_X1 U5358 ( .A(n4708), .B(n4707), .Z(n4709) );
  AOI22_X1 U5359 ( .A1(n6877), .A2(\adder_stage2[0][8] ), .B1(n4840), .B2(
        n4709), .ZN(n4710) );
  INV_X1 U5360 ( .A(n4710), .ZN(n9896) );
  OAI21_X1 U5361 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(n4718) );
  INV_X1 U5362 ( .A(n4714), .ZN(n4716) );
  NAND2_X1 U5363 ( .A1(n4716), .A2(n4715), .ZN(n4717) );
  XNOR2_X1 U5364 ( .A(n4718), .B(n4717), .ZN(n4719) );
  AOI22_X1 U5365 ( .A1(n7177), .A2(\adder_stage2[0][7] ), .B1(n4840), .B2(
        n4719), .ZN(n4720) );
  INV_X1 U5366 ( .A(n4720), .ZN(n9897) );
  BUF_X2 U5367 ( .A(n6352), .Z(n8294) );
  AOI22_X1 U5368 ( .A1(\x_mult_f_int[25][7] ), .A2(n8294), .B1(n7864), .B2(
        \x_mult_f[25][7] ), .ZN(n4721) );
  INV_X1 U5369 ( .A(n4721), .ZN(n9238) );
  BUF_X2 U5370 ( .A(n5767), .Z(n6272) );
  AOI22_X1 U5371 ( .A1(n6273), .A2(\x_mult_f[20][4] ), .B1(n6272), .B2(
        \x_mult_f_int[20][4] ), .ZN(n4722) );
  INV_X1 U5372 ( .A(n4722), .ZN(n9179) );
  NOR2_X1 U5373 ( .A1(\adder_stage1[8][1] ), .A2(\adder_stage1[9][1] ), .ZN(
        n4777) );
  INV_X1 U5374 ( .A(n4777), .ZN(n4723) );
  NAND2_X1 U5375 ( .A1(\adder_stage1[8][1] ), .A2(\adder_stage1[9][1] ), .ZN(
        n4775) );
  NAND2_X1 U5376 ( .A1(n4723), .A2(n4775), .ZN(n4724) );
  NAND2_X1 U5377 ( .A1(\adder_stage1[8][0] ), .A2(\adder_stage1[9][0] ), .ZN(
        n4776) );
  XOR2_X1 U5378 ( .A(n4724), .B(n4776), .Z(n4725) );
  AOI22_X1 U5379 ( .A1(n6273), .A2(\adder_stage2[4][1] ), .B1(n6272), .B2(
        n4725), .ZN(n4726) );
  INV_X1 U5380 ( .A(n4726), .ZN(n9835) );
  OR2_X1 U5381 ( .A1(\adder_stage1[8][0] ), .A2(\adder_stage1[9][0] ), .ZN(
        n4727) );
  AND2_X1 U5382 ( .A1(n4727), .A2(n4776), .ZN(n4728) );
  AOI22_X1 U5383 ( .A1(n6273), .A2(\adder_stage2[4][0] ), .B1(n6272), .B2(
        n4728), .ZN(n4729) );
  INV_X1 U5384 ( .A(n4729), .ZN(n9836) );
  BUF_X2 U5385 ( .A(n4645), .Z(n8311) );
  AOI22_X1 U5386 ( .A1(\x_mult_f_int[10][11] ), .A2(n8311), .B1(n8313), .B2(
        \x_mult_f[10][11] ), .ZN(n4730) );
  INV_X1 U5387 ( .A(n4730), .ZN(n9044) );
  AOI22_X1 U5388 ( .A1(\x_mult_f_int[10][8] ), .A2(n8311), .B1(n7640), .B2(
        \x_mult_f[10][8] ), .ZN(n4731) );
  INV_X1 U5389 ( .A(n4731), .ZN(n9047) );
  AOI22_X1 U5390 ( .A1(\x_mult_f_int[10][7] ), .A2(n8311), .B1(n8313), .B2(
        \x_mult_f[10][7] ), .ZN(n4732) );
  INV_X1 U5391 ( .A(n4732), .ZN(n9048) );
  AOI22_X1 U5392 ( .A1(\x_mult_f_int[10][6] ), .A2(n8311), .B1(n8325), .B2(
        \x_mult_f[10][6] ), .ZN(n4733) );
  INV_X1 U5393 ( .A(n4733), .ZN(n9049) );
  AOI22_X1 U5394 ( .A1(\x_mult_f_int[10][9] ), .A2(n8311), .B1(n8330), .B2(
        \x_mult_f[10][9] ), .ZN(n4734) );
  INV_X1 U5395 ( .A(n4734), .ZN(n9046) );
  AOI22_X1 U5396 ( .A1(\x_mult_f_int[10][10] ), .A2(n8311), .B1(n8328), .B2(
        \x_mult_f[10][10] ), .ZN(n4735) );
  INV_X1 U5397 ( .A(n4735), .ZN(n9045) );
  INV_X2 U5398 ( .A(n3408), .ZN(n8398) );
  AOI22_X1 U5399 ( .A1(\x_mult_f_int[26][9] ), .A2(n6626), .B1(n8398), .B2(
        \x_mult_f[26][9] ), .ZN(n4736) );
  INV_X1 U5400 ( .A(n4736), .ZN(n9250) );
  INV_X2 U5401 ( .A(n3408), .ZN(n8401) );
  AOI22_X1 U5402 ( .A1(\x_mult_f_int[26][11] ), .A2(n8235), .B1(n8401), .B2(
        \x_mult_f[26][11] ), .ZN(n4737) );
  INV_X1 U5403 ( .A(n4737), .ZN(n9248) );
  AOI22_X1 U5404 ( .A1(\x_mult_f_int[26][10] ), .A2(n7971), .B1(n8401), .B2(
        \x_mult_f[26][10] ), .ZN(n4738) );
  INV_X1 U5405 ( .A(n4738), .ZN(n9249) );
  INV_X2 U5406 ( .A(n6720), .ZN(n7640) );
  OR2_X1 U5407 ( .A1(\adder_stage1[0][0] ), .A2(\adder_stage1[1][0] ), .ZN(
        n4739) );
  AND2_X1 U5408 ( .A1(n4739), .A2(n4745), .ZN(n4740) );
  AOI22_X1 U5409 ( .A1(n7640), .A2(\adder_stage2[0][0] ), .B1(n4840), .B2(
        n4740), .ZN(n4741) );
  INV_X1 U5410 ( .A(n4741), .ZN(n9904) );
  INV_X1 U5411 ( .A(n4742), .ZN(n4744) );
  NAND2_X1 U5412 ( .A1(n4744), .A2(n4743), .ZN(n4746) );
  XOR2_X1 U5413 ( .A(n4746), .B(n4745), .Z(n4747) );
  AOI22_X1 U5414 ( .A1(n7640), .A2(\adder_stage2[0][1] ), .B1(n4840), .B2(
        n4747), .ZN(n4748) );
  INV_X1 U5415 ( .A(n4748), .ZN(n9903) );
  INV_X1 U5416 ( .A(n4749), .ZN(n4761) );
  OAI21_X1 U5417 ( .B1(n4761), .B2(n4757), .A(n4758), .ZN(n4754) );
  INV_X1 U5418 ( .A(n4750), .ZN(n4752) );
  NAND2_X1 U5419 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  XNOR2_X1 U5420 ( .A(n4754), .B(n4753), .ZN(n4755) );
  AOI22_X1 U5421 ( .A1(n7640), .A2(\adder_stage2[0][3] ), .B1(n4840), .B2(
        n4755), .ZN(n4756) );
  INV_X1 U5422 ( .A(n4756), .ZN(n9901) );
  INV_X1 U5423 ( .A(n4757), .ZN(n4759) );
  NAND2_X1 U5424 ( .A1(n4759), .A2(n4758), .ZN(n4760) );
  XOR2_X1 U5425 ( .A(n4761), .B(n4760), .Z(n4762) );
  AOI22_X1 U5426 ( .A1(n7640), .A2(\adder_stage2[0][2] ), .B1(n4840), .B2(
        n4762), .ZN(n4763) );
  INV_X1 U5427 ( .A(n4763), .ZN(n9902) );
  NAND2_X1 U5428 ( .A1(n4765), .A2(n4764), .ZN(n4766) );
  XNOR2_X1 U5429 ( .A(n4767), .B(n4766), .ZN(n4768) );
  AOI22_X1 U5430 ( .A1(n7640), .A2(\adder_stage2[0][4] ), .B1(n4840), .B2(
        n4768), .ZN(n4769) );
  INV_X1 U5431 ( .A(n4769), .ZN(n9900) );
  INV_X2 U5432 ( .A(n4990), .ZN(n6877) );
  AOI22_X1 U5433 ( .A1(n6877), .A2(\x_mult_f[4][3] ), .B1(n4840), .B2(
        \x_mult_f_int[4][3] ), .ZN(n4770) );
  INV_X1 U5434 ( .A(n4770), .ZN(n8977) );
  AOI22_X1 U5435 ( .A1(\x_mult_f_int[11][10] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][10] ), .ZN(n4772) );
  INV_X1 U5436 ( .A(n4772), .ZN(n9058) );
  AOI22_X1 U5437 ( .A1(\x_mult_f_int[11][11] ), .A2(n8314), .B1(n8427), .B2(
        \x_mult_f[11][11] ), .ZN(n4773) );
  INV_X1 U5438 ( .A(n4773), .ZN(n9057) );
  AOI22_X1 U5439 ( .A1(\x_mult_f_int[11][12] ), .A2(n8314), .B1(n8409), .B2(
        \x_mult_f[11][12] ), .ZN(n4774) );
  INV_X1 U5440 ( .A(n4774), .ZN(n9056) );
  NOR2_X1 U5441 ( .A1(\adder_stage1[8][2] ), .A2(\adder_stage1[9][2] ), .ZN(
        n4832) );
  NOR2_X1 U5442 ( .A1(n4832), .A2(n4800), .ZN(n4779) );
  OAI21_X1 U5443 ( .B1(n4777), .B2(n4776), .A(n4775), .ZN(n4799) );
  NAND2_X1 U5444 ( .A1(\adder_stage1[8][2] ), .A2(\adder_stage1[9][2] ), .ZN(
        n4833) );
  NAND2_X1 U5445 ( .A1(\adder_stage1[8][3] ), .A2(\adder_stage1[9][3] ), .ZN(
        n4801) );
  OAI21_X1 U5446 ( .B1(n4800), .B2(n4833), .A(n4801), .ZN(n4778) );
  INV_X1 U5447 ( .A(n4794), .ZN(n4814) );
  NOR2_X1 U5448 ( .A1(\adder_stage1[8][4] ), .A2(\adder_stage1[9][4] ), .ZN(
        n4783) );
  INV_X1 U5449 ( .A(n4783), .ZN(n4813) );
  NAND2_X1 U5450 ( .A1(\adder_stage1[9][4] ), .A2(\adder_stage1[8][4] ), .ZN(
        n4811) );
  NAND2_X1 U5451 ( .A1(n4813), .A2(n4811), .ZN(n4780) );
  XNOR2_X1 U5452 ( .A(n4814), .B(n4780), .ZN(n4781) );
  AOI22_X1 U5453 ( .A1(n8273), .A2(\adder_stage2[4][4] ), .B1(n6272), .B2(
        n4781), .ZN(n4782) );
  INV_X1 U5454 ( .A(n4782), .ZN(n9832) );
  NOR2_X1 U5455 ( .A1(\adder_stage1[8][5] ), .A2(\adder_stage1[9][5] ), .ZN(
        n4815) );
  NOR2_X1 U5456 ( .A1(n4783), .A2(n4815), .ZN(n4788) );
  NAND2_X1 U5457 ( .A1(\adder_stage1[8][5] ), .A2(\adder_stage1[9][5] ), .ZN(
        n4816) );
  OAI21_X1 U5458 ( .B1(n4815), .B2(n4811), .A(n4816), .ZN(n4790) );
  AOI21_X1 U5459 ( .B1(n4814), .B2(n4788), .A(n4790), .ZN(n4824) );
  NOR2_X1 U5460 ( .A1(\adder_stage1[8][6] ), .A2(\adder_stage1[9][6] ), .ZN(
        n4823) );
  INV_X1 U5461 ( .A(n4823), .ZN(n4784) );
  NAND2_X1 U5462 ( .A1(\adder_stage1[8][6] ), .A2(\adder_stage1[9][6] ), .ZN(
        n4822) );
  NAND2_X1 U5463 ( .A1(n4784), .A2(n4822), .ZN(n4785) );
  XOR2_X1 U5464 ( .A(n4824), .B(n4785), .Z(n4786) );
  AOI22_X1 U5465 ( .A1(n7669), .A2(\adder_stage2[4][6] ), .B1(n6272), .B2(
        n4786), .ZN(n4787) );
  INV_X1 U5466 ( .A(n4787), .ZN(n9830) );
  NOR2_X1 U5467 ( .A1(\adder_stage1[8][7] ), .A2(\adder_stage1[9][7] ), .ZN(
        n4825) );
  NOR2_X1 U5468 ( .A1(n4823), .A2(n4825), .ZN(n4791) );
  NAND2_X1 U5469 ( .A1(n4788), .A2(n4791), .ZN(n4793) );
  NAND2_X1 U5470 ( .A1(\adder_stage1[8][7] ), .A2(\adder_stage1[9][7] ), .ZN(
        n4826) );
  OAI21_X1 U5471 ( .B1(n4825), .B2(n4822), .A(n4826), .ZN(n4789) );
  AOI21_X1 U5472 ( .B1(n4791), .B2(n4790), .A(n4789), .ZN(n4792) );
  OAI21_X1 U5473 ( .B1(n4794), .B2(n4793), .A(n4792), .ZN(n5374) );
  INV_X1 U5474 ( .A(n5374), .ZN(n5997) );
  NOR2_X1 U5475 ( .A1(\adder_stage1[8][8] ), .A2(\adder_stage1[9][8] ), .ZN(
        n4807) );
  NAND2_X1 U5476 ( .A1(\adder_stage1[8][8] ), .A2(\adder_stage1[9][8] ), .ZN(
        n5367) );
  OAI21_X1 U5477 ( .B1(n5997), .B2(n4807), .A(n5367), .ZN(n4796) );
  OR2_X1 U5478 ( .A1(\adder_stage1[8][9] ), .A2(\adder_stage1[9][9] ), .ZN(
        n5371) );
  NAND2_X1 U5479 ( .A1(\adder_stage1[8][9] ), .A2(\adder_stage1[9][9] ), .ZN(
        n5368) );
  NAND2_X1 U5480 ( .A1(n5371), .A2(n5368), .ZN(n4795) );
  XNOR2_X1 U5481 ( .A(n4796), .B(n4795), .ZN(n4797) );
  AOI22_X1 U5482 ( .A1(n8338), .A2(\adder_stage2[4][9] ), .B1(n6272), .B2(
        n4797), .ZN(n4798) );
  INV_X1 U5483 ( .A(n4798), .ZN(n9827) );
  INV_X1 U5484 ( .A(n4799), .ZN(n4836) );
  OAI21_X1 U5485 ( .B1(n4836), .B2(n4832), .A(n4833), .ZN(n4804) );
  INV_X1 U5486 ( .A(n4800), .ZN(n4802) );
  NAND2_X1 U5487 ( .A1(n4802), .A2(n4801), .ZN(n4803) );
  XNOR2_X1 U5488 ( .A(n4804), .B(n4803), .ZN(n4805) );
  AOI22_X1 U5489 ( .A1(n7864), .A2(\adder_stage2[4][3] ), .B1(n6272), .B2(
        n4805), .ZN(n4806) );
  INV_X1 U5490 ( .A(n4806), .ZN(n9833) );
  INV_X1 U5491 ( .A(n4807), .ZN(n5366) );
  NAND2_X1 U5492 ( .A1(n5366), .A2(n5367), .ZN(n4808) );
  XOR2_X1 U5493 ( .A(n5997), .B(n4808), .Z(n4809) );
  AOI22_X1 U5494 ( .A1(n7864), .A2(\adder_stage2[4][8] ), .B1(n6272), .B2(
        n4809), .ZN(n4810) );
  INV_X1 U5495 ( .A(n4810), .ZN(n9828) );
  INV_X1 U5496 ( .A(n4811), .ZN(n4812) );
  AOI21_X1 U5497 ( .B1(n4814), .B2(n4813), .A(n4812), .ZN(n4819) );
  INV_X1 U5498 ( .A(n4815), .ZN(n4817) );
  NAND2_X1 U5499 ( .A1(n4817), .A2(n4816), .ZN(n4818) );
  XOR2_X1 U5500 ( .A(n4819), .B(n4818), .Z(n4820) );
  AOI22_X1 U5501 ( .A1(n8336), .A2(\adder_stage2[4][5] ), .B1(n6272), .B2(
        n4820), .ZN(n4821) );
  INV_X1 U5502 ( .A(n4821), .ZN(n9831) );
  OAI21_X1 U5503 ( .B1(n4824), .B2(n4823), .A(n4822), .ZN(n4829) );
  INV_X1 U5504 ( .A(n4825), .ZN(n4827) );
  NAND2_X1 U5505 ( .A1(n4827), .A2(n4826), .ZN(n4828) );
  XNOR2_X1 U5506 ( .A(n4829), .B(n4828), .ZN(n4830) );
  AOI22_X1 U5507 ( .A1(n8306), .A2(\adder_stage2[4][7] ), .B1(n6272), .B2(
        n4830), .ZN(n4831) );
  INV_X1 U5508 ( .A(n4831), .ZN(n9829) );
  INV_X1 U5509 ( .A(n4832), .ZN(n4834) );
  NAND2_X1 U5510 ( .A1(n4834), .A2(n4833), .ZN(n4835) );
  XOR2_X1 U5511 ( .A(n4836), .B(n4835), .Z(n4837) );
  AOI22_X1 U5512 ( .A1(n8336), .A2(\adder_stage2[4][2] ), .B1(n6272), .B2(
        n4837), .ZN(n4838) );
  INV_X1 U5513 ( .A(n4838), .ZN(n9834) );
  INV_X2 U5514 ( .A(n4990), .ZN(n8245) );
  AOI22_X1 U5515 ( .A1(n8245), .A2(\x_mult_f[4][5] ), .B1(n4840), .B2(
        \x_mult_f_int[4][5] ), .ZN(n4839) );
  INV_X1 U5516 ( .A(n4839), .ZN(n8975) );
  AOI22_X1 U5517 ( .A1(n8245), .A2(\x_mult_f[4][4] ), .B1(n4840), .B2(
        \x_mult_f_int[4][4] ), .ZN(n4841) );
  INV_X1 U5518 ( .A(n4841), .ZN(n8976) );
  BUF_X2 U5519 ( .A(n4894), .Z(n8304) );
  AOI22_X1 U5520 ( .A1(\x_mult_f_int[6][11] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[6][11] ), .ZN(n4842) );
  INV_X1 U5521 ( .A(n4842), .ZN(n8988) );
  NOR2_X1 U5522 ( .A1(n4843), .A2(n4846), .ZN(n7378) );
  NOR2_X1 U5523 ( .A1(\x_mult_f[26][6] ), .A2(\x_mult_f[27][6] ), .ZN(n7387)
         );
  NOR2_X1 U5524 ( .A1(\x_mult_f[26][7] ), .A2(\x_mult_f[27][7] ), .ZN(n7380)
         );
  NOR2_X1 U5525 ( .A1(n7387), .A2(n7380), .ZN(n4848) );
  NAND2_X1 U5526 ( .A1(n7378), .A2(n4848), .ZN(n4850) );
  OAI21_X1 U5527 ( .B1(n4846), .B2(n4845), .A(n4844), .ZN(n7377) );
  NAND2_X1 U5528 ( .A1(\x_mult_f[26][6] ), .A2(\x_mult_f[27][6] ), .ZN(n7388)
         );
  NAND2_X1 U5529 ( .A1(\x_mult_f[26][7] ), .A2(\x_mult_f[27][7] ), .ZN(n7381)
         );
  OAI21_X1 U5530 ( .B1(n7380), .B2(n7388), .A(n7381), .ZN(n4847) );
  AOI21_X1 U5531 ( .B1(n4848), .B2(n7377), .A(n4847), .ZN(n4849) );
  OAI21_X1 U5532 ( .B1(n4851), .B2(n4850), .A(n4849), .ZN(n7425) );
  OR2_X1 U5533 ( .A1(\x_mult_f[26][11] ), .A2(\x_mult_f[27][11] ), .ZN(n7428)
         );
  NAND2_X1 U5534 ( .A1(n7425), .A2(n7428), .ZN(n4858) );
  OR2_X1 U5535 ( .A1(\x_mult_f[26][8] ), .A2(\x_mult_f[27][8] ), .ZN(n7373) );
  OR2_X1 U5536 ( .A1(\x_mult_f[26][9] ), .A2(\x_mult_f[27][9] ), .ZN(n5686) );
  AND2_X1 U5537 ( .A1(n7373), .A2(n5686), .ZN(n7413) );
  OR2_X1 U5538 ( .A1(\x_mult_f[26][10] ), .A2(\x_mult_f[27][10] ), .ZN(n7415)
         );
  NAND2_X1 U5539 ( .A1(n7413), .A2(n7415), .ZN(n7420) );
  NAND2_X1 U5540 ( .A1(\x_mult_f[26][8] ), .A2(\x_mult_f[27][8] ), .ZN(n7372)
         );
  INV_X1 U5541 ( .A(n7372), .ZN(n5684) );
  NAND2_X1 U5542 ( .A1(\x_mult_f[26][9] ), .A2(\x_mult_f[27][9] ), .ZN(n5685)
         );
  INV_X1 U5543 ( .A(n5685), .ZN(n4852) );
  AOI21_X1 U5544 ( .B1(n5684), .B2(n5686), .A(n4852), .ZN(n7423) );
  INV_X1 U5545 ( .A(n7423), .ZN(n4856) );
  INV_X1 U5546 ( .A(n7415), .ZN(n7422) );
  INV_X1 U5547 ( .A(n7428), .ZN(n4853) );
  NOR2_X1 U5548 ( .A1(n7422), .A2(n4853), .ZN(n4855) );
  NAND2_X1 U5549 ( .A1(\x_mult_f[26][10] ), .A2(\x_mult_f[27][10] ), .ZN(n7421) );
  NAND2_X1 U5550 ( .A1(\x_mult_f[26][11] ), .A2(\x_mult_f[27][11] ), .ZN(n7427) );
  OAI21_X1 U5551 ( .B1(n7421), .B2(n4853), .A(n7427), .ZN(n4854) );
  AOI21_X1 U5552 ( .B1(n4856), .B2(n4855), .A(n4854), .ZN(n4857) );
  OAI21_X1 U5553 ( .B1(n4858), .B2(n7420), .A(n4857), .ZN(n8181) );
  OR2_X1 U5554 ( .A1(\x_mult_f[26][12] ), .A2(\x_mult_f[27][12] ), .ZN(n8179)
         );
  NAND2_X1 U5555 ( .A1(\x_mult_f[26][12] ), .A2(\x_mult_f[27][12] ), .ZN(n8178) );
  INV_X1 U5556 ( .A(n8178), .ZN(n4859) );
  AOI21_X1 U5557 ( .B1(n8181), .B2(n8179), .A(n4859), .ZN(n4866) );
  NOR2_X1 U5558 ( .A1(\x_mult_f[26][13] ), .A2(\x_mult_f[27][13] ), .ZN(n4862)
         );
  NAND2_X1 U5559 ( .A1(\x_mult_f[26][13] ), .A2(\x_mult_f[27][13] ), .ZN(n4863) );
  OAI21_X1 U5560 ( .B1(n4866), .B2(n4862), .A(n4863), .ZN(n7766) );
  BUF_X2 U5561 ( .A(n4645), .Z(n7819) );
  AOI22_X1 U5562 ( .A1(n4860), .A2(n7819), .B1(n8176), .B2(
        \adder_stage1[13][14] ), .ZN(n4861) );
  INV_X1 U5563 ( .A(n4861), .ZN(n9938) );
  INV_X1 U5564 ( .A(n4862), .ZN(n4864) );
  NAND2_X1 U5565 ( .A1(n4864), .A2(n4863), .ZN(n4865) );
  XOR2_X1 U5566 ( .A(n4866), .B(n4865), .Z(n4867) );
  AOI22_X1 U5567 ( .A1(n4867), .A2(n7819), .B1(n7669), .B2(
        \adder_stage1[13][13] ), .ZN(n4868) );
  INV_X1 U5568 ( .A(n4868), .ZN(n9939) );
  AOI22_X1 U5569 ( .A1(\x_mult_f_int[27][7] ), .A2(n7819), .B1(n7864), .B2(
        \x_mult_f[27][7] ), .ZN(n4869) );
  INV_X1 U5570 ( .A(n4869), .ZN(n9266) );
  AOI22_X1 U5571 ( .A1(\x_mult_f_int[27][6] ), .A2(n7819), .B1(n7864), .B2(
        \x_mult_f[27][6] ), .ZN(n4870) );
  INV_X1 U5572 ( .A(n4870), .ZN(n9267) );
  INV_X1 U5573 ( .A(n4871), .ZN(n4873) );
  NAND2_X1 U5574 ( .A1(n4873), .A2(n4872), .ZN(n4874) );
  XOR2_X1 U5575 ( .A(n4875), .B(n4874), .Z(n4876) );
  AOI22_X1 U5576 ( .A1(n7074), .A2(\adder_stage4[0][2] ), .B1(n6272), .B2(
        n4876), .ZN(n4877) );
  INV_X1 U5577 ( .A(n4877), .ZN(n9685) );
  INV_X1 U5578 ( .A(n4878), .ZN(n4880) );
  NAND2_X1 U5579 ( .A1(n4880), .A2(n4879), .ZN(n4881) );
  XOR2_X1 U5580 ( .A(n4881), .B(n6089), .Z(n4882) );
  AOI22_X1 U5581 ( .A1(n6854), .A2(\adder_stage4[0][1] ), .B1(n6036), .B2(
        n4882), .ZN(n4883) );
  INV_X1 U5582 ( .A(n4883), .ZN(n9686) );
  FA_X1 U5583 ( .A(\x_mult_f[10][14] ), .B(\x_mult_f[11][14] ), .CI(n4884), 
        .CO(n7701), .S(n4885) );
  AOI22_X1 U5584 ( .A1(n4885), .A2(n7819), .B1(n8313), .B2(
        \adder_stage1[5][14] ), .ZN(n4886) );
  INV_X1 U5585 ( .A(n4886), .ZN(n10072) );
  OAI21_X1 U5586 ( .B1(n4889), .B2(n4888), .A(n4887), .ZN(n8256) );
  OR2_X1 U5587 ( .A1(\adder_stage2[4][16] ), .A2(\adder_stage2[5][16] ), .ZN(
        n8254) );
  NAND2_X1 U5588 ( .A1(\adder_stage2[4][16] ), .A2(\adder_stage2[5][16] ), 
        .ZN(n8253) );
  INV_X1 U5589 ( .A(n8253), .ZN(n5492) );
  AOI21_X1 U5590 ( .B1(n8256), .B2(n8254), .A(n5492), .ZN(n4891) );
  OR2_X1 U5591 ( .A1(\adder_stage2[4][17] ), .A2(\adder_stage2[5][17] ), .ZN(
        n5491) );
  NAND2_X1 U5592 ( .A1(\adder_stage2[4][17] ), .A2(\adder_stage2[5][17] ), 
        .ZN(n5489) );
  NAND2_X1 U5593 ( .A1(n5491), .A2(n5489), .ZN(n4890) );
  XOR2_X1 U5594 ( .A(n4891), .B(n4890), .Z(n4892) );
  AOI22_X1 U5595 ( .A1(n4892), .A2(n8332), .B1(n8306), .B2(
        \adder_stage3[2][17] ), .ZN(n4893) );
  INV_X1 U5596 ( .A(n4893), .ZN(n9712) );
  AOI22_X1 U5597 ( .A1(\x_mult_f_int[6][7] ), .A2(n8334), .B1(n8306), .B2(
        \x_mult_f[6][7] ), .ZN(n4895) );
  INV_X1 U5598 ( .A(n4895), .ZN(n8992) );
  AOI22_X1 U5599 ( .A1(\x_mult_f_int[6][9] ), .A2(n8304), .B1(n8306), .B2(
        \x_mult_f[6][9] ), .ZN(n4896) );
  INV_X1 U5600 ( .A(n4896), .ZN(n8990) );
  AOI22_X1 U5601 ( .A1(\x_mult_f_int[6][8] ), .A2(n8304), .B1(n8306), .B2(
        \x_mult_f[6][8] ), .ZN(n4897) );
  INV_X1 U5602 ( .A(n4897), .ZN(n8991) );
  AOI22_X1 U5603 ( .A1(\x_mult_f_int[7][13] ), .A2(n8332), .B1(n8306), .B2(
        \x_mult_f[7][13] ), .ZN(n4898) );
  INV_X1 U5604 ( .A(n4898), .ZN(n9000) );
  AOI22_X1 U5605 ( .A1(\x_mult_f_int[6][6] ), .A2(n7919), .B1(n8306), .B2(
        \x_mult_f[6][6] ), .ZN(n4899) );
  INV_X1 U5606 ( .A(n4899), .ZN(n8993) );
  AOI22_X1 U5607 ( .A1(\x_mult_f_int[6][10] ), .A2(n8304), .B1(n8306), .B2(
        \x_mult_f[6][10] ), .ZN(n4900) );
  INV_X1 U5608 ( .A(n4900), .ZN(n8989) );
  BUF_X2 U5609 ( .A(n6352), .Z(n8117) );
  OR2_X1 U5610 ( .A1(\adder_stage1[4][0] ), .A2(\adder_stage1[5][0] ), .ZN(
        n4901) );
  AND2_X1 U5611 ( .A1(n4901), .A2(n4923), .ZN(n4902) );
  AOI22_X1 U5612 ( .A1(n8118), .A2(\adder_stage2[2][0] ), .B1(n8117), .B2(
        n4902), .ZN(n4903) );
  INV_X1 U5613 ( .A(n4903), .ZN(n9870) );
  AOI22_X1 U5614 ( .A1(n8118), .A2(\x_mult_f[12][5] ), .B1(n8117), .B2(
        \x_mult_f_int[12][5] ), .ZN(n4904) );
  INV_X1 U5615 ( .A(n4904), .ZN(n9077) );
  INV_X1 U5616 ( .A(n4905), .ZN(n4912) );
  INV_X1 U5617 ( .A(n4911), .ZN(n4906) );
  NAND2_X1 U5618 ( .A1(n4906), .A2(n4910), .ZN(n4907) );
  XOR2_X1 U5619 ( .A(n4912), .B(n4907), .Z(n4908) );
  AOI22_X1 U5620 ( .A1(n8118), .A2(\adder_stage2[2][2] ), .B1(n8117), .B2(
        n4908), .ZN(n4909) );
  INV_X1 U5621 ( .A(n4909), .ZN(n9868) );
  OAI21_X1 U5622 ( .B1(n4912), .B2(n4911), .A(n4910), .ZN(n4917) );
  INV_X1 U5623 ( .A(n4913), .ZN(n4915) );
  NAND2_X1 U5624 ( .A1(n4915), .A2(n4914), .ZN(n4916) );
  XNOR2_X1 U5625 ( .A(n4917), .B(n4916), .ZN(n4918) );
  AOI22_X1 U5626 ( .A1(n8118), .A2(\adder_stage2[2][3] ), .B1(n8117), .B2(
        n4918), .ZN(n4919) );
  INV_X1 U5627 ( .A(n4919), .ZN(n9867) );
  INV_X1 U5628 ( .A(n4920), .ZN(n4922) );
  NAND2_X1 U5629 ( .A1(n4922), .A2(n4921), .ZN(n4924) );
  XOR2_X1 U5630 ( .A(n4924), .B(n4923), .Z(n4925) );
  AOI22_X1 U5631 ( .A1(n8118), .A2(\adder_stage2[2][1] ), .B1(n8117), .B2(
        n4925), .ZN(n4926) );
  INV_X1 U5632 ( .A(n4926), .ZN(n9869) );
  INV_X1 U5633 ( .A(n4927), .ZN(n8110) );
  INV_X1 U5634 ( .A(n4928), .ZN(n8109) );
  NAND2_X1 U5635 ( .A1(n8109), .A2(n8107), .ZN(n4929) );
  XNOR2_X1 U5636 ( .A(n8110), .B(n4929), .ZN(n4930) );
  AOI22_X1 U5637 ( .A1(n8118), .A2(\adder_stage2[2][4] ), .B1(n8117), .B2(
        n4930), .ZN(n4931) );
  INV_X1 U5638 ( .A(n4931), .ZN(n9866) );
  INV_X2 U5639 ( .A(n3407), .ZN(n8309) );
  AOI22_X1 U5640 ( .A1(\x_mult_f_int[8][6] ), .A2(n7507), .B1(n8309), .B2(
        \x_mult_f[8][6] ), .ZN(n4932) );
  INV_X1 U5641 ( .A(n4932), .ZN(n9021) );
  AOI22_X1 U5642 ( .A1(\x_mult_f_int[8][7] ), .A2(n6875), .B1(n8309), .B2(
        \x_mult_f[8][7] ), .ZN(n4933) );
  INV_X1 U5643 ( .A(n4933), .ZN(n9020) );
  INV_X2 U5644 ( .A(n4990), .ZN(n7041) );
  NOR2_X1 U5645 ( .A1(\x_mult_f[6][2] ), .A2(\x_mult_f[7][2] ), .ZN(n4960) );
  NOR2_X1 U5646 ( .A1(\x_mult_f[6][3] ), .A2(\x_mult_f[7][3] ), .ZN(n4943) );
  NOR2_X1 U5647 ( .A1(n4960), .A2(n4943), .ZN(n4935) );
  NOR2_X1 U5648 ( .A1(\x_mult_f[6][1] ), .A2(\x_mult_f[7][1] ), .ZN(n4953) );
  NAND2_X1 U5649 ( .A1(\x_mult_f[7][0] ), .A2(\x_mult_f[6][0] ), .ZN(n4956) );
  NAND2_X1 U5650 ( .A1(\x_mult_f[7][1] ), .A2(\x_mult_f[6][1] ), .ZN(n4954) );
  OAI21_X1 U5651 ( .B1(n4953), .B2(n4956), .A(n4954), .ZN(n4942) );
  NAND2_X1 U5652 ( .A1(\x_mult_f[6][2] ), .A2(\x_mult_f[7][2] ), .ZN(n4961) );
  NAND2_X1 U5653 ( .A1(\x_mult_f[6][3] ), .A2(\x_mult_f[7][3] ), .ZN(n4944) );
  OAI21_X1 U5654 ( .B1(n4943), .B2(n4961), .A(n4944), .ZN(n4934) );
  AOI21_X1 U5655 ( .B1(n4935), .B2(n4942), .A(n4934), .ZN(n5463) );
  INV_X1 U5656 ( .A(n5463), .ZN(n6749) );
  NOR2_X1 U5657 ( .A1(\x_mult_f[6][4] ), .A2(\x_mult_f[7][4] ), .ZN(n5455) );
  INV_X1 U5658 ( .A(n5455), .ZN(n4974) );
  NAND2_X1 U5659 ( .A1(\x_mult_f[6][4] ), .A2(\x_mult_f[7][4] ), .ZN(n5457) );
  INV_X1 U5660 ( .A(n5457), .ZN(n4936) );
  AOI21_X1 U5661 ( .B1(n6749), .B2(n4974), .A(n4936), .ZN(n4939) );
  NOR2_X1 U5662 ( .A1(\x_mult_f[6][5] ), .A2(\x_mult_f[7][5] ), .ZN(n5458) );
  INV_X1 U5663 ( .A(n5458), .ZN(n4937) );
  NAND2_X1 U5664 ( .A1(\x_mult_f[6][5] ), .A2(\x_mult_f[7][5] ), .ZN(n5456) );
  NAND2_X1 U5665 ( .A1(n4937), .A2(n5456), .ZN(n4938) );
  XOR2_X1 U5666 ( .A(n4939), .B(n4938), .Z(n4940) );
  AOI22_X1 U5667 ( .A1(n7041), .A2(\adder_stage1[3][5] ), .B1(n8189), .B2(
        n4940), .ZN(n4941) );
  INV_X1 U5668 ( .A(n4941), .ZN(n10115) );
  INV_X1 U5669 ( .A(n4942), .ZN(n4964) );
  OAI21_X1 U5670 ( .B1(n4964), .B2(n4960), .A(n4961), .ZN(n4947) );
  INV_X1 U5671 ( .A(n4943), .ZN(n4945) );
  NAND2_X1 U5672 ( .A1(n4945), .A2(n4944), .ZN(n4946) );
  XNOR2_X1 U5673 ( .A(n4947), .B(n4946), .ZN(n4948) );
  AOI22_X1 U5674 ( .A1(n7041), .A2(\adder_stage1[3][3] ), .B1(n8189), .B2(
        n4948), .ZN(n4949) );
  INV_X1 U5675 ( .A(n4949), .ZN(n10117) );
  OR2_X1 U5676 ( .A1(\x_mult_f[6][0] ), .A2(\x_mult_f[7][0] ), .ZN(n4950) );
  AND2_X1 U5677 ( .A1(n4950), .A2(n4956), .ZN(n4951) );
  AOI22_X1 U5678 ( .A1(n7041), .A2(\adder_stage1[3][0] ), .B1(n8189), .B2(
        n4951), .ZN(n4952) );
  INV_X1 U5679 ( .A(n4952), .ZN(n10120) );
  INV_X1 U5680 ( .A(n4953), .ZN(n4955) );
  NAND2_X1 U5681 ( .A1(n4955), .A2(n4954), .ZN(n4957) );
  XOR2_X1 U5682 ( .A(n4957), .B(n4956), .Z(n4958) );
  AOI22_X1 U5683 ( .A1(n7041), .A2(\adder_stage1[3][1] ), .B1(n8189), .B2(
        n4958), .ZN(n4959) );
  INV_X1 U5684 ( .A(n4959), .ZN(n10119) );
  INV_X1 U5685 ( .A(n4960), .ZN(n4962) );
  NAND2_X1 U5686 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  XOR2_X1 U5687 ( .A(n4964), .B(n4963), .Z(n4965) );
  AOI22_X1 U5688 ( .A1(n7041), .A2(\adder_stage1[3][2] ), .B1(n8189), .B2(
        n4965), .ZN(n4966) );
  INV_X1 U5689 ( .A(n4966), .ZN(n10118) );
  NOR2_X1 U5690 ( .A1(\adder_stage1[2][2] ), .A2(\adder_stage1[3][2] ), .ZN(
        n7214) );
  NOR2_X1 U5691 ( .A1(\adder_stage1[2][3] ), .A2(\adder_stage1[3][3] ), .ZN(
        n7184) );
  NOR2_X1 U5692 ( .A1(n7214), .A2(n7184), .ZN(n4968) );
  NOR2_X1 U5693 ( .A1(\adder_stage1[2][1] ), .A2(\adder_stage1[3][1] ), .ZN(
        n7232) );
  NAND2_X1 U5694 ( .A1(\adder_stage1[2][1] ), .A2(\adder_stage1[3][1] ), .ZN(
        n7233) );
  OAI21_X1 U5695 ( .B1(n7232), .B2(n7238), .A(n7233), .ZN(n7183) );
  NAND2_X1 U5696 ( .A1(\adder_stage1[2][2] ), .A2(\adder_stage1[3][2] ), .ZN(
        n7215) );
  NAND2_X1 U5697 ( .A1(\adder_stage1[2][3] ), .A2(\adder_stage1[3][3] ), .ZN(
        n7185) );
  OAI21_X1 U5698 ( .B1(n7184), .B2(n7215), .A(n7185), .ZN(n4967) );
  AOI21_X1 U5699 ( .B1(n4968), .B2(n7183), .A(n4967), .ZN(n4986) );
  INV_X1 U5700 ( .A(n4986), .ZN(n7224) );
  NOR2_X1 U5701 ( .A1(\adder_stage1[2][4] ), .A2(\adder_stage1[3][4] ), .ZN(
        n7179) );
  NOR2_X1 U5702 ( .A1(\adder_stage1[2][5] ), .A2(\adder_stage1[3][5] ), .ZN(
        n7225) );
  NOR2_X1 U5703 ( .A1(n7179), .A2(n7225), .ZN(n4978) );
  NAND2_X1 U5704 ( .A1(\adder_stage1[2][4] ), .A2(\adder_stage1[3][4] ), .ZN(
        n7221) );
  NAND2_X1 U5705 ( .A1(\adder_stage1[2][5] ), .A2(\adder_stage1[3][5] ), .ZN(
        n7226) );
  OAI21_X1 U5706 ( .B1(n7225), .B2(n7221), .A(n7226), .ZN(n4982) );
  AOI21_X1 U5707 ( .B1(n7224), .B2(n4978), .A(n4982), .ZN(n7175) );
  NOR2_X1 U5708 ( .A1(\adder_stage1[2][6] ), .A2(\adder_stage1[3][6] ), .ZN(
        n7171) );
  NAND2_X1 U5709 ( .A1(\adder_stage1[2][6] ), .A2(\adder_stage1[3][6] ), .ZN(
        n7172) );
  OAI21_X1 U5710 ( .B1(n7175), .B2(n7171), .A(n7172), .ZN(n4971) );
  NOR2_X1 U5711 ( .A1(\adder_stage1[2][7] ), .A2(\adder_stage1[3][7] ), .ZN(
        n4980) );
  INV_X1 U5712 ( .A(n4980), .ZN(n4969) );
  NAND2_X1 U5713 ( .A1(\adder_stage1[2][7] ), .A2(\adder_stage1[3][7] ), .ZN(
        n4979) );
  NAND2_X1 U5714 ( .A1(n4969), .A2(n4979), .ZN(n4970) );
  XNOR2_X1 U5715 ( .A(n4971), .B(n4970), .ZN(n4972) );
  AOI22_X1 U5716 ( .A1(n7041), .A2(\adder_stage2[1][7] ), .B1(n8189), .B2(
        n4972), .ZN(n4973) );
  INV_X1 U5717 ( .A(n4973), .ZN(n9880) );
  NAND2_X1 U5718 ( .A1(n4974), .A2(n5457), .ZN(n4975) );
  XNOR2_X1 U5719 ( .A(n6749), .B(n4975), .ZN(n4976) );
  AOI22_X1 U5720 ( .A1(n7041), .A2(\adder_stage1[3][4] ), .B1(n8189), .B2(
        n4976), .ZN(n4977) );
  INV_X1 U5721 ( .A(n4977), .ZN(n10116) );
  NOR2_X1 U5722 ( .A1(n7171), .A2(n4980), .ZN(n4983) );
  NAND2_X1 U5723 ( .A1(n4978), .A2(n4983), .ZN(n4985) );
  OAI21_X1 U5724 ( .B1(n4980), .B2(n7172), .A(n4979), .ZN(n4981) );
  AOI21_X1 U5725 ( .B1(n4983), .B2(n4982), .A(n4981), .ZN(n4984) );
  OAI21_X1 U5726 ( .B1(n4986), .B2(n4985), .A(n4984), .ZN(n4995) );
  INV_X1 U5727 ( .A(n4995), .ZN(n5011) );
  NAND2_X1 U5728 ( .A1(n3484), .A2(n3457), .ZN(n5000) );
  NAND2_X1 U5729 ( .A1(\adder_stage1[2][8] ), .A2(\adder_stage1[3][8] ), .ZN(
        n5001) );
  NAND2_X1 U5730 ( .A1(n5000), .A2(n5001), .ZN(n4987) );
  XOR2_X1 U5731 ( .A(n5011), .B(n4987), .Z(n4988) );
  AOI22_X1 U5732 ( .A1(n6877), .A2(\adder_stage2[1][8] ), .B1(n8189), .B2(
        n4988), .ZN(n4989) );
  INV_X1 U5733 ( .A(n4989), .ZN(n9879) );
  INV_X2 U5734 ( .A(n4990), .ZN(n7177) );
  OR2_X1 U5735 ( .A1(\adder_stage1[2][9] ), .A2(\adder_stage1[3][9] ), .ZN(
        n5004) );
  NAND2_X1 U5736 ( .A1(n5004), .A2(n5000), .ZN(n5010) );
  NOR2_X1 U5737 ( .A1(\adder_stage1[2][10] ), .A2(\adder_stage1[3][10] ), .ZN(
        n5012) );
  NOR2_X1 U5738 ( .A1(n5010), .A2(n5012), .ZN(n4994) );
  INV_X1 U5739 ( .A(n5001), .ZN(n4992) );
  NAND2_X1 U5740 ( .A1(\adder_stage1[2][9] ), .A2(\adder_stage1[3][9] ), .ZN(
        n5003) );
  INV_X1 U5741 ( .A(n5003), .ZN(n4991) );
  AOI21_X1 U5742 ( .B1(n5004), .B2(n4992), .A(n4991), .ZN(n5009) );
  NAND2_X1 U5743 ( .A1(\adder_stage1[2][10] ), .A2(\adder_stage1[3][10] ), 
        .ZN(n5013) );
  OAI21_X1 U5744 ( .B1(n5009), .B2(n5012), .A(n5013), .ZN(n4993) );
  AOI21_X1 U5745 ( .B1(n4995), .B2(n4994), .A(n4993), .ZN(n6284) );
  NOR2_X1 U5746 ( .A1(\adder_stage1[2][11] ), .A2(\adder_stage1[3][11] ), .ZN(
        n6283) );
  INV_X1 U5747 ( .A(n6283), .ZN(n4996) );
  NAND2_X1 U5748 ( .A1(\adder_stage1[2][11] ), .A2(\adder_stage1[3][11] ), 
        .ZN(n6282) );
  NAND2_X1 U5749 ( .A1(n4996), .A2(n6282), .ZN(n4997) );
  XOR2_X1 U5750 ( .A(n6284), .B(n4997), .Z(n4998) );
  AOI22_X1 U5751 ( .A1(n7177), .A2(\adder_stage2[1][11] ), .B1(n8189), .B2(
        n4998), .ZN(n4999) );
  INV_X1 U5752 ( .A(n4999), .ZN(n9876) );
  INV_X1 U5753 ( .A(n5000), .ZN(n5002) );
  OAI21_X1 U5754 ( .B1(n5011), .B2(n5002), .A(n5001), .ZN(n5006) );
  NAND2_X1 U5755 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  XNOR2_X1 U5756 ( .A(n5006), .B(n5005), .ZN(n5007) );
  AOI22_X1 U5757 ( .A1(n8245), .A2(\adder_stage2[1][9] ), .B1(n8189), .B2(
        n5007), .ZN(n5008) );
  INV_X1 U5758 ( .A(n5008), .ZN(n9878) );
  OAI21_X1 U5759 ( .B1(n5011), .B2(n5010), .A(n5009), .ZN(n5016) );
  INV_X1 U5760 ( .A(n5012), .ZN(n5014) );
  NAND2_X1 U5761 ( .A1(n5014), .A2(n5013), .ZN(n5015) );
  XNOR2_X1 U5762 ( .A(n5016), .B(n5015), .ZN(n5017) );
  AOI22_X1 U5763 ( .A1(n7177), .A2(\adder_stage2[1][10] ), .B1(n8189), .B2(
        n5017), .ZN(n5018) );
  INV_X1 U5764 ( .A(n5018), .ZN(n9877) );
  NOR2_X1 U5765 ( .A1(\adder_stage2[6][2] ), .A2(\adder_stage2[7][2] ), .ZN(
        n7080) );
  NOR2_X1 U5766 ( .A1(\adder_stage2[6][3] ), .A2(\adder_stage2[7][3] ), .ZN(
        n7082) );
  NOR2_X1 U5767 ( .A1(n7080), .A2(n7082), .ZN(n5020) );
  NOR2_X1 U5768 ( .A1(\adder_stage2[6][1] ), .A2(\adder_stage2[7][1] ), .ZN(
        n6135) );
  NAND2_X1 U5769 ( .A1(\adder_stage2[6][0] ), .A2(\adder_stage2[7][0] ), .ZN(
        n6178) );
  NAND2_X1 U5770 ( .A1(\adder_stage2[6][1] ), .A2(\adder_stage2[7][1] ), .ZN(
        n6136) );
  OAI21_X1 U5771 ( .B1(n6135), .B2(n6178), .A(n6136), .ZN(n6130) );
  NAND2_X1 U5772 ( .A1(\adder_stage2[6][2] ), .A2(\adder_stage2[7][2] ), .ZN(
        n7079) );
  NAND2_X1 U5773 ( .A1(\adder_stage2[6][3] ), .A2(\adder_stage2[7][3] ), .ZN(
        n7083) );
  OAI21_X1 U5774 ( .B1(n7082), .B2(n7079), .A(n7083), .ZN(n5019) );
  AOI21_X1 U5775 ( .B1(n5020), .B2(n6130), .A(n5019), .ZN(n7100) );
  NOR2_X1 U5776 ( .A1(\adder_stage2[6][4] ), .A2(\adder_stage2[7][4] ), .ZN(
        n7101) );
  NOR2_X1 U5777 ( .A1(\adder_stage2[6][5] ), .A2(\adder_stage2[7][5] ), .ZN(
        n7103) );
  NOR2_X1 U5778 ( .A1(n7101), .A2(n7103), .ZN(n7252) );
  NOR2_X1 U5779 ( .A1(\adder_stage2[6][6] ), .A2(\adder_stage2[7][6] ), .ZN(
        n7268) );
  NOR2_X1 U5780 ( .A1(\adder_stage2[6][7] ), .A2(\adder_stage2[7][7] ), .ZN(
        n7270) );
  NOR2_X1 U5781 ( .A1(n7268), .A2(n7270), .ZN(n5022) );
  NAND2_X1 U5782 ( .A1(n7252), .A2(n5022), .ZN(n5024) );
  NAND2_X1 U5783 ( .A1(\adder_stage2[6][4] ), .A2(\adder_stage2[7][4] ), .ZN(
        n7118) );
  NAND2_X1 U5784 ( .A1(\adder_stage2[6][5] ), .A2(\adder_stage2[7][5] ), .ZN(
        n7104) );
  OAI21_X1 U5785 ( .B1(n7103), .B2(n7118), .A(n7104), .ZN(n7251) );
  NAND2_X1 U5786 ( .A1(\adder_stage2[6][6] ), .A2(\adder_stage2[7][6] ), .ZN(
        n7267) );
  NAND2_X1 U5787 ( .A1(\adder_stage2[6][7] ), .A2(\adder_stage2[7][7] ), .ZN(
        n7271) );
  OAI21_X1 U5788 ( .B1(n7270), .B2(n7267), .A(n7271), .ZN(n5021) );
  AOI21_X1 U5789 ( .B1(n5022), .B2(n7251), .A(n5021), .ZN(n5023) );
  OAI21_X1 U5790 ( .B1(n7100), .B2(n5024), .A(n5023), .ZN(n6487) );
  NOR2_X1 U5791 ( .A1(\adder_stage2[6][8] ), .A2(\adder_stage2[7][8] ), .ZN(
        n8099) );
  NOR2_X1 U5792 ( .A1(\adder_stage2[6][9] ), .A2(\adder_stage2[7][9] ), .ZN(
        n7279) );
  NOR2_X1 U5793 ( .A1(n8099), .A2(n7279), .ZN(n6488) );
  NOR2_X1 U5794 ( .A1(\adder_stage2[6][10] ), .A2(\adder_stage2[7][10] ), .ZN(
        n6492) );
  NOR2_X1 U5795 ( .A1(\adder_stage2[6][11] ), .A2(\adder_stage2[7][11] ), .ZN(
        n6494) );
  NOR2_X1 U5796 ( .A1(n6492), .A2(n6494), .ZN(n5026) );
  NAND2_X1 U5797 ( .A1(n6488), .A2(n5026), .ZN(n7259) );
  NOR2_X1 U5798 ( .A1(\adder_stage2[6][12] ), .A2(\adder_stage2[7][12] ), .ZN(
        n7260) );
  NOR2_X1 U5799 ( .A1(n7259), .A2(n7260), .ZN(n6466) );
  OR2_X1 U5800 ( .A1(\adder_stage2[6][13] ), .A2(\adder_stage2[7][13] ), .ZN(
        n6471) );
  NAND3_X1 U5801 ( .A1(n6487), .A2(n6466), .A3(n6471), .ZN(n5029) );
  NAND2_X1 U5802 ( .A1(\adder_stage2[6][8] ), .A2(\adder_stage2[7][8] ), .ZN(
        n8100) );
  NAND2_X1 U5803 ( .A1(\adder_stage2[6][9] ), .A2(\adder_stage2[7][9] ), .ZN(
        n7280) );
  OAI21_X1 U5804 ( .B1(n7279), .B2(n8100), .A(n7280), .ZN(n6489) );
  NAND2_X1 U5805 ( .A1(\adder_stage2[6][10] ), .A2(\adder_stage2[7][10] ), 
        .ZN(n6921) );
  NAND2_X1 U5806 ( .A1(\adder_stage2[6][11] ), .A2(\adder_stage2[7][11] ), 
        .ZN(n6495) );
  OAI21_X1 U5807 ( .B1(n6494), .B2(n6921), .A(n6495), .ZN(n5025) );
  AOI21_X1 U5808 ( .B1(n5026), .B2(n6489), .A(n5025), .ZN(n7258) );
  NAND2_X1 U5809 ( .A1(\adder_stage2[6][12] ), .A2(\adder_stage2[7][12] ), 
        .ZN(n7261) );
  OAI21_X1 U5810 ( .B1(n7258), .B2(n7260), .A(n7261), .ZN(n6467) );
  NAND2_X1 U5811 ( .A1(\adder_stage2[6][13] ), .A2(\adder_stage2[7][13] ), 
        .ZN(n6470) );
  INV_X1 U5812 ( .A(n6470), .ZN(n5027) );
  AOI21_X1 U5813 ( .B1(n6467), .B2(n6471), .A(n5027), .ZN(n5028) );
  NAND2_X1 U5814 ( .A1(n5029), .A2(n5028), .ZN(n6939) );
  OR2_X1 U5815 ( .A1(\adder_stage2[6][14] ), .A2(\adder_stage2[7][14] ), .ZN(
        n6937) );
  NAND2_X1 U5816 ( .A1(\adder_stage2[6][14] ), .A2(\adder_stage2[7][14] ), 
        .ZN(n6936) );
  INV_X1 U5817 ( .A(n6936), .ZN(n5030) );
  AOI21_X1 U5818 ( .B1(n6939), .B2(n6937), .A(n5030), .ZN(n6484) );
  NOR2_X1 U5819 ( .A1(\adder_stage2[6][15] ), .A2(\adder_stage2[7][15] ), .ZN(
        n6480) );
  NAND2_X1 U5820 ( .A1(\adder_stage2[6][15] ), .A2(\adder_stage2[7][15] ), 
        .ZN(n6481) );
  OAI21_X1 U5821 ( .B1(n6484), .B2(n6480), .A(n6481), .ZN(n8263) );
  OR2_X1 U5822 ( .A1(\adder_stage2[6][16] ), .A2(\adder_stage2[7][16] ), .ZN(
        n8261) );
  OR2_X1 U5823 ( .A1(\adder_stage2[6][17] ), .A2(\adder_stage2[7][17] ), .ZN(
        n5069) );
  AND2_X1 U5824 ( .A1(n8261), .A2(n5069), .ZN(n5074) );
  NOR2_X1 U5825 ( .A1(\adder_stage2[6][18] ), .A2(\adder_stage2[7][18] ), .ZN(
        n5032) );
  INV_X1 U5826 ( .A(n5032), .ZN(n5078) );
  AND2_X1 U5827 ( .A1(n5074), .A2(n5078), .ZN(n7753) );
  NAND2_X1 U5828 ( .A1(\adder_stage2[6][16] ), .A2(\adder_stage2[7][16] ), 
        .ZN(n8260) );
  INV_X1 U5829 ( .A(n8260), .ZN(n5067) );
  NAND2_X1 U5830 ( .A1(\adder_stage2[6][17] ), .A2(\adder_stage2[7][17] ), 
        .ZN(n5068) );
  INV_X1 U5831 ( .A(n5068), .ZN(n5031) );
  AOI21_X1 U5832 ( .B1(n5067), .B2(n5069), .A(n5031), .ZN(n5075) );
  NAND2_X1 U5833 ( .A1(\adder_stage2[6][18] ), .A2(\adder_stage2[7][18] ), 
        .ZN(n5077) );
  OAI21_X1 U5834 ( .B1(n5075), .B2(n5032), .A(n5077), .ZN(n7758) );
  AOI21_X1 U5835 ( .B1(n8263), .B2(n7753), .A(n7758), .ZN(n5034) );
  OR2_X1 U5836 ( .A1(\adder_stage2[6][19] ), .A2(\adder_stage2[7][19] ), .ZN(
        n7757) );
  NAND2_X1 U5837 ( .A1(\adder_stage2[6][19] ), .A2(\adder_stage2[7][19] ), 
        .ZN(n7755) );
  NAND2_X1 U5838 ( .A1(n7757), .A2(n7755), .ZN(n5033) );
  XOR2_X1 U5839 ( .A(n5034), .B(n5033), .Z(n5035) );
  BUF_X2 U5840 ( .A(n6352), .Z(n7962) );
  AOI22_X1 U5841 ( .A1(n5035), .A2(n7962), .B1(n7972), .B2(
        \adder_stage3[3][19] ), .ZN(n5036) );
  INV_X1 U5842 ( .A(n5036), .ZN(n9689) );
  BUF_X2 U5843 ( .A(n6352), .Z(n8301) );
  AOI22_X1 U5844 ( .A1(\x_mult_f_int[2][11] ), .A2(n8301), .B1(n8340), .B2(
        \x_mult_f[2][11] ), .ZN(n5037) );
  INV_X1 U5845 ( .A(n5037), .ZN(n8945) );
  INV_X2 U5846 ( .A(n3445), .ZN(n8434) );
  AOI22_X1 U5847 ( .A1(\x_mult_f_int[2][6] ), .A2(n8301), .B1(n8434), .B2(
        \x_mult_f[2][6] ), .ZN(n5038) );
  INV_X1 U5848 ( .A(n5038), .ZN(n8950) );
  AOI22_X1 U5849 ( .A1(\x_mult_f_int[2][10] ), .A2(n8301), .B1(n8434), .B2(
        \x_mult_f[2][10] ), .ZN(n5039) );
  INV_X1 U5850 ( .A(n5039), .ZN(n8946) );
  AOI22_X1 U5851 ( .A1(\x_mult_f_int[2][7] ), .A2(n8301), .B1(n8434), .B2(
        \x_mult_f[2][7] ), .ZN(n5040) );
  INV_X1 U5852 ( .A(n5040), .ZN(n8949) );
  AOI22_X1 U5853 ( .A1(\x_mult_f_int[2][9] ), .A2(n8301), .B1(n8434), .B2(
        \x_mult_f[2][9] ), .ZN(n5041) );
  INV_X1 U5854 ( .A(n5041), .ZN(n8947) );
  AOI22_X1 U5855 ( .A1(\x_mult_f_int[2][8] ), .A2(n8301), .B1(n8434), .B2(
        \x_mult_f[2][8] ), .ZN(n5042) );
  INV_X1 U5856 ( .A(n5042), .ZN(n8948) );
  AOI21_X1 U5857 ( .B1(n8110), .B2(n5044), .A(n5043), .ZN(n5051) );
  INV_X1 U5858 ( .A(n5050), .ZN(n5045) );
  NAND2_X1 U5859 ( .A1(n5045), .A2(n5049), .ZN(n5046) );
  XOR2_X1 U5860 ( .A(n5051), .B(n5046), .Z(n5047) );
  AOI22_X1 U5861 ( .A1(n7074), .A2(\adder_stage2[2][6] ), .B1(n8117), .B2(
        n5047), .ZN(n5048) );
  INV_X1 U5862 ( .A(n5048), .ZN(n9864) );
  OAI21_X1 U5863 ( .B1(n5051), .B2(n5050), .A(n5049), .ZN(n5056) );
  INV_X1 U5864 ( .A(n5052), .ZN(n5054) );
  NAND2_X1 U5865 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  XNOR2_X1 U5866 ( .A(n5056), .B(n5055), .ZN(n5057) );
  AOI22_X1 U5867 ( .A1(n7074), .A2(\adder_stage2[2][7] ), .B1(n8117), .B2(
        n5057), .ZN(n5058) );
  INV_X1 U5868 ( .A(n5058), .ZN(n9863) );
  OAI21_X1 U5869 ( .B1(n7049), .B2(n5059), .A(n7046), .ZN(n5063) );
  NAND2_X1 U5870 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  XNOR2_X1 U5871 ( .A(n5063), .B(n5062), .ZN(n5064) );
  AOI22_X1 U5872 ( .A1(n7074), .A2(\adder_stage2[2][12] ), .B1(n8117), .B2(
        n5064), .ZN(n5065) );
  INV_X1 U5873 ( .A(n5065), .ZN(n9858) );
  AOI22_X1 U5874 ( .A1(\x_mult_f_int[8][12] ), .A2(n7962), .B1(n8323), .B2(
        \x_mult_f[8][12] ), .ZN(n5066) );
  INV_X1 U5875 ( .A(n5066), .ZN(n9015) );
  AOI21_X1 U5876 ( .B1(n8263), .B2(n8261), .A(n5067), .ZN(n5071) );
  NAND2_X1 U5877 ( .A1(n5069), .A2(n5068), .ZN(n5070) );
  XOR2_X1 U5878 ( .A(n5071), .B(n5070), .Z(n5072) );
  AOI22_X1 U5879 ( .A1(n5072), .A2(n7962), .B1(n8434), .B2(
        \adder_stage3[3][17] ), .ZN(n5073) );
  INV_X1 U5880 ( .A(n5073), .ZN(n9691) );
  NAND2_X1 U5881 ( .A1(n8263), .A2(n5074), .ZN(n5076) );
  NAND2_X1 U5882 ( .A1(n5076), .A2(n5075), .ZN(n5080) );
  NAND2_X1 U5883 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  XNOR2_X1 U5884 ( .A(n5080), .B(n5079), .ZN(n5081) );
  AOI22_X1 U5885 ( .A1(n5081), .A2(n7962), .B1(n8434), .B2(
        \adder_stage3[3][18] ), .ZN(n5082) );
  INV_X1 U5886 ( .A(n5082), .ZN(n9690) );
  BUF_X2 U5887 ( .A(n6352), .Z(n7155) );
  NAND2_X1 U5888 ( .A1(n5087), .A2(n5086), .ZN(n5088) );
  XNOR2_X1 U5889 ( .A(n5089), .B(n5088), .ZN(n5090) );
  AOI22_X1 U5890 ( .A1(n8057), .A2(\adder_stage1[6][12] ), .B1(n7155), .B2(
        n5090), .ZN(n5091) );
  INV_X1 U5891 ( .A(n5091), .ZN(n10058) );
  NAND2_X1 U5892 ( .A1(n5097), .A2(n5092), .ZN(n5093) );
  XNOR2_X1 U5893 ( .A(n5098), .B(n5093), .ZN(n5094) );
  AOI22_X1 U5894 ( .A1(n8088), .A2(\adder_stage1[6][10] ), .B1(n7155), .B2(
        n5094), .ZN(n5095) );
  INV_X1 U5895 ( .A(n5095), .ZN(n10060) );
  NAND2_X1 U5896 ( .A1(n3506), .A2(n5100), .ZN(n5101) );
  XOR2_X1 U5897 ( .A(n5102), .B(n5101), .Z(n5103) );
  AOI22_X1 U5898 ( .A1(n8336), .A2(\adder_stage1[6][11] ), .B1(n7155), .B2(
        n5103), .ZN(n5104) );
  INV_X1 U5899 ( .A(n5104), .ZN(n10059) );
  AOI22_X1 U5900 ( .A1(\x_mult_f_int[12][6] ), .A2(n6272), .B1(n7855), .B2(
        \x_mult_f[12][6] ), .ZN(n5105) );
  INV_X1 U5901 ( .A(n5105), .ZN(n9076) );
  AOI22_X1 U5902 ( .A1(\x_mult_f_int[12][7] ), .A2(n6609), .B1(n7855), .B2(
        \x_mult_f[12][7] ), .ZN(n5106) );
  INV_X1 U5903 ( .A(n5106), .ZN(n9075) );
  OR2_X1 U5904 ( .A1(\x_mult_f[2][11] ), .A2(\x_mult_f[3][11] ), .ZN(n7941) );
  NAND2_X1 U5905 ( .A1(n7938), .A2(n7941), .ZN(n5114) );
  NAND2_X1 U5906 ( .A1(n5107), .A2(n5108), .ZN(n7933) );
  INV_X1 U5907 ( .A(n7936), .ZN(n5112) );
  INV_X1 U5908 ( .A(n5108), .ZN(n7935) );
  INV_X1 U5909 ( .A(n7941), .ZN(n5109) );
  NOR2_X1 U5910 ( .A1(n7935), .A2(n5109), .ZN(n5111) );
  NAND2_X1 U5911 ( .A1(\x_mult_f[2][11] ), .A2(\x_mult_f[3][11] ), .ZN(n7940)
         );
  OAI21_X1 U5912 ( .B1(n7934), .B2(n5109), .A(n7940), .ZN(n5110) );
  AOI21_X1 U5913 ( .B1(n5112), .B2(n5111), .A(n5110), .ZN(n5113) );
  OAI21_X1 U5914 ( .B1(n5114), .B2(n7933), .A(n5113), .ZN(n8052) );
  OR2_X1 U5915 ( .A1(\x_mult_f[2][12] ), .A2(\x_mult_f[3][12] ), .ZN(n8050) );
  NAND2_X1 U5916 ( .A1(\x_mult_f[2][12] ), .A2(\x_mult_f[3][12] ), .ZN(n8049)
         );
  INV_X1 U5917 ( .A(n8049), .ZN(n5115) );
  AOI21_X1 U5918 ( .B1(n8052), .B2(n8050), .A(n5115), .ZN(n5516) );
  NOR2_X1 U5919 ( .A1(\x_mult_f[2][13] ), .A2(\x_mult_f[3][13] ), .ZN(n5515)
         );
  INV_X1 U5920 ( .A(n5515), .ZN(n5116) );
  NAND2_X1 U5921 ( .A1(\x_mult_f[2][13] ), .A2(\x_mult_f[3][13] ), .ZN(n5514)
         );
  NAND2_X1 U5922 ( .A1(n5116), .A2(n5514), .ZN(n5117) );
  XOR2_X1 U5923 ( .A(n5516), .B(n5117), .Z(n5118) );
  INV_X2 U5924 ( .A(n3408), .ZN(n8319) );
  AOI22_X1 U5925 ( .A1(n5118), .A2(n7962), .B1(n8319), .B2(
        \adder_stage1[1][13] ), .ZN(n5119) );
  INV_X1 U5926 ( .A(n5119), .ZN(n10139) );
  AOI22_X1 U5927 ( .A1(\x_mult_f_int[3][6] ), .A2(n7962), .B1(n8319), .B2(
        \x_mult_f[3][6] ), .ZN(n5120) );
  INV_X1 U5928 ( .A(n5120), .ZN(n8964) );
  AOI22_X1 U5929 ( .A1(\x_mult_f_int[26][6] ), .A2(n8251), .B1(n8398), .B2(
        \x_mult_f[26][6] ), .ZN(n5121) );
  INV_X1 U5930 ( .A(n5121), .ZN(n9253) );
  AOI22_X1 U5931 ( .A1(\x_mult_f_int[26][8] ), .A2(n8216), .B1(n8398), .B2(
        \x_mult_f[26][8] ), .ZN(n5122) );
  INV_X1 U5932 ( .A(n5122), .ZN(n9251) );
  AOI22_X1 U5933 ( .A1(\x_mult_f_int[26][7] ), .A2(n8265), .B1(n8398), .B2(
        \x_mult_f[26][7] ), .ZN(n5123) );
  INV_X1 U5934 ( .A(n5123), .ZN(n9252) );
  BUF_X1 U5935 ( .A(n5124), .Z(n5384) );
  AOI22_X1 U5936 ( .A1(\x_mult_f_int[17][11] ), .A2(n7507), .B1(n8296), .B2(
        \x_mult_f[17][11] ), .ZN(n5125) );
  INV_X1 U5937 ( .A(n5125), .ZN(n9130) );
  AOI22_X1 U5938 ( .A1(\x_mult_f_int[17][8] ), .A2(n8024), .B1(n8325), .B2(
        \x_mult_f[17][8] ), .ZN(n5126) );
  INV_X1 U5939 ( .A(n5126), .ZN(n9133) );
  AOI22_X1 U5940 ( .A1(\x_mult_f_int[17][9] ), .A2(n8189), .B1(n8330), .B2(
        \x_mult_f[17][9] ), .ZN(n5127) );
  INV_X1 U5941 ( .A(n5127), .ZN(n9132) );
  AOI22_X1 U5942 ( .A1(\x_mult_f_int[17][6] ), .A2(n8301), .B1(n8328), .B2(
        \x_mult_f[17][6] ), .ZN(n5128) );
  INV_X1 U5943 ( .A(n5128), .ZN(n9135) );
  AOI22_X1 U5944 ( .A1(\x_mult_f_int[17][10] ), .A2(n4257), .B1(n8313), .B2(
        \x_mult_f[17][10] ), .ZN(n5129) );
  INV_X1 U5945 ( .A(n5129), .ZN(n9131) );
  AOI22_X1 U5946 ( .A1(\x_mult_f_int[17][7] ), .A2(n6036), .B1(n8434), .B2(
        \x_mult_f[17][7] ), .ZN(n5130) );
  INV_X1 U5947 ( .A(n5130), .ZN(n9134) );
  OR2_X1 U5948 ( .A1(\x_mult_f[22][8] ), .A2(\x_mult_f[23][8] ), .ZN(n7111) );
  OR2_X1 U5949 ( .A1(\x_mult_f[22][9] ), .A2(\x_mult_f[23][9] ), .ZN(n7113) );
  AND2_X1 U5950 ( .A1(n7111), .A2(n7113), .ZN(n6907) );
  OR2_X1 U5951 ( .A1(\x_mult_f[22][10] ), .A2(\x_mult_f[23][10] ), .ZN(n6911)
         );
  AND2_X1 U5952 ( .A1(n6907), .A2(n6911), .ZN(n5140) );
  NOR2_X1 U5953 ( .A1(\x_mult_f[22][2] ), .A2(\x_mult_f[23][2] ), .ZN(n6639)
         );
  NOR2_X1 U5954 ( .A1(\x_mult_f[22][3] ), .A2(\x_mult_f[23][3] ), .ZN(n6258)
         );
  NOR2_X1 U5955 ( .A1(n6639), .A2(n6258), .ZN(n5132) );
  NOR2_X1 U5956 ( .A1(\x_mult_f[22][1] ), .A2(\x_mult_f[23][1] ), .ZN(n6332)
         );
  NAND2_X1 U5957 ( .A1(\x_mult_f[22][0] ), .A2(\x_mult_f[23][0] ), .ZN(n7803)
         );
  NAND2_X1 U5958 ( .A1(\x_mult_f[22][1] ), .A2(\x_mult_f[23][1] ), .ZN(n6333)
         );
  OAI21_X1 U5959 ( .B1(n6332), .B2(n7803), .A(n6333), .ZN(n6257) );
  NAND2_X1 U5960 ( .A1(\x_mult_f[22][2] ), .A2(\x_mult_f[23][2] ), .ZN(n6640)
         );
  NAND2_X1 U5961 ( .A1(\x_mult_f[22][3] ), .A2(\x_mult_f[23][3] ), .ZN(n6259)
         );
  OAI21_X1 U5962 ( .B1(n6258), .B2(n6640), .A(n6259), .ZN(n5131) );
  AOI21_X1 U5963 ( .B1(n5132), .B2(n6257), .A(n5131), .ZN(n6527) );
  NOR2_X1 U5964 ( .A1(\x_mult_f[22][4] ), .A2(\x_mult_f[23][4] ), .ZN(n6528)
         );
  NOR2_X1 U5965 ( .A1(\x_mult_f[22][5] ), .A2(\x_mult_f[23][5] ), .ZN(n6530)
         );
  NOR2_X1 U5966 ( .A1(n6528), .A2(n6530), .ZN(n6559) );
  NOR2_X1 U5967 ( .A1(\x_mult_f[22][6] ), .A2(\x_mult_f[23][6] ), .ZN(n6900)
         );
  NOR2_X1 U5968 ( .A1(\x_mult_f[22][7] ), .A2(\x_mult_f[23][7] ), .ZN(n6560)
         );
  NOR2_X1 U5969 ( .A1(n6900), .A2(n6560), .ZN(n5134) );
  NAND2_X1 U5970 ( .A1(n6559), .A2(n5134), .ZN(n5136) );
  NAND2_X1 U5971 ( .A1(\x_mult_f[22][4] ), .A2(\x_mult_f[23][4] ), .ZN(n8162)
         );
  NAND2_X1 U5972 ( .A1(\x_mult_f[22][5] ), .A2(\x_mult_f[23][5] ), .ZN(n6531)
         );
  OAI21_X1 U5973 ( .B1(n6530), .B2(n8162), .A(n6531), .ZN(n6558) );
  NAND2_X1 U5974 ( .A1(\x_mult_f[22][6] ), .A2(\x_mult_f[23][6] ), .ZN(n6901)
         );
  NAND2_X1 U5975 ( .A1(\x_mult_f[22][7] ), .A2(\x_mult_f[23][7] ), .ZN(n6561)
         );
  OAI21_X1 U5976 ( .B1(n6560), .B2(n6901), .A(n6561), .ZN(n5133) );
  AOI21_X1 U5977 ( .B1(n5134), .B2(n6558), .A(n5133), .ZN(n5135) );
  OAI21_X1 U5978 ( .B1(n6527), .B2(n5136), .A(n5135), .ZN(n6918) );
  NAND2_X1 U5979 ( .A1(\x_mult_f[22][8] ), .A2(\x_mult_f[23][8] ), .ZN(n6916)
         );
  INV_X1 U5980 ( .A(n6916), .ZN(n7110) );
  NAND2_X1 U5981 ( .A1(\x_mult_f[22][9] ), .A2(\x_mult_f[23][9] ), .ZN(n7112)
         );
  INV_X1 U5982 ( .A(n7112), .ZN(n5137) );
  AOI21_X1 U5983 ( .B1(n7110), .B2(n7113), .A(n5137), .ZN(n6908) );
  INV_X1 U5984 ( .A(n6911), .ZN(n5138) );
  NAND2_X1 U5985 ( .A1(\x_mult_f[22][10] ), .A2(\x_mult_f[23][10] ), .ZN(n6910) );
  OAI21_X1 U5986 ( .B1(n6908), .B2(n5138), .A(n6910), .ZN(n5139) );
  AOI21_X1 U5987 ( .B1(n5140), .B2(n3433), .A(n5139), .ZN(n6463) );
  NOR2_X1 U5988 ( .A1(\x_mult_f[22][11] ), .A2(\x_mult_f[23][11] ), .ZN(n6459)
         );
  NAND2_X1 U5989 ( .A1(\x_mult_f[22][11] ), .A2(\x_mult_f[23][11] ), .ZN(n6460) );
  OAI21_X1 U5990 ( .B1(n3432), .B2(n6459), .A(n6460), .ZN(n6932) );
  OR2_X1 U5991 ( .A1(\x_mult_f[22][12] ), .A2(\x_mult_f[23][12] ), .ZN(n6930)
         );
  NAND2_X1 U5992 ( .A1(\x_mult_f[22][12] ), .A2(\x_mult_f[23][12] ), .ZN(n6929) );
  INV_X1 U5993 ( .A(n6929), .ZN(n5141) );
  AOI21_X1 U5994 ( .B1(n6932), .B2(n6930), .A(n5141), .ZN(n5159) );
  NOR2_X1 U5995 ( .A1(\x_mult_f[22][13] ), .A2(\x_mult_f[23][13] ), .ZN(n5158)
         );
  INV_X1 U5996 ( .A(n5158), .ZN(n5142) );
  NAND2_X1 U5997 ( .A1(\x_mult_f[22][13] ), .A2(\x_mult_f[23][13] ), .ZN(n5157) );
  NAND2_X1 U5998 ( .A1(n5142), .A2(n5157), .ZN(n5143) );
  XOR2_X1 U5999 ( .A(n5159), .B(n5143), .Z(n5144) );
  AOI22_X1 U6000 ( .A1(n5144), .A2(n8209), .B1(n7698), .B2(
        \adder_stage1[11][13] ), .ZN(n5145) );
  INV_X1 U6001 ( .A(n5145), .ZN(n9973) );
  AND2_X1 U6002 ( .A1(n5147), .A2(n5146), .ZN(n6630) );
  OR2_X1 U6003 ( .A1(\x_mult_f[20][13] ), .A2(\x_mult_f[21][13] ), .ZN(n6633)
         );
  AND2_X1 U6004 ( .A1(n6630), .A2(n6633), .ZN(n5148) );
  NAND2_X1 U6005 ( .A1(n5148), .A2(n6631), .ZN(n5154) );
  OAI21_X1 U6006 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n6629) );
  NAND2_X1 U6007 ( .A1(\x_mult_f[20][13] ), .A2(\x_mult_f[21][13] ), .ZN(n6632) );
  INV_X1 U6008 ( .A(n6632), .ZN(n5152) );
  AOI21_X1 U6009 ( .B1(n6629), .B2(n6633), .A(n5152), .ZN(n5153) );
  NAND2_X1 U6010 ( .A1(n5154), .A2(n5153), .ZN(n7778) );
  INV_X2 U6011 ( .A(n8004), .ZN(n8328) );
  AOI22_X1 U6012 ( .A1(n5155), .A2(n6307), .B1(n8328), .B2(
        \adder_stage1[10][14] ), .ZN(n5156) );
  INV_X1 U6013 ( .A(n5156), .ZN(n9989) );
  OAI21_X1 U6014 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(n7731) );
  AOI22_X1 U6015 ( .A1(n5160), .A2(n4840), .B1(n8309), .B2(
        \adder_stage1[11][14] ), .ZN(n5161) );
  INV_X1 U6016 ( .A(n5161), .ZN(n9972) );
  AOI22_X1 U6017 ( .A1(n7556), .A2(\x_mult_f[13][2] ), .B1(n7155), .B2(
        \x_mult_f_int[13][2] ), .ZN(n5162) );
  INV_X1 U6018 ( .A(n5162), .ZN(n9094) );
  AOI22_X1 U6019 ( .A1(n7556), .A2(\x_mult_f[13][4] ), .B1(n7155), .B2(
        \x_mult_f_int[13][4] ), .ZN(n5163) );
  INV_X1 U6020 ( .A(n5163), .ZN(n9092) );
  AOI22_X1 U6021 ( .A1(n7556), .A2(\x_mult_f[13][5] ), .B1(n7155), .B2(
        \x_mult_f_int[13][5] ), .ZN(n5164) );
  INV_X1 U6022 ( .A(n5164), .ZN(n9091) );
  AOI22_X1 U6023 ( .A1(\x_mult_f_int[23][7] ), .A2(n5175), .B1(n8428), .B2(
        \x_mult_f[23][7] ), .ZN(n5165) );
  INV_X1 U6024 ( .A(n5165), .ZN(n9218) );
  AOI22_X1 U6025 ( .A1(\x_mult_f_int[23][9] ), .A2(n5175), .B1(n8319), .B2(
        \x_mult_f[23][9] ), .ZN(n5166) );
  INV_X1 U6026 ( .A(n5166), .ZN(n9216) );
  AOI22_X1 U6027 ( .A1(\x_mult_f_int[23][8] ), .A2(n5175), .B1(n8401), .B2(
        \x_mult_f[23][8] ), .ZN(n5167) );
  INV_X1 U6028 ( .A(n5167), .ZN(n9217) );
  AOI22_X1 U6029 ( .A1(\x_mult_f_int[23][6] ), .A2(n5175), .B1(n8398), .B2(
        \x_mult_f[23][6] ), .ZN(n5168) );
  INV_X1 U6030 ( .A(n5168), .ZN(n9219) );
  AOI22_X1 U6031 ( .A1(\x_mult_f_int[23][10] ), .A2(n5175), .B1(n7698), .B2(
        \x_mult_f[23][10] ), .ZN(n5169) );
  INV_X1 U6032 ( .A(n5169), .ZN(n9215) );
  INV_X2 U6033 ( .A(n8004), .ZN(n8325) );
  AOI22_X1 U6034 ( .A1(\x_mult_f_int[21][11] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][11] ), .ZN(n5170) );
  INV_X1 U6035 ( .A(n5170), .ZN(n9186) );
  AOI22_X1 U6036 ( .A1(\x_mult_f_int[21][8] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][8] ), .ZN(n5171) );
  INV_X1 U6037 ( .A(n5171), .ZN(n9189) );
  AOI22_X1 U6038 ( .A1(\x_mult_f_int[21][9] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][9] ), .ZN(n5172) );
  INV_X1 U6039 ( .A(n5172), .ZN(n9188) );
  AOI22_X1 U6040 ( .A1(\x_mult_f_int[21][10] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][10] ), .ZN(n5173) );
  INV_X1 U6041 ( .A(n5173), .ZN(n9187) );
  AOI22_X1 U6042 ( .A1(\x_mult_f_int[21][7] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][7] ), .ZN(n5174) );
  INV_X1 U6043 ( .A(n5174), .ZN(n9190) );
  AOI22_X1 U6044 ( .A1(\x_mult_f_int[21][6] ), .A2(n6636), .B1(n8325), .B2(
        \x_mult_f[21][6] ), .ZN(n5176) );
  INV_X1 U6045 ( .A(n5176), .ZN(n9191) );
  INV_X2 U6046 ( .A(n8004), .ZN(n8330) );
  AOI22_X1 U6047 ( .A1(\x_mult_f_int[23][11] ), .A2(n5175), .B1(n8330), .B2(
        \x_mult_f[23][11] ), .ZN(n5177) );
  INV_X1 U6048 ( .A(n5177), .ZN(n9214) );
  AOI22_X1 U6049 ( .A1(\x_mult_f_int[12][12] ), .A2(n8311), .B1(n7855), .B2(
        \x_mult_f[12][12] ), .ZN(n5178) );
  INV_X1 U6050 ( .A(n5178), .ZN(n9070) );
  AOI22_X1 U6051 ( .A1(n8398), .A2(\x_mult_f[13][3] ), .B1(n7155), .B2(
        \x_mult_f_int[13][3] ), .ZN(n5179) );
  INV_X1 U6052 ( .A(n5179), .ZN(n9093) );
  AOI22_X1 U6053 ( .A1(n8398), .A2(\x_mult_f[13][0] ), .B1(n7155), .B2(
        \x_mult_f_int[13][0] ), .ZN(n5180) );
  INV_X1 U6054 ( .A(n5180), .ZN(n9353) );
  AOI22_X1 U6055 ( .A1(\x_mult_f_int[29][7] ), .A2(n4311), .B1(n8340), .B2(
        \x_mult_f[29][7] ), .ZN(n5182) );
  INV_X1 U6056 ( .A(n5182), .ZN(n9294) );
  AOI22_X1 U6057 ( .A1(\x_mult_f_int[29][9] ), .A2(n8054), .B1(n8340), .B2(
        \x_mult_f[29][9] ), .ZN(n5183) );
  INV_X1 U6058 ( .A(n5183), .ZN(n9292) );
  AOI22_X1 U6059 ( .A1(\x_mult_f_int[29][8] ), .A2(n6636), .B1(n8340), .B2(
        \x_mult_f[29][8] ), .ZN(n5184) );
  INV_X1 U6060 ( .A(n5184), .ZN(n9293) );
  NOR2_X1 U6061 ( .A1(\adder_stage2[0][2] ), .A2(\adder_stage2[1][2] ), .ZN(
        n6429) );
  NOR2_X1 U6062 ( .A1(\adder_stage2[0][3] ), .A2(\adder_stage2[1][3] ), .ZN(
        n6412) );
  NOR2_X1 U6063 ( .A1(n6429), .A2(n6412), .ZN(n5186) );
  NOR2_X1 U6064 ( .A1(\adder_stage2[0][1] ), .A2(\adder_stage2[1][1] ), .ZN(
        n6419) );
  NAND2_X1 U6065 ( .A1(\adder_stage2[0][0] ), .A2(\adder_stage2[1][0] ), .ZN(
        n6425) );
  NAND2_X1 U6066 ( .A1(\adder_stage2[0][1] ), .A2(\adder_stage2[1][1] ), .ZN(
        n6420) );
  OAI21_X1 U6067 ( .B1(n6419), .B2(n6425), .A(n6420), .ZN(n6411) );
  NAND2_X1 U6068 ( .A1(\adder_stage2[0][2] ), .A2(\adder_stage2[1][2] ), .ZN(
        n6430) );
  NAND2_X1 U6069 ( .A1(\adder_stage2[0][3] ), .A2(\adder_stage2[1][3] ), .ZN(
        n6413) );
  OAI21_X1 U6070 ( .B1(n6412), .B2(n6430), .A(n6413), .ZN(n5185) );
  AOI21_X1 U6071 ( .B1(n5186), .B2(n6411), .A(n5185), .ZN(n6265) );
  NOR2_X1 U6072 ( .A1(\adder_stage2[0][4] ), .A2(\adder_stage2[1][4] ), .ZN(
        n6266) );
  NOR2_X1 U6073 ( .A1(\adder_stage2[0][5] ), .A2(\adder_stage2[1][5] ), .ZN(
        n8229) );
  NOR2_X1 U6074 ( .A1(n6266), .A2(n8229), .ZN(n7517) );
  NOR2_X1 U6075 ( .A1(\adder_stage2[0][6] ), .A2(\adder_stage2[1][6] ), .ZN(
        n7527) );
  NOR2_X1 U6076 ( .A1(\adder_stage2[0][7] ), .A2(\adder_stage2[1][7] ), .ZN(
        n7518) );
  NOR2_X1 U6077 ( .A1(n7527), .A2(n7518), .ZN(n5188) );
  NAND2_X1 U6078 ( .A1(n7517), .A2(n5188), .ZN(n5190) );
  NAND2_X1 U6079 ( .A1(\adder_stage2[0][4] ), .A2(\adder_stage2[1][4] ), .ZN(
        n8225) );
  NAND2_X1 U6080 ( .A1(\adder_stage2[0][5] ), .A2(\adder_stage2[1][5] ), .ZN(
        n8230) );
  OAI21_X1 U6081 ( .B1(n8229), .B2(n8225), .A(n8230), .ZN(n7516) );
  NAND2_X1 U6082 ( .A1(\adder_stage2[0][6] ), .A2(\adder_stage2[1][6] ), .ZN(
        n7528) );
  NAND2_X1 U6083 ( .A1(\adder_stage2[0][7] ), .A2(\adder_stage2[1][7] ), .ZN(
        n7519) );
  OAI21_X1 U6084 ( .B1(n7518), .B2(n7528), .A(n7519), .ZN(n5187) );
  AOI21_X1 U6085 ( .B1(n5188), .B2(n7516), .A(n5187), .ZN(n5189) );
  OAI21_X1 U6086 ( .B1(n6265), .B2(n5190), .A(n5189), .ZN(n6344) );
  NOR2_X1 U6087 ( .A1(\adder_stage2[0][8] ), .A2(\adder_stage2[1][8] ), .ZN(
        n7509) );
  NOR2_X1 U6088 ( .A1(\adder_stage2[0][9] ), .A2(\adder_stage2[1][9] ), .ZN(
        n6345) );
  NOR2_X1 U6089 ( .A1(n7509), .A2(n6345), .ZN(n7197) );
  NOR2_X1 U6090 ( .A1(\adder_stage2[0][10] ), .A2(\adder_stage2[1][10] ), .ZN(
        n7201) );
  NOR2_X1 U6091 ( .A1(\adder_stage2[0][11] ), .A2(\adder_stage2[1][11] ), .ZN(
        n7203) );
  NOR2_X1 U6092 ( .A1(n7201), .A2(n7203), .ZN(n5192) );
  NAND2_X1 U6093 ( .A1(n7197), .A2(n5192), .ZN(n7243) );
  NOR2_X1 U6094 ( .A1(\adder_stage2[0][12] ), .A2(\adder_stage2[1][12] ), .ZN(
        n7244) );
  NOR2_X1 U6095 ( .A1(n7243), .A2(n7244), .ZN(n5194) );
  NAND2_X1 U6096 ( .A1(\adder_stage2[0][8] ), .A2(\adder_stage2[1][8] ), .ZN(
        n7510) );
  NAND2_X1 U6097 ( .A1(\adder_stage2[0][9] ), .A2(\adder_stage2[1][9] ), .ZN(
        n6346) );
  OAI21_X1 U6098 ( .B1(n6345), .B2(n7510), .A(n6346), .ZN(n7198) );
  NAND2_X1 U6099 ( .A1(\adder_stage2[0][10] ), .A2(\adder_stage2[1][10] ), 
        .ZN(n7635) );
  NAND2_X1 U6100 ( .A1(\adder_stage2[0][11] ), .A2(\adder_stage2[1][11] ), 
        .ZN(n7204) );
  OAI21_X1 U6101 ( .B1(n7203), .B2(n7635), .A(n7204), .ZN(n5191) );
  AOI21_X1 U6102 ( .B1(n5192), .B2(n7198), .A(n5191), .ZN(n7242) );
  NAND2_X1 U6103 ( .A1(\adder_stage2[0][12] ), .A2(\adder_stage2[1][12] ), 
        .ZN(n7245) );
  OAI21_X1 U6104 ( .B1(n7242), .B2(n7244), .A(n7245), .ZN(n5193) );
  AOI21_X1 U6105 ( .B1(n6344), .B2(n5194), .A(n5193), .ZN(n7168) );
  NOR2_X1 U6106 ( .A1(\adder_stage2[0][13] ), .A2(\adder_stage2[1][13] ), .ZN(
        n7164) );
  NAND2_X1 U6107 ( .A1(\adder_stage2[0][13] ), .A2(\adder_stage2[1][13] ), 
        .ZN(n7165) );
  OAI21_X1 U6108 ( .B1(n7168), .B2(n7164), .A(n7165), .ZN(n7194) );
  OR2_X1 U6109 ( .A1(\adder_stage2[0][14] ), .A2(\adder_stage2[1][14] ), .ZN(
        n7192) );
  NAND2_X1 U6110 ( .A1(\adder_stage2[0][14] ), .A2(\adder_stage2[1][14] ), 
        .ZN(n7191) );
  INV_X1 U6111 ( .A(n7191), .ZN(n5195) );
  AOI21_X1 U6112 ( .B1(n7194), .B2(n7192), .A(n5195), .ZN(n8239) );
  OR2_X1 U6113 ( .A1(\adder_stage2[0][16] ), .A2(\adder_stage2[1][16] ), .ZN(
        n8241) );
  NOR2_X1 U6114 ( .A1(\adder_stage2[0][15] ), .A2(\adder_stage2[1][15] ), .ZN(
        n8238) );
  INV_X1 U6115 ( .A(n8238), .ZN(n7210) );
  NAND2_X1 U6116 ( .A1(n8241), .A2(n7210), .ZN(n5207) );
  INV_X1 U6117 ( .A(n5207), .ZN(n5196) );
  NOR2_X1 U6118 ( .A1(\adder_stage2[0][17] ), .A2(\adder_stage2[1][17] ), .ZN(
        n5199) );
  INV_X1 U6119 ( .A(n5199), .ZN(n5210) );
  NAND2_X1 U6120 ( .A1(n5196), .A2(n5210), .ZN(n7135) );
  NAND2_X1 U6121 ( .A1(\adder_stage2[0][15] ), .A2(\adder_stage2[1][15] ), 
        .ZN(n8237) );
  INV_X1 U6122 ( .A(n8237), .ZN(n5198) );
  NAND2_X1 U6123 ( .A1(\adder_stage2[0][16] ), .A2(\adder_stage2[1][16] ), 
        .ZN(n8240) );
  INV_X1 U6124 ( .A(n8240), .ZN(n5197) );
  AOI21_X1 U6125 ( .B1(n8241), .B2(n5198), .A(n5197), .ZN(n5206) );
  NAND2_X1 U6126 ( .A1(\adder_stage2[0][17] ), .A2(\adder_stage2[1][17] ), 
        .ZN(n5209) );
  OAI21_X1 U6127 ( .B1(n5206), .B2(n5199), .A(n5209), .ZN(n5200) );
  INV_X1 U6128 ( .A(n5200), .ZN(n7140) );
  OAI21_X1 U6129 ( .B1(n8239), .B2(n7135), .A(n7140), .ZN(n5202) );
  OR2_X1 U6130 ( .A1(\adder_stage2[0][18] ), .A2(\adder_stage2[1][18] ), .ZN(
        n7137) );
  NAND2_X1 U6131 ( .A1(\adder_stage2[0][18] ), .A2(\adder_stage2[1][18] ), 
        .ZN(n7138) );
  NAND2_X1 U6132 ( .A1(n7137), .A2(n7138), .ZN(n5201) );
  XNOR2_X1 U6133 ( .A(n5202), .B(n5201), .ZN(n5203) );
  AOI22_X1 U6134 ( .A1(n5203), .A2(n7570), .B1(n8328), .B2(
        \adder_stage3[0][18] ), .ZN(n5204) );
  INV_X1 U6135 ( .A(n5204), .ZN(n9751) );
  AOI22_X1 U6136 ( .A1(\x_mult_f_int[29][6] ), .A2(n7155), .B1(n8434), .B2(
        \x_mult_f[29][6] ), .ZN(n5205) );
  INV_X1 U6137 ( .A(n5205), .ZN(n9295) );
  OAI21_X1 U6138 ( .B1(n8239), .B2(n5207), .A(n5206), .ZN(n5208) );
  INV_X1 U6139 ( .A(n5208), .ZN(n5212) );
  NAND2_X1 U6140 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  XOR2_X1 U6141 ( .A(n5212), .B(n5211), .Z(n5213) );
  AOI22_X1 U6142 ( .A1(n5213), .A2(n8272), .B1(n8328), .B2(
        \adder_stage3[0][17] ), .ZN(n5214) );
  INV_X1 U6143 ( .A(n5214), .ZN(n9752) );
  AOI22_X1 U6144 ( .A1(n8401), .A2(\x_mult_f[13][1] ), .B1(n7155), .B2(
        \x_mult_f_int[13][1] ), .ZN(n5215) );
  INV_X1 U6145 ( .A(n5215), .ZN(n9352) );
  AOI22_X1 U6146 ( .A1(\x_mult_f_int[18][9] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][9] ), .ZN(n5216) );
  INV_X1 U6147 ( .A(n5216), .ZN(n9146) );
  AOI22_X1 U6148 ( .A1(\x_mult_f_int[18][10] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][10] ), .ZN(n5217) );
  INV_X1 U6149 ( .A(n5217), .ZN(n9145) );
  NOR2_X1 U6150 ( .A1(\x_mult_f[16][2] ), .A2(\x_mult_f[17][2] ), .ZN(n5323)
         );
  NOR2_X1 U6151 ( .A1(\x_mult_f[16][3] ), .A2(\x_mult_f[17][3] ), .ZN(n5299)
         );
  NOR2_X1 U6152 ( .A1(n5323), .A2(n5299), .ZN(n5219) );
  NOR2_X1 U6153 ( .A1(\x_mult_f[16][1] ), .A2(\x_mult_f[17][1] ), .ZN(n5307)
         );
  NAND2_X1 U6154 ( .A1(\x_mult_f[16][0] ), .A2(\x_mult_f[17][0] ), .ZN(n5310)
         );
  NAND2_X1 U6155 ( .A1(\x_mult_f[16][1] ), .A2(\x_mult_f[17][1] ), .ZN(n5308)
         );
  OAI21_X1 U6156 ( .B1(n5307), .B2(n5310), .A(n5308), .ZN(n5298) );
  NAND2_X1 U6157 ( .A1(\x_mult_f[16][2] ), .A2(\x_mult_f[17][2] ), .ZN(n5324)
         );
  NAND2_X1 U6158 ( .A1(\x_mult_f[16][3] ), .A2(\x_mult_f[17][3] ), .ZN(n5300)
         );
  OAI21_X1 U6159 ( .B1(n5299), .B2(n5324), .A(n5300), .ZN(n5218) );
  AOI21_X1 U6160 ( .B1(n5219), .B2(n5298), .A(n5218), .ZN(n5252) );
  NOR2_X1 U6161 ( .A1(\x_mult_f[16][4] ), .A2(\x_mult_f[17][4] ), .ZN(n5253)
         );
  NOR2_X1 U6162 ( .A1(\x_mult_f[16][5] ), .A2(\x_mult_f[17][5] ), .ZN(n5277)
         );
  NOR2_X1 U6163 ( .A1(n5253), .A2(n5277), .ZN(n5264) );
  NOR2_X1 U6164 ( .A1(\x_mult_f[16][6] ), .A2(\x_mult_f[17][6] ), .ZN(n5316)
         );
  NOR2_X1 U6165 ( .A1(\x_mult_f[16][7] ), .A2(\x_mult_f[17][7] ), .ZN(n5265)
         );
  NOR2_X1 U6166 ( .A1(n5316), .A2(n5265), .ZN(n5221) );
  NAND2_X1 U6167 ( .A1(n5264), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6168 ( .A1(\x_mult_f[16][4] ), .A2(\x_mult_f[17][4] ), .ZN(n5273)
         );
  NAND2_X1 U6169 ( .A1(\x_mult_f[16][5] ), .A2(\x_mult_f[17][5] ), .ZN(n5278)
         );
  OAI21_X1 U6170 ( .B1(n5277), .B2(n5273), .A(n5278), .ZN(n5263) );
  NAND2_X1 U6171 ( .A1(\x_mult_f[16][6] ), .A2(\x_mult_f[17][6] ), .ZN(n5317)
         );
  NAND2_X1 U6172 ( .A1(\x_mult_f[16][7] ), .A2(\x_mult_f[17][7] ), .ZN(n5266)
         );
  OAI21_X1 U6173 ( .B1(n5265), .B2(n5317), .A(n5266), .ZN(n5220) );
  AOI21_X1 U6174 ( .B1(n5221), .B2(n5263), .A(n5220), .ZN(n5222) );
  OAI21_X1 U6175 ( .B1(n5252), .B2(n5223), .A(n5222), .ZN(n5352) );
  OR2_X1 U6176 ( .A1(\x_mult_f[16][8] ), .A2(\x_mult_f[17][8] ), .ZN(n8017) );
  OR2_X1 U6177 ( .A1(\x_mult_f[16][9] ), .A2(\x_mult_f[17][9] ), .ZN(n8020) );
  AND2_X1 U6178 ( .A1(n8017), .A2(n8020), .ZN(n5353) );
  OR2_X1 U6179 ( .A1(\x_mult_f[16][10] ), .A2(\x_mult_f[17][10] ), .ZN(n5357)
         );
  AND2_X1 U6180 ( .A1(n5353), .A2(n5357), .ZN(n5227) );
  NAND2_X1 U6181 ( .A1(\x_mult_f[16][8] ), .A2(\x_mult_f[17][8] ), .ZN(n5248)
         );
  INV_X1 U6182 ( .A(n5248), .ZN(n8016) );
  NAND2_X1 U6183 ( .A1(\x_mult_f[16][9] ), .A2(\x_mult_f[17][9] ), .ZN(n8019)
         );
  INV_X1 U6184 ( .A(n8019), .ZN(n5224) );
  AOI21_X1 U6185 ( .B1(n8016), .B2(n8020), .A(n5224), .ZN(n5354) );
  INV_X1 U6186 ( .A(n5357), .ZN(n5225) );
  NAND2_X1 U6187 ( .A1(\x_mult_f[16][10] ), .A2(\x_mult_f[17][10] ), .ZN(n5356) );
  OAI21_X1 U6188 ( .B1(n5354), .B2(n5225), .A(n5356), .ZN(n5226) );
  AOI21_X1 U6189 ( .B1(n5352), .B2(n5227), .A(n5226), .ZN(n5349) );
  NOR2_X1 U6190 ( .A1(\x_mult_f[16][11] ), .A2(\x_mult_f[17][11] ), .ZN(n5345)
         );
  NAND2_X1 U6191 ( .A1(\x_mult_f[16][11] ), .A2(\x_mult_f[17][11] ), .ZN(n5346) );
  OAI21_X1 U6192 ( .B1(n3427), .B2(n5345), .A(n5346), .ZN(n6042) );
  OR2_X1 U6193 ( .A1(\x_mult_f[16][12] ), .A2(\x_mult_f[17][12] ), .ZN(n6040)
         );
  NAND2_X1 U6194 ( .A1(\x_mult_f[16][12] ), .A2(\x_mult_f[17][12] ), .ZN(n6039) );
  INV_X1 U6195 ( .A(n6039), .ZN(n5228) );
  AOI21_X1 U6196 ( .B1(n6042), .B2(n6040), .A(n5228), .ZN(n5237) );
  NOR2_X1 U6197 ( .A1(\x_mult_f[16][13] ), .A2(\x_mult_f[17][13] ), .ZN(n5233)
         );
  NAND2_X1 U6198 ( .A1(\x_mult_f[16][13] ), .A2(\x_mult_f[17][13] ), .ZN(n5234) );
  OAI21_X1 U6199 ( .B1(n5237), .B2(n5233), .A(n5234), .ZN(n7692) );
  AOI22_X1 U6200 ( .A1(n5229), .A2(n8304), .B1(n8319), .B2(
        \adder_stage1[8][14] ), .ZN(n5230) );
  INV_X1 U6201 ( .A(n5230), .ZN(n10022) );
  AOI22_X1 U6202 ( .A1(\x_mult_f_int[18][12] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][12] ), .ZN(n5231) );
  INV_X1 U6203 ( .A(n5231), .ZN(n9143) );
  AOI22_X1 U6204 ( .A1(\x_mult_f_int[18][13] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][13] ), .ZN(n5232) );
  INV_X1 U6205 ( .A(n5232), .ZN(n9142) );
  INV_X1 U6206 ( .A(n5233), .ZN(n5235) );
  NAND2_X1 U6207 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  XOR2_X1 U6208 ( .A(n5237), .B(n5236), .Z(n5238) );
  AOI22_X1 U6209 ( .A1(n5238), .A2(n8332), .B1(n8319), .B2(
        \adder_stage1[8][13] ), .ZN(n5239) );
  INV_X1 U6210 ( .A(n5239), .ZN(n10023) );
  AOI22_X1 U6211 ( .A1(\x_mult_f_int[18][11] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][11] ), .ZN(n5240) );
  INV_X1 U6212 ( .A(n5240), .ZN(n9144) );
  AOI22_X1 U6213 ( .A1(n7556), .A2(\x_mult_f[2][3] ), .B1(n8054), .B2(
        \x_mult_f_int[2][3] ), .ZN(n5241) );
  INV_X1 U6214 ( .A(n5241), .ZN(n8953) );
  AOI22_X1 U6215 ( .A1(n7556), .A2(\x_mult_f[2][1] ), .B1(n8054), .B2(
        \x_mult_f_int[2][1] ), .ZN(n5242) );
  INV_X1 U6216 ( .A(n5242), .ZN(n9330) );
  AOI22_X1 U6217 ( .A1(n7556), .A2(\x_mult_f[2][4] ), .B1(n8054), .B2(
        \x_mult_f_int[2][4] ), .ZN(n5243) );
  INV_X1 U6218 ( .A(n5243), .ZN(n8952) );
  BUF_X2 U6219 ( .A(n4444), .Z(n7919) );
  AOI22_X1 U6220 ( .A1(n7920), .A2(\x_mult_f[18][3] ), .B1(n7919), .B2(
        \x_mult_f_int[18][3] ), .ZN(n5244) );
  INV_X1 U6221 ( .A(n5244), .ZN(n9152) );
  AOI22_X1 U6222 ( .A1(n7920), .A2(\x_mult_f[18][0] ), .B1(n7919), .B2(
        \x_mult_f_int[18][0] ), .ZN(n5245) );
  INV_X1 U6223 ( .A(n5245), .ZN(n9363) );
  AOI22_X1 U6224 ( .A1(n7920), .A2(\x_mult_f[18][1] ), .B1(n7919), .B2(
        \x_mult_f_int[18][1] ), .ZN(n5246) );
  INV_X1 U6225 ( .A(n5246), .ZN(n9362) );
  BUF_X2 U6226 ( .A(n5767), .Z(n8024) );
  NAND2_X1 U6227 ( .A1(n8017), .A2(n5248), .ZN(n5249) );
  XNOR2_X1 U6228 ( .A(n8018), .B(n5249), .ZN(n5250) );
  AOI22_X1 U6229 ( .A1(n7920), .A2(\adder_stage1[8][8] ), .B1(n8024), .B2(
        n5250), .ZN(n5251) );
  INV_X1 U6230 ( .A(n5251), .ZN(n10028) );
  INV_X1 U6231 ( .A(n5252), .ZN(n5276) );
  INV_X1 U6232 ( .A(n5253), .ZN(n5275) );
  NAND2_X1 U6233 ( .A1(n5275), .A2(n5273), .ZN(n5254) );
  XNOR2_X1 U6234 ( .A(n5276), .B(n5254), .ZN(n5255) );
  AOI22_X1 U6235 ( .A1(n7920), .A2(\adder_stage1[8][4] ), .B1(n8024), .B2(
        n5255), .ZN(n5256) );
  INV_X1 U6236 ( .A(n5256), .ZN(n10032) );
  AOI22_X1 U6237 ( .A1(n7614), .A2(\x_mult_f[18][4] ), .B1(n8024), .B2(
        \x_mult_f_int[18][4] ), .ZN(n5257) );
  INV_X1 U6238 ( .A(n5257), .ZN(n9151) );
  AOI22_X1 U6239 ( .A1(n7920), .A2(\x_mult_f[18][2] ), .B1(n7919), .B2(
        \x_mult_f_int[18][2] ), .ZN(n5258) );
  INV_X1 U6240 ( .A(n5258), .ZN(n9153) );
  AOI22_X1 U6241 ( .A1(n7920), .A2(\x_mult_f[19][2] ), .B1(n7919), .B2(
        \x_mult_f_int[19][2] ), .ZN(n5259) );
  INV_X1 U6242 ( .A(n5259), .ZN(n9167) );
  OR2_X1 U6243 ( .A1(\x_mult_f[16][0] ), .A2(\x_mult_f[17][0] ), .ZN(n5260) );
  AND2_X1 U6244 ( .A1(n5260), .A2(n5310), .ZN(n5261) );
  AOI22_X1 U6245 ( .A1(n7920), .A2(\adder_stage1[8][0] ), .B1(n8024), .B2(
        n5261), .ZN(n5262) );
  INV_X1 U6246 ( .A(n5262), .ZN(n10036) );
  AOI21_X1 U6247 ( .B1(n5276), .B2(n5264), .A(n5263), .ZN(n5320) );
  OAI21_X1 U6248 ( .B1(n5320), .B2(n5316), .A(n5317), .ZN(n5269) );
  INV_X1 U6249 ( .A(n5265), .ZN(n5267) );
  NAND2_X1 U6250 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6251 ( .A(n5269), .B(n5268), .ZN(n5270) );
  AOI22_X1 U6252 ( .A1(n7920), .A2(\adder_stage1[8][7] ), .B1(n8024), .B2(
        n5270), .ZN(n5271) );
  INV_X1 U6253 ( .A(n5271), .ZN(n10029) );
  AOI22_X1 U6254 ( .A1(n7920), .A2(\x_mult_f[19][5] ), .B1(n7919), .B2(
        \x_mult_f_int[19][5] ), .ZN(n5272) );
  INV_X1 U6255 ( .A(n5272), .ZN(n9164) );
  INV_X1 U6256 ( .A(n5273), .ZN(n5274) );
  AOI21_X1 U6257 ( .B1(n5276), .B2(n5275), .A(n5274), .ZN(n5281) );
  INV_X1 U6258 ( .A(n5277), .ZN(n5279) );
  NAND2_X1 U6259 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  XOR2_X1 U6260 ( .A(n5281), .B(n5280), .Z(n5282) );
  AOI22_X1 U6261 ( .A1(n7614), .A2(\adder_stage1[8][5] ), .B1(n8024), .B2(
        n5282), .ZN(n5283) );
  INV_X1 U6262 ( .A(n5283), .ZN(n10031) );
  NOR2_X1 U6263 ( .A1(\x_mult_f[18][2] ), .A2(\x_mult_f[19][2] ), .ZN(n5851)
         );
  NOR2_X1 U6264 ( .A1(n5851), .A2(n5853), .ZN(n5285) );
  NOR2_X1 U6265 ( .A1(\x_mult_f[18][1] ), .A2(\x_mult_f[19][1] ), .ZN(n5771)
         );
  NAND2_X1 U6266 ( .A1(\x_mult_f[18][0] ), .A2(\x_mult_f[19][0] ), .ZN(n5774)
         );
  NAND2_X1 U6267 ( .A1(\x_mult_f[18][1] ), .A2(\x_mult_f[19][1] ), .ZN(n5772)
         );
  OAI21_X1 U6268 ( .B1(n5771), .B2(n5774), .A(n5772), .ZN(n5792) );
  NAND2_X1 U6269 ( .A1(\x_mult_f[18][2] ), .A2(\x_mult_f[19][2] ), .ZN(n5850)
         );
  NAND2_X1 U6270 ( .A1(\x_mult_f[18][3] ), .A2(\x_mult_f[19][3] ), .ZN(n5854)
         );
  OAI21_X1 U6271 ( .B1(n5853), .B2(n5850), .A(n5854), .ZN(n5284) );
  NOR2_X1 U6272 ( .A1(\x_mult_f[18][4] ), .A2(\x_mult_f[19][4] ), .ZN(n5783)
         );
  NOR2_X1 U6273 ( .A1(\x_mult_f[18][5] ), .A2(\x_mult_f[19][5] ), .ZN(n5785)
         );
  NOR2_X1 U6274 ( .A1(n5783), .A2(n5785), .ZN(n5900) );
  NOR2_X1 U6275 ( .A1(\x_mult_f[18][6] ), .A2(\x_mult_f[19][6] ), .ZN(n5907)
         );
  NOR2_X1 U6276 ( .A1(\x_mult_f[18][7] ), .A2(\x_mult_f[19][7] ), .ZN(n5909)
         );
  NOR2_X1 U6277 ( .A1(n5907), .A2(n5909), .ZN(n5287) );
  NAND2_X1 U6278 ( .A1(n5900), .A2(n5287), .ZN(n5289) );
  NAND2_X1 U6279 ( .A1(\x_mult_f[18][4] ), .A2(\x_mult_f[19][4] ), .ZN(n5860)
         );
  NAND2_X1 U6280 ( .A1(\x_mult_f[18][5] ), .A2(\x_mult_f[19][5] ), .ZN(n5786)
         );
  OAI21_X1 U6281 ( .B1(n5785), .B2(n5860), .A(n5786), .ZN(n5899) );
  NAND2_X1 U6282 ( .A1(\x_mult_f[18][6] ), .A2(\x_mult_f[19][6] ), .ZN(n5906)
         );
  NAND2_X1 U6283 ( .A1(\x_mult_f[18][7] ), .A2(\x_mult_f[19][7] ), .ZN(n5910)
         );
  OAI21_X1 U6284 ( .B1(n5909), .B2(n5906), .A(n5910), .ZN(n5286) );
  AOI21_X1 U6285 ( .B1(n5287), .B2(n5899), .A(n5286), .ZN(n5288) );
  OAI21_X1 U6286 ( .B1(n5782), .B2(n5289), .A(n5288), .ZN(n5934) );
  OR2_X1 U6287 ( .A1(\x_mult_f[18][8] ), .A2(\x_mult_f[19][8] ), .ZN(n5932) );
  NAND2_X1 U6288 ( .A1(\x_mult_f[18][8] ), .A2(\x_mult_f[19][8] ), .ZN(n5931)
         );
  INV_X1 U6289 ( .A(n5931), .ZN(n5290) );
  OR2_X1 U6290 ( .A1(\x_mult_f[18][10] ), .A2(\x_mult_f[19][10] ), .ZN(n5335)
         );
  NOR2_X1 U6291 ( .A1(\x_mult_f[18][9] ), .A2(\x_mult_f[19][9] ), .ZN(n5333)
         );
  INV_X1 U6292 ( .A(n5333), .ZN(n5341) );
  NAND2_X1 U6293 ( .A1(n5335), .A2(n5341), .ZN(n5709) );
  NAND2_X1 U6294 ( .A1(\x_mult_f[18][9] ), .A2(\x_mult_f[19][9] ), .ZN(n5340)
         );
  INV_X1 U6295 ( .A(n5340), .ZN(n5292) );
  NAND2_X1 U6296 ( .A1(\x_mult_f[18][10] ), .A2(\x_mult_f[19][10] ), .ZN(n5334) );
  INV_X1 U6297 ( .A(n5334), .ZN(n5291) );
  AOI21_X1 U6298 ( .B1(n5335), .B2(n5292), .A(n5291), .ZN(n5715) );
  OAI21_X1 U6299 ( .B1(n7912), .B2(n5709), .A(n5715), .ZN(n5293) );
  INV_X1 U6300 ( .A(n5293), .ZN(n5295) );
  NOR2_X1 U6301 ( .A1(\x_mult_f[18][11] ), .A2(\x_mult_f[19][11] ), .ZN(n5714)
         );
  INV_X1 U6302 ( .A(n5714), .ZN(n5710) );
  NAND2_X1 U6303 ( .A1(\x_mult_f[18][11] ), .A2(\x_mult_f[19][11] ), .ZN(n5713) );
  NAND2_X1 U6304 ( .A1(n5710), .A2(n5713), .ZN(n5294) );
  XOR2_X1 U6305 ( .A(n5295), .B(n5294), .Z(n5296) );
  AOI22_X1 U6306 ( .A1(n7920), .A2(\adder_stage1[9][11] ), .B1(n7919), .B2(
        n5296), .ZN(n5297) );
  INV_X1 U6307 ( .A(n5297), .ZN(n10008) );
  INV_X1 U6308 ( .A(n5298), .ZN(n5327) );
  OAI21_X1 U6309 ( .B1(n5327), .B2(n5323), .A(n5324), .ZN(n5303) );
  INV_X1 U6310 ( .A(n5299), .ZN(n5301) );
  NAND2_X1 U6311 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  XNOR2_X1 U6312 ( .A(n5303), .B(n5302), .ZN(n5304) );
  AOI22_X1 U6313 ( .A1(n7920), .A2(\adder_stage1[8][3] ), .B1(n8024), .B2(
        n5304), .ZN(n5305) );
  INV_X1 U6314 ( .A(n5305), .ZN(n10033) );
  AOI22_X1 U6315 ( .A1(n7920), .A2(\x_mult_f[19][1] ), .B1(n7919), .B2(
        \x_mult_f_int[19][1] ), .ZN(n5306) );
  INV_X1 U6316 ( .A(n5306), .ZN(n9364) );
  INV_X1 U6317 ( .A(n5307), .ZN(n5309) );
  NAND2_X1 U6318 ( .A1(n5309), .A2(n5308), .ZN(n5311) );
  XOR2_X1 U6319 ( .A(n5311), .B(n5310), .Z(n5312) );
  AOI22_X1 U6320 ( .A1(n6273), .A2(\adder_stage1[8][1] ), .B1(n8024), .B2(
        n5312), .ZN(n5313) );
  INV_X1 U6321 ( .A(n5313), .ZN(n10035) );
  AOI22_X1 U6322 ( .A1(n7920), .A2(\x_mult_f[19][3] ), .B1(n7919), .B2(
        \x_mult_f_int[19][3] ), .ZN(n5314) );
  INV_X1 U6323 ( .A(n5314), .ZN(n9166) );
  AOI22_X1 U6324 ( .A1(n7920), .A2(\x_mult_f[19][4] ), .B1(n7919), .B2(
        \x_mult_f_int[19][4] ), .ZN(n5315) );
  INV_X1 U6325 ( .A(n5315), .ZN(n9165) );
  INV_X1 U6326 ( .A(n5316), .ZN(n5318) );
  NAND2_X1 U6327 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  XOR2_X1 U6328 ( .A(n5320), .B(n5319), .Z(n5321) );
  AOI22_X1 U6329 ( .A1(n7920), .A2(\adder_stage1[8][6] ), .B1(n8024), .B2(
        n5321), .ZN(n5322) );
  INV_X1 U6330 ( .A(n5322), .ZN(n10030) );
  INV_X1 U6331 ( .A(n5323), .ZN(n5325) );
  NAND2_X1 U6332 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  XOR2_X1 U6333 ( .A(n5327), .B(n5326), .Z(n5328) );
  AOI22_X1 U6334 ( .A1(n7525), .A2(\adder_stage1[8][2] ), .B1(n8024), .B2(
        n5328), .ZN(n5329) );
  INV_X1 U6335 ( .A(n5329), .ZN(n10034) );
  AOI22_X1 U6336 ( .A1(n7614), .A2(\x_mult_f[18][5] ), .B1(n8024), .B2(
        \x_mult_f_int[18][5] ), .ZN(n5330) );
  INV_X1 U6337 ( .A(n5330), .ZN(n9150) );
  AOI22_X1 U6338 ( .A1(n7920), .A2(\x_mult_f[19][0] ), .B1(n7919), .B2(
        \x_mult_f_int[19][0] ), .ZN(n5331) );
  INV_X1 U6339 ( .A(n5331), .ZN(n9365) );
  OAI21_X1 U6340 ( .B1(n7912), .B2(n5333), .A(n5340), .ZN(n5337) );
  NAND2_X1 U6341 ( .A1(n5335), .A2(n5334), .ZN(n5336) );
  XNOR2_X1 U6342 ( .A(n5337), .B(n5336), .ZN(n5338) );
  AOI22_X1 U6343 ( .A1(n8097), .A2(\adder_stage1[9][10] ), .B1(n7919), .B2(
        n5338), .ZN(n5339) );
  INV_X1 U6344 ( .A(n5339), .ZN(n10009) );
  NAND2_X1 U6345 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  XOR2_X1 U6346 ( .A(n7912), .B(n5342), .Z(n5343) );
  AOI22_X1 U6347 ( .A1(n8097), .A2(\adder_stage1[9][9] ), .B1(n7919), .B2(
        n5343), .ZN(n5344) );
  INV_X1 U6348 ( .A(n5344), .ZN(n10010) );
  INV_X2 U6349 ( .A(n3407), .ZN(n8168) );
  INV_X1 U6350 ( .A(n5345), .ZN(n5347) );
  NAND2_X1 U6351 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  XOR2_X1 U6352 ( .A(n5349), .B(n5348), .Z(n5350) );
  AOI22_X1 U6353 ( .A1(n8168), .A2(\adder_stage1[8][11] ), .B1(n8024), .B2(
        n5350), .ZN(n5351) );
  INV_X1 U6354 ( .A(n5351), .ZN(n10025) );
  NAND2_X1 U6355 ( .A1(n8018), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6356 ( .A1(n5355), .A2(n5354), .ZN(n5359) );
  NAND2_X1 U6357 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  XNOR2_X1 U6358 ( .A(n5359), .B(n5358), .ZN(n5360) );
  AOI22_X1 U6359 ( .A1(n8168), .A2(\adder_stage1[8][10] ), .B1(n8024), .B2(
        n5360), .ZN(n5361) );
  INV_X1 U6360 ( .A(n5361), .ZN(n10026) );
  AOI22_X1 U6361 ( .A1(\x_mult_f_int[8][10] ), .A2(n6279), .B1(n8309), .B2(
        \x_mult_f[8][10] ), .ZN(n5362) );
  INV_X1 U6362 ( .A(n5362), .ZN(n9017) );
  AOI22_X1 U6363 ( .A1(\x_mult_f_int[8][9] ), .A2(n6279), .B1(n8309), .B2(
        \x_mult_f[8][9] ), .ZN(n5363) );
  INV_X1 U6364 ( .A(n5363), .ZN(n9018) );
  OR2_X1 U6365 ( .A1(\adder_stage1[8][12] ), .A2(\adder_stage1[9][12] ), .ZN(
        n5985) );
  NOR2_X1 U6366 ( .A1(\adder_stage1[8][11] ), .A2(\adder_stage1[9][11] ), .ZN(
        n5983) );
  INV_X1 U6367 ( .A(n5983), .ZN(n5991) );
  NAND2_X1 U6368 ( .A1(n5985), .A2(n5991), .ZN(n8201) );
  INV_X1 U6369 ( .A(n8201), .ZN(n5364) );
  NOR2_X1 U6370 ( .A1(\adder_stage1[8][13] ), .A2(\adder_stage1[9][13] ), .ZN(
        n5377) );
  INV_X1 U6371 ( .A(n5377), .ZN(n8205) );
  NAND2_X1 U6372 ( .A1(n5364), .A2(n8205), .ZN(n8091) );
  INV_X1 U6373 ( .A(n8091), .ZN(n5365) );
  NOR2_X1 U6374 ( .A1(\adder_stage1[8][14] ), .A2(\adder_stage1[9][14] ), .ZN(
        n5379) );
  INV_X1 U6375 ( .A(n5379), .ZN(n8093) );
  AND2_X1 U6376 ( .A1(n5365), .A2(n8093), .ZN(n5382) );
  NAND2_X1 U6377 ( .A1(n5366), .A2(n5371), .ZN(n5996) );
  NOR2_X1 U6378 ( .A1(\adder_stage1[8][10] ), .A2(\adder_stage1[9][10] ), .ZN(
        n5998) );
  NOR2_X1 U6379 ( .A1(n5996), .A2(n5998), .ZN(n5373) );
  INV_X1 U6380 ( .A(n5367), .ZN(n5370) );
  INV_X1 U6381 ( .A(n5368), .ZN(n5369) );
  AOI21_X1 U6382 ( .B1(n5371), .B2(n5370), .A(n5369), .ZN(n5995) );
  NAND2_X1 U6383 ( .A1(\adder_stage1[8][10] ), .A2(\adder_stage1[9][10] ), 
        .ZN(n5999) );
  OAI21_X1 U6384 ( .B1(n5995), .B2(n5998), .A(n5999), .ZN(n5372) );
  INV_X1 U6385 ( .A(n8202), .ZN(n5381) );
  NAND2_X1 U6386 ( .A1(\adder_stage1[8][11] ), .A2(\adder_stage1[9][11] ), 
        .ZN(n5990) );
  INV_X1 U6387 ( .A(n5990), .ZN(n5376) );
  NAND2_X1 U6388 ( .A1(\adder_stage1[8][12] ), .A2(\adder_stage1[9][12] ), 
        .ZN(n5984) );
  INV_X1 U6389 ( .A(n5984), .ZN(n5375) );
  AOI21_X1 U6390 ( .B1(n5985), .B2(n5376), .A(n5375), .ZN(n8200) );
  NAND2_X1 U6391 ( .A1(\adder_stage1[8][13] ), .A2(\adder_stage1[9][13] ), 
        .ZN(n8204) );
  OAI21_X1 U6392 ( .B1(n8200), .B2(n5377), .A(n8204), .ZN(n5378) );
  INV_X1 U6393 ( .A(n5378), .ZN(n8090) );
  NAND2_X1 U6394 ( .A1(\adder_stage1[8][14] ), .A2(\adder_stage1[9][14] ), 
        .ZN(n8092) );
  OAI21_X1 U6395 ( .B1(n8090), .B2(n5379), .A(n8092), .ZN(n5380) );
  AOI21_X1 U6396 ( .B1(n5382), .B2(n5381), .A(n5380), .ZN(n5383) );
  INV_X1 U6397 ( .A(n5383), .ZN(n7774) );
  AOI22_X1 U6398 ( .A1(n5385), .A2(n6636), .B1(n8309), .B2(
        \adder_stage2[4][15] ), .ZN(n5386) );
  INV_X1 U6399 ( .A(n5386), .ZN(n9821) );
  AOI22_X1 U6400 ( .A1(\x_mult_f_int[22][6] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][6] ), .ZN(n5387) );
  INV_X1 U6401 ( .A(n5387), .ZN(n9205) );
  AOI22_X1 U6402 ( .A1(\x_mult_f_int[22][7] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][7] ), .ZN(n5388) );
  INV_X1 U6403 ( .A(n5388), .ZN(n9204) );
  AOI22_X1 U6404 ( .A1(\x_mult_f_int[22][10] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][10] ), .ZN(n5389) );
  INV_X1 U6405 ( .A(n5389), .ZN(n9201) );
  AOI22_X1 U6406 ( .A1(\x_mult_f_int[22][11] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][11] ), .ZN(n5390) );
  INV_X1 U6407 ( .A(n5390), .ZN(n9200) );
  AOI22_X1 U6408 ( .A1(\x_mult_f_int[22][9] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][9] ), .ZN(n5391) );
  INV_X1 U6409 ( .A(n5391), .ZN(n9202) );
  AOI22_X1 U6410 ( .A1(\x_mult_f_int[22][8] ), .A2(n6636), .B1(n8330), .B2(
        \x_mult_f[22][8] ), .ZN(n5392) );
  INV_X1 U6411 ( .A(n5392), .ZN(n9203) );
  AOI22_X1 U6412 ( .A1(n8398), .A2(\x_mult_f[2][2] ), .B1(n8054), .B2(
        \x_mult_f_int[2][2] ), .ZN(n5393) );
  INV_X1 U6413 ( .A(n5393), .ZN(n8954) );
  AOI22_X1 U6414 ( .A1(n8401), .A2(\x_mult_f[2][0] ), .B1(n8054), .B2(
        \x_mult_f_int[2][0] ), .ZN(n5394) );
  INV_X1 U6415 ( .A(n5394), .ZN(n9331) );
  AOI22_X1 U6416 ( .A1(\x_mult_f_int[18][7] ), .A2(n6636), .B1(n7855), .B2(
        \x_mult_f[18][7] ), .ZN(n5395) );
  INV_X1 U6417 ( .A(n5395), .ZN(n9148) );
  AOI22_X1 U6418 ( .A1(\x_mult_f_int[18][8] ), .A2(n6636), .B1(n8313), .B2(
        \x_mult_f[18][8] ), .ZN(n5396) );
  INV_X1 U6419 ( .A(n5396), .ZN(n9147) );
  AOI22_X1 U6420 ( .A1(\x_mult_f_int[19][11] ), .A2(n5175), .B1(n8336), .B2(
        \x_mult_f[19][11] ), .ZN(n5397) );
  INV_X1 U6421 ( .A(n5397), .ZN(n9158) );
  AOI22_X1 U6422 ( .A1(\x_mult_f_int[18][6] ), .A2(n5175), .B1(n7864), .B2(
        \x_mult_f[18][6] ), .ZN(n5398) );
  INV_X1 U6423 ( .A(n5398), .ZN(n9149) );
  INV_X1 U6424 ( .A(n5399), .ZN(n5402) );
  NOR3_X1 U6425 ( .A1(n7049), .A2(n5402), .A3(n5400), .ZN(n5405) );
  OAI21_X1 U6426 ( .B1(n5403), .B2(n5402), .A(n5401), .ZN(n5404) );
  OR2_X1 U6427 ( .A1(n5405), .A2(n5404), .ZN(n7675) );
  AOI22_X1 U6428 ( .A1(n5407), .A2(n7819), .B1(n8340), .B2(
        \adder_stage2[2][15] ), .ZN(n5408) );
  INV_X1 U6429 ( .A(n5408), .ZN(n9855) );
  AOI22_X1 U6430 ( .A1(\x_mult_f_int[15][7] ), .A2(n8294), .B1(n7622), .B2(
        \x_mult_f[15][7] ), .ZN(n5409) );
  INV_X1 U6431 ( .A(n5409), .ZN(n9117) );
  OR2_X1 U6432 ( .A1(\adder_stage1[6][12] ), .A2(\adder_stage1[7][12] ), .ZN(
        n5868) );
  NOR2_X1 U6433 ( .A1(\adder_stage1[6][11] ), .A2(\adder_stage1[7][11] ), .ZN(
        n5866) );
  INV_X1 U6434 ( .A(n5866), .ZN(n5778) );
  NAND2_X1 U6435 ( .A1(n5868), .A2(n5778), .ZN(n5970) );
  INV_X1 U6436 ( .A(n5970), .ZN(n5410) );
  NOR2_X1 U6437 ( .A1(\adder_stage1[6][13] ), .A2(\adder_stage1[7][13] ), .ZN(
        n5429) );
  INV_X1 U6438 ( .A(n5429), .ZN(n5973) );
  NAND2_X1 U6439 ( .A1(n5410), .A2(n5973), .ZN(n8192) );
  INV_X1 U6440 ( .A(n8192), .ZN(n5411) );
  OR2_X1 U6441 ( .A1(\adder_stage1[6][14] ), .A2(\adder_stage1[7][14] ), .ZN(
        n8195) );
  AND2_X1 U6442 ( .A1(n5411), .A2(n8195), .ZN(n5434) );
  NOR2_X1 U6443 ( .A1(n5412), .A2(n5416), .ZN(n5419) );
  NAND2_X1 U6444 ( .A1(n5413), .A2(n5419), .ZN(n5421) );
  OAI21_X1 U6445 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5417) );
  AOI21_X1 U6446 ( .B1(n5419), .B2(n5418), .A(n5417), .ZN(n5420) );
  OAI21_X1 U6447 ( .B1(n5422), .B2(n5421), .A(n5420), .ZN(n5916) );
  NOR2_X1 U6448 ( .A1(\adder_stage1[6][8] ), .A2(\adder_stage1[7][8] ), .ZN(
        n5917) );
  INV_X1 U6449 ( .A(n5917), .ZN(n5964) );
  NAND2_X1 U6450 ( .A1(n3485), .A2(n3458), .ZN(n5919) );
  NAND2_X1 U6451 ( .A1(n5964), .A2(n5919), .ZN(n5955) );
  NOR2_X1 U6452 ( .A1(\adder_stage1[6][10] ), .A2(\adder_stage1[7][10] ), .ZN(
        n5956) );
  NOR2_X1 U6453 ( .A1(n5955), .A2(n5956), .ZN(n5426) );
  NAND2_X1 U6454 ( .A1(\adder_stage1[7][8] ), .A2(\adder_stage1[6][8] ), .ZN(
        n5963) );
  INV_X1 U6455 ( .A(n5963), .ZN(n5424) );
  NAND2_X1 U6456 ( .A1(\adder_stage1[7][9] ), .A2(\adder_stage1[6][9] ), .ZN(
        n5918) );
  INV_X1 U6457 ( .A(n5918), .ZN(n5423) );
  AOI21_X1 U6458 ( .B1(n5424), .B2(n5919), .A(n5423), .ZN(n5954) );
  NAND2_X1 U6459 ( .A1(\adder_stage1[6][10] ), .A2(\adder_stage1[7][10] ), 
        .ZN(n5957) );
  OAI21_X1 U6460 ( .B1(n5954), .B2(n5956), .A(n5957), .ZN(n5425) );
  INV_X1 U6461 ( .A(n8193), .ZN(n5433) );
  NAND2_X1 U6462 ( .A1(\adder_stage1[6][11] ), .A2(\adder_stage1[7][11] ), 
        .ZN(n5865) );
  INV_X1 U6463 ( .A(n5865), .ZN(n5428) );
  NAND2_X1 U6464 ( .A1(\adder_stage1[6][12] ), .A2(\adder_stage1[7][12] ), 
        .ZN(n5867) );
  INV_X1 U6465 ( .A(n5867), .ZN(n5427) );
  AOI21_X1 U6466 ( .B1(n5868), .B2(n5428), .A(n5427), .ZN(n5969) );
  NAND2_X1 U6467 ( .A1(\adder_stage1[6][13] ), .A2(\adder_stage1[7][13] ), 
        .ZN(n5972) );
  OAI21_X1 U6468 ( .B1(n5969), .B2(n5429), .A(n5972), .ZN(n5430) );
  INV_X1 U6469 ( .A(n5430), .ZN(n8191) );
  INV_X1 U6470 ( .A(n8195), .ZN(n5431) );
  NAND2_X1 U6471 ( .A1(\adder_stage1[6][14] ), .A2(\adder_stage1[7][14] ), 
        .ZN(n8194) );
  OAI21_X1 U6472 ( .B1(n8191), .B2(n5431), .A(n8194), .ZN(n5432) );
  AOI21_X1 U6473 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5435) );
  INV_X1 U6474 ( .A(n5435), .ZN(n7800) );
  AOI22_X1 U6475 ( .A1(n5436), .A2(n8332), .B1(n7669), .B2(
        \adder_stage2[3][15] ), .ZN(n5437) );
  INV_X1 U6476 ( .A(n5437), .ZN(n9838) );
  AOI21_X1 U6477 ( .B1(n8070), .B2(n5439), .A(n5438), .ZN(n5443) );
  NAND2_X1 U6478 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  XOR2_X1 U6479 ( .A(n5443), .B(n5442), .Z(n5444) );
  AOI22_X1 U6480 ( .A1(n5444), .A2(n7819), .B1(n8434), .B2(
        \adder_stage1[5][13] ), .ZN(n5445) );
  INV_X1 U6481 ( .A(n5445), .ZN(n10073) );
  AOI22_X1 U6482 ( .A1(\x_mult_f_int[15][9] ), .A2(n8294), .B1(n8427), .B2(
        \x_mult_f[15][9] ), .ZN(n5446) );
  INV_X1 U6483 ( .A(n5446), .ZN(n9115) );
  INV_X2 U6484 ( .A(n8045), .ZN(n8296) );
  AOI22_X1 U6485 ( .A1(\x_mult_f_int[15][10] ), .A2(n8294), .B1(n8296), .B2(
        \x_mult_f[15][10] ), .ZN(n5447) );
  INV_X1 U6486 ( .A(n5447), .ZN(n9114) );
  AOI22_X1 U6487 ( .A1(\x_mult_f_int[7][9] ), .A2(n8332), .B1(n8296), .B2(
        \x_mult_f[7][9] ), .ZN(n5448) );
  INV_X1 U6488 ( .A(n5448), .ZN(n9004) );
  AOI22_X1 U6489 ( .A1(\x_mult_f_int[7][8] ), .A2(n8153), .B1(n8296), .B2(
        \x_mult_f[7][8] ), .ZN(n5450) );
  INV_X1 U6490 ( .A(n5450), .ZN(n9005) );
  AOI22_X1 U6491 ( .A1(\x_mult_f_int[7][7] ), .A2(n7507), .B1(n8296), .B2(
        \x_mult_f[7][7] ), .ZN(n5451) );
  INV_X1 U6492 ( .A(n5451), .ZN(n9006) );
  AOI22_X1 U6493 ( .A1(\x_mult_f_int[7][11] ), .A2(n8175), .B1(n8296), .B2(
        \x_mult_f[7][11] ), .ZN(n5452) );
  INV_X1 U6494 ( .A(n5452), .ZN(n9002) );
  AOI22_X1 U6495 ( .A1(\x_mult_f_int[7][12] ), .A2(n7450), .B1(n8296), .B2(
        \x_mult_f[7][12] ), .ZN(n5453) );
  INV_X1 U6496 ( .A(n5453), .ZN(n9001) );
  AOI22_X1 U6497 ( .A1(\x_mult_f_int[7][10] ), .A2(n5707), .B1(n8296), .B2(
        \x_mult_f[7][10] ), .ZN(n5454) );
  INV_X1 U6498 ( .A(n5454), .ZN(n9003) );
  OR2_X1 U6499 ( .A1(\x_mult_f[6][8] ), .A2(\x_mult_f[7][8] ), .ZN(n6742) );
  OR2_X1 U6500 ( .A1(\x_mult_f[6][9] ), .A2(\x_mult_f[7][9] ), .ZN(n6733) );
  AND2_X1 U6501 ( .A1(n6742), .A2(n6733), .ZN(n6817) );
  OR2_X1 U6502 ( .A1(\x_mult_f[6][10] ), .A2(\x_mult_f[7][10] ), .ZN(n6821) );
  AND2_X1 U6503 ( .A1(n6817), .A2(n6821), .ZN(n5467) );
  NOR2_X1 U6504 ( .A1(n5455), .A2(n5458), .ZN(n6748) );
  NOR2_X1 U6505 ( .A1(\x_mult_f[6][6] ), .A2(\x_mult_f[7][6] ), .ZN(n6810) );
  NOR2_X1 U6506 ( .A1(\x_mult_f[6][7] ), .A2(\x_mult_f[7][7] ), .ZN(n6750) );
  NOR2_X1 U6507 ( .A1(n6810), .A2(n6750), .ZN(n5460) );
  NAND2_X1 U6508 ( .A1(n6748), .A2(n5460), .ZN(n5462) );
  OAI21_X1 U6509 ( .B1(n5458), .B2(n5457), .A(n5456), .ZN(n6747) );
  NAND2_X1 U6510 ( .A1(\x_mult_f[6][6] ), .A2(\x_mult_f[7][6] ), .ZN(n6811) );
  NAND2_X1 U6511 ( .A1(\x_mult_f[6][7] ), .A2(\x_mult_f[7][7] ), .ZN(n6751) );
  OAI21_X1 U6512 ( .B1(n6750), .B2(n6811), .A(n6751), .ZN(n5459) );
  AOI21_X1 U6513 ( .B1(n5460), .B2(n6747), .A(n5459), .ZN(n5461) );
  OAI21_X1 U6514 ( .B1(n5463), .B2(n5462), .A(n5461), .ZN(n6744) );
  NAND2_X1 U6515 ( .A1(\x_mult_f[6][8] ), .A2(\x_mult_f[7][8] ), .ZN(n6741) );
  INV_X1 U6516 ( .A(n6741), .ZN(n6731) );
  NAND2_X1 U6517 ( .A1(\x_mult_f[6][9] ), .A2(\x_mult_f[7][9] ), .ZN(n6732) );
  INV_X1 U6518 ( .A(n6732), .ZN(n5464) );
  AOI21_X1 U6519 ( .B1(n6731), .B2(n6733), .A(n5464), .ZN(n6818) );
  INV_X1 U6520 ( .A(n6821), .ZN(n5465) );
  NAND2_X1 U6521 ( .A1(\x_mult_f[6][10] ), .A2(\x_mult_f[7][10] ), .ZN(n6820)
         );
  OAI21_X1 U6522 ( .B1(n6818), .B2(n5465), .A(n6820), .ZN(n5466) );
  AOI21_X1 U6523 ( .B1(n5467), .B2(n3441), .A(n5466), .ZN(n6761) );
  NOR2_X1 U6524 ( .A1(\x_mult_f[6][11] ), .A2(\x_mult_f[7][11] ), .ZN(n6757)
         );
  NAND2_X1 U6525 ( .A1(\x_mult_f[6][11] ), .A2(\x_mult_f[7][11] ), .ZN(n6758)
         );
  OAI21_X1 U6526 ( .B1(n3440), .B2(n6757), .A(n6758), .ZN(n6716) );
  OR2_X1 U6527 ( .A1(\x_mult_f[6][12] ), .A2(\x_mult_f[7][12] ), .ZN(n6714) );
  NAND2_X1 U6528 ( .A1(\x_mult_f[6][12] ), .A2(\x_mult_f[7][12] ), .ZN(n6713)
         );
  INV_X1 U6529 ( .A(n6713), .ZN(n5468) );
  AOI21_X1 U6530 ( .B1(n6716), .B2(n6714), .A(n5468), .ZN(n6294) );
  NOR2_X1 U6531 ( .A1(\x_mult_f[6][13] ), .A2(\x_mult_f[7][13] ), .ZN(n6290)
         );
  NAND2_X1 U6532 ( .A1(\x_mult_f[6][13] ), .A2(\x_mult_f[7][13] ), .ZN(n6291)
         );
  OAI21_X1 U6533 ( .B1(n6294), .B2(n6290), .A(n6291), .ZN(n7822) );
  AOI22_X1 U6534 ( .A1(n5469), .A2(n6875), .B1(n8296), .B2(
        \adder_stage1[3][14] ), .ZN(n5470) );
  INV_X1 U6535 ( .A(n5470), .ZN(n10106) );
  AOI22_X1 U6536 ( .A1(\x_mult_f_int[15][8] ), .A2(n8294), .B1(n8296), .B2(
        \x_mult_f[15][8] ), .ZN(n5471) );
  INV_X1 U6537 ( .A(n5471), .ZN(n9116) );
  AOI22_X1 U6538 ( .A1(\x_mult_f_int[7][6] ), .A2(n8311), .B1(n8296), .B2(
        \x_mult_f[7][6] ), .ZN(n5472) );
  INV_X1 U6539 ( .A(n5472), .ZN(n9007) );
  NAND2_X1 U6540 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  XNOR2_X1 U6541 ( .A(n5476), .B(n5475), .ZN(n5477) );
  AOI22_X1 U6542 ( .A1(n7669), .A2(\adder_stage3[2][4] ), .B1(n7927), .B2(
        n5477), .ZN(n5478) );
  INV_X1 U6543 ( .A(n5478), .ZN(n9725) );
  OAI21_X1 U6544 ( .B1(n5481), .B2(n5480), .A(n5479), .ZN(n5486) );
  INV_X1 U6545 ( .A(n5482), .ZN(n5484) );
  NAND2_X1 U6546 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  XNOR2_X1 U6547 ( .A(n5486), .B(n5485), .ZN(n5487) );
  AOI22_X1 U6548 ( .A1(n8273), .A2(\adder_stage3[2][3] ), .B1(n7927), .B2(
        n5487), .ZN(n5488) );
  INV_X1 U6549 ( .A(n5488), .ZN(n9726) );
  AND2_X1 U6550 ( .A1(n8254), .A2(n5491), .ZN(n5499) );
  NAND2_X1 U6551 ( .A1(n8256), .A2(n5499), .ZN(n5493) );
  INV_X1 U6552 ( .A(n5489), .ZN(n5490) );
  AOI21_X1 U6553 ( .B1(n5492), .B2(n5491), .A(n5490), .ZN(n5502) );
  NAND2_X1 U6554 ( .A1(n5493), .A2(n5502), .ZN(n5495) );
  NOR2_X1 U6555 ( .A1(\adder_stage2[4][18] ), .A2(\adder_stage2[5][18] ), .ZN(
        n5501) );
  INV_X1 U6556 ( .A(n5501), .ZN(n5498) );
  NAND2_X1 U6557 ( .A1(\adder_stage2[4][18] ), .A2(\adder_stage2[5][18] ), 
        .ZN(n5500) );
  NAND2_X1 U6558 ( .A1(n5498), .A2(n5500), .ZN(n5494) );
  XNOR2_X1 U6559 ( .A(n5495), .B(n5494), .ZN(n5496) );
  AOI22_X1 U6560 ( .A1(n5496), .A2(n7819), .B1(n8306), .B2(
        \adder_stage3[2][18] ), .ZN(n5497) );
  INV_X1 U6561 ( .A(n5497), .ZN(n9711) );
  AND2_X1 U6562 ( .A1(n5499), .A2(n5498), .ZN(n7783) );
  OAI21_X1 U6563 ( .B1(n5502), .B2(n5501), .A(n5500), .ZN(n7788) );
  AOI21_X1 U6564 ( .B1(n8256), .B2(n7783), .A(n7788), .ZN(n5504) );
  OR2_X1 U6565 ( .A1(\adder_stage2[4][19] ), .A2(\adder_stage2[5][19] ), .ZN(
        n7787) );
  NAND2_X1 U6566 ( .A1(\adder_stage2[4][19] ), .A2(\adder_stage2[5][19] ), 
        .ZN(n7785) );
  NAND2_X1 U6567 ( .A1(n7787), .A2(n7785), .ZN(n5503) );
  XOR2_X1 U6568 ( .A(n5504), .B(n5503), .Z(n5505) );
  AOI22_X1 U6569 ( .A1(n5505), .A2(n6279), .B1(n8306), .B2(
        \adder_stage3[2][19] ), .ZN(n5506) );
  INV_X1 U6570 ( .A(n5506), .ZN(n9710) );
  AOI22_X1 U6571 ( .A1(n8401), .A2(\x_mult_f[0][5] ), .B1(n8281), .B2(
        \x_mult_f_int[0][5] ), .ZN(n5507) );
  INV_X1 U6572 ( .A(n5507), .ZN(n8923) );
  BUF_X2 U6573 ( .A(n6352), .Z(n8087) );
  AOI22_X1 U6574 ( .A1(n8088), .A2(\x_mult_f[9][4] ), .B1(n8087), .B2(
        \x_mult_f_int[9][4] ), .ZN(n5508) );
  INV_X1 U6575 ( .A(n5508), .ZN(n9037) );
  AOI22_X1 U6576 ( .A1(n8088), .A2(\x_mult_f[9][2] ), .B1(n8087), .B2(
        \x_mult_f_int[9][2] ), .ZN(n5509) );
  INV_X1 U6577 ( .A(n5509), .ZN(n9039) );
  AOI22_X1 U6578 ( .A1(n8088), .A2(\x_mult_f[9][3] ), .B1(n8087), .B2(
        \x_mult_f_int[9][3] ), .ZN(n5510) );
  INV_X1 U6579 ( .A(n5510), .ZN(n9038) );
  INV_X2 U6580 ( .A(n3408), .ZN(n8428) );
  AOI22_X1 U6581 ( .A1(\x_mult_f_int[3][10] ), .A2(n7962), .B1(n8428), .B2(
        \x_mult_f[3][10] ), .ZN(n5511) );
  INV_X1 U6582 ( .A(n5511), .ZN(n8960) );
  AOI22_X1 U6583 ( .A1(\x_mult_f_int[30][9] ), .A2(n8024), .B1(n8428), .B2(
        \x_mult_f[30][9] ), .ZN(n5512) );
  INV_X1 U6584 ( .A(n5512), .ZN(n9306) );
  AOI22_X1 U6585 ( .A1(\x_mult_f_int[3][12] ), .A2(n8301), .B1(n8428), .B2(
        \x_mult_f[3][12] ), .ZN(n5513) );
  INV_X1 U6586 ( .A(n5513), .ZN(n8958) );
  OAI21_X1 U6587 ( .B1(n5516), .B2(n5515), .A(n5514), .ZN(n7722) );
  AOI22_X1 U6588 ( .A1(n5517), .A2(n7962), .B1(n8428), .B2(
        \adder_stage1[1][14] ), .ZN(n5518) );
  INV_X1 U6589 ( .A(n5518), .ZN(n10138) );
  AOI22_X1 U6590 ( .A1(\x_mult_f_int[3][8] ), .A2(n7962), .B1(n8428), .B2(
        \x_mult_f[3][8] ), .ZN(n5519) );
  INV_X1 U6591 ( .A(n5519), .ZN(n8962) );
  AOI22_X1 U6592 ( .A1(\x_mult_f_int[3][9] ), .A2(n7962), .B1(n8428), .B2(
        \x_mult_f[3][9] ), .ZN(n5520) );
  INV_X1 U6593 ( .A(n5520), .ZN(n8961) );
  AOI22_X1 U6594 ( .A1(\x_mult_f_int[3][11] ), .A2(n8301), .B1(n8428), .B2(
        \x_mult_f[3][11] ), .ZN(n5521) );
  INV_X1 U6595 ( .A(n5521), .ZN(n8959) );
  AOI22_X1 U6596 ( .A1(\x_mult_f_int[30][6] ), .A2(n7819), .B1(n8319), .B2(
        \x_mult_f[30][6] ), .ZN(n5522) );
  INV_X1 U6597 ( .A(n5522), .ZN(n9309) );
  AOI22_X1 U6598 ( .A1(\x_mult_f_int[30][8] ), .A2(n7507), .B1(n8428), .B2(
        \x_mult_f[30][8] ), .ZN(n5523) );
  INV_X1 U6599 ( .A(n5523), .ZN(n9307) );
  AOI22_X1 U6600 ( .A1(\x_mult_f_int[3][7] ), .A2(n7962), .B1(n8428), .B2(
        \x_mult_f[3][7] ), .ZN(n5524) );
  INV_X1 U6601 ( .A(n5524), .ZN(n8963) );
  AOI22_X1 U6602 ( .A1(\x_mult_f_int[13][11] ), .A2(n8078), .B1(n7864), .B2(
        \x_mult_f[13][11] ), .ZN(n5525) );
  INV_X1 U6603 ( .A(n5525), .ZN(n9085) );
  AOI22_X1 U6604 ( .A1(\x_mult_f_int[14][11] ), .A2(n8334), .B1(n8296), .B2(
        \x_mult_f[14][11] ), .ZN(n5526) );
  INV_X1 U6605 ( .A(n5526), .ZN(n9099) );
  AOI22_X1 U6606 ( .A1(\x_mult_f_int[14][10] ), .A2(n8334), .B1(n7622), .B2(
        \x_mult_f[14][10] ), .ZN(n5527) );
  INV_X1 U6607 ( .A(n5527), .ZN(n9100) );
  NOR2_X1 U6608 ( .A1(\x_mult_f[8][2] ), .A2(\x_mult_f[9][2] ), .ZN(n7542) );
  NOR2_X1 U6609 ( .A1(\x_mult_f[8][3] ), .A2(\x_mult_f[9][3] ), .ZN(n7535) );
  NOR2_X1 U6610 ( .A1(n7542), .A2(n7535), .ZN(n5529) );
  NOR2_X1 U6611 ( .A1(\x_mult_f[8][1] ), .A2(\x_mult_f[9][1] ), .ZN(n7549) );
  NAND2_X1 U6612 ( .A1(\x_mult_f[8][0] ), .A2(\x_mult_f[9][0] ), .ZN(n7552) );
  NAND2_X1 U6613 ( .A1(\x_mult_f[8][1] ), .A2(\x_mult_f[9][1] ), .ZN(n7550) );
  OAI21_X1 U6614 ( .B1(n7549), .B2(n7552), .A(n7550), .ZN(n7534) );
  NAND2_X1 U6615 ( .A1(\x_mult_f[8][2] ), .A2(\x_mult_f[9][2] ), .ZN(n7543) );
  NAND2_X1 U6616 ( .A1(\x_mult_f[8][3] ), .A2(\x_mult_f[9][3] ), .ZN(n7536) );
  OAI21_X1 U6617 ( .B1(n7535), .B2(n7543), .A(n7536), .ZN(n5528) );
  AOI21_X1 U6618 ( .B1(n5529), .B2(n7534), .A(n5528), .ZN(n5572) );
  NOR2_X1 U6619 ( .A1(\x_mult_f[8][4] ), .A2(\x_mult_f[9][4] ), .ZN(n6363) );
  NOR2_X1 U6620 ( .A1(\x_mult_f[8][5] ), .A2(\x_mult_f[9][5] ), .ZN(n6365) );
  NOR2_X1 U6621 ( .A1(n6363), .A2(n6365), .ZN(n5574) );
  NOR2_X1 U6622 ( .A1(\x_mult_f[8][6] ), .A2(\x_mult_f[9][6] ), .ZN(n6356) );
  NOR2_X1 U6623 ( .A1(\x_mult_f[8][7] ), .A2(\x_mult_f[9][7] ), .ZN(n5575) );
  NOR2_X1 U6624 ( .A1(n6356), .A2(n5575), .ZN(n5531) );
  NAND2_X1 U6625 ( .A1(n5574), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U6626 ( .A1(\x_mult_f[8][4] ), .A2(\x_mult_f[9][4] ), .ZN(n6373) );
  NAND2_X1 U6627 ( .A1(\x_mult_f[8][5] ), .A2(\x_mult_f[9][5] ), .ZN(n6366) );
  OAI21_X1 U6628 ( .B1(n6365), .B2(n6373), .A(n6366), .ZN(n5573) );
  NAND2_X1 U6629 ( .A1(\x_mult_f[8][6] ), .A2(\x_mult_f[9][6] ), .ZN(n6357) );
  NAND2_X1 U6630 ( .A1(\x_mult_f[8][7] ), .A2(\x_mult_f[9][7] ), .ZN(n5576) );
  OAI21_X1 U6631 ( .B1(n5575), .B2(n6357), .A(n5576), .ZN(n5530) );
  AOI21_X1 U6632 ( .B1(n5531), .B2(n5573), .A(n5530), .ZN(n5532) );
  OAI21_X1 U6633 ( .B1(n5572), .B2(n5533), .A(n5532), .ZN(n5557) );
  OR2_X1 U6634 ( .A1(\x_mult_f[8][8] ), .A2(\x_mult_f[9][8] ), .ZN(n5555) );
  NAND2_X1 U6635 ( .A1(\x_mult_f[8][8] ), .A2(\x_mult_f[9][8] ), .ZN(n5554) );
  INV_X1 U6636 ( .A(n5554), .ZN(n5534) );
  OR2_X1 U6637 ( .A1(\x_mult_f[8][10] ), .A2(\x_mult_f[9][10] ), .ZN(n5562) );
  NOR2_X1 U6638 ( .A1(\x_mult_f[8][9] ), .A2(\x_mult_f[9][9] ), .ZN(n5560) );
  INV_X1 U6639 ( .A(n5560), .ZN(n5568) );
  NAND2_X1 U6640 ( .A1(n5562), .A2(n5568), .ZN(n5543) );
  NOR2_X1 U6641 ( .A1(n5727), .A2(n5543), .ZN(n5538) );
  NAND2_X1 U6642 ( .A1(\x_mult_f[8][9] ), .A2(\x_mult_f[9][9] ), .ZN(n5567) );
  INV_X1 U6643 ( .A(n5567), .ZN(n5536) );
  NAND2_X1 U6644 ( .A1(\x_mult_f[8][10] ), .A2(\x_mult_f[9][10] ), .ZN(n5561)
         );
  INV_X1 U6645 ( .A(n5561), .ZN(n5535) );
  AOI21_X1 U6646 ( .B1(n5562), .B2(n5536), .A(n5535), .ZN(n5548) );
  INV_X1 U6647 ( .A(n5548), .ZN(n5537) );
  NOR2_X1 U6648 ( .A1(n5538), .A2(n5537), .ZN(n5540) );
  NOR2_X1 U6649 ( .A1(\x_mult_f[8][11] ), .A2(\x_mult_f[9][11] ), .ZN(n5547)
         );
  INV_X1 U6650 ( .A(n5547), .ZN(n5544) );
  NAND2_X1 U6651 ( .A1(\x_mult_f[8][11] ), .A2(\x_mult_f[9][11] ), .ZN(n5546)
         );
  NAND2_X1 U6652 ( .A1(n5544), .A2(n5546), .ZN(n5539) );
  XOR2_X1 U6653 ( .A(n5540), .B(n5539), .Z(n5541) );
  AOI22_X1 U6654 ( .A1(n8057), .A2(\adder_stage1[4][11] ), .B1(n8087), .B2(
        n5541), .ZN(n5542) );
  INV_X1 U6655 ( .A(n5542), .ZN(n10092) );
  INV_X1 U6656 ( .A(n5543), .ZN(n5545) );
  NAND2_X1 U6657 ( .A1(n5545), .A2(n5544), .ZN(n5729) );
  OAI21_X1 U6658 ( .B1(n5548), .B2(n5547), .A(n5546), .ZN(n5549) );
  INV_X1 U6659 ( .A(n5549), .ZN(n5732) );
  OAI21_X1 U6660 ( .B1(n3414), .B2(n5729), .A(n5732), .ZN(n5551) );
  OR2_X1 U6661 ( .A1(\x_mult_f[8][12] ), .A2(\x_mult_f[9][12] ), .ZN(n5728) );
  NAND2_X1 U6662 ( .A1(\x_mult_f[8][12] ), .A2(\x_mult_f[9][12] ), .ZN(n5730)
         );
  NAND2_X1 U6663 ( .A1(n5728), .A2(n5730), .ZN(n5550) );
  XNOR2_X1 U6664 ( .A(n5551), .B(n5550), .ZN(n5552) );
  AOI22_X1 U6665 ( .A1(n8057), .A2(\adder_stage1[4][12] ), .B1(n8087), .B2(
        n5552), .ZN(n5553) );
  INV_X1 U6666 ( .A(n5553), .ZN(n10091) );
  INV_X2 U6667 ( .A(n3409), .ZN(n7622) );
  NAND2_X1 U6668 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  XNOR2_X1 U6669 ( .A(n5557), .B(n5556), .ZN(n5558) );
  AOI22_X1 U6670 ( .A1(n7622), .A2(\adder_stage1[4][8] ), .B1(n8087), .B2(
        n5558), .ZN(n5559) );
  INV_X1 U6671 ( .A(n5559), .ZN(n10095) );
  OAI21_X1 U6672 ( .B1(n3414), .B2(n5560), .A(n5567), .ZN(n5564) );
  NAND2_X1 U6673 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  XNOR2_X1 U6674 ( .A(n5564), .B(n5563), .ZN(n5565) );
  AOI22_X1 U6675 ( .A1(n7622), .A2(\adder_stage1[4][10] ), .B1(n8087), .B2(
        n5565), .ZN(n5566) );
  INV_X1 U6676 ( .A(n5566), .ZN(n10093) );
  NAND2_X1 U6677 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  XOR2_X1 U6678 ( .A(n3414), .B(n5569), .Z(n5570) );
  AOI22_X1 U6679 ( .A1(n7622), .A2(\adder_stage1[4][9] ), .B1(n8087), .B2(
        n5570), .ZN(n5571) );
  INV_X1 U6680 ( .A(n5571), .ZN(n10094) );
  INV_X1 U6681 ( .A(n5572), .ZN(n6376) );
  AOI21_X1 U6682 ( .B1(n6376), .B2(n5574), .A(n5573), .ZN(n6360) );
  OAI21_X1 U6683 ( .B1(n6360), .B2(n6356), .A(n6357), .ZN(n5579) );
  INV_X1 U6684 ( .A(n5575), .ZN(n5577) );
  NAND2_X1 U6685 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  XNOR2_X1 U6686 ( .A(n5579), .B(n5578), .ZN(n5580) );
  AOI22_X1 U6687 ( .A1(n7622), .A2(\adder_stage1[4][7] ), .B1(n8087), .B2(
        n5580), .ZN(n5581) );
  INV_X1 U6688 ( .A(n5581), .ZN(n10096) );
  OAI21_X1 U6689 ( .B1(n5584), .B2(n5583), .A(n5582), .ZN(n8419) );
  OR2_X1 U6690 ( .A1(\adder_stage2[2][16] ), .A2(\adder_stage2[3][16] ), .ZN(
        n8248) );
  NAND2_X1 U6691 ( .A1(\adder_stage2[2][16] ), .A2(\adder_stage2[3][16] ), 
        .ZN(n8247) );
  INV_X1 U6692 ( .A(n8247), .ZN(n7739) );
  AOI21_X1 U6693 ( .B1(n8419), .B2(n8248), .A(n7739), .ZN(n5586) );
  OR2_X1 U6694 ( .A1(\adder_stage2[2][17] ), .A2(\adder_stage2[3][17] ), .ZN(
        n7738) );
  NAND2_X1 U6695 ( .A1(\adder_stage2[2][17] ), .A2(\adder_stage2[3][17] ), 
        .ZN(n7736) );
  NAND2_X1 U6696 ( .A1(n7738), .A2(n7736), .ZN(n5585) );
  XOR2_X1 U6697 ( .A(n5586), .B(n5585), .Z(n5587) );
  AOI22_X1 U6698 ( .A1(n5587), .A2(n7507), .B1(n7972), .B2(
        \adder_stage3[1][17] ), .ZN(n5588) );
  INV_X1 U6699 ( .A(n5588), .ZN(n9731) );
  OR2_X1 U6700 ( .A1(\x_mult_f[0][0] ), .A2(\x_mult_f[1][0] ), .ZN(n5589) );
  AND2_X1 U6701 ( .A1(n5589), .A2(n5667), .ZN(n5590) );
  AOI22_X1 U6702 ( .A1(n8245), .A2(\adder_stage1[0][0] ), .B1(n5707), .B2(
        n5590), .ZN(n5591) );
  INV_X1 U6703 ( .A(n5591), .ZN(n10169) );
  INV_X2 U6704 ( .A(n3408), .ZN(n7959) );
  BUF_X2 U6705 ( .A(n7343), .Z(n8175) );
  AOI22_X1 U6706 ( .A1(n7959), .A2(\x_mult_f[31][1] ), .B1(n8175), .B2(
        \x_mult_f_int[31][1] ), .ZN(n5592) );
  INV_X1 U6707 ( .A(n5592), .ZN(n9388) );
  INV_X1 U6708 ( .A(n5593), .ZN(n5595) );
  NAND2_X1 U6709 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  XOR2_X1 U6710 ( .A(n5596), .B(n5631), .Z(n5597) );
  AOI22_X1 U6711 ( .A1(n7952), .A2(\adder_stage1[14][1] ), .B1(n7507), .B2(
        n5597), .ZN(n5598) );
  INV_X1 U6712 ( .A(n5598), .ZN(n9934) );
  AOI22_X1 U6713 ( .A1(n7959), .A2(\x_mult_f[31][4] ), .B1(n8175), .B2(
        \x_mult_f_int[31][4] ), .ZN(n5599) );
  INV_X1 U6714 ( .A(n5599), .ZN(n9323) );
  AOI22_X1 U6715 ( .A1(n7959), .A2(\x_mult_f[31][2] ), .B1(n8175), .B2(
        \x_mult_f_int[31][2] ), .ZN(n5600) );
  INV_X1 U6716 ( .A(n5600), .ZN(n9325) );
  AOI22_X1 U6717 ( .A1(n7959), .A2(\x_mult_f[31][5] ), .B1(n8175), .B2(
        \x_mult_f_int[31][5] ), .ZN(n5601) );
  INV_X1 U6718 ( .A(n5601), .ZN(n9322) );
  INV_X1 U6719 ( .A(n5602), .ZN(n5610) );
  INV_X1 U6720 ( .A(n5609), .ZN(n5603) );
  NAND2_X1 U6721 ( .A1(n5603), .A2(n5608), .ZN(n5604) );
  XOR2_X1 U6722 ( .A(n5610), .B(n5604), .Z(n5605) );
  AOI22_X1 U6723 ( .A1(n7952), .A2(\adder_stage1[14][2] ), .B1(n8301), .B2(
        n5605), .ZN(n5606) );
  INV_X1 U6724 ( .A(n5606), .ZN(n9933) );
  AOI22_X1 U6725 ( .A1(n7959), .A2(\x_mult_f[31][3] ), .B1(n8175), .B2(
        \x_mult_f_int[31][3] ), .ZN(n5607) );
  INV_X1 U6726 ( .A(n5607), .ZN(n9324) );
  OAI21_X1 U6727 ( .B1(n5610), .B2(n5609), .A(n5608), .ZN(n5615) );
  INV_X1 U6728 ( .A(n5611), .ZN(n5613) );
  NAND2_X1 U6729 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  XNOR2_X1 U6730 ( .A(n5615), .B(n5614), .ZN(n5616) );
  AOI22_X1 U6731 ( .A1(n7952), .A2(\adder_stage1[14][3] ), .B1(n6272), .B2(
        n5616), .ZN(n5617) );
  INV_X1 U6732 ( .A(n5617), .ZN(n9932) );
  OR2_X1 U6733 ( .A1(\x_mult_f[30][8] ), .A2(\x_mult_f[31][8] ), .ZN(n7368) );
  OR2_X1 U6734 ( .A1(\x_mult_f[30][9] ), .A2(\x_mult_f[31][9] ), .ZN(n7352) );
  AND2_X1 U6735 ( .A1(n7368), .A2(n7352), .ZN(n7395) );
  NOR2_X1 U6736 ( .A1(n5618), .A2(n7444), .ZN(n7359) );
  NOR2_X1 U6737 ( .A1(\x_mult_f[30][6] ), .A2(\x_mult_f[31][6] ), .ZN(n7433)
         );
  NOR2_X1 U6738 ( .A1(\x_mult_f[30][7] ), .A2(\x_mult_f[31][7] ), .ZN(n7360)
         );
  NOR2_X1 U6739 ( .A1(n7433), .A2(n7360), .ZN(n5621) );
  NAND2_X1 U6740 ( .A1(n7359), .A2(n5621), .ZN(n7348) );
  INV_X1 U6741 ( .A(n7348), .ZN(n5619) );
  OR2_X1 U6742 ( .A1(\x_mult_f[30][10] ), .A2(\x_mult_f[31][10] ), .ZN(n7399)
         );
  NAND2_X1 U6743 ( .A1(n5619), .A2(n7399), .ZN(n5622) );
  NAND2_X1 U6744 ( .A1(\x_mult_f[30][5] ), .A2(\x_mult_f[31][5] ), .ZN(n7445)
         );
  OAI21_X1 U6745 ( .B1(n7444), .B2(n7440), .A(n7445), .ZN(n7358) );
  NAND2_X1 U6746 ( .A1(\x_mult_f[30][6] ), .A2(\x_mult_f[31][6] ), .ZN(n7434)
         );
  NAND2_X1 U6747 ( .A1(\x_mult_f[30][7] ), .A2(\x_mult_f[31][7] ), .ZN(n7361)
         );
  OAI21_X1 U6748 ( .B1(n7360), .B2(n7434), .A(n7361), .ZN(n5620) );
  AOI21_X1 U6749 ( .B1(n5621), .B2(n7358), .A(n5620), .ZN(n7347) );
  OAI22_X1 U6750 ( .A1(n5622), .A2(n7349), .B1(n7347), .B2(n5624), .ZN(n5626)
         );
  NAND2_X1 U6751 ( .A1(\x_mult_f[30][8] ), .A2(\x_mult_f[31][8] ), .ZN(n7367)
         );
  INV_X1 U6752 ( .A(n7367), .ZN(n7350) );
  NAND2_X1 U6753 ( .A1(\x_mult_f[30][9] ), .A2(\x_mult_f[31][9] ), .ZN(n7351)
         );
  INV_X1 U6754 ( .A(n7351), .ZN(n5623) );
  AOI21_X1 U6755 ( .B1(n7350), .B2(n7352), .A(n5623), .ZN(n7396) );
  INV_X1 U6756 ( .A(n7399), .ZN(n5624) );
  NAND2_X1 U6757 ( .A1(\x_mult_f[30][10] ), .A2(\x_mult_f[31][10] ), .ZN(n7398) );
  OAI21_X1 U6758 ( .B1(n7396), .B2(n5624), .A(n7398), .ZN(n5625) );
  AOI21_X1 U6759 ( .B1(n5626), .B2(n7395), .A(n5625), .ZN(n7326) );
  NOR2_X1 U6760 ( .A1(\x_mult_f[30][11] ), .A2(\x_mult_f[31][11] ), .ZN(n7325)
         );
  INV_X1 U6761 ( .A(n7325), .ZN(n5627) );
  NAND2_X1 U6762 ( .A1(\x_mult_f[30][11] ), .A2(\x_mult_f[31][11] ), .ZN(n7324) );
  NAND2_X1 U6763 ( .A1(n5627), .A2(n7324), .ZN(n5628) );
  XOR2_X1 U6764 ( .A(n7326), .B(n5628), .Z(n5629) );
  AOI22_X1 U6765 ( .A1(n7959), .A2(\adder_stage1[15][11] ), .B1(n6036), .B2(
        n5629), .ZN(n5630) );
  INV_X1 U6766 ( .A(n5630), .ZN(n9907) );
  OR2_X1 U6767 ( .A1(\x_mult_f[28][0] ), .A2(\x_mult_f[29][0] ), .ZN(n5632) );
  AND2_X1 U6768 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  AOI22_X1 U6769 ( .A1(n7952), .A2(\adder_stage1[14][0] ), .B1(n8175), .B2(
        n5633), .ZN(n5634) );
  INV_X1 U6770 ( .A(n5634), .ZN(n9935) );
  NOR2_X1 U6771 ( .A1(\x_mult_f[24][5] ), .A2(\x_mult_f[25][5] ), .ZN(n6022)
         );
  NOR2_X1 U6772 ( .A1(n5635), .A2(n6022), .ZN(n6010) );
  NOR2_X1 U6773 ( .A1(\x_mult_f[24][6] ), .A2(\x_mult_f[25][6] ), .ZN(n6029)
         );
  NOR2_X1 U6774 ( .A1(\x_mult_f[24][7] ), .A2(\x_mult_f[25][7] ), .ZN(n6011)
         );
  NOR2_X1 U6775 ( .A1(n6029), .A2(n6011), .ZN(n5637) );
  NAND2_X1 U6776 ( .A1(n6010), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U6777 ( .A1(\x_mult_f[24][5] ), .A2(\x_mult_f[25][5] ), .ZN(n6023)
         );
  OAI21_X1 U6778 ( .B1(n6022), .B2(n6018), .A(n6023), .ZN(n6009) );
  NAND2_X1 U6779 ( .A1(\x_mult_f[24][6] ), .A2(\x_mult_f[25][6] ), .ZN(n6030)
         );
  NAND2_X1 U6780 ( .A1(\x_mult_f[24][7] ), .A2(\x_mult_f[25][7] ), .ZN(n6012)
         );
  OAI21_X1 U6781 ( .B1(n6011), .B2(n6030), .A(n6012), .ZN(n5636) );
  AOI21_X1 U6782 ( .B1(n5637), .B2(n6009), .A(n5636), .ZN(n5638) );
  OAI21_X1 U6783 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n7452) );
  OR2_X1 U6784 ( .A1(\x_mult_f[24][8] ), .A2(\x_mult_f[25][8] ), .ZN(n7454) );
  OR2_X1 U6785 ( .A1(\x_mult_f[24][9] ), .A2(\x_mult_f[25][9] ), .ZN(n7456) );
  AND2_X1 U6786 ( .A1(n7454), .A2(n7456), .ZN(n7461) );
  OR2_X1 U6787 ( .A1(\x_mult_f[24][10] ), .A2(\x_mult_f[25][10] ), .ZN(n7465)
         );
  AND2_X1 U6788 ( .A1(n7461), .A2(n7465), .ZN(n5644) );
  NAND2_X1 U6789 ( .A1(\x_mult_f[24][8] ), .A2(\x_mult_f[25][8] ), .ZN(n6005)
         );
  INV_X1 U6790 ( .A(n6005), .ZN(n7453) );
  NAND2_X1 U6791 ( .A1(\x_mult_f[24][9] ), .A2(\x_mult_f[25][9] ), .ZN(n7455)
         );
  INV_X1 U6792 ( .A(n7455), .ZN(n5641) );
  AOI21_X1 U6793 ( .B1(n7453), .B2(n7456), .A(n5641), .ZN(n7462) );
  INV_X1 U6794 ( .A(n7465), .ZN(n5642) );
  NAND2_X1 U6795 ( .A1(\x_mult_f[24][10] ), .A2(\x_mult_f[25][10] ), .ZN(n7464) );
  OAI21_X1 U6796 ( .B1(n7462), .B2(n5642), .A(n7464), .ZN(n5643) );
  AOI21_X1 U6797 ( .B1(n3435), .B2(n5644), .A(n5643), .ZN(n6455) );
  NOR2_X1 U6798 ( .A1(\x_mult_f[24][11] ), .A2(\x_mult_f[25][11] ), .ZN(n6454)
         );
  INV_X1 U6799 ( .A(n6454), .ZN(n5645) );
  NAND2_X1 U6800 ( .A1(\x_mult_f[24][11] ), .A2(\x_mult_f[25][11] ), .ZN(n6453) );
  NAND2_X1 U6801 ( .A1(n5645), .A2(n6453), .ZN(n5646) );
  XOR2_X1 U6802 ( .A(n6455), .B(n5646), .Z(n5647) );
  AOI22_X1 U6803 ( .A1(n8176), .A2(\adder_stage1[12][11] ), .B1(n8175), .B2(
        n5647), .ZN(n5648) );
  INV_X1 U6804 ( .A(n5648), .ZN(n9958) );
  AOI22_X1 U6805 ( .A1(n8176), .A2(\x_mult_f[25][1] ), .B1(n8209), .B2(
        \x_mult_f_int[25][1] ), .ZN(n5649) );
  INV_X1 U6806 ( .A(n5649), .ZN(n9376) );
  AOI22_X1 U6807 ( .A1(n7959), .A2(\x_mult_f[27][2] ), .B1(n8175), .B2(
        \x_mult_f_int[27][2] ), .ZN(n5650) );
  INV_X1 U6808 ( .A(n5650), .ZN(n9271) );
  AOI22_X1 U6809 ( .A1(n7177), .A2(\x_mult_f[27][1] ), .B1(n8024), .B2(
        \x_mult_f_int[27][1] ), .ZN(n5651) );
  INV_X1 U6810 ( .A(n5651), .ZN(n9380) );
  AOI22_X1 U6811 ( .A1(n8176), .A2(\x_mult_f[25][0] ), .B1(n7507), .B2(
        \x_mult_f_int[25][0] ), .ZN(n5652) );
  INV_X1 U6812 ( .A(n5652), .ZN(n9377) );
  AOI22_X1 U6813 ( .A1(n7928), .A2(\x_mult_f[27][4] ), .B1(n8175), .B2(
        \x_mult_f_int[27][4] ), .ZN(n5653) );
  INV_X1 U6814 ( .A(n5653), .ZN(n9269) );
  AOI22_X1 U6815 ( .A1(n7920), .A2(\x_mult_f[27][0] ), .B1(n8235), .B2(
        \x_mult_f_int[27][0] ), .ZN(n5654) );
  INV_X1 U6816 ( .A(n5654), .ZN(n9381) );
  AOI22_X1 U6817 ( .A1(n7614), .A2(\x_mult_f[27][3] ), .B1(n8175), .B2(
        \x_mult_f_int[27][3] ), .ZN(n5655) );
  INV_X1 U6818 ( .A(n5655), .ZN(n9270) );
  INV_X1 U6819 ( .A(n5656), .ZN(n5680) );
  OAI21_X1 U6820 ( .B1(n5680), .B2(n5676), .A(n5677), .ZN(n5661) );
  INV_X1 U6821 ( .A(n5657), .ZN(n5659) );
  NAND2_X1 U6822 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  XNOR2_X1 U6823 ( .A(n5661), .B(n5660), .ZN(n5662) );
  AOI22_X1 U6824 ( .A1(n6854), .A2(\adder_stage1[0][3] ), .B1(n5707), .B2(
        n5662), .ZN(n5663) );
  INV_X1 U6825 ( .A(n5663), .ZN(n10166) );
  INV_X1 U6826 ( .A(n5664), .ZN(n5666) );
  NAND2_X1 U6827 ( .A1(n5666), .A2(n5665), .ZN(n5668) );
  XOR2_X1 U6828 ( .A(n5668), .B(n5667), .Z(n5669) );
  AOI22_X1 U6829 ( .A1(n6854), .A2(\adder_stage1[0][1] ), .B1(n5707), .B2(
        n5669), .ZN(n5670) );
  INV_X1 U6830 ( .A(n5670), .ZN(n10168) );
  NAND2_X1 U6831 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  XNOR2_X1 U6832 ( .A(n5693), .B(n5673), .ZN(n5674) );
  AOI22_X1 U6833 ( .A1(n6854), .A2(\adder_stage1[0][4] ), .B1(n5707), .B2(
        n5674), .ZN(n5675) );
  INV_X1 U6834 ( .A(n5675), .ZN(n10165) );
  INV_X1 U6835 ( .A(n5676), .ZN(n5678) );
  NAND2_X1 U6836 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  XOR2_X1 U6837 ( .A(n5680), .B(n5679), .Z(n5681) );
  AOI22_X1 U6838 ( .A1(n6854), .A2(\adder_stage1[0][2] ), .B1(n5707), .B2(
        n5681), .ZN(n5682) );
  INV_X1 U6839 ( .A(n5682), .ZN(n10167) );
  AOI22_X1 U6840 ( .A1(n7556), .A2(\x_mult_f[2][5] ), .B1(n5707), .B2(
        \x_mult_f_int[2][5] ), .ZN(n5683) );
  INV_X1 U6841 ( .A(n5683), .ZN(n8951) );
  AOI21_X1 U6842 ( .B1(n7425), .B2(n7373), .A(n5684), .ZN(n5688) );
  NAND2_X1 U6843 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  XOR2_X1 U6844 ( .A(n5688), .B(n5687), .Z(n5689) );
  AOI22_X1 U6845 ( .A1(n7640), .A2(\adder_stage1[13][9] ), .B1(n7570), .B2(
        n5689), .ZN(n5690) );
  INV_X1 U6846 ( .A(n5690), .ZN(n9943) );
  AOI21_X1 U6847 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n5700) );
  INV_X1 U6848 ( .A(n5699), .ZN(n5694) );
  NAND2_X1 U6849 ( .A1(n5694), .A2(n5698), .ZN(n5695) );
  XOR2_X1 U6850 ( .A(n5700), .B(n5695), .Z(n5696) );
  AOI22_X1 U6851 ( .A1(n7074), .A2(\adder_stage1[0][6] ), .B1(n5707), .B2(
        n5696), .ZN(n5697) );
  INV_X1 U6852 ( .A(n5697), .ZN(n10163) );
  OAI21_X1 U6853 ( .B1(n5700), .B2(n5699), .A(n5698), .ZN(n5705) );
  INV_X1 U6854 ( .A(n5701), .ZN(n5703) );
  NAND2_X1 U6855 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  XNOR2_X1 U6856 ( .A(n5705), .B(n5704), .ZN(n5706) );
  AOI22_X1 U6857 ( .A1(n7074), .A2(\adder_stage1[0][7] ), .B1(n5707), .B2(
        n5706), .ZN(n5708) );
  INV_X1 U6858 ( .A(n5708), .ZN(n10162) );
  INV_X1 U6859 ( .A(n5709), .ZN(n5711) );
  NAND2_X1 U6860 ( .A1(n5711), .A2(n5710), .ZN(n7911) );
  NOR2_X1 U6861 ( .A1(\x_mult_f[18][12] ), .A2(\x_mult_f[19][12] ), .ZN(n7913)
         );
  OR2_X1 U6862 ( .A1(n7911), .A2(n7913), .ZN(n5712) );
  NOR2_X1 U6863 ( .A1(n5712), .A2(n7912), .ZN(n5718) );
  OAI21_X1 U6864 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5716) );
  INV_X1 U6865 ( .A(n5716), .ZN(n7910) );
  NAND2_X1 U6866 ( .A1(\x_mult_f[18][12] ), .A2(\x_mult_f[19][12] ), .ZN(n7914) );
  OAI21_X1 U6867 ( .B1(n7910), .B2(n7913), .A(n7914), .ZN(n5717) );
  NOR2_X1 U6868 ( .A1(n5718), .A2(n5717), .ZN(n7340) );
  NOR2_X1 U6869 ( .A1(\x_mult_f[18][13] ), .A2(\x_mult_f[19][13] ), .ZN(n7336)
         );
  NAND2_X1 U6870 ( .A1(\x_mult_f[18][13] ), .A2(\x_mult_f[19][13] ), .ZN(n7337) );
  OAI21_X1 U6871 ( .B1(n7340), .B2(n7336), .A(n7337), .ZN(n7500) );
  INV_X2 U6872 ( .A(n3407), .ZN(n7698) );
  AOI22_X1 U6873 ( .A1(n5719), .A2(n8314), .B1(n7698), .B2(
        \adder_stage1[9][14] ), .ZN(n5720) );
  INV_X1 U6874 ( .A(n5720), .ZN(n10005) );
  AOI22_X1 U6875 ( .A1(\x_mult_f_int[9][7] ), .A2(n6307), .B1(n7698), .B2(
        \x_mult_f[9][7] ), .ZN(n5721) );
  INV_X1 U6876 ( .A(n5721), .ZN(n9034) );
  AOI22_X1 U6877 ( .A1(\x_mult_f_int[9][8] ), .A2(n6875), .B1(n7698), .B2(
        \x_mult_f[9][8] ), .ZN(n5722) );
  INV_X1 U6878 ( .A(n5722), .ZN(n9033) );
  AOI22_X1 U6879 ( .A1(\x_mult_f_int[19][6] ), .A2(n7862), .B1(n7698), .B2(
        \x_mult_f[19][6] ), .ZN(n5723) );
  INV_X1 U6880 ( .A(n5723), .ZN(n9163) );
  AOI22_X1 U6881 ( .A1(\x_mult_f_int[9][6] ), .A2(n6307), .B1(n7698), .B2(
        \x_mult_f[9][6] ), .ZN(n5724) );
  INV_X1 U6882 ( .A(n5724), .ZN(n9035) );
  AOI22_X1 U6883 ( .A1(\x_mult_f_int[19][7] ), .A2(n8153), .B1(n7698), .B2(
        \x_mult_f[19][7] ), .ZN(n5725) );
  INV_X1 U6884 ( .A(n5725), .ZN(n9162) );
  AOI22_X1 U6885 ( .A1(\x_mult_f_int[19][10] ), .A2(n7971), .B1(n8313), .B2(
        \x_mult_f[19][10] ), .ZN(n5726) );
  INV_X1 U6886 ( .A(n5726), .ZN(n9159) );
  INV_X1 U6887 ( .A(n5727), .ZN(n5735) );
  INV_X1 U6888 ( .A(n5728), .ZN(n5731) );
  NOR2_X1 U6889 ( .A1(n5729), .A2(n5731), .ZN(n5734) );
  OAI21_X1 U6890 ( .B1(n5732), .B2(n5731), .A(n5730), .ZN(n5733) );
  AOI21_X1 U6891 ( .B1(n5735), .B2(n5734), .A(n5733), .ZN(n6057) );
  NOR2_X1 U6892 ( .A1(\x_mult_f[8][13] ), .A2(\x_mult_f[9][13] ), .ZN(n6056)
         );
  INV_X1 U6893 ( .A(n6056), .ZN(n5736) );
  NAND2_X1 U6894 ( .A1(\x_mult_f[8][13] ), .A2(\x_mult_f[9][13] ), .ZN(n6055)
         );
  NAND2_X1 U6895 ( .A1(n5736), .A2(n6055), .ZN(n5737) );
  XOR2_X1 U6896 ( .A(n3413), .B(n5737), .Z(n5738) );
  AOI22_X1 U6897 ( .A1(n5738), .A2(n6307), .B1(n8319), .B2(
        \adder_stage1[4][13] ), .ZN(n5739) );
  INV_X1 U6898 ( .A(n5739), .ZN(n10090) );
  BUF_X2 U6899 ( .A(n5767), .Z(n6036) );
  AOI22_X1 U6900 ( .A1(n7556), .A2(\x_mult_f[0][0] ), .B1(n6036), .B2(
        \x_mult_f_int[0][0] ), .ZN(n5740) );
  INV_X1 U6901 ( .A(n5740), .ZN(n9327) );
  AOI22_X1 U6902 ( .A1(n7556), .A2(\x_mult_f[0][1] ), .B1(n6036), .B2(
        \x_mult_f_int[0][1] ), .ZN(n5741) );
  INV_X1 U6903 ( .A(n5741), .ZN(n9326) );
  AOI22_X1 U6904 ( .A1(n7525), .A2(\x_mult_f[0][3] ), .B1(n6036), .B2(
        \x_mult_f_int[0][3] ), .ZN(n5742) );
  INV_X1 U6905 ( .A(n5742), .ZN(n8925) );
  AOI22_X1 U6906 ( .A1(n7556), .A2(\x_mult_f[0][4] ), .B1(n6036), .B2(
        \x_mult_f_int[0][4] ), .ZN(n5743) );
  INV_X1 U6907 ( .A(n5743), .ZN(n8924) );
  AOI22_X1 U6908 ( .A1(n7177), .A2(\x_mult_f[1][0] ), .B1(n6036), .B2(
        \x_mult_f_int[1][0] ), .ZN(n5744) );
  INV_X1 U6909 ( .A(n5744), .ZN(n9329) );
  AOI22_X1 U6910 ( .A1(n7177), .A2(\x_mult_f[1][1] ), .B1(n6036), .B2(
        \x_mult_f_int[1][1] ), .ZN(n5745) );
  INV_X1 U6911 ( .A(n5745), .ZN(n9328) );
  AOI22_X1 U6912 ( .A1(n8168), .A2(\x_mult_f[1][2] ), .B1(n6036), .B2(
        \x_mult_f_int[1][2] ), .ZN(n5746) );
  INV_X1 U6913 ( .A(n5746), .ZN(n8940) );
  BUF_X2 U6914 ( .A(n6238), .Z(n5981) );
  AOI22_X1 U6915 ( .A1(n7920), .A2(\x_mult_f[14][2] ), .B1(n5981), .B2(
        \x_mult_f_int[14][2] ), .ZN(n5747) );
  INV_X1 U6916 ( .A(n5747), .ZN(n9108) );
  AOI22_X1 U6917 ( .A1(n6273), .A2(\x_mult_f[20][1] ), .B1(n6036), .B2(
        \x_mult_f_int[20][1] ), .ZN(n5748) );
  INV_X1 U6918 ( .A(n5748), .ZN(n9366) );
  AOI22_X1 U6919 ( .A1(n6273), .A2(\x_mult_f[20][0] ), .B1(n6036), .B2(
        \x_mult_f_int[20][0] ), .ZN(n5749) );
  INV_X1 U6920 ( .A(n5749), .ZN(n9367) );
  AOI22_X1 U6921 ( .A1(n7525), .A2(\x_mult_f[14][3] ), .B1(n5981), .B2(
        \x_mult_f_int[14][3] ), .ZN(n5750) );
  INV_X1 U6922 ( .A(n5750), .ZN(n9107) );
  AOI22_X1 U6923 ( .A1(n7959), .A2(\x_mult_f[1][3] ), .B1(n6036), .B2(
        \x_mult_f_int[1][3] ), .ZN(n5751) );
  INV_X1 U6924 ( .A(n5751), .ZN(n8939) );
  AOI22_X1 U6925 ( .A1(n6273), .A2(\x_mult_f[14][4] ), .B1(n5981), .B2(
        \x_mult_f_int[14][4] ), .ZN(n5752) );
  INV_X1 U6926 ( .A(n5752), .ZN(n9106) );
  AOI22_X1 U6927 ( .A1(n7920), .A2(\x_mult_f[14][5] ), .B1(n5981), .B2(
        \x_mult_f_int[14][5] ), .ZN(n5753) );
  INV_X1 U6928 ( .A(n5753), .ZN(n9105) );
  AOI22_X1 U6929 ( .A1(n7928), .A2(\x_mult_f[1][4] ), .B1(n6036), .B2(
        \x_mult_f_int[1][4] ), .ZN(n5754) );
  INV_X1 U6930 ( .A(n5754), .ZN(n8938) );
  AOI22_X1 U6931 ( .A1(n8176), .A2(\x_mult_f[1][5] ), .B1(n6036), .B2(
        \x_mult_f_int[1][5] ), .ZN(n5755) );
  INV_X1 U6932 ( .A(n5755), .ZN(n8937) );
  AOI22_X1 U6933 ( .A1(n6273), .A2(\x_mult_f[21][5] ), .B1(n6036), .B2(
        \x_mult_f_int[21][5] ), .ZN(n5756) );
  INV_X1 U6934 ( .A(n5756), .ZN(n9192) );
  INV_X1 U6935 ( .A(n5757), .ZN(n5946) );
  AOI21_X1 U6936 ( .B1(n5946), .B2(n5759), .A(n5758), .ZN(n5928) );
  OAI21_X1 U6937 ( .B1(n5928), .B2(n5924), .A(n5925), .ZN(n5764) );
  INV_X1 U6938 ( .A(n5760), .ZN(n5762) );
  NAND2_X1 U6939 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  XNOR2_X1 U6940 ( .A(n5764), .B(n5763), .ZN(n5765) );
  AOI22_X1 U6941 ( .A1(n8336), .A2(\adder_stage1[6][7] ), .B1(n5981), .B2(
        n5765), .ZN(n5766) );
  INV_X1 U6942 ( .A(n5766), .ZN(n10063) );
  BUF_X2 U6943 ( .A(n5767), .Z(n8209) );
  OR2_X1 U6944 ( .A1(\x_mult_f[18][0] ), .A2(\x_mult_f[19][0] ), .ZN(n5768) );
  AND2_X1 U6945 ( .A1(n5768), .A2(n5774), .ZN(n5769) );
  AOI22_X1 U6946 ( .A1(n8097), .A2(\adder_stage1[9][0] ), .B1(n8209), .B2(
        n5769), .ZN(n5770) );
  INV_X1 U6947 ( .A(n5770), .ZN(n10019) );
  INV_X1 U6948 ( .A(n5771), .ZN(n5773) );
  NAND2_X1 U6949 ( .A1(n5773), .A2(n5772), .ZN(n5775) );
  XOR2_X1 U6950 ( .A(n5775), .B(n5774), .Z(n5776) );
  AOI22_X1 U6951 ( .A1(n8097), .A2(\adder_stage1[9][1] ), .B1(n8209), .B2(
        n5776), .ZN(n5777) );
  INV_X1 U6952 ( .A(n5777), .ZN(n10018) );
  NAND2_X1 U6953 ( .A1(n5778), .A2(n5865), .ZN(n5779) );
  XOR2_X1 U6954 ( .A(n8193), .B(n5779), .Z(n5780) );
  AOI22_X1 U6955 ( .A1(n8057), .A2(\adder_stage2[3][11] ), .B1(n8281), .B2(
        n5780), .ZN(n5781) );
  INV_X1 U6956 ( .A(n5781), .ZN(n9842) );
  INV_X1 U6957 ( .A(n5782), .ZN(n5901) );
  INV_X1 U6958 ( .A(n5783), .ZN(n5861) );
  INV_X1 U6959 ( .A(n5860), .ZN(n5784) );
  AOI21_X1 U6960 ( .B1(n5901), .B2(n5861), .A(n5784), .ZN(n5789) );
  INV_X1 U6961 ( .A(n5785), .ZN(n5787) );
  NAND2_X1 U6962 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XOR2_X1 U6963 ( .A(n5789), .B(n5788), .Z(n5790) );
  AOI22_X1 U6964 ( .A1(n8097), .A2(\adder_stage1[9][5] ), .B1(n8209), .B2(
        n5790), .ZN(n5791) );
  INV_X1 U6965 ( .A(n5791), .ZN(n10014) );
  INV_X1 U6966 ( .A(n5792), .ZN(n5852) );
  INV_X1 U6967 ( .A(n5851), .ZN(n5793) );
  NAND2_X1 U6968 ( .A1(n5793), .A2(n5850), .ZN(n5794) );
  XOR2_X1 U6969 ( .A(n5852), .B(n5794), .Z(n5795) );
  AOI22_X1 U6970 ( .A1(n8097), .A2(\adder_stage1[9][2] ), .B1(n8209), .B2(
        n5795), .ZN(n5796) );
  INV_X1 U6971 ( .A(n5796), .ZN(n10017) );
  INV_X1 U6972 ( .A(n5797), .ZN(n5799) );
  NAND2_X1 U6973 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  XOR2_X1 U6974 ( .A(n5801), .B(n5800), .Z(n5802) );
  AOI22_X1 U6975 ( .A1(n7855), .A2(\adder_stage1[7][6] ), .B1(n8292), .B2(
        n5802), .ZN(n5803) );
  INV_X1 U6976 ( .A(n5803), .ZN(n10047) );
  INV_X1 U6977 ( .A(n5804), .ZN(n5814) );
  INV_X1 U6978 ( .A(n5813), .ZN(n5805) );
  AOI21_X1 U6979 ( .B1(n5816), .B2(n5814), .A(n5805), .ZN(n5810) );
  INV_X1 U6980 ( .A(n5806), .ZN(n5808) );
  NAND2_X1 U6981 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XOR2_X1 U6982 ( .A(n5810), .B(n5809), .Z(n5811) );
  AOI22_X1 U6983 ( .A1(n6854), .A2(\adder_stage1[7][5] ), .B1(n6626), .B2(
        n5811), .ZN(n5812) );
  INV_X1 U6984 ( .A(n5812), .ZN(n10048) );
  NAND2_X1 U6985 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  XNOR2_X1 U6986 ( .A(n5816), .B(n5815), .ZN(n5817) );
  AOI22_X1 U6987 ( .A1(n8118), .A2(\adder_stage1[7][4] ), .B1(n8153), .B2(
        n5817), .ZN(n5818) );
  INV_X1 U6988 ( .A(n5818), .ZN(n10049) );
  INV_X1 U6989 ( .A(n5819), .ZN(n5831) );
  OAI21_X1 U6990 ( .B1(n5831), .B2(n5827), .A(n5828), .ZN(n5824) );
  INV_X1 U6991 ( .A(n5820), .ZN(n5822) );
  NAND2_X1 U6992 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U6993 ( .A(n5824), .B(n5823), .ZN(n5825) );
  AOI22_X1 U6994 ( .A1(n7074), .A2(\adder_stage1[7][3] ), .B1(n5981), .B2(
        n5825), .ZN(n5826) );
  INV_X1 U6995 ( .A(n5826), .ZN(n10050) );
  INV_X1 U6996 ( .A(n5827), .ZN(n5829) );
  NAND2_X1 U6997 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  XOR2_X1 U6998 ( .A(n5831), .B(n5830), .Z(n5832) );
  NAND2_X1 U6999 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XNOR2_X1 U7000 ( .A(n5837), .B(n5836), .ZN(n5838) );
  AOI22_X1 U7001 ( .A1(n8057), .A2(\adder_stage1[6][8] ), .B1(n5981), .B2(
        n5838), .ZN(n5839) );
  INV_X1 U7002 ( .A(n5839), .ZN(n10062) );
  INV_X1 U7003 ( .A(n5840), .ZN(n5842) );
  NAND2_X1 U7004 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  XOR2_X1 U7005 ( .A(n5843), .B(n5846), .Z(n5844) );
  AOI22_X1 U7006 ( .A1(n8057), .A2(\adder_stage1[7][1] ), .B1(n6626), .B2(
        n5844), .ZN(n5845) );
  INV_X1 U7007 ( .A(n5845), .ZN(n10052) );
  OR2_X1 U7008 ( .A1(\x_mult_f[14][0] ), .A2(\x_mult_f[15][0] ), .ZN(n5847) );
  AND2_X1 U7009 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  AOI22_X1 U7010 ( .A1(n7041), .A2(\adder_stage1[7][0] ), .B1(n8153), .B2(
        n5848), .ZN(n5849) );
  INV_X1 U7011 ( .A(n5849), .ZN(n10053) );
  OAI21_X1 U7012 ( .B1(n5852), .B2(n5851), .A(n5850), .ZN(n5857) );
  INV_X1 U7013 ( .A(n5853), .ZN(n5855) );
  NAND2_X1 U7014 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  XNOR2_X1 U7015 ( .A(n5857), .B(n5856), .ZN(n5858) );
  AOI22_X1 U7016 ( .A1(n8097), .A2(\adder_stage1[9][3] ), .B1(n8209), .B2(
        n5858), .ZN(n5859) );
  INV_X1 U7017 ( .A(n5859), .ZN(n10016) );
  NAND2_X1 U7018 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  XNOR2_X1 U7019 ( .A(n5901), .B(n5862), .ZN(n5863) );
  AOI22_X1 U7020 ( .A1(n8097), .A2(\adder_stage1[9][4] ), .B1(n8209), .B2(
        n5863), .ZN(n5864) );
  INV_X1 U7021 ( .A(n5864), .ZN(n10015) );
  OAI21_X1 U7022 ( .B1(n8193), .B2(n5866), .A(n5865), .ZN(n5870) );
  NAND2_X1 U7023 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U7024 ( .A(n5870), .B(n5869), .ZN(n5871) );
  AOI22_X1 U7025 ( .A1(n7525), .A2(\adder_stage2[3][12] ), .B1(n8292), .B2(
        n5871), .ZN(n5872) );
  INV_X1 U7026 ( .A(n5872), .ZN(n9841) );
  INV_X1 U7027 ( .A(n5873), .ZN(n5875) );
  NAND2_X1 U7028 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  XOR2_X1 U7029 ( .A(n5877), .B(n5876), .Z(n5878) );
  AOI22_X1 U7030 ( .A1(n7698), .A2(\adder_stage1[6][9] ), .B1(n5981), .B2(
        n5878), .ZN(n5879) );
  INV_X1 U7031 ( .A(n5879), .ZN(n10061) );
  INV_X1 U7032 ( .A(n5880), .ZN(n5896) );
  OAI21_X1 U7033 ( .B1(n5896), .B2(n5892), .A(n5893), .ZN(n5885) );
  INV_X1 U7034 ( .A(n5881), .ZN(n5883) );
  NAND2_X1 U7035 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  XNOR2_X1 U7036 ( .A(n5885), .B(n5884), .ZN(n5886) );
  AOI22_X1 U7037 ( .A1(n8168), .A2(\adder_stage1[6][3] ), .B1(n5981), .B2(
        n5886), .ZN(n5887) );
  INV_X1 U7038 ( .A(n5887), .ZN(n10067) );
  INV_X1 U7039 ( .A(n5888), .ZN(n5945) );
  NAND2_X1 U7040 ( .A1(n5945), .A2(n5943), .ZN(n5889) );
  XNOR2_X1 U7041 ( .A(n5946), .B(n5889), .ZN(n5890) );
  AOI22_X1 U7042 ( .A1(n7556), .A2(\adder_stage1[6][4] ), .B1(n5981), .B2(
        n5890), .ZN(n5891) );
  INV_X1 U7043 ( .A(n5891), .ZN(n10066) );
  INV_X1 U7044 ( .A(n5892), .ZN(n5894) );
  NAND2_X1 U7045 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  XOR2_X1 U7046 ( .A(n5896), .B(n5895), .Z(n5897) );
  AOI22_X1 U7047 ( .A1(n8097), .A2(\adder_stage1[6][2] ), .B1(n5981), .B2(
        n5897), .ZN(n5898) );
  INV_X1 U7048 ( .A(n5898), .ZN(n10068) );
  AOI21_X1 U7049 ( .B1(n5901), .B2(n5900), .A(n5899), .ZN(n5908) );
  INV_X1 U7050 ( .A(n5907), .ZN(n5902) );
  NAND2_X1 U7051 ( .A1(n5902), .A2(n5906), .ZN(n5903) );
  XOR2_X1 U7052 ( .A(n5908), .B(n5903), .Z(n5904) );
  AOI22_X1 U7053 ( .A1(n8097), .A2(\adder_stage1[9][6] ), .B1(n8209), .B2(
        n5904), .ZN(n5905) );
  INV_X1 U7054 ( .A(n5905), .ZN(n10013) );
  OAI21_X1 U7055 ( .B1(n5908), .B2(n5907), .A(n5906), .ZN(n5913) );
  INV_X1 U7056 ( .A(n5909), .ZN(n5911) );
  NAND2_X1 U7057 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  XNOR2_X1 U7058 ( .A(n5913), .B(n5912), .ZN(n5914) );
  AOI22_X1 U7059 ( .A1(n8097), .A2(\adder_stage1[9][7] ), .B1(n8209), .B2(
        n5914), .ZN(n5915) );
  INV_X1 U7060 ( .A(n5915), .ZN(n10012) );
  INV_X1 U7061 ( .A(n5916), .ZN(n5966) );
  OAI21_X1 U7062 ( .B1(n5966), .B2(n5917), .A(n5963), .ZN(n5921) );
  NAND2_X1 U7063 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  XNOR2_X1 U7064 ( .A(n5921), .B(n5920), .ZN(n5922) );
  AOI22_X1 U7065 ( .A1(n8325), .A2(\adder_stage2[3][9] ), .B1(n7627), .B2(
        n5922), .ZN(n5923) );
  INV_X1 U7066 ( .A(n5923), .ZN(n9844) );
  INV_X1 U7067 ( .A(n5924), .ZN(n5926) );
  NAND2_X1 U7068 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  XOR2_X1 U7069 ( .A(n5928), .B(n5927), .Z(n5929) );
  AOI22_X1 U7070 ( .A1(n7855), .A2(\adder_stage1[6][6] ), .B1(n5981), .B2(
        n5929), .ZN(n5930) );
  INV_X1 U7071 ( .A(n5930), .ZN(n10064) );
  NAND2_X1 U7072 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  XNOR2_X1 U7073 ( .A(n5934), .B(n5933), .ZN(n5935) );
  AOI22_X1 U7074 ( .A1(n8097), .A2(\adder_stage1[9][8] ), .B1(n8209), .B2(
        n5935), .ZN(n5936) );
  INV_X1 U7075 ( .A(n5936), .ZN(n10011) );
  INV_X1 U7076 ( .A(n5937), .ZN(n5939) );
  NAND2_X1 U7077 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  XOR2_X1 U7078 ( .A(n5940), .B(n5978), .Z(n5941) );
  AOI22_X1 U7079 ( .A1(n7855), .A2(\adder_stage1[6][1] ), .B1(n5981), .B2(
        n5941), .ZN(n5942) );
  INV_X1 U7080 ( .A(n5942), .ZN(n10069) );
  INV_X1 U7081 ( .A(n5943), .ZN(n5944) );
  AOI21_X1 U7082 ( .B1(n5946), .B2(n5945), .A(n5944), .ZN(n5951) );
  INV_X1 U7083 ( .A(n5947), .ZN(n5949) );
  NAND2_X1 U7084 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  XOR2_X1 U7085 ( .A(n5951), .B(n5950), .Z(n5952) );
  AOI22_X1 U7086 ( .A1(n7041), .A2(\adder_stage1[6][5] ), .B1(n5981), .B2(
        n5952), .ZN(n5953) );
  INV_X1 U7087 ( .A(n5953), .ZN(n10065) );
  OAI21_X1 U7088 ( .B1(n5966), .B2(n5955), .A(n5954), .ZN(n5960) );
  INV_X1 U7089 ( .A(n5956), .ZN(n5958) );
  NAND2_X1 U7090 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7091 ( .A(n5960), .B(n5959), .ZN(n5961) );
  AOI22_X1 U7092 ( .A1(n6273), .A2(\adder_stage2[3][10] ), .B1(n5981), .B2(
        n5961), .ZN(n5962) );
  INV_X1 U7093 ( .A(n5962), .ZN(n9843) );
  NAND2_X1 U7094 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  XOR2_X1 U7095 ( .A(n5966), .B(n5965), .Z(n5967) );
  AOI22_X1 U7096 ( .A1(n8330), .A2(\adder_stage2[3][8] ), .B1(n6279), .B2(
        n5967), .ZN(n5968) );
  INV_X1 U7097 ( .A(n5968), .ZN(n9845) );
  OAI21_X1 U7098 ( .B1(n8193), .B2(n5970), .A(n5969), .ZN(n5971) );
  INV_X1 U7099 ( .A(n5971), .ZN(n5975) );
  NAND2_X1 U7100 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  XOR2_X1 U7101 ( .A(n5975), .B(n5974), .Z(n5976) );
  AOI22_X1 U7102 ( .A1(n7920), .A2(\adder_stage2[3][13] ), .B1(n6626), .B2(
        n5976), .ZN(n5977) );
  INV_X1 U7103 ( .A(n5977), .ZN(n9840) );
  OR2_X1 U7104 ( .A1(\x_mult_f[12][0] ), .A2(\x_mult_f[13][0] ), .ZN(n5979) );
  AND2_X1 U7105 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  AOI22_X1 U7106 ( .A1(n8057), .A2(\adder_stage1[6][0] ), .B1(n5981), .B2(
        n5980), .ZN(n5982) );
  INV_X1 U7107 ( .A(n5982), .ZN(n10070) );
  OAI21_X1 U7108 ( .B1(n8202), .B2(n5983), .A(n5990), .ZN(n5987) );
  NAND2_X1 U7109 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  XNOR2_X1 U7110 ( .A(n5987), .B(n5986), .ZN(n5988) );
  AOI22_X1 U7111 ( .A1(n8306), .A2(\adder_stage2[4][12] ), .B1(n8209), .B2(
        n5988), .ZN(n5989) );
  INV_X1 U7112 ( .A(n5989), .ZN(n9824) );
  NAND2_X1 U7113 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  XOR2_X1 U7114 ( .A(n8202), .B(n5992), .Z(n5993) );
  AOI22_X1 U7115 ( .A1(n8313), .A2(\adder_stage2[4][11] ), .B1(n8209), .B2(
        n5993), .ZN(n5994) );
  INV_X1 U7116 ( .A(n5994), .ZN(n9825) );
  OAI21_X1 U7117 ( .B1(n5997), .B2(n5996), .A(n5995), .ZN(n6002) );
  INV_X1 U7118 ( .A(n5998), .ZN(n6000) );
  NAND2_X1 U7119 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  XNOR2_X1 U7120 ( .A(n6002), .B(n6001), .ZN(n6003) );
  AOI22_X1 U7121 ( .A1(n8168), .A2(\adder_stage2[4][10] ), .B1(n8209), .B2(
        n6003), .ZN(n6004) );
  INV_X1 U7122 ( .A(n6004), .ZN(n9826) );
  NAND2_X1 U7123 ( .A1(n7454), .A2(n6005), .ZN(n6006) );
  XNOR2_X1 U7124 ( .A(n3435), .B(n6006), .ZN(n6007) );
  AOI22_X1 U7125 ( .A1(n8057), .A2(\adder_stage1[12][8] ), .B1(n8105), .B2(
        n6007), .ZN(n6008) );
  INV_X1 U7126 ( .A(n6008), .ZN(n9961) );
  AOI21_X1 U7127 ( .B1(n6021), .B2(n6010), .A(n6009), .ZN(n6033) );
  OAI21_X1 U7128 ( .B1(n6033), .B2(n6029), .A(n6030), .ZN(n6015) );
  INV_X1 U7129 ( .A(n6011), .ZN(n6013) );
  NAND2_X1 U7130 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  XNOR2_X1 U7131 ( .A(n6015), .B(n6014), .ZN(n6016) );
  AOI22_X1 U7132 ( .A1(n7041), .A2(\adder_stage1[12][7] ), .B1(n8209), .B2(
        n6016), .ZN(n6017) );
  INV_X1 U7133 ( .A(n6017), .ZN(n9962) );
  INV_X1 U7134 ( .A(n6018), .ZN(n6019) );
  AOI21_X1 U7135 ( .B1(n6021), .B2(n6020), .A(n6019), .ZN(n6026) );
  INV_X1 U7136 ( .A(n6022), .ZN(n6024) );
  NAND2_X1 U7137 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  XOR2_X1 U7138 ( .A(n6026), .B(n6025), .Z(n6027) );
  AOI22_X1 U7139 ( .A1(n7669), .A2(\adder_stage1[12][5] ), .B1(n6036), .B2(
        n6027), .ZN(n6028) );
  INV_X1 U7140 ( .A(n6028), .ZN(n9964) );
  INV_X1 U7141 ( .A(n6029), .ZN(n6031) );
  NAND2_X1 U7142 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  XOR2_X1 U7143 ( .A(n6033), .B(n6032), .Z(n6034) );
  AOI22_X1 U7144 ( .A1(n6854), .A2(\adder_stage1[12][6] ), .B1(n4645), .B2(
        n6034), .ZN(n6035) );
  INV_X1 U7145 ( .A(n6035), .ZN(n9963) );
  AOI22_X1 U7146 ( .A1(n8398), .A2(\x_mult_f[0][2] ), .B1(n6036), .B2(
        \x_mult_f_int[0][2] ), .ZN(n6037) );
  INV_X1 U7147 ( .A(n6037), .ZN(n8926) );
  BUF_X2 U7148 ( .A(n4671), .Z(n7507) );
  AOI22_X1 U7149 ( .A1(n8168), .A2(\x_mult_f[17][3] ), .B1(n7507), .B2(
        \x_mult_f_int[17][3] ), .ZN(n6038) );
  INV_X1 U7150 ( .A(n6038), .ZN(n9138) );
  NAND2_X1 U7151 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  XNOR2_X1 U7152 ( .A(n6042), .B(n6041), .ZN(n6043) );
  AOI22_X1 U7153 ( .A1(n8168), .A2(\adder_stage1[8][12] ), .B1(n7507), .B2(
        n6043), .ZN(n6044) );
  INV_X1 U7154 ( .A(n6044), .ZN(n10024) );
  AOI22_X1 U7155 ( .A1(n8168), .A2(\x_mult_f[17][4] ), .B1(n7507), .B2(
        \x_mult_f_int[17][4] ), .ZN(n6045) );
  INV_X1 U7156 ( .A(n6045), .ZN(n9137) );
  AOI22_X1 U7157 ( .A1(n8168), .A2(\x_mult_f[17][1] ), .B1(n7507), .B2(
        \x_mult_f_int[17][1] ), .ZN(n6046) );
  INV_X1 U7158 ( .A(n6046), .ZN(n9360) );
  AOI22_X1 U7159 ( .A1(n8168), .A2(\x_mult_f[16][1] ), .B1(n7507), .B2(
        \x_mult_f_int[16][1] ), .ZN(n6047) );
  INV_X1 U7160 ( .A(n6047), .ZN(n9358) );
  AOI22_X1 U7161 ( .A1(n8168), .A2(\x_mult_f[17][2] ), .B1(n7507), .B2(
        \x_mult_f_int[17][2] ), .ZN(n6048) );
  INV_X1 U7162 ( .A(n6048), .ZN(n9139) );
  AOI22_X1 U7163 ( .A1(n8168), .A2(\x_mult_f[17][5] ), .B1(n7507), .B2(
        \x_mult_f_int[17][5] ), .ZN(n6049) );
  INV_X1 U7164 ( .A(n6049), .ZN(n9136) );
  AOI22_X1 U7165 ( .A1(n8168), .A2(\x_mult_f[17][0] ), .B1(n7507), .B2(
        \x_mult_f_int[17][0] ), .ZN(n6050) );
  INV_X1 U7166 ( .A(n6050), .ZN(n9361) );
  AOI22_X1 U7167 ( .A1(n8168), .A2(\x_mult_f[16][0] ), .B1(n7507), .B2(
        \x_mult_f_int[16][0] ), .ZN(n6051) );
  INV_X1 U7168 ( .A(n6051), .ZN(n9359) );
  AOI22_X1 U7169 ( .A1(n7959), .A2(\x_mult_f[28][3] ), .B1(n5707), .B2(
        \x_mult_f_int[28][3] ), .ZN(n6052) );
  INV_X1 U7170 ( .A(n6052), .ZN(n9284) );
  AOI22_X1 U7171 ( .A1(n7928), .A2(\x_mult_f[28][1] ), .B1(n8078), .B2(
        \x_mult_f_int[28][1] ), .ZN(n6053) );
  INV_X1 U7172 ( .A(n6053), .ZN(n9382) );
  AOI22_X1 U7173 ( .A1(n8057), .A2(\x_mult_f[28][2] ), .B1(n4444), .B2(
        \x_mult_f_int[28][2] ), .ZN(n6054) );
  INV_X1 U7174 ( .A(n6054), .ZN(n9285) );
  OAI21_X1 U7175 ( .B1(n6057), .B2(n6056), .A(n6055), .ZN(n7749) );
  AOI22_X1 U7176 ( .A1(n6058), .A2(n7155), .B1(n8306), .B2(
        \adder_stage1[4][14] ), .ZN(n6059) );
  INV_X1 U7177 ( .A(n6059), .ZN(n10089) );
  INV_X1 U7178 ( .A(n6060), .ZN(n6061) );
  AOI21_X1 U7179 ( .B1(n3422), .B2(n6062), .A(n6061), .ZN(n6070) );
  NOR2_X1 U7180 ( .A1(\x_mult_f[0][13] ), .A2(\x_mult_f[1][13] ), .ZN(n6069)
         );
  INV_X1 U7181 ( .A(n6069), .ZN(n6064) );
  NAND2_X1 U7182 ( .A1(\x_mult_f[0][13] ), .A2(\x_mult_f[1][13] ), .ZN(n6068)
         );
  NAND2_X1 U7183 ( .A1(n6064), .A2(n6068), .ZN(n6065) );
  XOR2_X1 U7184 ( .A(n6070), .B(n6065), .Z(n6066) );
  AOI22_X1 U7185 ( .A1(n6066), .A2(n8054), .B1(n8340), .B2(
        \adder_stage1[0][13] ), .ZN(n6067) );
  INV_X1 U7186 ( .A(n6067), .ZN(n10156) );
  OAI21_X1 U7187 ( .B1(n3431), .B2(n6069), .A(n6068), .ZN(n7727) );
  AOI22_X1 U7188 ( .A1(n6071), .A2(n4311), .B1(n7669), .B2(
        \adder_stage1[0][14] ), .ZN(n6072) );
  INV_X1 U7189 ( .A(n6072), .ZN(n10155) );
  OAI21_X1 U7190 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(n6080) );
  INV_X1 U7191 ( .A(n6076), .ZN(n6078) );
  NAND2_X1 U7192 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  XNOR2_X1 U7193 ( .A(n6080), .B(n6079), .ZN(n6081) );
  AOI22_X1 U7194 ( .A1(n7614), .A2(\adder_stage1[10][7] ), .B1(n4444), .B2(
        n6081), .ZN(n6082) );
  INV_X1 U7195 ( .A(n6082), .ZN(n9996) );
  NAND2_X1 U7196 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  XNOR2_X1 U7197 ( .A(n6086), .B(n6085), .ZN(n6087) );
  AOI22_X1 U7198 ( .A1(n7614), .A2(\adder_stage1[10][8] ), .B1(n4444), .B2(
        n6087), .ZN(n6088) );
  INV_X1 U7199 ( .A(n6088), .ZN(n9995) );
  OR2_X1 U7200 ( .A1(\adder_stage3[0][0] ), .A2(\adder_stage3[1][0] ), .ZN(
        n6090) );
  AND2_X1 U7201 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  AOI22_X1 U7202 ( .A1(n7622), .A2(\adder_stage4[0][0] ), .B1(n7507), .B2(
        n6091), .ZN(n6092) );
  INV_X1 U7203 ( .A(n6092), .ZN(n9687) );
  BUF_X2 U7204 ( .A(n4444), .Z(n6609) );
  NOR2_X1 U7205 ( .A1(\adder_stage1[10][2] ), .A2(\adder_stage1[11][2] ), .ZN(
        n6229) );
  NOR2_X1 U7206 ( .A1(\adder_stage1[10][3] ), .A2(\adder_stage1[11][3] ), .ZN(
        n6231) );
  NOR2_X1 U7207 ( .A1(n6229), .A2(n6231), .ZN(n6095) );
  NOR2_X1 U7208 ( .A1(\adder_stage1[10][1] ), .A2(\adder_stage1[11][1] ), .ZN(
        n6218) );
  NAND2_X1 U7209 ( .A1(\adder_stage1[10][0] ), .A2(\adder_stage1[11][0] ), 
        .ZN(n6224) );
  NAND2_X1 U7210 ( .A1(\adder_stage1[10][1] ), .A2(\adder_stage1[11][1] ), 
        .ZN(n6219) );
  OAI21_X1 U7211 ( .B1(n6218), .B2(n6224), .A(n6219), .ZN(n6213) );
  NAND2_X1 U7212 ( .A1(\adder_stage1[10][2] ), .A2(\adder_stage1[11][2] ), 
        .ZN(n6228) );
  NAND2_X1 U7213 ( .A1(\adder_stage1[10][3] ), .A2(\adder_stage1[11][3] ), 
        .ZN(n6232) );
  OAI21_X1 U7214 ( .B1(n6231), .B2(n6228), .A(n6232), .ZN(n6094) );
  AOI21_X1 U7215 ( .B1(n6095), .B2(n6213), .A(n6094), .ZN(n6106) );
  INV_X1 U7216 ( .A(n6106), .ZN(n6122) );
  NOR2_X1 U7217 ( .A1(\adder_stage1[10][4] ), .A2(\adder_stage1[11][4] ), .ZN(
        n6110) );
  NOR2_X1 U7218 ( .A1(\adder_stage1[10][5] ), .A2(\adder_stage1[11][5] ), .ZN(
        n6112) );
  NOR2_X1 U7219 ( .A1(n6110), .A2(n6112), .ZN(n6100) );
  NAND2_X1 U7220 ( .A1(\adder_stage1[10][4] ), .A2(\adder_stage1[11][4] ), 
        .ZN(n6119) );
  NAND2_X1 U7221 ( .A1(\adder_stage1[10][5] ), .A2(\adder_stage1[11][5] ), 
        .ZN(n6113) );
  OAI21_X1 U7222 ( .B1(n6112), .B2(n6119), .A(n6113), .ZN(n6102) );
  AOI21_X1 U7223 ( .B1(n6122), .B2(n6100), .A(n6102), .ZN(n6170) );
  NOR2_X1 U7224 ( .A1(\adder_stage1[10][6] ), .A2(\adder_stage1[11][6] ), .ZN(
        n6169) );
  INV_X1 U7225 ( .A(n6169), .ZN(n6096) );
  NAND2_X1 U7226 ( .A1(\adder_stage1[10][6] ), .A2(\adder_stage1[11][6] ), 
        .ZN(n6168) );
  NAND2_X1 U7227 ( .A1(n6096), .A2(n6168), .ZN(n6097) );
  XOR2_X1 U7228 ( .A(n6170), .B(n6097), .Z(n6098) );
  AOI22_X1 U7229 ( .A1(n8168), .A2(\adder_stage2[5][6] ), .B1(n6609), .B2(
        n6098), .ZN(n6099) );
  INV_X1 U7230 ( .A(n6099), .ZN(n9813) );
  NOR2_X1 U7231 ( .A1(\adder_stage1[10][7] ), .A2(\adder_stage1[11][7] ), .ZN(
        n6171) );
  NOR2_X1 U7232 ( .A1(n6169), .A2(n6171), .ZN(n6103) );
  NAND2_X1 U7233 ( .A1(n6100), .A2(n6103), .ZN(n6105) );
  NAND2_X1 U7234 ( .A1(\adder_stage1[10][7] ), .A2(\adder_stage1[11][7] ), 
        .ZN(n6172) );
  OAI21_X1 U7235 ( .B1(n6171), .B2(n6168), .A(n6172), .ZN(n6101) );
  AOI21_X1 U7236 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(n6104) );
  OAI21_X1 U7237 ( .B1(n6106), .B2(n6105), .A(n6104), .ZN(n6149) );
  INV_X1 U7238 ( .A(n6149), .ZN(n6242) );
  NOR2_X1 U7239 ( .A1(\adder_stage1[10][8] ), .A2(\adder_stage1[11][8] ), .ZN(
        n6125) );
  INV_X1 U7240 ( .A(n6125), .ZN(n6141) );
  NAND2_X1 U7241 ( .A1(\adder_stage1[10][8] ), .A2(\adder_stage1[11][8] ), 
        .ZN(n6142) );
  NAND2_X1 U7242 ( .A1(n6141), .A2(n6142), .ZN(n6107) );
  XOR2_X1 U7243 ( .A(n6242), .B(n6107), .Z(n6108) );
  AOI22_X1 U7244 ( .A1(n6854), .A2(\adder_stage2[5][8] ), .B1(n6609), .B2(
        n6108), .ZN(n6109) );
  INV_X1 U7245 ( .A(n6109), .ZN(n9811) );
  INV_X1 U7246 ( .A(n6110), .ZN(n6120) );
  INV_X1 U7247 ( .A(n6119), .ZN(n6111) );
  AOI21_X1 U7248 ( .B1(n6122), .B2(n6120), .A(n6111), .ZN(n6116) );
  INV_X1 U7249 ( .A(n6112), .ZN(n6114) );
  NAND2_X1 U7250 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  XOR2_X1 U7251 ( .A(n6116), .B(n6115), .Z(n6117) );
  AOI22_X1 U7252 ( .A1(n8118), .A2(\adder_stage2[5][5] ), .B1(n6609), .B2(
        n6117), .ZN(n6118) );
  INV_X1 U7253 ( .A(n6118), .ZN(n9814) );
  NAND2_X1 U7254 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  XNOR2_X1 U7255 ( .A(n6122), .B(n6121), .ZN(n6123) );
  AOI22_X1 U7256 ( .A1(n7074), .A2(\adder_stage2[5][4] ), .B1(n6609), .B2(
        n6123), .ZN(n6124) );
  INV_X1 U7257 ( .A(n6124), .ZN(n9815) );
  BUF_X2 U7258 ( .A(n4645), .Z(n8216) );
  OAI21_X1 U7259 ( .B1(n6242), .B2(n6125), .A(n6142), .ZN(n6127) );
  OR2_X1 U7260 ( .A1(\adder_stage1[10][9] ), .A2(\adder_stage1[11][9] ), .ZN(
        n6146) );
  NAND2_X1 U7261 ( .A1(\adder_stage1[10][9] ), .A2(\adder_stage1[11][9] ), 
        .ZN(n6143) );
  NAND2_X1 U7262 ( .A1(n6146), .A2(n6143), .ZN(n6126) );
  XNOR2_X1 U7263 ( .A(n6127), .B(n6126), .ZN(n6128) );
  AOI22_X1 U7264 ( .A1(n8336), .A2(\adder_stage2[5][9] ), .B1(n8216), .B2(
        n6128), .ZN(n6129) );
  INV_X1 U7265 ( .A(n6129), .ZN(n9810) );
  BUF_X2 U7266 ( .A(n6238), .Z(n6626) );
  INV_X1 U7267 ( .A(n6130), .ZN(n7081) );
  INV_X1 U7268 ( .A(n7080), .ZN(n6131) );
  NAND2_X1 U7269 ( .A1(n6131), .A2(n7079), .ZN(n6132) );
  XOR2_X1 U7270 ( .A(n7081), .B(n6132), .Z(n6133) );
  AOI22_X1 U7271 ( .A1(n8057), .A2(\adder_stage3[3][2] ), .B1(n6626), .B2(
        n6133), .ZN(n6134) );
  INV_X1 U7272 ( .A(n6134), .ZN(n9706) );
  INV_X1 U7273 ( .A(n6135), .ZN(n6137) );
  NAND2_X1 U7274 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  XOR2_X1 U7275 ( .A(n6138), .B(n6178), .Z(n6139) );
  AOI22_X1 U7276 ( .A1(n8088), .A2(\adder_stage3[3][1] ), .B1(n6626), .B2(
        n6139), .ZN(n6140) );
  INV_X1 U7277 ( .A(n6140), .ZN(n9707) );
  NAND2_X1 U7278 ( .A1(n6141), .A2(n6146), .ZN(n6241) );
  NOR2_X1 U7279 ( .A1(\adder_stage1[10][10] ), .A2(\adder_stage1[11][10] ), 
        .ZN(n6243) );
  NOR2_X1 U7280 ( .A1(n6241), .A2(n6243), .ZN(n6148) );
  INV_X1 U7281 ( .A(n6142), .ZN(n6145) );
  INV_X1 U7282 ( .A(n6143), .ZN(n6144) );
  AOI21_X1 U7283 ( .B1(n6146), .B2(n6145), .A(n6144), .ZN(n6240) );
  NAND2_X1 U7284 ( .A1(\adder_stage1[10][10] ), .A2(\adder_stage1[11][10] ), 
        .ZN(n6244) );
  OAI21_X1 U7285 ( .B1(n6240), .B2(n6243), .A(n6244), .ZN(n6147) );
  AOI21_X1 U7286 ( .B1(n6149), .B2(n6148), .A(n6147), .ZN(n6156) );
  NOR2_X1 U7287 ( .A1(\adder_stage1[10][11] ), .A2(\adder_stage1[11][11] ), 
        .ZN(n6155) );
  INV_X1 U7288 ( .A(n6155), .ZN(n6150) );
  NAND2_X1 U7289 ( .A1(\adder_stage1[10][11] ), .A2(\adder_stage1[11][11] ), 
        .ZN(n6154) );
  NAND2_X1 U7290 ( .A1(n6150), .A2(n6154), .ZN(n6151) );
  XOR2_X1 U7291 ( .A(n3437), .B(n6151), .Z(n6152) );
  AOI22_X1 U7292 ( .A1(n8168), .A2(\adder_stage2[5][11] ), .B1(n8216), .B2(
        n6152), .ZN(n6153) );
  INV_X1 U7293 ( .A(n6153), .ZN(n9808) );
  OAI21_X1 U7294 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(n6163) );
  OR2_X1 U7295 ( .A1(\adder_stage1[10][12] ), .A2(\adder_stage1[11][12] ), 
        .ZN(n6162) );
  NAND2_X1 U7296 ( .A1(\adder_stage1[10][12] ), .A2(\adder_stage1[11][12] ), 
        .ZN(n6160) );
  NAND2_X1 U7297 ( .A1(n6162), .A2(n6160), .ZN(n6157) );
  XNOR2_X1 U7298 ( .A(n6163), .B(n6157), .ZN(n6158) );
  AOI22_X1 U7299 ( .A1(n6877), .A2(\adder_stage2[5][12] ), .B1(n8216), .B2(
        n6158), .ZN(n6159) );
  INV_X1 U7300 ( .A(n6159), .ZN(n9807) );
  INV_X1 U7301 ( .A(n6160), .ZN(n6161) );
  AOI21_X1 U7302 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n7159) );
  NOR2_X1 U7303 ( .A1(\adder_stage1[10][13] ), .A2(\adder_stage1[11][13] ), 
        .ZN(n7158) );
  INV_X1 U7304 ( .A(n7158), .ZN(n6164) );
  NAND2_X1 U7305 ( .A1(\adder_stage1[10][13] ), .A2(\adder_stage1[11][13] ), 
        .ZN(n7157) );
  NAND2_X1 U7306 ( .A1(n6164), .A2(n7157), .ZN(n6165) );
  XOR2_X1 U7307 ( .A(n3436), .B(n6165), .Z(n6166) );
  AOI22_X1 U7308 ( .A1(n8273), .A2(\adder_stage2[5][13] ), .B1(n8216), .B2(
        n6166), .ZN(n6167) );
  INV_X1 U7309 ( .A(n6167), .ZN(n9806) );
  OAI21_X1 U7310 ( .B1(n6170), .B2(n6169), .A(n6168), .ZN(n6175) );
  INV_X1 U7311 ( .A(n6171), .ZN(n6173) );
  NAND2_X1 U7312 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  XNOR2_X1 U7313 ( .A(n6175), .B(n6174), .ZN(n6176) );
  AOI22_X1 U7314 ( .A1(n7525), .A2(\adder_stage2[5][7] ), .B1(n6609), .B2(
        n6176), .ZN(n6177) );
  INV_X1 U7315 ( .A(n6177), .ZN(n9812) );
  OR2_X1 U7316 ( .A1(\adder_stage2[6][0] ), .A2(\adder_stage2[7][0] ), .ZN(
        n6179) );
  AND2_X1 U7317 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  AOI22_X1 U7318 ( .A1(n8057), .A2(\adder_stage3[3][0] ), .B1(n6626), .B2(
        n6180), .ZN(n6181) );
  INV_X1 U7319 ( .A(n6181), .ZN(n9708) );
  NOR2_X1 U7320 ( .A1(n6182), .A2(n6185), .ZN(n6684) );
  NOR2_X1 U7321 ( .A1(\adder_stage3[2][6] ), .A2(\adder_stage3[3][6] ), .ZN(
        n8284) );
  NOR2_X1 U7322 ( .A1(\adder_stage3[2][7] ), .A2(\adder_stage3[3][7] ), .ZN(
        n8286) );
  NOR2_X1 U7323 ( .A1(n8284), .A2(n8286), .ZN(n6187) );
  NAND2_X1 U7324 ( .A1(n6684), .A2(n6187), .ZN(n6189) );
  OAI21_X1 U7325 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(n6683) );
  NAND2_X1 U7326 ( .A1(\adder_stage3[2][6] ), .A2(\adder_stage3[3][6] ), .ZN(
        n8283) );
  NAND2_X1 U7327 ( .A1(\adder_stage3[2][7] ), .A2(\adder_stage3[3][7] ), .ZN(
        n8287) );
  OAI21_X1 U7328 ( .B1(n8286), .B2(n8283), .A(n8287), .ZN(n6186) );
  AOI21_X1 U7329 ( .B1(n6187), .B2(n6683), .A(n6186), .ZN(n6188) );
  OAI21_X1 U7330 ( .B1(n6190), .B2(n6189), .A(n6188), .ZN(n6650) );
  NOR2_X1 U7331 ( .A1(\adder_stage3[2][8] ), .A2(\adder_stage3[3][8] ), .ZN(
        n6677) );
  NOR2_X1 U7332 ( .A1(\adder_stage3[2][9] ), .A2(\adder_stage3[3][9] ), .ZN(
        n6651) );
  NOR2_X1 U7333 ( .A1(n6677), .A2(n6651), .ZN(n6658) );
  NOR2_X1 U7334 ( .A1(\adder_stage3[3][11] ), .A2(\adder_stage3[2][11] ), .ZN(
        n6664) );
  NOR2_X1 U7335 ( .A1(\adder_stage3[2][10] ), .A2(\adder_stage3[3][10] ), .ZN(
        n6662) );
  NOR2_X1 U7336 ( .A1(n6664), .A2(n6662), .ZN(n6192) );
  NAND2_X1 U7337 ( .A1(n6658), .A2(n6192), .ZN(n6691) );
  NOR2_X1 U7338 ( .A1(\adder_stage3[2][12] ), .A2(\adder_stage3[3][12] ), .ZN(
        n6693) );
  NOR2_X1 U7339 ( .A1(n6691), .A2(n6693), .ZN(n6194) );
  NAND2_X1 U7340 ( .A1(\adder_stage3[2][8] ), .A2(\adder_stage3[3][8] ), .ZN(
        n6678) );
  NAND2_X1 U7341 ( .A1(\adder_stage3[2][9] ), .A2(\adder_stage3[3][9] ), .ZN(
        n6652) );
  OAI21_X1 U7342 ( .B1(n6651), .B2(n6678), .A(n6652), .ZN(n6659) );
  NAND2_X1 U7343 ( .A1(\adder_stage3[2][10] ), .A2(\adder_stage3[3][10] ), 
        .ZN(n6671) );
  NAND2_X1 U7344 ( .A1(\adder_stage3[2][11] ), .A2(\adder_stage3[3][11] ), 
        .ZN(n6665) );
  OAI21_X1 U7345 ( .B1(n6664), .B2(n6671), .A(n6665), .ZN(n6191) );
  AOI21_X1 U7346 ( .B1(n6192), .B2(n6659), .A(n6191), .ZN(n6690) );
  NAND2_X1 U7347 ( .A1(\adder_stage3[2][12] ), .A2(\adder_stage3[3][12] ), 
        .ZN(n6694) );
  OAI21_X1 U7348 ( .B1(n6690), .B2(n6693), .A(n6694), .ZN(n6193) );
  AOI21_X1 U7349 ( .B1(n6650), .B2(n6194), .A(n6193), .ZN(n6210) );
  NOR2_X1 U7350 ( .A1(\adder_stage3[2][13] ), .A2(\adder_stage3[3][13] ), .ZN(
        n6206) );
  NAND2_X1 U7351 ( .A1(\adder_stage3[2][13] ), .A2(\adder_stage3[3][13] ), 
        .ZN(n6207) );
  OAI21_X1 U7352 ( .B1(n6210), .B2(n6206), .A(n6207), .ZN(n6253) );
  OR2_X1 U7353 ( .A1(\adder_stage3[2][14] ), .A2(\adder_stage3[3][14] ), .ZN(
        n6251) );
  NAND2_X1 U7354 ( .A1(\adder_stage3[2][14] ), .A2(\adder_stage3[3][14] ), 
        .ZN(n6250) );
  INV_X1 U7355 ( .A(n6250), .ZN(n6195) );
  AOI21_X1 U7356 ( .B1(n6253), .B2(n6251), .A(n6195), .ZN(n6202) );
  NOR2_X1 U7357 ( .A1(\adder_stage3[2][15] ), .A2(\adder_stage3[3][15] ), .ZN(
        n6201) );
  INV_X1 U7358 ( .A(n6201), .ZN(n6196) );
  NAND2_X1 U7359 ( .A1(\adder_stage3[2][15] ), .A2(\adder_stage3[3][15] ), 
        .ZN(n6200) );
  NAND2_X1 U7360 ( .A1(n6196), .A2(n6200), .ZN(n6197) );
  XOR2_X1 U7361 ( .A(n6202), .B(n6197), .Z(n6198) );
  AOI22_X1 U7362 ( .A1(n8088), .A2(\adder_stage4[1][15] ), .B1(n6626), .B2(
        n6198), .ZN(n6199) );
  INV_X1 U7363 ( .A(n6199), .ZN(n9651) );
  OAI21_X1 U7364 ( .B1(n6202), .B2(n6201), .A(n6200), .ZN(n8137) );
  OR2_X1 U7365 ( .A1(\adder_stage3[2][16] ), .A2(\adder_stage3[3][16] ), .ZN(
        n8136) );
  NAND2_X1 U7366 ( .A1(\adder_stage3[2][16] ), .A2(\adder_stage3[3][16] ), 
        .ZN(n6446) );
  NAND2_X1 U7367 ( .A1(n8136), .A2(n6446), .ZN(n6203) );
  XNOR2_X1 U7368 ( .A(n8137), .B(n6203), .ZN(n6204) );
  AOI22_X1 U7369 ( .A1(n8057), .A2(\adder_stage4[1][16] ), .B1(n6626), .B2(
        n6204), .ZN(n6205) );
  INV_X1 U7370 ( .A(n6205), .ZN(n9650) );
  INV_X1 U7371 ( .A(n6206), .ZN(n6208) );
  NAND2_X1 U7372 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  XOR2_X1 U7373 ( .A(n6210), .B(n6209), .Z(n6211) );
  AOI22_X1 U7374 ( .A1(n8057), .A2(\adder_stage4[1][13] ), .B1(n6626), .B2(
        n6211), .ZN(n6212) );
  INV_X1 U7375 ( .A(n6212), .ZN(n9653) );
  INV_X1 U7376 ( .A(n6213), .ZN(n6230) );
  INV_X1 U7377 ( .A(n6229), .ZN(n6214) );
  NAND2_X1 U7378 ( .A1(n6214), .A2(n6228), .ZN(n6215) );
  XOR2_X1 U7379 ( .A(n6230), .B(n6215), .Z(n6216) );
  AOI22_X1 U7380 ( .A1(n7041), .A2(\adder_stage2[5][2] ), .B1(n6609), .B2(
        n6216), .ZN(n6217) );
  INV_X1 U7381 ( .A(n6217), .ZN(n9817) );
  INV_X1 U7382 ( .A(n6218), .ZN(n6220) );
  NAND2_X1 U7383 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  XOR2_X1 U7384 ( .A(n6221), .B(n6224), .Z(n6222) );
  AOI22_X1 U7385 ( .A1(n8338), .A2(\adder_stage2[5][1] ), .B1(n6609), .B2(
        n6222), .ZN(n6223) );
  INV_X1 U7386 ( .A(n6223), .ZN(n9818) );
  OR2_X1 U7387 ( .A1(\adder_stage1[10][0] ), .A2(\adder_stage1[11][0] ), .ZN(
        n6225) );
  AND2_X1 U7388 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  AOI22_X1 U7389 ( .A1(n8325), .A2(\adder_stage2[5][0] ), .B1(n6609), .B2(
        n6226), .ZN(n6227) );
  INV_X1 U7390 ( .A(n6227), .ZN(n9819) );
  OAI21_X1 U7391 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(n6235) );
  INV_X1 U7392 ( .A(n6231), .ZN(n6233) );
  NAND2_X1 U7393 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  XNOR2_X1 U7394 ( .A(n6235), .B(n6234), .ZN(n6236) );
  AOI22_X1 U7395 ( .A1(n8330), .A2(\adder_stage2[5][3] ), .B1(n6609), .B2(
        n6236), .ZN(n6237) );
  INV_X1 U7396 ( .A(n6237), .ZN(n9816) );
  BUF_X2 U7397 ( .A(n4645), .Z(n8265) );
  AOI22_X1 U7398 ( .A1(n7928), .A2(\x_mult_f[29][1] ), .B1(n8265), .B2(
        \x_mult_f_int[29][1] ), .ZN(n6239) );
  INV_X1 U7399 ( .A(n6239), .ZN(n9384) );
  OAI21_X1 U7400 ( .B1(n6242), .B2(n6241), .A(n6240), .ZN(n6247) );
  INV_X1 U7401 ( .A(n6243), .ZN(n6245) );
  NAND2_X1 U7402 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  XNOR2_X1 U7403 ( .A(n6247), .B(n6246), .ZN(n6248) );
  AOI22_X1 U7404 ( .A1(n8168), .A2(\adder_stage2[5][10] ), .B1(n8216), .B2(
        n6248), .ZN(n6249) );
  INV_X1 U7405 ( .A(n6249), .ZN(n9809) );
  NAND2_X1 U7406 ( .A1(n6251), .A2(n6250), .ZN(n6252) );
  XNOR2_X1 U7407 ( .A(n6253), .B(n6252), .ZN(n6254) );
  AOI22_X1 U7408 ( .A1(n7855), .A2(\adder_stage4[1][14] ), .B1(n6626), .B2(
        n6254), .ZN(n6255) );
  INV_X1 U7409 ( .A(n6255), .ZN(n9652) );
  AOI22_X1 U7410 ( .A1(n7928), .A2(\x_mult_f[29][2] ), .B1(n8265), .B2(
        \x_mult_f_int[29][2] ), .ZN(n6256) );
  INV_X1 U7411 ( .A(n6256), .ZN(n9299) );
  INV_X1 U7412 ( .A(n6257), .ZN(n6643) );
  OAI21_X1 U7413 ( .B1(n6643), .B2(n6639), .A(n6640), .ZN(n6262) );
  INV_X1 U7414 ( .A(n6258), .ZN(n6260) );
  NAND2_X1 U7415 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  XNOR2_X1 U7416 ( .A(n6262), .B(n6261), .ZN(n6263) );
  AOI22_X1 U7417 ( .A1(n8176), .A2(\adder_stage1[11][3] ), .B1(n8265), .B2(
        n6263), .ZN(n6264) );
  INV_X1 U7418 ( .A(n6264), .ZN(n9983) );
  BUF_X2 U7419 ( .A(n6352), .Z(n8235) );
  INV_X1 U7420 ( .A(n6265), .ZN(n8228) );
  INV_X1 U7421 ( .A(n6266), .ZN(n8227) );
  NAND2_X1 U7422 ( .A1(n8227), .A2(n8225), .ZN(n6267) );
  XNOR2_X1 U7423 ( .A(n8228), .B(n6267), .ZN(n6268) );
  AOI22_X1 U7424 ( .A1(n8245), .A2(\adder_stage3[0][4] ), .B1(n8235), .B2(
        n6268), .ZN(n6269) );
  INV_X1 U7425 ( .A(n6269), .ZN(n9765) );
  AOI22_X1 U7426 ( .A1(n6273), .A2(\x_mult_f[20][2] ), .B1(n6272), .B2(
        \x_mult_f_int[20][2] ), .ZN(n6270) );
  INV_X1 U7427 ( .A(n6270), .ZN(n9181) );
  AOI22_X1 U7428 ( .A1(n6273), .A2(\x_mult_f[20][5] ), .B1(n6272), .B2(
        \x_mult_f_int[20][5] ), .ZN(n6271) );
  INV_X1 U7429 ( .A(n6271), .ZN(n9178) );
  AOI22_X1 U7430 ( .A1(n6273), .A2(\x_mult_f[20][3] ), .B1(n6272), .B2(
        \x_mult_f_int[20][3] ), .ZN(n6274) );
  INV_X1 U7431 ( .A(n6274), .ZN(n9180) );
  OAI21_X1 U7432 ( .B1(n6277), .B2(n6276), .A(n6275), .ZN(n7925) );
  OR2_X1 U7433 ( .A1(\x_mult_f[28][12] ), .A2(\x_mult_f[29][12] ), .ZN(n7923)
         );
  NAND2_X1 U7434 ( .A1(\x_mult_f[28][12] ), .A2(\x_mult_f[29][12] ), .ZN(n7922) );
  INV_X1 U7435 ( .A(n7922), .ZN(n6278) );
  AOI21_X1 U7436 ( .B1(n7925), .B2(n7923), .A(n6278), .ZN(n7296) );
  NOR2_X1 U7437 ( .A1(\x_mult_f[28][13] ), .A2(\x_mult_f[29][13] ), .ZN(n7292)
         );
  NAND2_X1 U7438 ( .A1(\x_mult_f[28][13] ), .A2(\x_mult_f[29][13] ), .ZN(n7293) );
  OAI21_X1 U7439 ( .B1(n3426), .B2(n7292), .A(n7293), .ZN(n7704) );
  AOI22_X1 U7440 ( .A1(n6280), .A2(n7507), .B1(n8434), .B2(
        \adder_stage1[14][14] ), .ZN(n6281) );
  INV_X1 U7441 ( .A(n6281), .ZN(n9921) );
  OAI21_X1 U7442 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(n8187) );
  OR2_X1 U7443 ( .A1(\adder_stage1[2][12] ), .A2(\adder_stage1[3][12] ), .ZN(
        n8185) );
  NAND2_X1 U7444 ( .A1(\adder_stage1[2][12] ), .A2(\adder_stage1[3][12] ), 
        .ZN(n8184) );
  INV_X1 U7445 ( .A(n8184), .ZN(n6285) );
  AOI21_X1 U7446 ( .B1(n8187), .B2(n8185), .A(n6285), .ZN(n7039) );
  NOR2_X1 U7447 ( .A1(\adder_stage1[2][13] ), .A2(\adder_stage1[3][13] ), .ZN(
        n7035) );
  NAND2_X1 U7448 ( .A1(\adder_stage1[2][13] ), .A2(\adder_stage1[3][13] ), 
        .ZN(n7036) );
  OAI21_X1 U7449 ( .B1(n7039), .B2(n7035), .A(n7036), .ZN(n7032) );
  OR2_X1 U7450 ( .A1(\adder_stage1[2][14] ), .A2(\adder_stage1[3][14] ), .ZN(
        n7030) );
  NAND2_X1 U7451 ( .A1(\adder_stage1[2][14] ), .A2(\adder_stage1[3][14] ), 
        .ZN(n7029) );
  INV_X1 U7452 ( .A(n7029), .ZN(n6286) );
  XOR2_X1 U7453 ( .A(\adder_stage1[3][15] ), .B(\adder_stage1[2][15] ), .Z(
        n6287) );
  AOI22_X1 U7454 ( .A1(n6288), .A2(n6875), .B1(n8309), .B2(
        \adder_stage2[1][15] ), .ZN(n6289) );
  INV_X1 U7455 ( .A(n6289), .ZN(n9872) );
  INV_X1 U7456 ( .A(n6290), .ZN(n6292) );
  NAND2_X1 U7457 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  XOR2_X1 U7458 ( .A(n6294), .B(n6293), .Z(n6295) );
  AOI22_X1 U7459 ( .A1(n6295), .A2(n8087), .B1(n7698), .B2(
        \adder_stage1[3][13] ), .ZN(n6296) );
  INV_X1 U7460 ( .A(n6296), .ZN(n10107) );
  OR2_X1 U7461 ( .A1(\x_mult_f[26][0] ), .A2(\x_mult_f[27][0] ), .ZN(n6297) );
  AND2_X1 U7462 ( .A1(n6297), .A2(n6303), .ZN(n6298) );
  AOI22_X1 U7463 ( .A1(n8168), .A2(\adder_stage1[13][0] ), .B1(n8265), .B2(
        n6298), .ZN(n6299) );
  INV_X1 U7464 ( .A(n6299), .ZN(n9952) );
  INV_X1 U7465 ( .A(n6300), .ZN(n6302) );
  NAND2_X1 U7466 ( .A1(n6302), .A2(n6301), .ZN(n6304) );
  XOR2_X1 U7467 ( .A(n6304), .B(n6303), .Z(n6305) );
  AOI22_X1 U7468 ( .A1(n8328), .A2(\adder_stage1[13][1] ), .B1(n8265), .B2(
        n6305), .ZN(n6306) );
  INV_X1 U7469 ( .A(n6306), .ZN(n9951) );
  AOI22_X1 U7470 ( .A1(\x_mult_f_int[9][14] ), .A2(n7507), .B1(n8309), .B2(
        \x_mult_f[9][14] ), .ZN(n6308) );
  INV_X1 U7471 ( .A(n6308), .ZN(n9027) );
  BUF_X2 U7472 ( .A(n4444), .Z(n8078) );
  INV_X1 U7473 ( .A(n6309), .ZN(n6311) );
  NAND2_X1 U7474 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  XOR2_X1 U7475 ( .A(n6313), .B(n6312), .Z(n6314) );
  AOI22_X1 U7476 ( .A1(n6877), .A2(\adder_stage1[5][9] ), .B1(n8078), .B2(
        n6314), .ZN(n6315) );
  INV_X1 U7477 ( .A(n6315), .ZN(n10077) );
  NOR2_X1 U7478 ( .A1(\adder_stage1[12][1] ), .A2(\adder_stage1[13][1] ), .ZN(
        n6954) );
  INV_X1 U7479 ( .A(n6954), .ZN(n6316) );
  NAND2_X1 U7480 ( .A1(\adder_stage1[12][1] ), .A2(\adder_stage1[13][1] ), 
        .ZN(n6952) );
  NAND2_X1 U7481 ( .A1(n6316), .A2(n6952), .ZN(n6317) );
  NAND2_X1 U7482 ( .A1(\adder_stage1[12][0] ), .A2(\adder_stage1[13][0] ), 
        .ZN(n6953) );
  XOR2_X1 U7483 ( .A(n6317), .B(n6953), .Z(n6318) );
  AOI22_X1 U7484 ( .A1(n6854), .A2(\adder_stage2[6][1] ), .B1(n6626), .B2(
        n6318), .ZN(n6319) );
  INV_X1 U7485 ( .A(n6319), .ZN(n9802) );
  NAND2_X1 U7486 ( .A1(n6325), .A2(n6320), .ZN(n6321) );
  XNOR2_X1 U7487 ( .A(n8070), .B(n6321), .ZN(n6322) );
  AOI22_X1 U7488 ( .A1(n7698), .A2(\adder_stage1[5][10] ), .B1(n8078), .B2(
        n6322), .ZN(n6323) );
  INV_X1 U7489 ( .A(n6323), .ZN(n10076) );
  AOI21_X1 U7490 ( .B1(n8070), .B2(n6325), .A(n6324), .ZN(n6329) );
  NAND2_X1 U7491 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  XOR2_X1 U7492 ( .A(n6329), .B(n6328), .Z(n6330) );
  AOI22_X1 U7493 ( .A1(n7640), .A2(\adder_stage1[5][11] ), .B1(n8078), .B2(
        n6330), .ZN(n6331) );
  INV_X1 U7494 ( .A(n6331), .ZN(n10075) );
  INV_X1 U7495 ( .A(n6332), .ZN(n6334) );
  NAND2_X1 U7496 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  XOR2_X1 U7497 ( .A(n6335), .B(n7803), .Z(n6336) );
  AOI22_X1 U7498 ( .A1(n8118), .A2(\adder_stage1[11][1] ), .B1(n8265), .B2(
        n6336), .ZN(n6337) );
  INV_X1 U7499 ( .A(n6337), .ZN(n9985) );
  NAND2_X1 U7500 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  XNOR2_X1 U7501 ( .A(n6341), .B(n6340), .ZN(n6342) );
  AOI22_X1 U7502 ( .A1(n7972), .A2(\adder_stage1[5][8] ), .B1(n8078), .B2(
        n6342), .ZN(n6343) );
  INV_X1 U7503 ( .A(n6343), .ZN(n10078) );
  INV_X1 U7504 ( .A(n6344), .ZN(n7513) );
  OAI21_X1 U7505 ( .B1(n7513), .B2(n7509), .A(n7510), .ZN(n6349) );
  INV_X1 U7506 ( .A(n6345), .ZN(n6347) );
  NAND2_X1 U7507 ( .A1(n6347), .A2(n6346), .ZN(n6348) );
  XNOR2_X1 U7508 ( .A(n6349), .B(n6348), .ZN(n6350) );
  AOI22_X1 U7509 ( .A1(n7640), .A2(\adder_stage3[0][9] ), .B1(n8235), .B2(
        n6350), .ZN(n6351) );
  INV_X1 U7510 ( .A(n6351), .ZN(n9760) );
  BUF_X2 U7511 ( .A(n6352), .Z(n7570) );
  OR2_X1 U7512 ( .A1(\x_mult_f[8][0] ), .A2(\x_mult_f[9][0] ), .ZN(n6353) );
  AND2_X1 U7513 ( .A1(n6353), .A2(n7552), .ZN(n6354) );
  AOI22_X1 U7514 ( .A1(n7640), .A2(\adder_stage1[4][0] ), .B1(n7570), .B2(
        n6354), .ZN(n6355) );
  INV_X1 U7515 ( .A(n6355), .ZN(n10103) );
  INV_X1 U7516 ( .A(n6356), .ZN(n6358) );
  NAND2_X1 U7517 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  XOR2_X1 U7518 ( .A(n6360), .B(n6359), .Z(n6361) );
  AOI22_X1 U7519 ( .A1(n7622), .A2(\adder_stage1[4][6] ), .B1(n7570), .B2(
        n6361), .ZN(n6362) );
  INV_X1 U7520 ( .A(n6362), .ZN(n10097) );
  INV_X1 U7521 ( .A(n6363), .ZN(n6374) );
  INV_X1 U7522 ( .A(n6373), .ZN(n6364) );
  AOI21_X1 U7523 ( .B1(n6376), .B2(n6374), .A(n6364), .ZN(n6369) );
  INV_X1 U7524 ( .A(n6365), .ZN(n6367) );
  NAND2_X1 U7525 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  XOR2_X1 U7526 ( .A(n6369), .B(n6368), .Z(n6370) );
  AOI22_X1 U7527 ( .A1(n7622), .A2(\adder_stage1[4][5] ), .B1(n7570), .B2(
        n6370), .ZN(n6371) );
  INV_X1 U7528 ( .A(n6371), .ZN(n10098) );
  AOI22_X1 U7529 ( .A1(n7525), .A2(\x_mult_f[11][5] ), .B1(n7570), .B2(
        \x_mult_f_int[11][5] ), .ZN(n6372) );
  INV_X1 U7530 ( .A(n6372), .ZN(n9063) );
  NAND2_X1 U7531 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  XNOR2_X1 U7532 ( .A(n6376), .B(n6375), .ZN(n6377) );
  AOI22_X1 U7533 ( .A1(n7622), .A2(\adder_stage1[4][4] ), .B1(n7570), .B2(
        n6377), .ZN(n6378) );
  INV_X1 U7534 ( .A(n6378), .ZN(n10099) );
  INV_X1 U7535 ( .A(n6379), .ZN(n6852) );
  AOI21_X1 U7536 ( .B1(n6852), .B2(n6381), .A(n6380), .ZN(n6400) );
  INV_X1 U7537 ( .A(n6399), .ZN(n6382) );
  NAND2_X1 U7538 ( .A1(n6382), .A2(n6398), .ZN(n6383) );
  XOR2_X1 U7539 ( .A(n6400), .B(n6383), .Z(n6384) );
  AOI22_X1 U7540 ( .A1(n6854), .A2(\adder_stage1[5][6] ), .B1(n8078), .B2(
        n6384), .ZN(n6385) );
  INV_X1 U7541 ( .A(n6385), .ZN(n10080) );
  AOI22_X1 U7542 ( .A1(n7525), .A2(\x_mult_f[11][4] ), .B1(n8078), .B2(
        \x_mult_f_int[11][4] ), .ZN(n6386) );
  INV_X1 U7543 ( .A(n6386), .ZN(n9064) );
  INV_X1 U7544 ( .A(n6387), .ZN(n6850) );
  INV_X1 U7545 ( .A(n6849), .ZN(n6388) );
  AOI21_X1 U7546 ( .B1(n6852), .B2(n6850), .A(n6388), .ZN(n6393) );
  INV_X1 U7547 ( .A(n6389), .ZN(n6391) );
  NAND2_X1 U7548 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  XOR2_X1 U7549 ( .A(n6393), .B(n6392), .Z(n6394) );
  AOI22_X1 U7550 ( .A1(n6854), .A2(\adder_stage1[5][5] ), .B1(n8078), .B2(
        n6394), .ZN(n6395) );
  INV_X1 U7551 ( .A(n6395), .ZN(n10081) );
  AOI22_X1 U7552 ( .A1(n7525), .A2(\x_mult_f[11][1] ), .B1(n8078), .B2(
        \x_mult_f_int[11][1] ), .ZN(n6396) );
  INV_X1 U7553 ( .A(n6396), .ZN(n9348) );
  AOI22_X1 U7554 ( .A1(n7525), .A2(\x_mult_f[11][2] ), .B1(n8078), .B2(
        \x_mult_f_int[11][2] ), .ZN(n6397) );
  INV_X1 U7555 ( .A(n6397), .ZN(n9066) );
  OAI21_X1 U7556 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6405) );
  INV_X1 U7557 ( .A(n6401), .ZN(n6403) );
  NAND2_X1 U7558 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  XNOR2_X1 U7559 ( .A(n6405), .B(n6404), .ZN(n6406) );
  AOI22_X1 U7560 ( .A1(n6854), .A2(\adder_stage1[5][7] ), .B1(n8078), .B2(
        n6406), .ZN(n6407) );
  INV_X1 U7561 ( .A(n6407), .ZN(n10079) );
  AOI22_X1 U7562 ( .A1(n7525), .A2(\x_mult_f[11][3] ), .B1(n8078), .B2(
        \x_mult_f_int[11][3] ), .ZN(n6408) );
  INV_X1 U7563 ( .A(n6408), .ZN(n9065) );
  AOI22_X1 U7564 ( .A1(n7525), .A2(\x_mult_f[11][0] ), .B1(n8078), .B2(
        \x_mult_f_int[11][0] ), .ZN(n6409) );
  INV_X1 U7565 ( .A(n6409), .ZN(n9349) );
  AOI22_X1 U7566 ( .A1(n7556), .A2(\x_mult_f[10][0] ), .B1(n7570), .B2(
        \x_mult_f_int[10][0] ), .ZN(n6410) );
  INV_X1 U7567 ( .A(n6410), .ZN(n9347) );
  INV_X1 U7568 ( .A(n6411), .ZN(n6433) );
  OAI21_X1 U7569 ( .B1(n6433), .B2(n6429), .A(n6430), .ZN(n6416) );
  INV_X1 U7570 ( .A(n6412), .ZN(n6414) );
  NAND2_X1 U7571 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  XNOR2_X1 U7572 ( .A(n6416), .B(n6415), .ZN(n6417) );
  AOI22_X1 U7573 ( .A1(n8325), .A2(\adder_stage3[0][3] ), .B1(n8235), .B2(
        n6417), .ZN(n6418) );
  INV_X1 U7574 ( .A(n6418), .ZN(n9766) );
  INV_X1 U7575 ( .A(n6419), .ZN(n6421) );
  NAND2_X1 U7576 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  XOR2_X1 U7577 ( .A(n6422), .B(n6425), .Z(n6423) );
  AOI22_X1 U7578 ( .A1(n8330), .A2(\adder_stage3[0][1] ), .B1(n8235), .B2(
        n6423), .ZN(n6424) );
  INV_X1 U7579 ( .A(n6424), .ZN(n9768) );
  OR2_X1 U7580 ( .A1(\adder_stage2[0][0] ), .A2(\adder_stage2[1][0] ), .ZN(
        n6426) );
  AND2_X1 U7581 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  AOI22_X1 U7582 ( .A1(n8118), .A2(\adder_stage3[0][0] ), .B1(n8235), .B2(
        n6427), .ZN(n6428) );
  INV_X1 U7583 ( .A(n6428), .ZN(n9769) );
  INV_X1 U7584 ( .A(n6429), .ZN(n6431) );
  NAND2_X1 U7585 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  XOR2_X1 U7586 ( .A(n6433), .B(n6432), .Z(n6434) );
  AOI22_X1 U7587 ( .A1(n6854), .A2(\adder_stage3[0][2] ), .B1(n8235), .B2(
        n6434), .ZN(n6435) );
  INV_X1 U7588 ( .A(n6435), .ZN(n9767) );
  AOI22_X1 U7589 ( .A1(\x_mult_f_int[28][8] ), .A2(n8258), .B1(n8338), .B2(
        \x_mult_f[28][8] ), .ZN(n6437) );
  INV_X1 U7590 ( .A(n6437), .ZN(n9279) );
  AOI22_X1 U7591 ( .A1(\x_mult_f_int[28][6] ), .A2(n7927), .B1(n8409), .B2(
        \x_mult_f[28][6] ), .ZN(n6438) );
  INV_X1 U7592 ( .A(n6438), .ZN(n9281) );
  AOI22_X1 U7593 ( .A1(\x_mult_f_int[28][7] ), .A2(n7450), .B1(n8340), .B2(
        \x_mult_f[28][7] ), .ZN(n6439) );
  INV_X1 U7594 ( .A(n6439), .ZN(n9280) );
  OR2_X1 U7595 ( .A1(\adder_stage3[2][0] ), .A2(\adder_stage3[3][0] ), .ZN(
        n6440) );
  AND2_X1 U7596 ( .A1(n6440), .A2(n8278), .ZN(n6441) );
  AOI22_X1 U7597 ( .A1(n7972), .A2(\adder_stage4[1][0] ), .B1(n8078), .B2(
        n6441), .ZN(n6442) );
  INV_X1 U7598 ( .A(n6442), .ZN(n9666) );
  AOI22_X1 U7599 ( .A1(\x_mult_f_int[14][9] ), .A2(n8334), .B1(n8340), .B2(
        \x_mult_f[14][9] ), .ZN(n6443) );
  INV_X1 U7600 ( .A(n6443), .ZN(n9101) );
  BUF_X2 U7601 ( .A(n4645), .Z(n8167) );
  AOI22_X1 U7602 ( .A1(n7928), .A2(\x_mult_f[29][3] ), .B1(n8167), .B2(
        \x_mult_f_int[29][3] ), .ZN(n6444) );
  INV_X1 U7603 ( .A(n6444), .ZN(n9298) );
  AOI22_X1 U7604 ( .A1(\x_mult_f_int[1][6] ), .A2(n5175), .B1(n8401), .B2(
        \x_mult_f[1][6] ), .ZN(n6445) );
  INV_X1 U7605 ( .A(n6445), .ZN(n8936) );
  OR2_X1 U7606 ( .A1(\adder_stage3[2][17] ), .A2(\adder_stage3[3][17] ), .ZN(
        n8139) );
  AND2_X1 U7607 ( .A1(n8136), .A2(n8139), .ZN(n7708) );
  NAND2_X1 U7608 ( .A1(n8137), .A2(n7708), .ZN(n6448) );
  INV_X1 U7609 ( .A(n6446), .ZN(n8135) );
  NAND2_X1 U7610 ( .A1(\adder_stage3[2][17] ), .A2(\adder_stage3[3][17] ), 
        .ZN(n8138) );
  INV_X1 U7611 ( .A(n8138), .ZN(n6447) );
  AOI21_X1 U7612 ( .B1(n8135), .B2(n8139), .A(n6447), .ZN(n7713) );
  NAND2_X1 U7613 ( .A1(n6448), .A2(n7713), .ZN(n6450) );
  OR2_X1 U7614 ( .A1(\adder_stage3[2][18] ), .A2(\adder_stage3[3][18] ), .ZN(
        n7710) );
  NAND2_X1 U7615 ( .A1(\adder_stage3[2][18] ), .A2(\adder_stage3[3][18] ), 
        .ZN(n7711) );
  NAND2_X1 U7616 ( .A1(n7710), .A2(n7711), .ZN(n6449) );
  XNOR2_X1 U7617 ( .A(n6450), .B(n6449), .ZN(n6451) );
  AOI22_X1 U7618 ( .A1(n6451), .A2(n8175), .B1(n8401), .B2(
        \adder_stage4[1][18] ), .ZN(n6452) );
  INV_X1 U7619 ( .A(n6452), .ZN(n9648) );
  OAI21_X1 U7620 ( .B1(n3434), .B2(n6454), .A(n6453), .ZN(n8173) );
  OR2_X1 U7621 ( .A1(\x_mult_f[24][12] ), .A2(\x_mult_f[25][12] ), .ZN(n8171)
         );
  NAND2_X1 U7622 ( .A1(\x_mult_f[24][12] ), .A2(\x_mult_f[25][12] ), .ZN(n8170) );
  INV_X1 U7623 ( .A(n8170), .ZN(n6456) );
  AOI21_X1 U7624 ( .B1(n8173), .B2(n8171), .A(n6456), .ZN(n7594) );
  NOR2_X1 U7625 ( .A1(\x_mult_f[24][13] ), .A2(\x_mult_f[25][13] ), .ZN(n7590)
         );
  NAND2_X1 U7626 ( .A1(\x_mult_f[24][13] ), .A2(\x_mult_f[25][13] ), .ZN(n7591) );
  OAI21_X1 U7627 ( .B1(n7594), .B2(n7590), .A(n7591), .ZN(n8030) );
  AOI22_X1 U7628 ( .A1(n6457), .A2(n6279), .B1(n8409), .B2(
        \adder_stage1[12][14] ), .ZN(n6458) );
  INV_X1 U7629 ( .A(n6458), .ZN(n9955) );
  INV_X1 U7630 ( .A(n6459), .ZN(n6461) );
  NAND2_X1 U7631 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  XOR2_X1 U7632 ( .A(n6463), .B(n6462), .Z(n6464) );
  AOI22_X1 U7633 ( .A1(n8296), .A2(\adder_stage1[11][11] ), .B1(n8265), .B2(
        n6464), .ZN(n6465) );
  INV_X1 U7634 ( .A(n6465), .ZN(n9975) );
  NAND2_X1 U7635 ( .A1(n6487), .A2(n6466), .ZN(n6469) );
  INV_X1 U7636 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U7637 ( .A1(n6469), .A2(n6468), .ZN(n6473) );
  NAND2_X1 U7638 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  XNOR2_X1 U7639 ( .A(n6473), .B(n6472), .ZN(n6474) );
  AOI22_X1 U7640 ( .A1(n8097), .A2(\adder_stage3[3][13] ), .B1(n8265), .B2(
        n6474), .ZN(n6475) );
  INV_X1 U7641 ( .A(n6475), .ZN(n9695) );
  NOR2_X1 U7642 ( .A1(\adder_stage1[14][1] ), .A2(\adder_stage1[15][1] ), .ZN(
        n6502) );
  INV_X1 U7643 ( .A(n6502), .ZN(n6476) );
  NAND2_X1 U7644 ( .A1(\adder_stage1[14][1] ), .A2(\adder_stage1[15][1] ), 
        .ZN(n6501) );
  NAND2_X1 U7645 ( .A1(n6476), .A2(n6501), .ZN(n6477) );
  NAND2_X1 U7646 ( .A1(\adder_stage1[14][0] ), .A2(\adder_stage1[15][0] ), 
        .ZN(n7096) );
  XOR2_X1 U7647 ( .A(n6477), .B(n7096), .Z(n6478) );
  AOI22_X1 U7648 ( .A1(n8245), .A2(\adder_stage2[7][1] ), .B1(n8216), .B2(
        n6478), .ZN(n6479) );
  INV_X1 U7649 ( .A(n6479), .ZN(n9785) );
  INV_X1 U7650 ( .A(n6480), .ZN(n6482) );
  NAND2_X1 U7651 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  XOR2_X1 U7652 ( .A(n6484), .B(n6483), .Z(n6485) );
  AOI22_X1 U7653 ( .A1(n8168), .A2(\adder_stage3[3][15] ), .B1(n8265), .B2(
        n6485), .ZN(n6486) );
  INV_X1 U7654 ( .A(n6486), .ZN(n9693) );
  INV_X1 U7655 ( .A(n6487), .ZN(n8103) );
  INV_X1 U7656 ( .A(n6488), .ZN(n6491) );
  INV_X1 U7657 ( .A(n6489), .ZN(n6490) );
  OAI21_X1 U7658 ( .B1(n8103), .B2(n6491), .A(n6490), .ZN(n6924) );
  INV_X1 U7659 ( .A(n6492), .ZN(n6922) );
  INV_X1 U7660 ( .A(n6921), .ZN(n6493) );
  AOI21_X1 U7661 ( .B1(n6924), .B2(n6922), .A(n6493), .ZN(n6498) );
  INV_X1 U7662 ( .A(n6494), .ZN(n6496) );
  NAND2_X1 U7663 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  XOR2_X1 U7664 ( .A(n6498), .B(n6497), .Z(n6499) );
  AOI22_X1 U7665 ( .A1(n8273), .A2(\adder_stage3[3][11] ), .B1(n8265), .B2(
        n6499), .ZN(n6500) );
  INV_X1 U7666 ( .A(n6500), .ZN(n9697) );
  NOR2_X1 U7667 ( .A1(\adder_stage1[14][2] ), .A2(\adder_stage1[15][2] ), .ZN(
        n6613) );
  NOR2_X1 U7668 ( .A1(n6613), .A2(n6615), .ZN(n6504) );
  OAI21_X1 U7669 ( .B1(n6502), .B2(n7096), .A(n6501), .ZN(n6537) );
  NAND2_X1 U7670 ( .A1(\adder_stage1[14][2] ), .A2(\adder_stage1[15][2] ), 
        .ZN(n6612) );
  NAND2_X1 U7671 ( .A1(\adder_stage1[14][3] ), .A2(\adder_stage1[15][3] ), 
        .ZN(n6616) );
  OAI21_X1 U7672 ( .B1(n6615), .B2(n6612), .A(n6616), .ZN(n6503) );
  AOI21_X1 U7673 ( .B1(n6504), .B2(n6537), .A(n6503), .ZN(n6517) );
  NOR2_X1 U7674 ( .A1(\adder_stage1[14][4] ), .A2(\adder_stage1[15][4] ), .ZN(
        n6518) );
  NOR2_X1 U7675 ( .A1(\adder_stage1[14][5] ), .A2(\adder_stage1[15][5] ), .ZN(
        n6520) );
  NOR2_X1 U7676 ( .A1(n6518), .A2(n6520), .ZN(n6543) );
  NOR2_X1 U7677 ( .A1(\adder_stage1[14][6] ), .A2(\adder_stage1[15][6] ), .ZN(
        n6578) );
  NOR2_X1 U7678 ( .A1(\adder_stage1[14][7] ), .A2(\adder_stage1[15][7] ), .ZN(
        n6580) );
  NOR2_X1 U7679 ( .A1(n6578), .A2(n6580), .ZN(n6506) );
  NAND2_X1 U7680 ( .A1(n6543), .A2(n6506), .ZN(n6508) );
  NAND2_X1 U7681 ( .A1(\adder_stage1[14][4] ), .A2(\adder_stage1[15][4] ), 
        .ZN(n6571) );
  NAND2_X1 U7682 ( .A1(\adder_stage1[14][5] ), .A2(\adder_stage1[15][5] ), 
        .ZN(n6521) );
  OAI21_X1 U7683 ( .B1(n6520), .B2(n6571), .A(n6521), .ZN(n6542) );
  NAND2_X1 U7684 ( .A1(\adder_stage1[14][6] ), .A2(\adder_stage1[15][6] ), 
        .ZN(n6577) );
  NAND2_X1 U7685 ( .A1(\adder_stage1[14][7] ), .A2(\adder_stage1[15][7] ), 
        .ZN(n6581) );
  OAI21_X1 U7686 ( .B1(n6580), .B2(n6577), .A(n6581), .ZN(n6505) );
  AOI21_X1 U7687 ( .B1(n6506), .B2(n6542), .A(n6505), .ZN(n6507) );
  OAI21_X1 U7688 ( .B1(n3428), .B2(n6508), .A(n6507), .ZN(n6548) );
  NOR2_X1 U7689 ( .A1(\adder_stage1[14][8] ), .A2(\adder_stage1[15][8] ), .ZN(
        n6596) );
  INV_X1 U7690 ( .A(n6596), .ZN(n6567) );
  OR2_X1 U7691 ( .A1(\adder_stage1[14][9] ), .A2(\adder_stage1[15][9] ), .ZN(
        n6599) );
  NAND2_X1 U7692 ( .A1(n6567), .A2(n6599), .ZN(n6550) );
  NOR2_X1 U7693 ( .A1(\adder_stage1[14][10] ), .A2(\adder_stage1[15][10] ), 
        .ZN(n6551) );
  NOR2_X1 U7694 ( .A1(n6550), .A2(n6551), .ZN(n6512) );
  NAND2_X1 U7695 ( .A1(\adder_stage1[14][8] ), .A2(\adder_stage1[15][8] ), 
        .ZN(n6595) );
  INV_X1 U7696 ( .A(n6595), .ZN(n6510) );
  NAND2_X1 U7697 ( .A1(\adder_stage1[14][9] ), .A2(\adder_stage1[15][9] ), 
        .ZN(n6598) );
  INV_X1 U7698 ( .A(n6598), .ZN(n6509) );
  AOI21_X1 U7699 ( .B1(n6599), .B2(n6510), .A(n6509), .ZN(n6549) );
  NAND2_X1 U7700 ( .A1(\adder_stage1[14][10] ), .A2(\adder_stage1[15][10] ), 
        .ZN(n6552) );
  OAI21_X1 U7701 ( .B1(n6549), .B2(n6551), .A(n6552), .ZN(n6511) );
  AOI21_X1 U7702 ( .B1(n6548), .B2(n6512), .A(n6511), .ZN(n6589) );
  NOR2_X1 U7703 ( .A1(\adder_stage1[14][11] ), .A2(\adder_stage1[15][11] ), 
        .ZN(n6588) );
  INV_X1 U7704 ( .A(n6588), .ZN(n6513) );
  NAND2_X1 U7705 ( .A1(\adder_stage1[14][11] ), .A2(\adder_stage1[15][11] ), 
        .ZN(n6587) );
  NAND2_X1 U7706 ( .A1(n6513), .A2(n6587), .ZN(n6514) );
  XOR2_X1 U7707 ( .A(n3429), .B(n6514), .Z(n6515) );
  AOI22_X1 U7708 ( .A1(n7614), .A2(\adder_stage2[7][11] ), .B1(n6609), .B2(
        n6515), .ZN(n6516) );
  INV_X1 U7709 ( .A(n6516), .ZN(n9775) );
  INV_X1 U7710 ( .A(n6517), .ZN(n6574) );
  INV_X1 U7711 ( .A(n6518), .ZN(n6572) );
  INV_X1 U7712 ( .A(n6571), .ZN(n6519) );
  AOI21_X1 U7713 ( .B1(n6574), .B2(n6572), .A(n6519), .ZN(n6524) );
  INV_X1 U7714 ( .A(n6520), .ZN(n6522) );
  NAND2_X1 U7715 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  XOR2_X1 U7716 ( .A(n6524), .B(n6523), .Z(n6525) );
  AOI22_X1 U7717 ( .A1(n7972), .A2(\adder_stage2[7][5] ), .B1(n8216), .B2(
        n6525), .ZN(n6526) );
  INV_X1 U7718 ( .A(n6526), .ZN(n9781) );
  INV_X1 U7719 ( .A(n6527), .ZN(n8165) );
  INV_X1 U7720 ( .A(n6528), .ZN(n8163) );
  INV_X1 U7721 ( .A(n8162), .ZN(n6529) );
  AOI21_X1 U7722 ( .B1(n8165), .B2(n8163), .A(n6529), .ZN(n6534) );
  INV_X1 U7723 ( .A(n6530), .ZN(n6532) );
  NAND2_X1 U7724 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  XOR2_X1 U7725 ( .A(n6534), .B(n6533), .Z(n6535) );
  AOI22_X1 U7726 ( .A1(n8313), .A2(\adder_stage1[11][5] ), .B1(n8265), .B2(
        n6535), .ZN(n6536) );
  INV_X1 U7727 ( .A(n6536), .ZN(n9981) );
  INV_X1 U7728 ( .A(n6537), .ZN(n6614) );
  INV_X1 U7729 ( .A(n6613), .ZN(n6538) );
  NAND2_X1 U7730 ( .A1(n6538), .A2(n6612), .ZN(n6539) );
  XOR2_X1 U7731 ( .A(n6614), .B(n6539), .Z(n6540) );
  AOI22_X1 U7732 ( .A1(n8434), .A2(\adder_stage2[7][2] ), .B1(n8216), .B2(
        n6540), .ZN(n6541) );
  INV_X1 U7733 ( .A(n6541), .ZN(n9784) );
  AOI21_X1 U7734 ( .B1(n6574), .B2(n6543), .A(n6542), .ZN(n6579) );
  INV_X1 U7735 ( .A(n6578), .ZN(n6544) );
  NAND2_X1 U7736 ( .A1(n6544), .A2(n6577), .ZN(n6545) );
  XOR2_X1 U7737 ( .A(n6579), .B(n6545), .Z(n6546) );
  AOI22_X1 U7738 ( .A1(n8325), .A2(\adder_stage2[7][6] ), .B1(n8216), .B2(
        n6546), .ZN(n6547) );
  INV_X1 U7739 ( .A(n6547), .ZN(n9780) );
  INV_X1 U7740 ( .A(n6548), .ZN(n6597) );
  OAI21_X1 U7741 ( .B1(n6597), .B2(n6550), .A(n6549), .ZN(n6555) );
  INV_X1 U7742 ( .A(n6551), .ZN(n6553) );
  NAND2_X1 U7743 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  XNOR2_X1 U7744 ( .A(n6555), .B(n6554), .ZN(n6556) );
  AOI22_X1 U7745 ( .A1(n8398), .A2(\adder_stage2[7][10] ), .B1(n6609), .B2(
        n6556), .ZN(n6557) );
  INV_X1 U7746 ( .A(n6557), .ZN(n9776) );
  AOI21_X1 U7747 ( .B1(n8165), .B2(n6559), .A(n6558), .ZN(n6904) );
  OAI21_X1 U7748 ( .B1(n6904), .B2(n6900), .A(n6901), .ZN(n6564) );
  INV_X1 U7749 ( .A(n6560), .ZN(n6562) );
  NAND2_X1 U7750 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  XNOR2_X1 U7751 ( .A(n6564), .B(n6563), .ZN(n6565) );
  AOI22_X1 U7752 ( .A1(n8296), .A2(\adder_stage1[11][7] ), .B1(n8265), .B2(
        n6565), .ZN(n6566) );
  INV_X1 U7753 ( .A(n6566), .ZN(n9979) );
  NAND2_X1 U7754 ( .A1(n6567), .A2(n6595), .ZN(n6568) );
  XOR2_X1 U7755 ( .A(n6597), .B(n6568), .Z(n6569) );
  AOI22_X1 U7756 ( .A1(n7640), .A2(\adder_stage2[7][8] ), .B1(n8216), .B2(
        n6569), .ZN(n6570) );
  INV_X1 U7757 ( .A(n6570), .ZN(n9778) );
  NAND2_X1 U7758 ( .A1(n6572), .A2(n6571), .ZN(n6573) );
  XNOR2_X1 U7759 ( .A(n6574), .B(n6573), .ZN(n6575) );
  AOI22_X1 U7760 ( .A1(n8176), .A2(\adder_stage2[7][4] ), .B1(n8216), .B2(
        n6575), .ZN(n6576) );
  INV_X1 U7761 ( .A(n6576), .ZN(n9782) );
  OAI21_X1 U7762 ( .B1(n6579), .B2(n6578), .A(n6577), .ZN(n6584) );
  INV_X1 U7763 ( .A(n6580), .ZN(n6582) );
  NAND2_X1 U7764 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  XNOR2_X1 U7765 ( .A(n6584), .B(n6583), .ZN(n6585) );
  AOI22_X1 U7766 ( .A1(n8296), .A2(\adder_stage2[7][7] ), .B1(n8216), .B2(
        n6585), .ZN(n6586) );
  INV_X1 U7767 ( .A(n6586), .ZN(n9779) );
  OAI21_X1 U7768 ( .B1(n6589), .B2(n6588), .A(n6587), .ZN(n6607) );
  OR2_X1 U7769 ( .A1(\adder_stage1[14][12] ), .A2(\adder_stage1[15][12] ), 
        .ZN(n6605) );
  NAND2_X1 U7770 ( .A1(\adder_stage1[14][12] ), .A2(\adder_stage1[15][12] ), 
        .ZN(n6604) );
  INV_X1 U7771 ( .A(n6604), .ZN(n6590) );
  AOI21_X1 U7772 ( .B1(n6607), .B2(n6605), .A(n6590), .ZN(n7565) );
  NOR2_X1 U7773 ( .A1(\adder_stage1[14][13] ), .A2(\adder_stage1[15][13] ), 
        .ZN(n7564) );
  INV_X1 U7774 ( .A(n7564), .ZN(n6591) );
  NAND2_X1 U7775 ( .A1(\adder_stage1[14][13] ), .A2(\adder_stage1[15][13] ), 
        .ZN(n7563) );
  NAND2_X1 U7776 ( .A1(n6591), .A2(n7563), .ZN(n6592) );
  XOR2_X1 U7777 ( .A(n7565), .B(n6592), .Z(n6593) );
  AOI22_X1 U7778 ( .A1(n8330), .A2(\adder_stage2[7][13] ), .B1(n6609), .B2(
        n6593), .ZN(n6594) );
  INV_X1 U7779 ( .A(n6594), .ZN(n9773) );
  OAI21_X1 U7780 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6601) );
  NAND2_X1 U7781 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  XNOR2_X1 U7782 ( .A(n6601), .B(n6600), .ZN(n6602) );
  AOI22_X1 U7783 ( .A1(n8313), .A2(\adder_stage2[7][9] ), .B1(n6609), .B2(
        n6602), .ZN(n6603) );
  INV_X1 U7784 ( .A(n6603), .ZN(n9777) );
  NAND2_X1 U7785 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  XNOR2_X1 U7786 ( .A(n6607), .B(n6606), .ZN(n6608) );
  AOI22_X1 U7787 ( .A1(n7177), .A2(\adder_stage2[7][12] ), .B1(n6609), .B2(
        n6608), .ZN(n6610) );
  INV_X1 U7788 ( .A(n6610), .ZN(n9774) );
  AOI22_X1 U7789 ( .A1(n8434), .A2(\x_mult_f[22][4] ), .B1(n6626), .B2(
        \x_mult_f_int[22][4] ), .ZN(n6611) );
  INV_X1 U7790 ( .A(n6611), .ZN(n9207) );
  OAI21_X1 U7791 ( .B1(n6614), .B2(n6613), .A(n6612), .ZN(n6619) );
  INV_X1 U7792 ( .A(n6615), .ZN(n6617) );
  NAND2_X1 U7793 ( .A1(n6617), .A2(n6616), .ZN(n6618) );
  XNOR2_X1 U7794 ( .A(n6619), .B(n6618), .ZN(n6620) );
  AOI22_X1 U7795 ( .A1(n8328), .A2(\adder_stage2[7][3] ), .B1(n8216), .B2(
        n6620), .ZN(n6621) );
  INV_X1 U7796 ( .A(n6621), .ZN(n9783) );
  AOI22_X1 U7797 ( .A1(n7074), .A2(\x_mult_f[22][2] ), .B1(n6626), .B2(
        \x_mult_f_int[22][2] ), .ZN(n6622) );
  INV_X1 U7798 ( .A(n6622), .ZN(n9209) );
  AOI22_X1 U7799 ( .A1(n8328), .A2(\x_mult_f[22][1] ), .B1(n6626), .B2(
        \x_mult_f_int[22][1] ), .ZN(n6623) );
  INV_X1 U7800 ( .A(n6623), .ZN(n9370) );
  AOI22_X1 U7801 ( .A1(n8296), .A2(\x_mult_f[22][0] ), .B1(n6626), .B2(
        \x_mult_f_int[22][0] ), .ZN(n6624) );
  INV_X1 U7802 ( .A(n6624), .ZN(n9371) );
  AOI22_X1 U7803 ( .A1(n8273), .A2(\x_mult_f[22][5] ), .B1(n6626), .B2(
        \x_mult_f_int[22][5] ), .ZN(n6625) );
  INV_X1 U7804 ( .A(n6625), .ZN(n9206) );
  AOI22_X1 U7805 ( .A1(n8273), .A2(\x_mult_f[22][3] ), .B1(n6626), .B2(
        \x_mult_f_int[22][3] ), .ZN(n6627) );
  INV_X1 U7806 ( .A(n6627), .ZN(n9208) );
  AOI22_X1 U7807 ( .A1(n8401), .A2(\x_mult_f[10][4] ), .B1(n7570), .B2(
        \x_mult_f_int[10][4] ), .ZN(n6628) );
  INV_X1 U7808 ( .A(n6628), .ZN(n9051) );
  AOI21_X1 U7809 ( .B1(n3410), .B2(n6630), .A(n6629), .ZN(n6635) );
  NAND2_X1 U7810 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  XOR2_X1 U7811 ( .A(n6635), .B(n6634), .Z(n6637) );
  AOI22_X1 U7812 ( .A1(n6637), .A2(n6636), .B1(n8328), .B2(
        \adder_stage1[10][13] ), .ZN(n6638) );
  INV_X1 U7813 ( .A(n6638), .ZN(n9990) );
  INV_X1 U7814 ( .A(n6639), .ZN(n6641) );
  NAND2_X1 U7815 ( .A1(n6641), .A2(n6640), .ZN(n6642) );
  XOR2_X1 U7816 ( .A(n6643), .B(n6642), .Z(n6644) );
  AOI22_X1 U7817 ( .A1(n7074), .A2(\adder_stage1[11][2] ), .B1(n8167), .B2(
        n6644), .ZN(n6645) );
  INV_X1 U7818 ( .A(n6645), .ZN(n9984) );
  AOI22_X1 U7819 ( .A1(\x_mult_f_int[30][7] ), .A2(n7507), .B1(n8428), .B2(
        \x_mult_f[30][7] ), .ZN(n6646) );
  INV_X1 U7820 ( .A(n6646), .ZN(n9308) );
  AOI22_X1 U7821 ( .A1(\x_mult_f_int[20][7] ), .A2(n6636), .B1(n8325), .B2(
        \x_mult_f[20][7] ), .ZN(n6647) );
  INV_X1 U7822 ( .A(n6647), .ZN(n9176) );
  AOI22_X1 U7823 ( .A1(\x_mult_f_int[20][6] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[20][6] ), .ZN(n6648) );
  INV_X1 U7824 ( .A(n6648), .ZN(n9177) );
  AOI22_X1 U7825 ( .A1(\x_mult_f_int[25][6] ), .A2(n8294), .B1(n8336), .B2(
        \x_mult_f[25][6] ), .ZN(n6649) );
  INV_X1 U7826 ( .A(n6649), .ZN(n9239) );
  BUF_X2 U7827 ( .A(n6238), .Z(n8292) );
  INV_X1 U7828 ( .A(n6650), .ZN(n6692) );
  OAI21_X1 U7829 ( .B1(n6692), .B2(n6677), .A(n6678), .ZN(n6655) );
  INV_X1 U7830 ( .A(n6651), .ZN(n6653) );
  NAND2_X1 U7831 ( .A1(n6653), .A2(n6652), .ZN(n6654) );
  XNOR2_X1 U7832 ( .A(n6655), .B(n6654), .ZN(n6656) );
  AOI22_X1 U7833 ( .A1(n8057), .A2(\adder_stage4[1][9] ), .B1(n8292), .B2(
        n6656), .ZN(n6657) );
  INV_X1 U7834 ( .A(n6657), .ZN(n9657) );
  INV_X1 U7835 ( .A(n6658), .ZN(n6661) );
  INV_X1 U7836 ( .A(n6659), .ZN(n6660) );
  OAI21_X1 U7837 ( .B1(n6692), .B2(n6661), .A(n6660), .ZN(n6674) );
  INV_X1 U7838 ( .A(n6662), .ZN(n6672) );
  INV_X1 U7839 ( .A(n6671), .ZN(n6663) );
  AOI21_X1 U7840 ( .B1(n6674), .B2(n6672), .A(n6663), .ZN(n6668) );
  INV_X1 U7841 ( .A(n6664), .ZN(n6666) );
  NAND2_X1 U7842 ( .A1(n6666), .A2(n6665), .ZN(n6667) );
  XOR2_X1 U7843 ( .A(n6668), .B(n6667), .Z(n6669) );
  AOI22_X1 U7844 ( .A1(n8057), .A2(\adder_stage4[1][11] ), .B1(n8292), .B2(
        n6669), .ZN(n6670) );
  INV_X1 U7845 ( .A(n6670), .ZN(n9655) );
  NAND2_X1 U7846 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  XNOR2_X1 U7847 ( .A(n6674), .B(n6673), .ZN(n6675) );
  AOI22_X1 U7848 ( .A1(n8336), .A2(\adder_stage4[1][10] ), .B1(n8292), .B2(
        n6675), .ZN(n6676) );
  INV_X1 U7849 ( .A(n6676), .ZN(n9656) );
  INV_X1 U7850 ( .A(n6677), .ZN(n6679) );
  NAND2_X1 U7851 ( .A1(n6679), .A2(n6678), .ZN(n6680) );
  XOR2_X1 U7852 ( .A(n6692), .B(n6680), .Z(n6681) );
  AOI22_X1 U7853 ( .A1(n8313), .A2(\adder_stage4[1][8] ), .B1(n8292), .B2(
        n6681), .ZN(n6682) );
  INV_X1 U7854 ( .A(n6682), .ZN(n9658) );
  AOI21_X1 U7855 ( .B1(n6685), .B2(n6684), .A(n6683), .ZN(n8285) );
  INV_X1 U7856 ( .A(n8284), .ZN(n6686) );
  NAND2_X1 U7857 ( .A1(n6686), .A2(n8283), .ZN(n6687) );
  XOR2_X1 U7858 ( .A(n8285), .B(n6687), .Z(n6688) );
  AOI22_X1 U7859 ( .A1(n8338), .A2(\adder_stage4[1][6] ), .B1(n8292), .B2(
        n6688), .ZN(n6689) );
  INV_X1 U7860 ( .A(n6689), .ZN(n9660) );
  OAI21_X1 U7861 ( .B1(n6692), .B2(n6691), .A(n6690), .ZN(n6697) );
  INV_X1 U7862 ( .A(n6693), .ZN(n6695) );
  NAND2_X1 U7863 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  XNOR2_X1 U7864 ( .A(n6697), .B(n6696), .ZN(n6698) );
  AOI22_X1 U7865 ( .A1(n8088), .A2(\adder_stage4[1][12] ), .B1(n8292), .B2(
        n6698), .ZN(n6699) );
  INV_X1 U7866 ( .A(n6699), .ZN(n9654) );
  AOI22_X1 U7867 ( .A1(\x_mult_f_int[15][12] ), .A2(n7862), .B1(n8296), .B2(
        \x_mult_f[15][12] ), .ZN(n6700) );
  INV_X1 U7868 ( .A(n6700), .ZN(n9112) );
  AOI22_X1 U7869 ( .A1(\x_mult_f_int[15][11] ), .A2(n6279), .B1(n8340), .B2(
        \x_mult_f[15][11] ), .ZN(n6701) );
  INV_X1 U7870 ( .A(n6701), .ZN(n9113) );
  AOI22_X1 U7871 ( .A1(n6877), .A2(\x_mult_f[7][4] ), .B1(n8189), .B2(
        \x_mult_f_int[7][4] ), .ZN(n6702) );
  INV_X1 U7872 ( .A(n6702), .ZN(n9009) );
  BUF_X2 U7873 ( .A(n6352), .Z(n7971) );
  NOR2_X1 U7874 ( .A1(\x_mult_f[4][2] ), .A2(\x_mult_f[5][2] ), .ZN(n6867) );
  NOR2_X1 U7875 ( .A1(n6867), .A2(n6869), .ZN(n6704) );
  NOR2_X1 U7876 ( .A1(\x_mult_f[4][1] ), .A2(\x_mult_f[5][1] ), .ZN(n6856) );
  NAND2_X1 U7877 ( .A1(\x_mult_f[4][0] ), .A2(\x_mult_f[5][0] ), .ZN(n6862) );
  NAND2_X1 U7878 ( .A1(\x_mult_f[4][1] ), .A2(\x_mult_f[5][1] ), .ZN(n6857) );
  OAI21_X1 U7879 ( .B1(n6856), .B2(n6862), .A(n6857), .ZN(n6844) );
  NAND2_X1 U7880 ( .A1(\x_mult_f[4][3] ), .A2(\x_mult_f[5][3] ), .ZN(n6870) );
  OAI21_X1 U7881 ( .B1(n6869), .B2(n6866), .A(n6870), .ZN(n6703) );
  NOR2_X1 U7882 ( .A1(\x_mult_f[4][4] ), .A2(\x_mult_f[5][4] ), .ZN(n6801) );
  NOR2_X1 U7883 ( .A1(\x_mult_f[4][5] ), .A2(\x_mult_f[5][5] ), .ZN(n6803) );
  NOR2_X1 U7884 ( .A1(n6801), .A2(n6803), .ZN(n6785) );
  NOR2_X1 U7885 ( .A1(\x_mult_f[4][6] ), .A2(\x_mult_f[5][6] ), .ZN(n6794) );
  NOR2_X1 U7886 ( .A1(\x_mult_f[4][7] ), .A2(\x_mult_f[5][7] ), .ZN(n6786) );
  NOR2_X1 U7887 ( .A1(n6794), .A2(n6786), .ZN(n6706) );
  NAND2_X1 U7888 ( .A1(n6785), .A2(n6706), .ZN(n6708) );
  NAND2_X1 U7889 ( .A1(\x_mult_f[4][4] ), .A2(\x_mult_f[5][4] ), .ZN(n6837) );
  NAND2_X1 U7890 ( .A1(\x_mult_f[4][5] ), .A2(\x_mult_f[5][5] ), .ZN(n6804) );
  OAI21_X1 U7891 ( .B1(n6803), .B2(n6837), .A(n6804), .ZN(n6784) );
  NAND2_X1 U7892 ( .A1(\x_mult_f[4][6] ), .A2(\x_mult_f[5][6] ), .ZN(n6795) );
  NAND2_X1 U7893 ( .A1(\x_mult_f[4][7] ), .A2(\x_mult_f[5][7] ), .ZN(n6787) );
  OAI21_X1 U7894 ( .B1(n6786), .B2(n6795), .A(n6787), .ZN(n6705) );
  AOI21_X1 U7895 ( .B1(n6706), .B2(n6784), .A(n6705), .ZN(n6707) );
  OAI21_X1 U7896 ( .B1(n6783), .B2(n6708), .A(n6707), .ZN(n6778) );
  OR2_X1 U7897 ( .A1(\x_mult_f[4][8] ), .A2(\x_mult_f[5][8] ), .ZN(n6776) );
  NAND2_X1 U7898 ( .A1(\x_mult_f[4][8] ), .A2(\x_mult_f[5][8] ), .ZN(n6775) );
  INV_X1 U7899 ( .A(n6775), .ZN(n6725) );
  AOI21_X1 U7900 ( .B1(n6721), .B2(n6776), .A(n6725), .ZN(n6710) );
  OR2_X1 U7901 ( .A1(\x_mult_f[4][9] ), .A2(\x_mult_f[5][9] ), .ZN(n6724) );
  NAND2_X1 U7902 ( .A1(\x_mult_f[4][9] ), .A2(\x_mult_f[5][9] ), .ZN(n6722) );
  NAND2_X1 U7903 ( .A1(n6724), .A2(n6722), .ZN(n6709) );
  XOR2_X1 U7904 ( .A(n6710), .B(n6709), .Z(n6711) );
  AOI22_X1 U7905 ( .A1(n7177), .A2(\adder_stage1[2][9] ), .B1(n7971), .B2(
        n6711), .ZN(n6712) );
  INV_X1 U7906 ( .A(n6712), .ZN(n10126) );
  NAND2_X1 U7907 ( .A1(n6714), .A2(n6713), .ZN(n6715) );
  XNOR2_X1 U7908 ( .A(n6716), .B(n6715), .ZN(n6717) );
  AOI22_X1 U7909 ( .A1(n6877), .A2(\adder_stage1[3][12] ), .B1(n7163), .B2(
        n6717), .ZN(n6718) );
  INV_X1 U7910 ( .A(n6718), .ZN(n10108) );
  AOI22_X1 U7911 ( .A1(n6877), .A2(\x_mult_f[7][5] ), .B1(n6036), .B2(
        \x_mult_f_int[7][5] ), .ZN(n6719) );
  INV_X1 U7912 ( .A(n6719), .ZN(n9008) );
  INV_X2 U7913 ( .A(n6720), .ZN(n7972) );
  AND2_X1 U7914 ( .A1(n6776), .A2(n6724), .ZN(n6764) );
  NAND2_X1 U7915 ( .A1(n6721), .A2(n6764), .ZN(n6726) );
  INV_X1 U7916 ( .A(n6722), .ZN(n6723) );
  AOI21_X1 U7917 ( .B1(n6725), .B2(n6724), .A(n6723), .ZN(n6768) );
  NAND2_X1 U7918 ( .A1(n6726), .A2(n6768), .ZN(n6728) );
  OR2_X1 U7919 ( .A1(\x_mult_f[4][10] ), .A2(\x_mult_f[5][10] ), .ZN(n6765) );
  NAND2_X1 U7920 ( .A1(\x_mult_f[4][10] ), .A2(\x_mult_f[5][10] ), .ZN(n6766)
         );
  NAND2_X1 U7921 ( .A1(n6765), .A2(n6766), .ZN(n6727) );
  XNOR2_X1 U7922 ( .A(n6728), .B(n6727), .ZN(n6729) );
  AOI22_X1 U7923 ( .A1(n7972), .A2(\adder_stage1[2][10] ), .B1(n7971), .B2(
        n6729), .ZN(n6730) );
  INV_X1 U7924 ( .A(n6730), .ZN(n10125) );
  AOI21_X1 U7925 ( .B1(n3441), .B2(n6742), .A(n6731), .ZN(n6735) );
  NAND2_X1 U7926 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  XOR2_X1 U7927 ( .A(n6735), .B(n6734), .Z(n6736) );
  AOI22_X1 U7928 ( .A1(n7041), .A2(\adder_stage1[3][9] ), .B1(n7507), .B2(
        n6736), .ZN(n6737) );
  INV_X1 U7929 ( .A(n6737), .ZN(n10111) );
  BUF_X2 U7930 ( .A(n5449), .Z(n6875) );
  AOI22_X1 U7931 ( .A1(n7972), .A2(\x_mult_f[6][5] ), .B1(n6875), .B2(
        \x_mult_f_int[6][5] ), .ZN(n6738) );
  INV_X1 U7932 ( .A(n6738), .ZN(n8994) );
  AOI22_X1 U7933 ( .A1(n7972), .A2(\x_mult_f[6][4] ), .B1(n6875), .B2(
        \x_mult_f_int[6][4] ), .ZN(n6739) );
  INV_X1 U7934 ( .A(n6739), .ZN(n8995) );
  AOI22_X1 U7935 ( .A1(n7972), .A2(\x_mult_f[6][3] ), .B1(n6875), .B2(
        \x_mult_f_int[6][3] ), .ZN(n6740) );
  INV_X1 U7936 ( .A(n6740), .ZN(n8996) );
  NAND2_X1 U7937 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  XNOR2_X1 U7938 ( .A(n3441), .B(n6743), .ZN(n6745) );
  AOI22_X1 U7939 ( .A1(n7041), .A2(\adder_stage1[3][8] ), .B1(n8024), .B2(
        n6745), .ZN(n6746) );
  INV_X1 U7940 ( .A(n6746), .ZN(n10112) );
  AOI21_X1 U7941 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n6814) );
  OAI21_X1 U7942 ( .B1(n6814), .B2(n6810), .A(n6811), .ZN(n6754) );
  INV_X1 U7943 ( .A(n6750), .ZN(n6752) );
  NAND2_X1 U7944 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  XNOR2_X1 U7945 ( .A(n6754), .B(n6753), .ZN(n6755) );
  AOI22_X1 U7946 ( .A1(n7041), .A2(\adder_stage1[3][7] ), .B1(n7163), .B2(
        n6755), .ZN(n6756) );
  INV_X1 U7947 ( .A(n6756), .ZN(n10113) );
  INV_X1 U7948 ( .A(n6757), .ZN(n6759) );
  NAND2_X1 U7949 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  XOR2_X1 U7950 ( .A(n6761), .B(n6760), .Z(n6762) );
  AOI22_X1 U7951 ( .A1(n6877), .A2(\adder_stage1[3][11] ), .B1(n7570), .B2(
        n6762), .ZN(n6763) );
  INV_X1 U7952 ( .A(n6763), .ZN(n10109) );
  AND2_X1 U7953 ( .A1(n6764), .A2(n6765), .ZN(n6770) );
  INV_X1 U7954 ( .A(n6765), .ZN(n6767) );
  OAI21_X1 U7955 ( .B1(n6768), .B2(n6767), .A(n6766), .ZN(n6769) );
  AOI21_X1 U7956 ( .B1(n6778), .B2(n6770), .A(n6769), .ZN(n7320) );
  NOR2_X1 U7957 ( .A1(\x_mult_f[4][11] ), .A2(\x_mult_f[5][11] ), .ZN(n7319)
         );
  INV_X1 U7958 ( .A(n7319), .ZN(n6771) );
  NAND2_X1 U7959 ( .A1(\x_mult_f[4][11] ), .A2(\x_mult_f[5][11] ), .ZN(n7318)
         );
  NAND2_X1 U7960 ( .A1(n6771), .A2(n7318), .ZN(n6772) );
  XOR2_X1 U7961 ( .A(n3412), .B(n6772), .Z(n6773) );
  AOI22_X1 U7962 ( .A1(n7972), .A2(\adder_stage1[2][11] ), .B1(n7971), .B2(
        n6773), .ZN(n6774) );
  INV_X1 U7963 ( .A(n6774), .ZN(n10124) );
  NAND2_X1 U7964 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  XNOR2_X1 U7965 ( .A(n6778), .B(n6777), .ZN(n6779) );
  AOI22_X1 U7966 ( .A1(n7177), .A2(\adder_stage1[2][8] ), .B1(n7971), .B2(
        n6779), .ZN(n6780) );
  INV_X1 U7967 ( .A(n6780), .ZN(n10127) );
  AOI22_X1 U7968 ( .A1(n7972), .A2(\x_mult_f[6][1] ), .B1(n6875), .B2(
        \x_mult_f_int[6][1] ), .ZN(n6781) );
  INV_X1 U7969 ( .A(n6781), .ZN(n9338) );
  AOI22_X1 U7970 ( .A1(n7972), .A2(\x_mult_f[6][2] ), .B1(n6875), .B2(
        \x_mult_f_int[6][2] ), .ZN(n6782) );
  INV_X1 U7971 ( .A(n6782), .ZN(n8997) );
  INV_X1 U7972 ( .A(n6783), .ZN(n6840) );
  AOI21_X1 U7973 ( .B1(n6840), .B2(n6785), .A(n6784), .ZN(n6798) );
  OAI21_X1 U7974 ( .B1(n6798), .B2(n6794), .A(n6795), .ZN(n6790) );
  INV_X1 U7975 ( .A(n6786), .ZN(n6788) );
  NAND2_X1 U7976 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  XNOR2_X1 U7977 ( .A(n6790), .B(n6789), .ZN(n6791) );
  AOI22_X1 U7978 ( .A1(n7177), .A2(\adder_stage1[2][7] ), .B1(n6875), .B2(
        n6791), .ZN(n6792) );
  INV_X1 U7979 ( .A(n6792), .ZN(n10128) );
  AOI22_X1 U7980 ( .A1(n7972), .A2(\x_mult_f[6][0] ), .B1(n6875), .B2(
        \x_mult_f_int[6][0] ), .ZN(n6793) );
  INV_X1 U7981 ( .A(n6793), .ZN(n9339) );
  INV_X1 U7982 ( .A(n6794), .ZN(n6796) );
  NAND2_X1 U7983 ( .A1(n6796), .A2(n6795), .ZN(n6797) );
  XOR2_X1 U7984 ( .A(n6798), .B(n6797), .Z(n6799) );
  AOI22_X1 U7985 ( .A1(n7177), .A2(\adder_stage1[2][6] ), .B1(n6875), .B2(
        n6799), .ZN(n6800) );
  INV_X1 U7986 ( .A(n6800), .ZN(n10129) );
  INV_X1 U7987 ( .A(n6801), .ZN(n6838) );
  INV_X1 U7988 ( .A(n6837), .ZN(n6802) );
  AOI21_X1 U7989 ( .B1(n6840), .B2(n6838), .A(n6802), .ZN(n6807) );
  INV_X1 U7990 ( .A(n6803), .ZN(n6805) );
  NAND2_X1 U7991 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  XOR2_X1 U7992 ( .A(n6807), .B(n6806), .Z(n6808) );
  AOI22_X1 U7993 ( .A1(n7177), .A2(\adder_stage1[2][5] ), .B1(n6875), .B2(
        n6808), .ZN(n6809) );
  INV_X1 U7994 ( .A(n6809), .ZN(n10130) );
  INV_X1 U7995 ( .A(n6810), .ZN(n6812) );
  NAND2_X1 U7996 ( .A1(n6812), .A2(n6811), .ZN(n6813) );
  XOR2_X1 U7997 ( .A(n6814), .B(n6813), .Z(n6815) );
  AOI22_X1 U7998 ( .A1(n7041), .A2(\adder_stage1[3][6] ), .B1(n7155), .B2(
        n6815), .ZN(n6816) );
  INV_X1 U7999 ( .A(n6816), .ZN(n10114) );
  NAND2_X1 U8000 ( .A1(n3441), .A2(n6817), .ZN(n6819) );
  NAND2_X1 U8001 ( .A1(n6819), .A2(n6818), .ZN(n6823) );
  NAND2_X1 U8002 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  XNOR2_X1 U8003 ( .A(n6823), .B(n6822), .ZN(n6824) );
  AOI22_X1 U8004 ( .A1(n6877), .A2(\adder_stage1[3][10] ), .B1(n8272), .B2(
        n6824), .ZN(n6825) );
  INV_X1 U8005 ( .A(n6825), .ZN(n10110) );
  AOI22_X1 U8006 ( .A1(n6877), .A2(\x_mult_f[5][4] ), .B1(n7971), .B2(
        \x_mult_f_int[5][4] ), .ZN(n6826) );
  INV_X1 U8007 ( .A(n6826), .ZN(n8981) );
  AOI22_X1 U8008 ( .A1(n6877), .A2(\x_mult_f[7][3] ), .B1(n6272), .B2(
        \x_mult_f_int[7][3] ), .ZN(n6827) );
  INV_X1 U8009 ( .A(n6827), .ZN(n9010) );
  AOI22_X1 U8010 ( .A1(n6877), .A2(\x_mult_f[7][2] ), .B1(n8209), .B2(
        \x_mult_f_int[7][2] ), .ZN(n6828) );
  INV_X1 U8011 ( .A(n6828), .ZN(n9011) );
  AOI22_X1 U8012 ( .A1(n6877), .A2(\x_mult_f[7][1] ), .B1(n8087), .B2(
        \x_mult_f_int[7][1] ), .ZN(n6829) );
  INV_X1 U8013 ( .A(n6829), .ZN(n9340) );
  AOI22_X1 U8014 ( .A1(n6877), .A2(\x_mult_f[7][0] ), .B1(n7919), .B2(
        \x_mult_f_int[7][0] ), .ZN(n6830) );
  INV_X1 U8015 ( .A(n6830), .ZN(n9341) );
  AOI22_X1 U8016 ( .A1(n6877), .A2(\x_mult_f[5][3] ), .B1(n7971), .B2(
        \x_mult_f_int[5][3] ), .ZN(n6831) );
  INV_X1 U8017 ( .A(n6831), .ZN(n8982) );
  AOI22_X1 U8018 ( .A1(n6877), .A2(\x_mult_f[5][5] ), .B1(n7971), .B2(
        \x_mult_f_int[5][5] ), .ZN(n6832) );
  INV_X1 U8019 ( .A(n6832), .ZN(n8980) );
  AOI22_X1 U8020 ( .A1(n8245), .A2(\x_mult_f[4][1] ), .B1(n7971), .B2(
        \x_mult_f_int[4][1] ), .ZN(n6833) );
  INV_X1 U8021 ( .A(n6833), .ZN(n9334) );
  AOI22_X1 U8022 ( .A1(n7972), .A2(\x_mult_f[5][2] ), .B1(n7971), .B2(
        \x_mult_f_int[5][2] ), .ZN(n6834) );
  INV_X1 U8023 ( .A(n6834), .ZN(n8983) );
  AOI22_X1 U8024 ( .A1(n7972), .A2(\x_mult_f[5][1] ), .B1(n7971), .B2(
        \x_mult_f_int[5][1] ), .ZN(n6835) );
  INV_X1 U8025 ( .A(n6835), .ZN(n9336) );
  AOI22_X1 U8026 ( .A1(n7972), .A2(\x_mult_f[5][0] ), .B1(n7971), .B2(
        \x_mult_f_int[5][0] ), .ZN(n6836) );
  INV_X1 U8027 ( .A(n6836), .ZN(n9337) );
  NAND2_X1 U8028 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  XNOR2_X1 U8029 ( .A(n6840), .B(n6839), .ZN(n6841) );
  AOI22_X1 U8030 ( .A1(n7177), .A2(\adder_stage1[2][4] ), .B1(n6875), .B2(
        n6841), .ZN(n6842) );
  INV_X1 U8031 ( .A(n6842), .ZN(n10131) );
  AOI22_X1 U8032 ( .A1(n7177), .A2(\x_mult_f[4][2] ), .B1(n7971), .B2(
        \x_mult_f_int[4][2] ), .ZN(n6843) );
  INV_X1 U8033 ( .A(n6843), .ZN(n8978) );
  INV_X1 U8034 ( .A(n6844), .ZN(n6868) );
  INV_X1 U8035 ( .A(n6867), .ZN(n6845) );
  NAND2_X1 U8036 ( .A1(n6845), .A2(n6866), .ZN(n6846) );
  XOR2_X1 U8037 ( .A(n6868), .B(n6846), .Z(n6847) );
  AOI22_X1 U8038 ( .A1(n7177), .A2(\adder_stage1[2][2] ), .B1(n6875), .B2(
        n6847), .ZN(n6848) );
  INV_X1 U8039 ( .A(n6848), .ZN(n10133) );
  NAND2_X1 U8040 ( .A1(n6850), .A2(n6849), .ZN(n6851) );
  XNOR2_X1 U8041 ( .A(n6852), .B(n6851), .ZN(n6853) );
  AOI22_X1 U8042 ( .A1(n6854), .A2(\adder_stage1[5][4] ), .B1(n7962), .B2(
        n6853), .ZN(n6855) );
  INV_X1 U8043 ( .A(n6855), .ZN(n10082) );
  INV_X1 U8044 ( .A(n6856), .ZN(n6858) );
  NAND2_X1 U8045 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  XOR2_X1 U8046 ( .A(n6859), .B(n6862), .Z(n6860) );
  AOI22_X1 U8047 ( .A1(n7177), .A2(\adder_stage1[2][1] ), .B1(n6875), .B2(
        n6860), .ZN(n6861) );
  INV_X1 U8048 ( .A(n6861), .ZN(n10134) );
  OR2_X1 U8049 ( .A1(\x_mult_f[4][0] ), .A2(\x_mult_f[5][0] ), .ZN(n6863) );
  AND2_X1 U8050 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  AOI22_X1 U8051 ( .A1(n7177), .A2(\adder_stage1[2][0] ), .B1(n6875), .B2(
        n6864), .ZN(n6865) );
  INV_X1 U8052 ( .A(n6865), .ZN(n10135) );
  OAI21_X1 U8053 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6873) );
  INV_X1 U8054 ( .A(n6869), .ZN(n6871) );
  NAND2_X1 U8055 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  XNOR2_X1 U8056 ( .A(n6873), .B(n6872), .ZN(n6874) );
  AOI22_X1 U8057 ( .A1(n7177), .A2(\adder_stage1[2][3] ), .B1(n6875), .B2(
        n6874), .ZN(n6876) );
  INV_X1 U8058 ( .A(n6876), .ZN(n10132) );
  AOI22_X1 U8059 ( .A1(n6877), .A2(\x_mult_f[4][0] ), .B1(n7971), .B2(
        \x_mult_f_int[4][0] ), .ZN(n6878) );
  INV_X1 U8060 ( .A(n6878), .ZN(n9335) );
  AND2_X1 U8061 ( .A1(n6879), .A2(n6883), .ZN(n8144) );
  NOR2_X1 U8062 ( .A1(\x_mult_f[14][12] ), .A2(\x_mult_f[15][12] ), .ZN(n6885)
         );
  INV_X1 U8063 ( .A(n6885), .ZN(n8149) );
  AND2_X1 U8064 ( .A1(n8144), .A2(n8149), .ZN(n6893) );
  OR2_X1 U8065 ( .A1(\x_mult_f[14][13] ), .A2(\x_mult_f[15][13] ), .ZN(n6895)
         );
  AND2_X1 U8066 ( .A1(n6893), .A2(n6895), .ZN(n6880) );
  NAND2_X1 U8067 ( .A1(n6880), .A2(n8145), .ZN(n6888) );
  INV_X1 U8068 ( .A(n6881), .ZN(n6882) );
  AOI21_X1 U8069 ( .B1(n6884), .B2(n6883), .A(n6882), .ZN(n8146) );
  NAND2_X1 U8070 ( .A1(\x_mult_f[14][12] ), .A2(\x_mult_f[15][12] ), .ZN(n8148) );
  OAI21_X1 U8071 ( .B1(n8146), .B2(n6885), .A(n8148), .ZN(n6892) );
  NAND2_X1 U8072 ( .A1(\x_mult_f[14][13] ), .A2(\x_mult_f[15][13] ), .ZN(n6894) );
  INV_X1 U8073 ( .A(n6894), .ZN(n6886) );
  AOI21_X1 U8074 ( .B1(n6892), .B2(n6895), .A(n6886), .ZN(n6887) );
  NAND2_X1 U8075 ( .A1(n6888), .A2(n6887), .ZN(n7770) );
  AOI22_X1 U8076 ( .A1(n6889), .A2(n8294), .B1(n7855), .B2(
        \adder_stage1[7][14] ), .ZN(n6890) );
  INV_X1 U8077 ( .A(n6890), .ZN(n10039) );
  AOI22_X1 U8078 ( .A1(\x_mult_f_int[15][6] ), .A2(n8294), .B1(n7855), .B2(
        \x_mult_f[15][6] ), .ZN(n6891) );
  INV_X1 U8079 ( .A(n6891), .ZN(n9118) );
  AOI21_X1 U8080 ( .B1(n8145), .B2(n6893), .A(n6892), .ZN(n6897) );
  NAND2_X1 U8081 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  XOR2_X1 U8082 ( .A(n6897), .B(n6896), .Z(n6898) );
  AOI22_X1 U8083 ( .A1(n6898), .A2(n8294), .B1(n7855), .B2(
        \adder_stage1[7][13] ), .ZN(n6899) );
  INV_X1 U8084 ( .A(n6899), .ZN(n10040) );
  INV_X1 U8085 ( .A(n6900), .ZN(n6902) );
  NAND2_X1 U8086 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  XOR2_X1 U8087 ( .A(n6904), .B(n6903), .Z(n6905) );
  AOI22_X1 U8088 ( .A1(n7041), .A2(\adder_stage1[11][6] ), .B1(n8167), .B2(
        n6905), .ZN(n6906) );
  INV_X1 U8089 ( .A(n6906), .ZN(n9980) );
  NAND2_X1 U8090 ( .A1(n3433), .A2(n6907), .ZN(n6909) );
  NAND2_X1 U8091 ( .A1(n6909), .A2(n6908), .ZN(n6913) );
  NAND2_X1 U8092 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  XNOR2_X1 U8093 ( .A(n6913), .B(n6912), .ZN(n6914) );
  AOI22_X1 U8094 ( .A1(n8340), .A2(\adder_stage1[11][10] ), .B1(n8167), .B2(
        n6914), .ZN(n6915) );
  INV_X1 U8095 ( .A(n6915), .ZN(n9976) );
  NAND2_X1 U8096 ( .A1(n7111), .A2(n6916), .ZN(n6917) );
  XNOR2_X1 U8097 ( .A(n3433), .B(n6917), .ZN(n6919) );
  AOI22_X1 U8098 ( .A1(n8313), .A2(\adder_stage1[11][8] ), .B1(n8167), .B2(
        n6919), .ZN(n6920) );
  INV_X1 U8099 ( .A(n6920), .ZN(n9978) );
  NAND2_X1 U8100 ( .A1(n6922), .A2(n6921), .ZN(n6923) );
  XNOR2_X1 U8101 ( .A(n6924), .B(n6923), .ZN(n6925) );
  AOI22_X1 U8102 ( .A1(n8340), .A2(\adder_stage3[3][10] ), .B1(n8167), .B2(
        n6925), .ZN(n6926) );
  INV_X1 U8103 ( .A(n6926), .ZN(n9698) );
  AOI22_X1 U8104 ( .A1(n8057), .A2(\x_mult_f[23][1] ), .B1(n8167), .B2(
        \x_mult_f_int[23][1] ), .ZN(n6927) );
  INV_X1 U8105 ( .A(n6927), .ZN(n9372) );
  AOI22_X1 U8106 ( .A1(n8434), .A2(\x_mult_f[23][0] ), .B1(n8167), .B2(
        \x_mult_f_int[23][0] ), .ZN(n6928) );
  INV_X1 U8107 ( .A(n6928), .ZN(n9373) );
  NAND2_X1 U8108 ( .A1(n6930), .A2(n6929), .ZN(n6931) );
  XNOR2_X1 U8109 ( .A(n6932), .B(n6931), .ZN(n6933) );
  AOI22_X1 U8110 ( .A1(n8273), .A2(\adder_stage1[11][12] ), .B1(n8167), .B2(
        n6933), .ZN(n6934) );
  INV_X1 U8111 ( .A(n6934), .ZN(n9974) );
  AOI22_X1 U8112 ( .A1(n8313), .A2(\x_mult_f[23][4] ), .B1(n8167), .B2(
        \x_mult_f_int[23][4] ), .ZN(n6935) );
  INV_X1 U8113 ( .A(n6935), .ZN(n9221) );
  NAND2_X1 U8114 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  XNOR2_X1 U8115 ( .A(n6939), .B(n6938), .ZN(n6940) );
  AOI22_X1 U8116 ( .A1(n8325), .A2(\adder_stage3[3][14] ), .B1(n8167), .B2(
        n6940), .ZN(n6941) );
  INV_X1 U8117 ( .A(n6941), .ZN(n9694) );
  AOI22_X1 U8118 ( .A1(n8296), .A2(\x_mult_f[23][2] ), .B1(n8167), .B2(
        \x_mult_f_int[23][2] ), .ZN(n6942) );
  INV_X1 U8119 ( .A(n6942), .ZN(n9223) );
  OR2_X1 U8120 ( .A1(\adder_stage1[12][0] ), .A2(\adder_stage1[13][0] ), .ZN(
        n6943) );
  AND2_X1 U8121 ( .A1(n6943), .A2(n6953), .ZN(n6944) );
  AOI22_X1 U8122 ( .A1(n7041), .A2(\adder_stage2[6][0] ), .B1(n8292), .B2(
        n6944), .ZN(n6945) );
  INV_X1 U8123 ( .A(n6945), .ZN(n9803) );
  INV_X1 U8124 ( .A(n6946), .ZN(n7606) );
  NAND2_X1 U8125 ( .A1(n7606), .A2(n7604), .ZN(n6947) );
  XNOR2_X1 U8126 ( .A(n7607), .B(n6947), .ZN(n6948) );
  AOI22_X1 U8127 ( .A1(n7614), .A2(\adder_stage1[10][4] ), .B1(n8292), .B2(
        n6948), .ZN(n6949) );
  INV_X1 U8128 ( .A(n6949), .ZN(n9999) );
  OR2_X1 U8129 ( .A1(\adder_stage1[12][12] ), .A2(\adder_stage1[13][12] ), 
        .ZN(n7665) );
  NOR2_X1 U8130 ( .A1(\adder_stage1[12][11] ), .A2(\adder_stage1[13][11] ), 
        .ZN(n7662) );
  INV_X1 U8131 ( .A(n7662), .ZN(n7624) );
  NAND2_X1 U8132 ( .A1(n7665), .A2(n7624), .ZN(n7643) );
  INV_X1 U8133 ( .A(n7643), .ZN(n6950) );
  NOR2_X1 U8134 ( .A1(\adder_stage1[12][13] ), .A2(\adder_stage1[13][13] ), 
        .ZN(n6967) );
  INV_X1 U8135 ( .A(n6967), .ZN(n7646) );
  NAND2_X1 U8136 ( .A1(n6950), .A2(n7646), .ZN(n7573) );
  INV_X1 U8137 ( .A(n7573), .ZN(n6951) );
  NOR2_X1 U8138 ( .A1(\adder_stage1[12][14] ), .A2(\adder_stage1[13][14] ), 
        .ZN(n6969) );
  INV_X1 U8139 ( .A(n6969), .ZN(n7575) );
  AND2_X1 U8140 ( .A1(n6951), .A2(n7575), .ZN(n6972) );
  NOR2_X1 U8141 ( .A1(\adder_stage1[12][2] ), .A2(\adder_stage1[13][2] ), .ZN(
        n7616) );
  NOR2_X1 U8142 ( .A1(n7616), .A2(n6987), .ZN(n6956) );
  OAI21_X1 U8143 ( .B1(n6954), .B2(n6953), .A(n6952), .ZN(n6986) );
  NAND2_X1 U8144 ( .A1(\adder_stage1[12][2] ), .A2(\adder_stage1[13][2] ), 
        .ZN(n7617) );
  NAND2_X1 U8145 ( .A1(\adder_stage1[12][3] ), .A2(\adder_stage1[13][3] ), 
        .ZN(n6988) );
  OAI21_X1 U8146 ( .B1(n6987), .B2(n7617), .A(n6988), .ZN(n6955) );
  NOR2_X1 U8147 ( .A1(\adder_stage1[12][4] ), .A2(\adder_stage1[13][4] ), .ZN(
        n6977) );
  NOR2_X1 U8148 ( .A1(\adder_stage1[12][5] ), .A2(\adder_stage1[13][5] ), .ZN(
        n6979) );
  NOR2_X1 U8149 ( .A1(n6977), .A2(n6979), .ZN(n7008) );
  NOR2_X1 U8150 ( .A1(\adder_stage1[12][7] ), .A2(\adder_stage1[13][7] ), .ZN(
        n7016) );
  NOR2_X1 U8151 ( .A1(\adder_stage1[12][6] ), .A2(\adder_stage1[13][6] ), .ZN(
        n7014) );
  NOR2_X1 U8152 ( .A1(n7016), .A2(n7014), .ZN(n6958) );
  NAND2_X1 U8153 ( .A1(n7008), .A2(n6958), .ZN(n6960) );
  NAND2_X1 U8154 ( .A1(\adder_stage1[12][4] ), .A2(\adder_stage1[13][4] ), 
        .ZN(n7023) );
  NAND2_X1 U8155 ( .A1(\adder_stage1[12][5] ), .A2(\adder_stage1[13][5] ), 
        .ZN(n6980) );
  OAI21_X1 U8156 ( .B1(n6979), .B2(n7023), .A(n6980), .ZN(n7007) );
  NAND2_X1 U8157 ( .A1(\adder_stage1[12][6] ), .A2(\adder_stage1[13][6] ), 
        .ZN(n7013) );
  NAND2_X1 U8158 ( .A1(\adder_stage1[12][7] ), .A2(\adder_stage1[13][7] ), 
        .ZN(n7017) );
  OAI21_X1 U8159 ( .B1(n7016), .B2(n7013), .A(n7017), .ZN(n6957) );
  AOI21_X1 U8160 ( .B1(n6958), .B2(n7007), .A(n6957), .ZN(n6959) );
  OAI21_X1 U8161 ( .B1(n6976), .B2(n6960), .A(n6959), .ZN(n6994) );
  NOR2_X1 U8162 ( .A1(\adder_stage1[12][8] ), .A2(\adder_stage1[13][8] ), .ZN(
        n7000) );
  INV_X1 U8163 ( .A(n7000), .ZN(n6995) );
  OR2_X1 U8164 ( .A1(\adder_stage1[12][9] ), .A2(\adder_stage1[13][9] ), .ZN(
        n7002) );
  NAND2_X1 U8165 ( .A1(n6995), .A2(n7002), .ZN(n7652) );
  NOR2_X1 U8166 ( .A1(\adder_stage1[12][10] ), .A2(\adder_stage1[13][10] ), 
        .ZN(n7654) );
  NOR2_X1 U8167 ( .A1(n7652), .A2(n7654), .ZN(n6964) );
  NAND2_X1 U8168 ( .A1(\adder_stage1[12][8] ), .A2(\adder_stage1[13][8] ), 
        .ZN(n6999) );
  INV_X1 U8169 ( .A(n6999), .ZN(n6962) );
  NAND2_X1 U8170 ( .A1(\adder_stage1[12][9] ), .A2(\adder_stage1[13][9] ), 
        .ZN(n7001) );
  INV_X1 U8171 ( .A(n7001), .ZN(n6961) );
  AOI21_X1 U8172 ( .B1(n7002), .B2(n6962), .A(n6961), .ZN(n7651) );
  NAND2_X1 U8173 ( .A1(\adder_stage1[12][10] ), .A2(\adder_stage1[13][10] ), 
        .ZN(n7655) );
  OAI21_X1 U8174 ( .B1(n7651), .B2(n7654), .A(n7655), .ZN(n6963) );
  INV_X1 U8175 ( .A(n7663), .ZN(n6971) );
  NAND2_X1 U8176 ( .A1(\adder_stage1[12][11] ), .A2(\adder_stage1[13][11] ), 
        .ZN(n7661) );
  INV_X1 U8177 ( .A(n7661), .ZN(n6966) );
  NAND2_X1 U8178 ( .A1(\adder_stage1[12][12] ), .A2(\adder_stage1[13][12] ), 
        .ZN(n7664) );
  INV_X1 U8179 ( .A(n7664), .ZN(n6965) );
  AOI21_X1 U8180 ( .B1(n7665), .B2(n6966), .A(n6965), .ZN(n7642) );
  NAND2_X1 U8181 ( .A1(\adder_stage1[12][13] ), .A2(\adder_stage1[13][13] ), 
        .ZN(n7645) );
  OAI21_X1 U8182 ( .B1(n7642), .B2(n6967), .A(n7645), .ZN(n6968) );
  INV_X1 U8183 ( .A(n6968), .ZN(n7572) );
  NAND2_X1 U8184 ( .A1(\adder_stage1[12][14] ), .A2(\adder_stage1[13][14] ), 
        .ZN(n7574) );
  OAI21_X1 U8185 ( .B1(n7572), .B2(n6969), .A(n7574), .ZN(n6970) );
  AOI21_X1 U8186 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6973) );
  INV_X1 U8187 ( .A(n6973), .ZN(n7902) );
  AOI22_X1 U8188 ( .A1(n6974), .A2(n8311), .B1(n8338), .B2(
        \adder_stage2[6][15] ), .ZN(n6975) );
  INV_X1 U8189 ( .A(n6975), .ZN(n9788) );
  INV_X2 U8190 ( .A(n3409), .ZN(n7669) );
  BUF_X2 U8191 ( .A(n6238), .Z(n7627) );
  INV_X1 U8192 ( .A(n6976), .ZN(n7026) );
  INV_X1 U8193 ( .A(n6977), .ZN(n7024) );
  INV_X1 U8194 ( .A(n7023), .ZN(n6978) );
  AOI21_X1 U8195 ( .B1(n7026), .B2(n7024), .A(n6978), .ZN(n6983) );
  INV_X1 U8196 ( .A(n6979), .ZN(n6981) );
  NAND2_X1 U8197 ( .A1(n6981), .A2(n6980), .ZN(n6982) );
  XOR2_X1 U8198 ( .A(n6983), .B(n6982), .Z(n6984) );
  AOI22_X1 U8199 ( .A1(n7669), .A2(\adder_stage2[6][5] ), .B1(n7627), .B2(
        n6984), .ZN(n6985) );
  INV_X1 U8200 ( .A(n6985), .ZN(n9798) );
  INV_X1 U8201 ( .A(n6986), .ZN(n7620) );
  OAI21_X1 U8202 ( .B1(n7620), .B2(n7616), .A(n7617), .ZN(n6991) );
  INV_X1 U8203 ( .A(n6987), .ZN(n6989) );
  NAND2_X1 U8204 ( .A1(n6989), .A2(n6988), .ZN(n6990) );
  XNOR2_X1 U8205 ( .A(n6991), .B(n6990), .ZN(n6992) );
  AOI22_X1 U8206 ( .A1(n7669), .A2(\adder_stage2[6][3] ), .B1(n7627), .B2(
        n6992), .ZN(n6993) );
  INV_X1 U8207 ( .A(n6993), .ZN(n9800) );
  INV_X1 U8208 ( .A(n6994), .ZN(n7653) );
  NAND2_X1 U8209 ( .A1(n6995), .A2(n6999), .ZN(n6996) );
  XOR2_X1 U8210 ( .A(n7653), .B(n6996), .Z(n6997) );
  AOI22_X1 U8211 ( .A1(n7669), .A2(\adder_stage2[6][8] ), .B1(n7627), .B2(
        n6997), .ZN(n6998) );
  INV_X1 U8212 ( .A(n6998), .ZN(n9795) );
  OAI21_X1 U8213 ( .B1(n7653), .B2(n7000), .A(n6999), .ZN(n7004) );
  NAND2_X1 U8214 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  XNOR2_X1 U8215 ( .A(n7004), .B(n7003), .ZN(n7005) );
  AOI22_X1 U8216 ( .A1(n7669), .A2(\adder_stage2[6][9] ), .B1(n7627), .B2(
        n7005), .ZN(n7006) );
  INV_X1 U8217 ( .A(n7006), .ZN(n9794) );
  AOI21_X1 U8218 ( .B1(n7026), .B2(n7008), .A(n7007), .ZN(n7015) );
  INV_X1 U8219 ( .A(n7014), .ZN(n7009) );
  NAND2_X1 U8220 ( .A1(n7009), .A2(n7013), .ZN(n7010) );
  XOR2_X1 U8221 ( .A(n7015), .B(n7010), .Z(n7011) );
  AOI22_X1 U8222 ( .A1(n7669), .A2(\adder_stage2[6][6] ), .B1(n7627), .B2(
        n7011), .ZN(n7012) );
  INV_X1 U8223 ( .A(n7012), .ZN(n9797) );
  OAI21_X1 U8224 ( .B1(n7015), .B2(n7014), .A(n7013), .ZN(n7020) );
  INV_X1 U8225 ( .A(n7016), .ZN(n7018) );
  NAND2_X1 U8226 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  XNOR2_X1 U8227 ( .A(n7020), .B(n7019), .ZN(n7021) );
  AOI22_X1 U8228 ( .A1(n7669), .A2(\adder_stage2[6][7] ), .B1(n7627), .B2(
        n7021), .ZN(n7022) );
  INV_X1 U8229 ( .A(n7022), .ZN(n9796) );
  NAND2_X1 U8230 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  XNOR2_X1 U8231 ( .A(n7026), .B(n7025), .ZN(n7027) );
  AOI22_X1 U8232 ( .A1(n7669), .A2(\adder_stage2[6][4] ), .B1(n7627), .B2(
        n7027), .ZN(n7028) );
  INV_X1 U8233 ( .A(n7028), .ZN(n9799) );
  NAND2_X1 U8234 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  XNOR2_X1 U8235 ( .A(n3421), .B(n7031), .ZN(n7033) );
  AOI22_X1 U8236 ( .A1(n7041), .A2(\adder_stage2[1][14] ), .B1(n8189), .B2(
        n7033), .ZN(n7034) );
  INV_X1 U8237 ( .A(n7034), .ZN(n9873) );
  INV_X1 U8238 ( .A(n7035), .ZN(n7037) );
  NAND2_X1 U8239 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  XOR2_X1 U8240 ( .A(n7039), .B(n7038), .Z(n7040) );
  AOI22_X1 U8241 ( .A1(n7041), .A2(\adder_stage2[1][13] ), .B1(n8189), .B2(
        n7040), .ZN(n7042) );
  INV_X1 U8242 ( .A(n7042), .ZN(n9874) );
  BUF_X2 U8243 ( .A(n4645), .Z(n8105) );
  AOI22_X1 U8244 ( .A1(n7928), .A2(\x_mult_f[29][0] ), .B1(n8105), .B2(
        \x_mult_f_int[29][0] ), .ZN(n7043) );
  INV_X1 U8245 ( .A(n7043), .ZN(n9385) );
  AOI22_X1 U8246 ( .A1(n7928), .A2(\x_mult_f[29][4] ), .B1(n8105), .B2(
        \x_mult_f_int[29][4] ), .ZN(n7044) );
  INV_X1 U8247 ( .A(n7044), .ZN(n9297) );
  AOI22_X1 U8248 ( .A1(n7855), .A2(\x_mult_f[26][3] ), .B1(n8105), .B2(
        \x_mult_f_int[26][3] ), .ZN(n7045) );
  INV_X1 U8249 ( .A(n7045), .ZN(n9256) );
  NAND2_X1 U8250 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  XOR2_X1 U8251 ( .A(n7049), .B(n7048), .Z(n7050) );
  AOI22_X1 U8252 ( .A1(n7074), .A2(\adder_stage2[2][11] ), .B1(n8117), .B2(
        n7050), .ZN(n7051) );
  INV_X1 U8253 ( .A(n7051), .ZN(n9859) );
  INV_X1 U8254 ( .A(n7052), .ZN(n7072) );
  OAI21_X1 U8255 ( .B1(n7072), .B2(n7053), .A(n7069), .ZN(n7057) );
  NAND2_X1 U8256 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  XNOR2_X1 U8257 ( .A(n7057), .B(n7056), .ZN(n7058) );
  AOI22_X1 U8258 ( .A1(n7074), .A2(\adder_stage2[2][9] ), .B1(n8117), .B2(
        n7058), .ZN(n7059) );
  INV_X1 U8259 ( .A(n7059), .ZN(n9861) );
  OAI21_X1 U8260 ( .B1(n7072), .B2(n7061), .A(n7060), .ZN(n7066) );
  INV_X1 U8261 ( .A(n7062), .ZN(n7064) );
  NAND2_X1 U8262 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  XNOR2_X1 U8263 ( .A(n7066), .B(n7065), .ZN(n7067) );
  AOI22_X1 U8264 ( .A1(n7074), .A2(\adder_stage2[2][10] ), .B1(n8117), .B2(
        n7067), .ZN(n7068) );
  INV_X1 U8265 ( .A(n7068), .ZN(n9860) );
  NAND2_X1 U8266 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  XOR2_X1 U8267 ( .A(n7072), .B(n7071), .Z(n7073) );
  AOI22_X1 U8268 ( .A1(n7074), .A2(\adder_stage2[2][8] ), .B1(n8117), .B2(
        n7073), .ZN(n7075) );
  INV_X1 U8269 ( .A(n7075), .ZN(n9862) );
  OR2_X1 U8270 ( .A1(\x_mult_f[20][0] ), .A2(\x_mult_f[21][0] ), .ZN(n7076) );
  AND2_X1 U8271 ( .A1(n7076), .A2(n7092), .ZN(n7077) );
  AOI22_X1 U8272 ( .A1(n8118), .A2(\adder_stage1[10][0] ), .B1(n8292), .B2(
        n7077), .ZN(n7078) );
  INV_X1 U8273 ( .A(n7078), .ZN(n10002) );
  OAI21_X1 U8274 ( .B1(n7081), .B2(n7080), .A(n7079), .ZN(n7086) );
  INV_X1 U8275 ( .A(n7082), .ZN(n7084) );
  NAND2_X1 U8276 ( .A1(n7084), .A2(n7083), .ZN(n7085) );
  XNOR2_X1 U8277 ( .A(n7086), .B(n7085), .ZN(n7087) );
  AOI22_X1 U8278 ( .A1(n8330), .A2(\adder_stage3[3][3] ), .B1(n7627), .B2(
        n7087), .ZN(n7088) );
  INV_X1 U8279 ( .A(n7088), .ZN(n9705) );
  INV_X1 U8280 ( .A(n7089), .ZN(n7091) );
  NAND2_X1 U8281 ( .A1(n7091), .A2(n7090), .ZN(n7093) );
  XOR2_X1 U8282 ( .A(n7093), .B(n7092), .Z(n7094) );
  AOI22_X1 U8283 ( .A1(n8434), .A2(\adder_stage1[10][1] ), .B1(n8292), .B2(
        n7094), .ZN(n7095) );
  INV_X1 U8284 ( .A(n7095), .ZN(n10001) );
  OR2_X1 U8285 ( .A1(\adder_stage1[14][0] ), .A2(\adder_stage1[15][0] ), .ZN(
        n7097) );
  AND2_X1 U8286 ( .A1(n7097), .A2(n7096), .ZN(n7098) );
  AOI22_X1 U8287 ( .A1(n8325), .A2(\adder_stage2[7][0] ), .B1(n7627), .B2(
        n7098), .ZN(n7099) );
  INV_X1 U8288 ( .A(n7099), .ZN(n9786) );
  INV_X1 U8289 ( .A(n7100), .ZN(n7253) );
  INV_X1 U8290 ( .A(n7101), .ZN(n7119) );
  INV_X1 U8291 ( .A(n7118), .ZN(n7102) );
  AOI21_X1 U8292 ( .B1(n7253), .B2(n7119), .A(n7102), .ZN(n7107) );
  INV_X1 U8293 ( .A(n7103), .ZN(n7105) );
  NAND2_X1 U8294 ( .A1(n7105), .A2(n7104), .ZN(n7106) );
  XOR2_X1 U8295 ( .A(n7107), .B(n7106), .Z(n7108) );
  AOI22_X1 U8296 ( .A1(n7959), .A2(\adder_stage3[3][5] ), .B1(n7627), .B2(
        n7108), .ZN(n7109) );
  INV_X1 U8297 ( .A(n7109), .ZN(n9703) );
  AOI21_X1 U8298 ( .B1(n3433), .B2(n7111), .A(n7110), .ZN(n7115) );
  NAND2_X1 U8299 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  XOR2_X1 U8300 ( .A(n7115), .B(n7114), .Z(n7116) );
  AOI22_X1 U8301 ( .A1(n8338), .A2(\adder_stage1[11][9] ), .B1(n7627), .B2(
        n7116), .ZN(n7117) );
  INV_X1 U8302 ( .A(n7117), .ZN(n9977) );
  NAND2_X1 U8303 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  XNOR2_X1 U8304 ( .A(n7253), .B(n7120), .ZN(n7121) );
  AOI22_X1 U8305 ( .A1(n7928), .A2(\adder_stage3[3][4] ), .B1(n7627), .B2(
        n7121), .ZN(n7122) );
  INV_X1 U8306 ( .A(n7122), .ZN(n9704) );
  AOI22_X1 U8307 ( .A1(\x_mult_f_int[31][11] ), .A2(n8304), .B1(n8325), .B2(
        \x_mult_f[31][11] ), .ZN(n7123) );
  INV_X1 U8308 ( .A(n7123), .ZN(n9318) );
  AOI22_X1 U8309 ( .A1(\x_mult_f_int[31][8] ), .A2(n8304), .B1(n8330), .B2(
        \x_mult_f[31][8] ), .ZN(n7124) );
  INV_X1 U8310 ( .A(n7124), .ZN(n9321) );
  AOI22_X1 U8311 ( .A1(\x_mult_f_int[31][10] ), .A2(n8304), .B1(n8328), .B2(
        \x_mult_f[31][10] ), .ZN(n7125) );
  INV_X1 U8312 ( .A(n7125), .ZN(n9319) );
  AOI22_X1 U8313 ( .A1(\x_mult_f_int[31][9] ), .A2(n8304), .B1(n7614), .B2(
        \x_mult_f[31][9] ), .ZN(n7126) );
  INV_X1 U8314 ( .A(n7126), .ZN(n9320) );
  AOI22_X1 U8315 ( .A1(n7952), .A2(\x_mult_f[29][5] ), .B1(n8105), .B2(
        \x_mult_f_int[29][5] ), .ZN(n7127) );
  INV_X1 U8316 ( .A(n7127), .ZN(n9296) );
  AOI22_X1 U8317 ( .A1(\x_mult_f_int[1][7] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[1][7] ), .ZN(n7128) );
  INV_X1 U8318 ( .A(n7128), .ZN(n8935) );
  AOI22_X1 U8319 ( .A1(\x_mult_f_int[29][11] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][11] ), .ZN(n7129) );
  INV_X1 U8320 ( .A(n7129), .ZN(n9290) );
  AOI22_X1 U8321 ( .A1(\x_mult_f_int[0][8] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[0][8] ), .ZN(n7130) );
  INV_X1 U8322 ( .A(n7130), .ZN(n8920) );
  AOI22_X1 U8323 ( .A1(\x_mult_f_int[0][6] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[0][6] ), .ZN(n7131) );
  INV_X1 U8324 ( .A(n7131), .ZN(n8922) );
  AOI22_X1 U8325 ( .A1(\x_mult_f_int[0][7] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[0][7] ), .ZN(n7132) );
  INV_X1 U8326 ( .A(n7132), .ZN(n8921) );
  AOI22_X1 U8327 ( .A1(\x_mult_f_int[1][11] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[1][11] ), .ZN(n7133) );
  INV_X1 U8328 ( .A(n7133), .ZN(n8931) );
  AOI22_X1 U8329 ( .A1(\x_mult_f_int[29][10] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][10] ), .ZN(n7134) );
  INV_X1 U8330 ( .A(n7134), .ZN(n9291) );
  INV_X1 U8331 ( .A(n7135), .ZN(n7136) );
  NAND2_X1 U8332 ( .A1(n7136), .A2(n7137), .ZN(n7143) );
  INV_X1 U8333 ( .A(n7137), .ZN(n7139) );
  OAI21_X1 U8334 ( .B1(n7140), .B2(n7139), .A(n7138), .ZN(n7141) );
  INV_X1 U8335 ( .A(n7141), .ZN(n7142) );
  OAI21_X1 U8336 ( .B1(n8239), .B2(n7143), .A(n7142), .ZN(n7144) );
  INV_X1 U8337 ( .A(n7144), .ZN(n8082) );
  NOR2_X1 U8338 ( .A1(\adder_stage2[0][19] ), .A2(\adder_stage2[1][19] ), .ZN(
        n8081) );
  INV_X1 U8339 ( .A(n8081), .ZN(n7145) );
  NAND2_X1 U8340 ( .A1(\adder_stage2[0][19] ), .A2(\adder_stage2[1][19] ), 
        .ZN(n8080) );
  NAND2_X1 U8341 ( .A1(n7145), .A2(n8080), .ZN(n7146) );
  XOR2_X1 U8342 ( .A(n8082), .B(n7146), .Z(n7147) );
  AOI22_X1 U8343 ( .A1(n7147), .A2(n8298), .B1(n8328), .B2(
        \adder_stage3[0][19] ), .ZN(n7148) );
  INV_X1 U8344 ( .A(n7148), .ZN(n9750) );
  AOI22_X1 U8345 ( .A1(\x_mult_f_int[27][8] ), .A2(n7819), .B1(n7864), .B2(
        \x_mult_f[27][8] ), .ZN(n7149) );
  INV_X1 U8346 ( .A(n7149), .ZN(n9265) );
  AOI22_X1 U8347 ( .A1(\x_mult_f_int[27][9] ), .A2(n7819), .B1(n7864), .B2(
        \x_mult_f[27][9] ), .ZN(n7150) );
  INV_X1 U8348 ( .A(n7150), .ZN(n9264) );
  AOI22_X1 U8349 ( .A1(n7074), .A2(\x_mult_f[12][4] ), .B1(n7155), .B2(
        \x_mult_f_int[12][4] ), .ZN(n7151) );
  INV_X1 U8350 ( .A(n7151), .ZN(n9078) );
  AOI22_X1 U8351 ( .A1(n6854), .A2(\x_mult_f[12][3] ), .B1(n7155), .B2(
        \x_mult_f_int[12][3] ), .ZN(n7152) );
  INV_X1 U8352 ( .A(n7152), .ZN(n9079) );
  AOI22_X1 U8353 ( .A1(n7525), .A2(\x_mult_f[12][1] ), .B1(n7155), .B2(
        \x_mult_f_int[12][1] ), .ZN(n7153) );
  INV_X1 U8354 ( .A(n7153), .ZN(n9350) );
  AOI22_X1 U8355 ( .A1(n7525), .A2(\x_mult_f[12][2] ), .B1(n7155), .B2(
        \x_mult_f_int[12][2] ), .ZN(n7154) );
  INV_X1 U8356 ( .A(n7154), .ZN(n9080) );
  AOI22_X1 U8357 ( .A1(n7525), .A2(\x_mult_f[12][0] ), .B1(n7155), .B2(
        \x_mult_f_int[12][0] ), .ZN(n7156) );
  INV_X1 U8358 ( .A(n7156), .ZN(n9351) );
  OAI21_X1 U8359 ( .B1(n7159), .B2(n7158), .A(n7157), .ZN(n8214) );
  OR2_X1 U8360 ( .A1(\adder_stage1[10][14] ), .A2(\adder_stage1[11][14] ), 
        .ZN(n8212) );
  NAND2_X1 U8361 ( .A1(n8214), .A2(n8212), .ZN(n7160) );
  NAND2_X1 U8362 ( .A1(\adder_stage1[10][14] ), .A2(\adder_stage1[11][14] ), 
        .ZN(n8211) );
  NAND2_X1 U8363 ( .A1(n7160), .A2(n8211), .ZN(n7994) );
  AOI22_X1 U8364 ( .A1(n7161), .A2(n6875), .B1(n8296), .B2(
        \adder_stage2[5][15] ), .ZN(n7162) );
  INV_X1 U8365 ( .A(n7162), .ZN(n9804) );
  INV_X1 U8366 ( .A(n7164), .ZN(n7166) );
  NAND2_X1 U8367 ( .A1(n7166), .A2(n7165), .ZN(n7167) );
  XOR2_X1 U8368 ( .A(n7168), .B(n7167), .Z(n7169) );
  AOI22_X1 U8369 ( .A1(n8245), .A2(\adder_stage3[0][13] ), .B1(n8024), .B2(
        n7169), .ZN(n7170) );
  INV_X1 U8370 ( .A(n7170), .ZN(n9756) );
  INV_X1 U8371 ( .A(n7171), .ZN(n7173) );
  NAND2_X1 U8372 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  XOR2_X1 U8373 ( .A(n7175), .B(n7174), .Z(n7176) );
  AOI22_X1 U8374 ( .A1(n7177), .A2(\adder_stage2[1][6] ), .B1(n6272), .B2(
        n7176), .ZN(n7178) );
  INV_X1 U8375 ( .A(n7178), .ZN(n9881) );
  INV_X1 U8376 ( .A(n7179), .ZN(n7223) );
  NAND2_X1 U8377 ( .A1(n7223), .A2(n7221), .ZN(n7180) );
  XNOR2_X1 U8378 ( .A(n7224), .B(n7180), .ZN(n7181) );
  AOI22_X1 U8379 ( .A1(n8245), .A2(\adder_stage2[1][4] ), .B1(n8209), .B2(
        n7181), .ZN(n7182) );
  INV_X1 U8380 ( .A(n7182), .ZN(n9883) );
  INV_X1 U8381 ( .A(n7183), .ZN(n7218) );
  OAI21_X1 U8382 ( .B1(n7218), .B2(n7214), .A(n7215), .ZN(n7188) );
  INV_X1 U8383 ( .A(n7184), .ZN(n7186) );
  NAND2_X1 U8384 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  XNOR2_X1 U8385 ( .A(n7188), .B(n7187), .ZN(n7189) );
  AOI22_X1 U8386 ( .A1(n8245), .A2(\adder_stage2[1][3] ), .B1(n6036), .B2(
        n7189), .ZN(n7190) );
  INV_X1 U8387 ( .A(n7190), .ZN(n9884) );
  NAND2_X1 U8388 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  XNOR2_X1 U8389 ( .A(n7194), .B(n7193), .ZN(n7195) );
  AOI22_X1 U8390 ( .A1(n8245), .A2(\adder_stage3[0][14] ), .B1(n8024), .B2(
        n7195), .ZN(n7196) );
  INV_X1 U8391 ( .A(n7196), .ZN(n9755) );
  INV_X1 U8392 ( .A(n7197), .ZN(n7200) );
  INV_X1 U8393 ( .A(n7198), .ZN(n7199) );
  OAI21_X1 U8394 ( .B1(n7513), .B2(n7200), .A(n7199), .ZN(n7638) );
  INV_X1 U8395 ( .A(n7201), .ZN(n7636) );
  INV_X1 U8396 ( .A(n7635), .ZN(n7202) );
  AOI21_X1 U8397 ( .B1(n7638), .B2(n7636), .A(n7202), .ZN(n7207) );
  INV_X1 U8398 ( .A(n7203), .ZN(n7205) );
  NAND2_X1 U8399 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  XOR2_X1 U8400 ( .A(n7207), .B(n7206), .Z(n7208) );
  AOI22_X1 U8401 ( .A1(n7640), .A2(\adder_stage3[0][11] ), .B1(n8117), .B2(
        n7208), .ZN(n7209) );
  INV_X1 U8402 ( .A(n7209), .ZN(n9758) );
  NAND2_X1 U8403 ( .A1(n7210), .A2(n8237), .ZN(n7211) );
  XOR2_X1 U8404 ( .A(n8239), .B(n7211), .Z(n7212) );
  AOI22_X1 U8405 ( .A1(n8245), .A2(\adder_stage3[0][15] ), .B1(n6036), .B2(
        n7212), .ZN(n7213) );
  INV_X1 U8406 ( .A(n7213), .ZN(n9754) );
  INV_X1 U8407 ( .A(n7214), .ZN(n7216) );
  NAND2_X1 U8408 ( .A1(n7216), .A2(n7215), .ZN(n7217) );
  XOR2_X1 U8409 ( .A(n7218), .B(n7217), .Z(n7219) );
  AOI22_X1 U8410 ( .A1(n8245), .A2(\adder_stage2[1][2] ), .B1(n6272), .B2(
        n7219), .ZN(n7220) );
  INV_X1 U8411 ( .A(n7220), .ZN(n9885) );
  INV_X1 U8412 ( .A(n7221), .ZN(n7222) );
  AOI21_X1 U8413 ( .B1(n7224), .B2(n7223), .A(n7222), .ZN(n7229) );
  INV_X1 U8414 ( .A(n7225), .ZN(n7227) );
  NAND2_X1 U8415 ( .A1(n7227), .A2(n7226), .ZN(n7228) );
  XOR2_X1 U8416 ( .A(n7229), .B(n7228), .Z(n7230) );
  AOI22_X1 U8417 ( .A1(n8245), .A2(\adder_stage2[1][5] ), .B1(n8209), .B2(
        n7230), .ZN(n7231) );
  INV_X1 U8418 ( .A(n7231), .ZN(n9882) );
  INV_X1 U8419 ( .A(n7232), .ZN(n7234) );
  NAND2_X1 U8420 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  XOR2_X1 U8421 ( .A(n7235), .B(n7238), .Z(n7236) );
  AOI22_X1 U8422 ( .A1(n8245), .A2(\adder_stage2[1][1] ), .B1(n6352), .B2(
        n7236), .ZN(n7237) );
  INV_X1 U8423 ( .A(n7237), .ZN(n9886) );
  OR2_X1 U8424 ( .A1(\adder_stage1[2][0] ), .A2(\adder_stage1[3][0] ), .ZN(
        n7239) );
  AND2_X1 U8425 ( .A1(n7239), .A2(n7238), .ZN(n7240) );
  AOI22_X1 U8426 ( .A1(n8245), .A2(\adder_stage2[1][0] ), .B1(n8235), .B2(
        n7240), .ZN(n7241) );
  INV_X1 U8427 ( .A(n7241), .ZN(n9887) );
  OAI21_X1 U8428 ( .B1(n7513), .B2(n7243), .A(n7242), .ZN(n7248) );
  INV_X1 U8429 ( .A(n7244), .ZN(n7246) );
  NAND2_X1 U8430 ( .A1(n7246), .A2(n7245), .ZN(n7247) );
  XNOR2_X1 U8431 ( .A(n7248), .B(n7247), .ZN(n7249) );
  AOI22_X1 U8432 ( .A1(n8245), .A2(\adder_stage3[0][12] ), .B1(n6636), .B2(
        n7249), .ZN(n7250) );
  INV_X1 U8433 ( .A(n7250), .ZN(n9757) );
  AOI21_X1 U8434 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(n7269) );
  INV_X1 U8435 ( .A(n7268), .ZN(n7254) );
  NAND2_X1 U8436 ( .A1(n7254), .A2(n7267), .ZN(n7255) );
  XOR2_X1 U8437 ( .A(n7269), .B(n7255), .Z(n7256) );
  AOI22_X1 U8438 ( .A1(n8273), .A2(\adder_stage3[3][6] ), .B1(n8105), .B2(
        n7256), .ZN(n7257) );
  INV_X1 U8439 ( .A(n7257), .ZN(n9702) );
  OAI21_X1 U8440 ( .B1(n8103), .B2(n7259), .A(n7258), .ZN(n7264) );
  INV_X1 U8441 ( .A(n7260), .ZN(n7262) );
  NAND2_X1 U8442 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  XNOR2_X1 U8443 ( .A(n7264), .B(n7263), .ZN(n7265) );
  AOI22_X1 U8444 ( .A1(n8434), .A2(\adder_stage3[3][12] ), .B1(n8105), .B2(
        n7265), .ZN(n7266) );
  INV_X1 U8445 ( .A(n7266), .ZN(n9696) );
  OAI21_X1 U8446 ( .B1(n7269), .B2(n7268), .A(n7267), .ZN(n7274) );
  INV_X1 U8447 ( .A(n7270), .ZN(n7272) );
  NAND2_X1 U8448 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  XNOR2_X1 U8449 ( .A(n7274), .B(n7273), .ZN(n7275) );
  AOI22_X1 U8450 ( .A1(n7928), .A2(\adder_stage3[3][7] ), .B1(n8105), .B2(
        n7275), .ZN(n7276) );
  INV_X1 U8451 ( .A(n7276), .ZN(n9701) );
  AOI22_X1 U8452 ( .A1(n7952), .A2(\x_mult_f[23][5] ), .B1(n8105), .B2(
        \x_mult_f_int[23][5] ), .ZN(n7277) );
  INV_X1 U8453 ( .A(n7277), .ZN(n9220) );
  AOI22_X1 U8454 ( .A1(n7959), .A2(\x_mult_f[23][3] ), .B1(n8105), .B2(
        \x_mult_f_int[23][3] ), .ZN(n7278) );
  INV_X1 U8455 ( .A(n7278), .ZN(n9222) );
  OAI21_X1 U8456 ( .B1(n8103), .B2(n8099), .A(n8100), .ZN(n7283) );
  INV_X1 U8457 ( .A(n7279), .ZN(n7281) );
  NAND2_X1 U8458 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  XNOR2_X1 U8459 ( .A(n7283), .B(n7282), .ZN(n7284) );
  AOI22_X1 U8460 ( .A1(n7556), .A2(\adder_stage3[3][9] ), .B1(n8105), .B2(
        n7284), .ZN(n7285) );
  INV_X1 U8461 ( .A(n7285), .ZN(n9699) );
  AOI22_X1 U8462 ( .A1(\x_mult_f_int[8][8] ), .A2(n6875), .B1(n8309), .B2(
        \x_mult_f[8][8] ), .ZN(n7286) );
  INV_X1 U8463 ( .A(n7286), .ZN(n9019) );
  AOI22_X1 U8464 ( .A1(\x_mult_f_int[8][11] ), .A2(n8294), .B1(n8309), .B2(
        \x_mult_f[8][11] ), .ZN(n7287) );
  INV_X1 U8465 ( .A(n7287), .ZN(n9016) );
  AOI22_X1 U8466 ( .A1(\x_mult_f_int[1][10] ), .A2(n8298), .B1(n8398), .B2(
        \x_mult_f[1][10] ), .ZN(n7288) );
  INV_X1 U8467 ( .A(n7288), .ZN(n8932) );
  AOI22_X1 U8468 ( .A1(\x_mult_f_int[1][8] ), .A2(n8298), .B1(n8398), .B2(
        \x_mult_f[1][8] ), .ZN(n7289) );
  INV_X1 U8469 ( .A(n7289), .ZN(n8934) );
  AOI22_X1 U8470 ( .A1(\x_mult_f_int[1][9] ), .A2(n8298), .B1(n8398), .B2(
        \x_mult_f[1][9] ), .ZN(n7290) );
  INV_X1 U8471 ( .A(n7290), .ZN(n8933) );
  AOI22_X1 U8472 ( .A1(\x_mult_f_int[8][13] ), .A2(n7507), .B1(n8323), .B2(
        \x_mult_f[8][13] ), .ZN(n7291) );
  INV_X1 U8473 ( .A(n7291), .ZN(n9014) );
  INV_X1 U8474 ( .A(n7292), .ZN(n7294) );
  NAND2_X1 U8475 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  XOR2_X1 U8476 ( .A(n7296), .B(n7295), .Z(n7297) );
  AOI22_X1 U8477 ( .A1(n7297), .A2(n8298), .B1(n8428), .B2(
        \adder_stage1[14][13] ), .ZN(n7298) );
  INV_X1 U8478 ( .A(n7298), .ZN(n9922) );
  AOI22_X1 U8479 ( .A1(\x_mult_f_int[12][8] ), .A2(n8105), .B1(n7855), .B2(
        \x_mult_f[12][8] ), .ZN(n7299) );
  INV_X1 U8480 ( .A(n7299), .ZN(n9074) );
  AOI22_X1 U8481 ( .A1(\x_mult_f_int[12][9] ), .A2(n8314), .B1(n7855), .B2(
        \x_mult_f[12][9] ), .ZN(n7300) );
  INV_X1 U8482 ( .A(n7300), .ZN(n9073) );
  AOI22_X1 U8483 ( .A1(\x_mult_f_int[12][10] ), .A2(n7819), .B1(n7855), .B2(
        \x_mult_f[12][10] ), .ZN(n7301) );
  INV_X1 U8484 ( .A(n7301), .ZN(n9072) );
  AOI22_X1 U8485 ( .A1(\x_mult_f_int[25][8] ), .A2(n4645), .B1(n8338), .B2(
        \x_mult_f[25][8] ), .ZN(n7302) );
  INV_X1 U8486 ( .A(n7302), .ZN(n9237) );
  AOI22_X1 U8487 ( .A1(\x_mult_f_int[27][10] ), .A2(n8167), .B1(n7864), .B2(
        \x_mult_f[27][10] ), .ZN(n7303) );
  INV_X1 U8488 ( .A(n7303), .ZN(n9263) );
  AOI22_X1 U8489 ( .A1(\x_mult_f_int[27][11] ), .A2(n8153), .B1(n7864), .B2(
        \x_mult_f[27][11] ), .ZN(n7304) );
  INV_X1 U8490 ( .A(n7304), .ZN(n9262) );
  AOI22_X1 U8491 ( .A1(\x_mult_f_int[12][11] ), .A2(n8314), .B1(n7855), .B2(
        \x_mult_f[12][11] ), .ZN(n7305) );
  INV_X1 U8492 ( .A(n7305), .ZN(n9071) );
  AOI22_X1 U8493 ( .A1(\x_mult_f_int[4][10] ), .A2(n5981), .B1(n8338), .B2(
        \x_mult_f[4][10] ), .ZN(n7306) );
  INV_X1 U8494 ( .A(n7306), .ZN(n8974) );
  AOI22_X1 U8495 ( .A1(\x_mult_f_int[4][11] ), .A2(n8258), .B1(n8338), .B2(
        \x_mult_f[4][11] ), .ZN(n7307) );
  INV_X1 U8496 ( .A(n7307), .ZN(n8973) );
  INV_X1 U8497 ( .A(n7308), .ZN(n7312) );
  NOR3_X1 U8498 ( .A1(n7310), .A2(n7312), .A3(n7309), .ZN(n7315) );
  OAI21_X1 U8499 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n7314) );
  OR2_X1 U8500 ( .A1(n7315), .A2(n7314), .ZN(n7884) );
  AOI22_X1 U8501 ( .A1(n7316), .A2(n7627), .B1(n8338), .B2(
        \adder_stage2[0][15] ), .ZN(n7317) );
  INV_X1 U8502 ( .A(n7317), .ZN(n9889) );
  OAI21_X1 U8503 ( .B1(n7320), .B2(n7319), .A(n7318), .ZN(n7969) );
  OR2_X1 U8504 ( .A1(\x_mult_f[4][12] ), .A2(\x_mult_f[5][12] ), .ZN(n7967) );
  NAND2_X1 U8505 ( .A1(\x_mult_f[4][12] ), .A2(\x_mult_f[5][12] ), .ZN(n7966)
         );
  INV_X1 U8506 ( .A(n7966), .ZN(n7321) );
  AOI21_X1 U8507 ( .B1(n7969), .B2(n7967), .A(n7321), .ZN(n8403) );
  NOR2_X1 U8508 ( .A1(\x_mult_f[4][13] ), .A2(\x_mult_f[5][13] ), .ZN(n8404)
         );
  NAND2_X1 U8509 ( .A1(\x_mult_f[4][13] ), .A2(\x_mult_f[5][13] ), .ZN(n8405)
         );
  OAI21_X1 U8510 ( .B1(n8403), .B2(n8404), .A(n8405), .ZN(n8044) );
  AOI22_X1 U8511 ( .A1(n7322), .A2(n8292), .B1(n8336), .B2(
        \adder_stage1[2][14] ), .ZN(n7323) );
  INV_X1 U8512 ( .A(n7323), .ZN(n10122) );
  OAI21_X1 U8513 ( .B1(n7326), .B2(n7325), .A(n7324), .ZN(n7957) );
  OR2_X1 U8514 ( .A1(\x_mult_f[30][12] ), .A2(\x_mult_f[31][12] ), .ZN(n7955)
         );
  NAND2_X1 U8515 ( .A1(\x_mult_f[30][12] ), .A2(\x_mult_f[31][12] ), .ZN(n7954) );
  INV_X1 U8516 ( .A(n7954), .ZN(n7327) );
  AOI21_X1 U8517 ( .B1(n7957), .B2(n7955), .A(n7327), .ZN(n8433) );
  NOR2_X1 U8518 ( .A1(\x_mult_f[30][13] ), .A2(\x_mult_f[31][13] ), .ZN(n8429)
         );
  NAND2_X1 U8519 ( .A1(\x_mult_f[30][13] ), .A2(\x_mult_f[31][13] ), .ZN(n8430) );
  OAI21_X1 U8520 ( .B1(n8433), .B2(n8429), .A(n8430), .ZN(n8127) );
  INV_X1 U8521 ( .A(n7328), .ZN(n7329) );
  AOI22_X1 U8522 ( .A1(n7329), .A2(n6626), .B1(n8319), .B2(
        \adder_stage1[15][20] ), .ZN(n7330) );
  INV_X1 U8523 ( .A(n7330), .ZN(n9905) );
  AOI22_X1 U8524 ( .A1(\x_mult_f_int[0][9] ), .A2(n8087), .B1(n8336), .B2(
        \x_mult_f[0][9] ), .ZN(n7331) );
  INV_X1 U8525 ( .A(n7331), .ZN(n8919) );
  AOI22_X1 U8526 ( .A1(\x_mult_f_int[0][10] ), .A2(n8167), .B1(n8336), .B2(
        \x_mult_f[0][10] ), .ZN(n7332) );
  INV_X1 U8527 ( .A(n7332), .ZN(n8918) );
  AOI22_X1 U8528 ( .A1(\x_mult_f_int[0][11] ), .A2(n7962), .B1(n8336), .B2(
        \x_mult_f[0][11] ), .ZN(n7333) );
  INV_X1 U8529 ( .A(n7333), .ZN(n8917) );
  AOI22_X1 U8530 ( .A1(n8328), .A2(\x_mult_f[8][0] ), .B1(n8087), .B2(
        \x_mult_f_int[8][0] ), .ZN(n7334) );
  INV_X1 U8531 ( .A(n7334), .ZN(n9343) );
  AOI22_X1 U8532 ( .A1(n8328), .A2(\x_mult_f[8][1] ), .B1(n8087), .B2(
        \x_mult_f_int[8][1] ), .ZN(n7335) );
  INV_X1 U8533 ( .A(n7335), .ZN(n9342) );
  INV_X1 U8534 ( .A(n7336), .ZN(n7338) );
  NAND2_X1 U8535 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
  XOR2_X1 U8536 ( .A(n7340), .B(n7339), .Z(n7341) );
  AOI22_X1 U8537 ( .A1(n7341), .A2(n6636), .B1(n7698), .B2(
        \adder_stage1[9][13] ), .ZN(n7342) );
  INV_X1 U8538 ( .A(n7342), .ZN(n10006) );
  BUF_X2 U8539 ( .A(n7343), .Z(n7450) );
  AOI22_X1 U8540 ( .A1(n8176), .A2(\x_mult_f[25][3] ), .B1(n7450), .B2(
        \x_mult_f_int[25][3] ), .ZN(n7344) );
  INV_X1 U8541 ( .A(n7344), .ZN(n9242) );
  AOI22_X1 U8542 ( .A1(n8176), .A2(\x_mult_f[25][5] ), .B1(n7450), .B2(
        \x_mult_f_int[25][5] ), .ZN(n7345) );
  INV_X1 U8543 ( .A(n7345), .ZN(n9240) );
  AOI22_X1 U8544 ( .A1(n8176), .A2(\x_mult_f[25][2] ), .B1(n7450), .B2(
        \x_mult_f_int[25][2] ), .ZN(n7346) );
  INV_X1 U8545 ( .A(n7346), .ZN(n9243) );
  OAI21_X1 U8546 ( .B1(n7349), .B2(n7348), .A(n7347), .ZN(n7394) );
  AOI21_X1 U8547 ( .B1(n7394), .B2(n7368), .A(n7350), .ZN(n7354) );
  NAND2_X1 U8548 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  XOR2_X1 U8549 ( .A(n7354), .B(n7353), .Z(n7355) );
  AOI22_X1 U8550 ( .A1(n7959), .A2(\adder_stage1[15][9] ), .B1(n7450), .B2(
        n7355), .ZN(n7356) );
  INV_X1 U8551 ( .A(n7356), .ZN(n9909) );
  AOI22_X1 U8552 ( .A1(n8176), .A2(\x_mult_f[25][4] ), .B1(n7450), .B2(
        \x_mult_f_int[25][4] ), .ZN(n7357) );
  INV_X1 U8553 ( .A(n7357), .ZN(n9241) );
  AOI21_X1 U8554 ( .B1(n7443), .B2(n7359), .A(n7358), .ZN(n7437) );
  OAI21_X1 U8555 ( .B1(n7437), .B2(n7433), .A(n7434), .ZN(n7364) );
  INV_X1 U8556 ( .A(n7360), .ZN(n7362) );
  NAND2_X1 U8557 ( .A1(n7362), .A2(n7361), .ZN(n7363) );
  XNOR2_X1 U8558 ( .A(n7364), .B(n7363), .ZN(n7365) );
  AOI22_X1 U8559 ( .A1(n7959), .A2(\adder_stage1[15][7] ), .B1(n7450), .B2(
        n7365), .ZN(n7366) );
  INV_X1 U8560 ( .A(n7366), .ZN(n9911) );
  NAND2_X1 U8561 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  XNOR2_X1 U8562 ( .A(n7394), .B(n7369), .ZN(n7370) );
  AOI22_X1 U8563 ( .A1(n7959), .A2(\adder_stage1[15][8] ), .B1(n7450), .B2(
        n7370), .ZN(n7371) );
  INV_X1 U8564 ( .A(n7371), .ZN(n9910) );
  NAND2_X1 U8565 ( .A1(n7373), .A2(n7372), .ZN(n7374) );
  XNOR2_X1 U8566 ( .A(n7425), .B(n7374), .ZN(n7375) );
  AOI22_X1 U8567 ( .A1(n8057), .A2(\adder_stage1[13][8] ), .B1(n7450), .B2(
        n7375), .ZN(n7376) );
  INV_X1 U8568 ( .A(n7376), .ZN(n9944) );
  AOI21_X1 U8569 ( .B1(n7379), .B2(n7378), .A(n7377), .ZN(n7391) );
  OAI21_X1 U8570 ( .B1(n7391), .B2(n7387), .A(n7388), .ZN(n7384) );
  INV_X1 U8571 ( .A(n7380), .ZN(n7382) );
  NAND2_X1 U8572 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  XNOR2_X1 U8573 ( .A(n7384), .B(n7383), .ZN(n7385) );
  AOI22_X1 U8574 ( .A1(n6854), .A2(\adder_stage1[13][7] ), .B1(n7450), .B2(
        n7385), .ZN(n7386) );
  INV_X1 U8575 ( .A(n7386), .ZN(n9945) );
  INV_X1 U8576 ( .A(n7387), .ZN(n7389) );
  NAND2_X1 U8577 ( .A1(n7389), .A2(n7388), .ZN(n7390) );
  XOR2_X1 U8578 ( .A(n7391), .B(n7390), .Z(n7392) );
  AOI22_X1 U8579 ( .A1(n8057), .A2(\adder_stage1[13][6] ), .B1(n7450), .B2(
        n7392), .ZN(n7393) );
  INV_X1 U8580 ( .A(n7393), .ZN(n9946) );
  NAND2_X1 U8581 ( .A1(n7395), .A2(n7394), .ZN(n7397) );
  NAND2_X1 U8582 ( .A1(n7397), .A2(n7396), .ZN(n7401) );
  NAND2_X1 U8583 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  XNOR2_X1 U8584 ( .A(n7401), .B(n7400), .ZN(n7402) );
  AOI22_X1 U8585 ( .A1(n7959), .A2(\adder_stage1[15][10] ), .B1(n7450), .B2(
        n7402), .ZN(n7403) );
  INV_X1 U8586 ( .A(n7403), .ZN(n9908) );
  INV_X1 U8587 ( .A(n7404), .ZN(n7948) );
  INV_X1 U8588 ( .A(n7947), .ZN(n7405) );
  AOI21_X1 U8589 ( .B1(n7950), .B2(n7948), .A(n7405), .ZN(n7410) );
  INV_X1 U8590 ( .A(n7406), .ZN(n7408) );
  NAND2_X1 U8591 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  XOR2_X1 U8592 ( .A(n7410), .B(n7409), .Z(n7411) );
  AOI22_X1 U8593 ( .A1(n7952), .A2(\adder_stage1[14][5] ), .B1(n7450), .B2(
        n7411), .ZN(n7412) );
  INV_X1 U8594 ( .A(n7412), .ZN(n9930) );
  NAND2_X1 U8595 ( .A1(n7425), .A2(n7413), .ZN(n7414) );
  NAND2_X1 U8596 ( .A1(n7414), .A2(n7423), .ZN(n7417) );
  NAND2_X1 U8597 ( .A1(n7415), .A2(n7421), .ZN(n7416) );
  XNOR2_X1 U8598 ( .A(n7417), .B(n7416), .ZN(n7418) );
  AOI22_X1 U8599 ( .A1(n7525), .A2(\adder_stage1[13][10] ), .B1(n7971), .B2(
        n7418), .ZN(n7419) );
  INV_X1 U8600 ( .A(n7419), .ZN(n9942) );
  INV_X1 U8601 ( .A(n7420), .ZN(n7426) );
  OAI21_X1 U8602 ( .B1(n7423), .B2(n7422), .A(n7421), .ZN(n7424) );
  AOI21_X1 U8603 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n7430) );
  NAND2_X1 U8604 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  XOR2_X1 U8605 ( .A(n7430), .B(n7429), .Z(n7431) );
  AOI22_X1 U8606 ( .A1(n6273), .A2(\adder_stage1[13][11] ), .B1(n8087), .B2(
        n7431), .ZN(n7432) );
  INV_X1 U8607 ( .A(n7432), .ZN(n9941) );
  INV_X1 U8608 ( .A(n7433), .ZN(n7435) );
  NAND2_X1 U8609 ( .A1(n7435), .A2(n7434), .ZN(n7436) );
  XOR2_X1 U8610 ( .A(n7437), .B(n7436), .Z(n7438) );
  AOI22_X1 U8611 ( .A1(n7959), .A2(\adder_stage1[15][6] ), .B1(n7450), .B2(
        n7438), .ZN(n7439) );
  INV_X1 U8612 ( .A(n7439), .ZN(n9912) );
  INV_X1 U8613 ( .A(n7440), .ZN(n7441) );
  AOI21_X1 U8614 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n7448) );
  INV_X1 U8615 ( .A(n7444), .ZN(n7446) );
  NAND2_X1 U8616 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  XOR2_X1 U8617 ( .A(n7448), .B(n7447), .Z(n7449) );
  AOI22_X1 U8618 ( .A1(n7928), .A2(\adder_stage1[15][5] ), .B1(n7450), .B2(
        n7449), .ZN(n7451) );
  INV_X1 U8619 ( .A(n7451), .ZN(n9913) );
  AOI21_X1 U8620 ( .B1(n3435), .B2(n7454), .A(n7453), .ZN(n7458) );
  NAND2_X1 U8621 ( .A1(n7456), .A2(n7455), .ZN(n7457) );
  XOR2_X1 U8622 ( .A(n7458), .B(n7457), .Z(n7459) );
  AOI22_X1 U8623 ( .A1(n8118), .A2(\adder_stage1[12][9] ), .B1(n8175), .B2(
        n7459), .ZN(n7460) );
  INV_X1 U8624 ( .A(n7460), .ZN(n9960) );
  NAND2_X1 U8625 ( .A1(n3435), .A2(n7461), .ZN(n7463) );
  NAND2_X1 U8626 ( .A1(n7463), .A2(n7462), .ZN(n7467) );
  NAND2_X1 U8627 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  XNOR2_X1 U8628 ( .A(n7467), .B(n7466), .ZN(n7468) );
  AOI22_X1 U8629 ( .A1(n7074), .A2(\adder_stage1[12][10] ), .B1(n8175), .B2(
        n7468), .ZN(n7469) );
  INV_X1 U8630 ( .A(n7469), .ZN(n9959) );
  OAI21_X1 U8631 ( .B1(n7472), .B2(n7471), .A(n7470), .ZN(n8270) );
  OR2_X1 U8632 ( .A1(\adder_stage3[0][16] ), .A2(\adder_stage3[1][16] ), .ZN(
        n8268) );
  NAND2_X1 U8633 ( .A1(\adder_stage3[0][16] ), .A2(\adder_stage3[1][16] ), 
        .ZN(n8267) );
  INV_X1 U8634 ( .A(n8267), .ZN(n7480) );
  AOI21_X1 U8635 ( .B1(n8270), .B2(n8268), .A(n7480), .ZN(n7474) );
  OR2_X1 U8636 ( .A1(\adder_stage3[0][17] ), .A2(\adder_stage3[1][17] ), .ZN(
        n7479) );
  NAND2_X1 U8637 ( .A1(\adder_stage3[0][17] ), .A2(\adder_stage3[1][17] ), 
        .ZN(n7477) );
  NAND2_X1 U8638 ( .A1(n7479), .A2(n7477), .ZN(n7473) );
  XOR2_X1 U8639 ( .A(n7474), .B(n7473), .Z(n7475) );
  AOI22_X1 U8640 ( .A1(n7475), .A2(n8301), .B1(n8313), .B2(
        \adder_stage4[0][17] ), .ZN(n7476) );
  INV_X1 U8641 ( .A(n7476), .ZN(n9670) );
  AND2_X1 U8642 ( .A1(n8268), .A2(n7479), .ZN(n7486) );
  OR2_X1 U8643 ( .A1(\adder_stage3[0][18] ), .A2(\adder_stage3[1][18] ), .ZN(
        n7490) );
  AND2_X1 U8644 ( .A1(n7486), .A2(n7490), .ZN(n7679) );
  INV_X1 U8645 ( .A(n7477), .ZN(n7478) );
  AOI21_X1 U8646 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7487) );
  INV_X1 U8647 ( .A(n7490), .ZN(n7481) );
  NAND2_X1 U8648 ( .A1(\adder_stage3[0][18] ), .A2(\adder_stage3[1][18] ), 
        .ZN(n7489) );
  OAI21_X1 U8649 ( .B1(n7487), .B2(n7481), .A(n7489), .ZN(n7684) );
  AOI21_X1 U8650 ( .B1(n8270), .B2(n7679), .A(n7684), .ZN(n7483) );
  OR2_X1 U8651 ( .A1(\adder_stage3[0][19] ), .A2(\adder_stage3[1][19] ), .ZN(
        n7683) );
  NAND2_X1 U8652 ( .A1(\adder_stage3[0][19] ), .A2(\adder_stage3[1][19] ), 
        .ZN(n7681) );
  NAND2_X1 U8653 ( .A1(n7683), .A2(n7681), .ZN(n7482) );
  XOR2_X1 U8654 ( .A(n7483), .B(n7482), .Z(n7484) );
  AOI22_X1 U8655 ( .A1(n7484), .A2(n7507), .B1(n8313), .B2(
        \adder_stage4[0][19] ), .ZN(n7485) );
  INV_X1 U8656 ( .A(n7485), .ZN(n9668) );
  NAND2_X1 U8657 ( .A1(n8270), .A2(n7486), .ZN(n7488) );
  NAND2_X1 U8658 ( .A1(n7488), .A2(n7487), .ZN(n7492) );
  NAND2_X1 U8659 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  XNOR2_X1 U8660 ( .A(n7492), .B(n7491), .ZN(n7493) );
  AOI22_X1 U8661 ( .A1(n7493), .A2(n8314), .B1(n8313), .B2(
        \adder_stage4[0][18] ), .ZN(n7494) );
  INV_X1 U8662 ( .A(n7494), .ZN(n9669) );
  AOI22_X1 U8663 ( .A1(\x_mult_f_int[19][9] ), .A2(n7962), .B1(n8330), .B2(
        \x_mult_f[19][9] ), .ZN(n7495) );
  INV_X1 U8664 ( .A(n7495), .ZN(n9160) );
  AOI22_X1 U8665 ( .A1(\x_mult_f_int[19][8] ), .A2(n7627), .B1(n8325), .B2(
        \x_mult_f[19][8] ), .ZN(n7496) );
  INV_X1 U8666 ( .A(n7496), .ZN(n9161) );
  AOI22_X1 U8667 ( .A1(\x_mult_f_int[28][13] ), .A2(n6609), .B1(n8434), .B2(
        \x_mult_f[28][13] ), .ZN(n7497) );
  INV_X1 U8668 ( .A(n7497), .ZN(n9274) );
  AOI22_X1 U8669 ( .A1(\x_mult_f_int[28][12] ), .A2(n6636), .B1(n7855), .B2(
        \x_mult_f[28][12] ), .ZN(n7498) );
  INV_X1 U8670 ( .A(n7498), .ZN(n9275) );
  AOI22_X1 U8671 ( .A1(\x_mult_f_int[28][11] ), .A2(n6636), .B1(n7622), .B2(
        \x_mult_f[28][11] ), .ZN(n7499) );
  INV_X1 U8672 ( .A(n7499), .ZN(n9276) );
  FA_X1 U8673 ( .A(\x_mult_f[18][14] ), .B(\x_mult_f[19][14] ), .CI(n7500), 
        .CO(n7696), .S(n5719) );
  INV_X1 U8674 ( .A(n7501), .ZN(n7502) );
  AOI22_X1 U8675 ( .A1(n7502), .A2(n4444), .B1(n7698), .B2(
        \adder_stage1[9][20] ), .ZN(n7503) );
  INV_X1 U8676 ( .A(n7503), .ZN(n10003) );
  AOI22_X1 U8677 ( .A1(n8309), .A2(\x_mult_f[16][4] ), .B1(n7507), .B2(
        \x_mult_f_int[16][4] ), .ZN(n7504) );
  INV_X1 U8678 ( .A(n7504), .ZN(n9127) );
  AOI22_X1 U8679 ( .A1(n7622), .A2(\x_mult_f[16][3] ), .B1(n7507), .B2(
        \x_mult_f_int[16][3] ), .ZN(n7505) );
  INV_X1 U8680 ( .A(n7505), .ZN(n9128) );
  AOI22_X1 U8681 ( .A1(n8176), .A2(\x_mult_f[16][5] ), .B1(n7507), .B2(
        \x_mult_f_int[16][5] ), .ZN(n7506) );
  INV_X1 U8682 ( .A(n7506), .ZN(n9126) );
  AOI22_X1 U8683 ( .A1(n8273), .A2(\x_mult_f[16][2] ), .B1(n7507), .B2(
        \x_mult_f_int[16][2] ), .ZN(n7508) );
  INV_X1 U8684 ( .A(n7508), .ZN(n9129) );
  INV_X1 U8685 ( .A(n7509), .ZN(n7511) );
  NAND2_X1 U8686 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  XOR2_X1 U8687 ( .A(n7513), .B(n7512), .Z(n7514) );
  AOI22_X1 U8688 ( .A1(n7640), .A2(\adder_stage3[0][8] ), .B1(n8235), .B2(
        n7514), .ZN(n7515) );
  INV_X1 U8689 ( .A(n7515), .ZN(n9761) );
  AOI21_X1 U8690 ( .B1(n8228), .B2(n7517), .A(n7516), .ZN(n7531) );
  OAI21_X1 U8691 ( .B1(n7531), .B2(n7527), .A(n7528), .ZN(n7522) );
  INV_X1 U8692 ( .A(n7518), .ZN(n7520) );
  NAND2_X1 U8693 ( .A1(n7520), .A2(n7519), .ZN(n7521) );
  XNOR2_X1 U8694 ( .A(n7522), .B(n7521), .ZN(n7523) );
  AOI22_X1 U8695 ( .A1(n7640), .A2(\adder_stage3[0][7] ), .B1(n8235), .B2(
        n7523), .ZN(n7524) );
  INV_X1 U8696 ( .A(n7524), .ZN(n9762) );
  AOI22_X1 U8697 ( .A1(n7525), .A2(\x_mult_f[10][1] ), .B1(n7570), .B2(
        \x_mult_f_int[10][1] ), .ZN(n7526) );
  INV_X1 U8698 ( .A(n7526), .ZN(n9346) );
  INV_X1 U8699 ( .A(n7527), .ZN(n7529) );
  NAND2_X1 U8700 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  XOR2_X1 U8701 ( .A(n7531), .B(n7530), .Z(n7532) );
  AOI22_X1 U8702 ( .A1(n7640), .A2(\adder_stage3[0][6] ), .B1(n8235), .B2(
        n7532), .ZN(n7533) );
  INV_X1 U8703 ( .A(n7533), .ZN(n9763) );
  INV_X1 U8704 ( .A(n7534), .ZN(n7546) );
  OAI21_X1 U8705 ( .B1(n7546), .B2(n7542), .A(n7543), .ZN(n7539) );
  INV_X1 U8706 ( .A(n7535), .ZN(n7537) );
  NAND2_X1 U8707 ( .A1(n7537), .A2(n7536), .ZN(n7538) );
  XNOR2_X1 U8708 ( .A(n7539), .B(n7538), .ZN(n7540) );
  AOI22_X1 U8709 ( .A1(n7622), .A2(\adder_stage1[4][3] ), .B1(n7570), .B2(
        n7540), .ZN(n7541) );
  INV_X1 U8710 ( .A(n7541), .ZN(n10100) );
  INV_X1 U8711 ( .A(n7542), .ZN(n7544) );
  NAND2_X1 U8712 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  XOR2_X1 U8713 ( .A(n7546), .B(n7545), .Z(n7547) );
  AOI22_X1 U8714 ( .A1(n7622), .A2(\adder_stage1[4][2] ), .B1(n7570), .B2(
        n7547), .ZN(n7548) );
  INV_X1 U8715 ( .A(n7548), .ZN(n10101) );
  INV_X1 U8716 ( .A(n7549), .ZN(n7551) );
  NAND2_X1 U8717 ( .A1(n7551), .A2(n7550), .ZN(n7553) );
  XOR2_X1 U8718 ( .A(n7553), .B(n7552), .Z(n7554) );
  AOI22_X1 U8719 ( .A1(n7622), .A2(\adder_stage1[4][1] ), .B1(n7570), .B2(
        n7554), .ZN(n7555) );
  INV_X1 U8720 ( .A(n7555), .ZN(n10102) );
  AOI22_X1 U8721 ( .A1(n7556), .A2(\x_mult_f[10][3] ), .B1(n7570), .B2(
        \x_mult_f_int[10][3] ), .ZN(n7557) );
  INV_X1 U8722 ( .A(n7557), .ZN(n9052) );
  AOI22_X1 U8723 ( .A1(n8330), .A2(\x_mult_f[8][3] ), .B1(n8235), .B2(
        \x_mult_f_int[8][3] ), .ZN(n7558) );
  INV_X1 U8724 ( .A(n7558), .ZN(n9024) );
  AOI22_X1 U8725 ( .A1(n8273), .A2(\x_mult_f[8][5] ), .B1(n8235), .B2(
        \x_mult_f_int[8][5] ), .ZN(n7559) );
  INV_X1 U8726 ( .A(n7559), .ZN(n9022) );
  AOI22_X1 U8727 ( .A1(n8088), .A2(\x_mult_f[8][4] ), .B1(n8235), .B2(
        \x_mult_f_int[8][4] ), .ZN(n7560) );
  INV_X1 U8728 ( .A(n7560), .ZN(n9023) );
  AOI22_X1 U8729 ( .A1(n7972), .A2(\x_mult_f[8][2] ), .B1(n8235), .B2(
        \x_mult_f_int[8][2] ), .ZN(n7561) );
  INV_X1 U8730 ( .A(n7561), .ZN(n9025) );
  AOI22_X1 U8731 ( .A1(n8398), .A2(\x_mult_f[10][5] ), .B1(n7570), .B2(
        \x_mult_f_int[10][5] ), .ZN(n7562) );
  INV_X1 U8732 ( .A(n7562), .ZN(n9050) );
  OAI21_X1 U8733 ( .B1(n7565), .B2(n7564), .A(n7563), .ZN(n8218) );
  OR2_X1 U8734 ( .A1(\adder_stage1[14][14] ), .A2(\adder_stage1[15][14] ), 
        .ZN(n8220) );
  NAND2_X1 U8735 ( .A1(\adder_stage1[14][14] ), .A2(\adder_stage1[15][14] ), 
        .ZN(n8219) );
  INV_X1 U8736 ( .A(n8219), .ZN(n7566) );
  XOR2_X1 U8737 ( .A(\adder_stage1[15][15] ), .B(\adder_stage1[14][15] ), .Z(
        n7567) );
  AOI22_X1 U8738 ( .A1(n7568), .A2(n8281), .B1(n8338), .B2(
        \adder_stage2[7][15] ), .ZN(n7569) );
  INV_X1 U8739 ( .A(n7569), .ZN(n9771) );
  AOI22_X1 U8740 ( .A1(n8401), .A2(\x_mult_f[10][2] ), .B1(n7570), .B2(
        \x_mult_f_int[10][2] ), .ZN(n7571) );
  INV_X1 U8741 ( .A(n7571), .ZN(n9053) );
  OAI21_X1 U8742 ( .B1(n7663), .B2(n7573), .A(n7572), .ZN(n7577) );
  NAND2_X1 U8743 ( .A1(n7575), .A2(n7574), .ZN(n7576) );
  XNOR2_X1 U8744 ( .A(n7577), .B(n7576), .ZN(n7578) );
  AOI22_X1 U8745 ( .A1(n7669), .A2(\adder_stage2[6][14] ), .B1(n8167), .B2(
        n7578), .ZN(n7579) );
  INV_X1 U8746 ( .A(n7579), .ZN(n9789) );
  AOI22_X1 U8747 ( .A1(\x_mult_f_int[30][11] ), .A2(n6875), .B1(n8296), .B2(
        \x_mult_f[30][11] ), .ZN(n7580) );
  INV_X1 U8748 ( .A(n7580), .ZN(n9304) );
  AOI22_X1 U8749 ( .A1(\x_mult_f_int[30][10] ), .A2(n8087), .B1(n7614), .B2(
        \x_mult_f[30][10] ), .ZN(n7581) );
  INV_X1 U8750 ( .A(n7581), .ZN(n9305) );
  AOI22_X1 U8751 ( .A1(\x_mult_f_int[14][7] ), .A2(n7862), .B1(n8313), .B2(
        \x_mult_f[14][7] ), .ZN(n7582) );
  INV_X1 U8752 ( .A(n7582), .ZN(n9103) );
  AOI22_X1 U8753 ( .A1(\x_mult_f_int[14][8] ), .A2(n7862), .B1(n8409), .B2(
        \x_mult_f[14][8] ), .ZN(n7583) );
  INV_X1 U8754 ( .A(n7583), .ZN(n9102) );
  AOI22_X1 U8755 ( .A1(\x_mult_f_int[14][6] ), .A2(n6279), .B1(n8427), .B2(
        \x_mult_f[14][6] ), .ZN(n7584) );
  INV_X1 U8756 ( .A(n7584), .ZN(n9104) );
  AOI22_X1 U8757 ( .A1(\x_mult_f_int[9][10] ), .A2(n7862), .B1(n7698), .B2(
        \x_mult_f[9][10] ), .ZN(n7585) );
  INV_X1 U8758 ( .A(n7585), .ZN(n9031) );
  AOI22_X1 U8759 ( .A1(\x_mult_f_int[9][11] ), .A2(n8311), .B1(n7698), .B2(
        \x_mult_f[9][11] ), .ZN(n7586) );
  INV_X1 U8760 ( .A(n7586), .ZN(n9030) );
  AOI22_X1 U8761 ( .A1(\x_mult_f_int[9][9] ), .A2(n5981), .B1(n7698), .B2(
        \x_mult_f[9][9] ), .ZN(n7587) );
  INV_X1 U8762 ( .A(n7587), .ZN(n9032) );
  AOI22_X1 U8763 ( .A1(\x_mult_f_int[28][9] ), .A2(n6279), .B1(n8309), .B2(
        \x_mult_f[28][9] ), .ZN(n7588) );
  INV_X1 U8764 ( .A(n7588), .ZN(n9278) );
  AOI22_X1 U8765 ( .A1(\x_mult_f_int[28][10] ), .A2(n7962), .B1(n8434), .B2(
        \x_mult_f[28][10] ), .ZN(n7589) );
  INV_X1 U8766 ( .A(n7589), .ZN(n9277) );
  INV_X1 U8767 ( .A(n7590), .ZN(n7592) );
  NAND2_X1 U8768 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  XOR2_X1 U8769 ( .A(n7594), .B(n7593), .Z(n7595) );
  AOI22_X1 U8770 ( .A1(n7595), .A2(n7862), .B1(n8336), .B2(
        \adder_stage1[12][13] ), .ZN(n7596) );
  INV_X1 U8771 ( .A(n7596), .ZN(n9956) );
  INV_X1 U8772 ( .A(n7597), .ZN(n8159) );
  OAI21_X1 U8773 ( .B1(n8159), .B2(n8155), .A(n8156), .ZN(n7602) );
  INV_X1 U8774 ( .A(n7598), .ZN(n7600) );
  NAND2_X1 U8775 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  XNOR2_X1 U8776 ( .A(n7602), .B(n7601), .ZN(n7603) );
  AOI22_X1 U8777 ( .A1(n7614), .A2(\adder_stage1[10][3] ), .B1(n8292), .B2(
        n7603), .ZN(n8892) );
  INV_X1 U8778 ( .A(n7604), .ZN(n7605) );
  AOI21_X1 U8779 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n7612) );
  INV_X1 U8780 ( .A(n7608), .ZN(n7610) );
  NAND2_X1 U8781 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  XOR2_X1 U8782 ( .A(n7612), .B(n7611), .Z(n7613) );
  AOI22_X1 U8783 ( .A1(n7614), .A2(\adder_stage1[10][5] ), .B1(n8292), .B2(
        n7613), .ZN(n7615) );
  INV_X1 U8784 ( .A(n7615), .ZN(n9998) );
  INV_X1 U8785 ( .A(n7616), .ZN(n7618) );
  NAND2_X1 U8786 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  XOR2_X1 U8787 ( .A(n7620), .B(n7619), .Z(n7621) );
  AOI22_X1 U8788 ( .A1(n7622), .A2(\adder_stage2[6][2] ), .B1(n7627), .B2(
        n7621), .ZN(n7623) );
  INV_X1 U8789 ( .A(n7623), .ZN(n9801) );
  NAND2_X1 U8790 ( .A1(n7624), .A2(n7661), .ZN(n7625) );
  XOR2_X1 U8791 ( .A(n7663), .B(n7625), .Z(n7626) );
  AOI22_X1 U8792 ( .A1(n7669), .A2(\adder_stage2[6][11] ), .B1(n7627), .B2(
        n7626), .ZN(n7628) );
  INV_X1 U8793 ( .A(n7628), .ZN(n9792) );
  AOI22_X1 U8794 ( .A1(\x_mult_f_int[20][10] ), .A2(n8153), .B1(n8323), .B2(
        \x_mult_f[20][10] ), .ZN(n7629) );
  INV_X1 U8795 ( .A(n7629), .ZN(n9173) );
  AOI22_X1 U8796 ( .A1(\x_mult_f_int[20][13] ), .A2(n5981), .B1(n8323), .B2(
        \x_mult_f[20][13] ), .ZN(n7630) );
  INV_X1 U8797 ( .A(n7630), .ZN(n9170) );
  AOI22_X1 U8798 ( .A1(\x_mult_f_int[20][9] ), .A2(n7927), .B1(n8323), .B2(
        \x_mult_f[20][9] ), .ZN(n7631) );
  INV_X1 U8799 ( .A(n7631), .ZN(n9174) );
  AOI22_X1 U8800 ( .A1(\x_mult_f_int[20][12] ), .A2(n8294), .B1(n8323), .B2(
        \x_mult_f[20][12] ), .ZN(n7632) );
  INV_X1 U8801 ( .A(n7632), .ZN(n9171) );
  AOI22_X1 U8802 ( .A1(\x_mult_f_int[20][8] ), .A2(n6307), .B1(n8323), .B2(
        \x_mult_f[20][8] ), .ZN(n7633) );
  INV_X1 U8803 ( .A(n7633), .ZN(n9175) );
  AOI22_X1 U8804 ( .A1(\x_mult_f_int[20][11] ), .A2(n7627), .B1(n8323), .B2(
        \x_mult_f[20][11] ), .ZN(n7634) );
  INV_X1 U8805 ( .A(n7634), .ZN(n9172) );
  NAND2_X1 U8806 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  XNOR2_X1 U8807 ( .A(n7638), .B(n7637), .ZN(n7639) );
  AOI22_X1 U8808 ( .A1(n7640), .A2(\adder_stage3[0][10] ), .B1(n8298), .B2(
        n7639), .ZN(n7641) );
  INV_X1 U8809 ( .A(n7641), .ZN(n9759) );
  OAI21_X1 U8810 ( .B1(n7663), .B2(n7643), .A(n7642), .ZN(n7644) );
  INV_X1 U8811 ( .A(n7644), .ZN(n7648) );
  NAND2_X1 U8812 ( .A1(n7646), .A2(n7645), .ZN(n7647) );
  XOR2_X1 U8813 ( .A(n7648), .B(n7647), .Z(n7649) );
  AOI22_X1 U8814 ( .A1(n7669), .A2(\adder_stage2[6][13] ), .B1(n8105), .B2(
        n7649), .ZN(n7650) );
  INV_X1 U8815 ( .A(n7650), .ZN(n9790) );
  OAI21_X1 U8816 ( .B1(n7653), .B2(n7652), .A(n7651), .ZN(n7658) );
  INV_X1 U8817 ( .A(n7654), .ZN(n7656) );
  NAND2_X1 U8818 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  XNOR2_X1 U8819 ( .A(n7658), .B(n7657), .ZN(n7659) );
  AOI22_X1 U8820 ( .A1(n7669), .A2(\adder_stage2[6][10] ), .B1(n8105), .B2(
        n7659), .ZN(n7660) );
  INV_X1 U8821 ( .A(n7660), .ZN(n9793) );
  OAI21_X1 U8822 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7667) );
  NAND2_X1 U8823 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  XNOR2_X1 U8824 ( .A(n7667), .B(n7666), .ZN(n7668) );
  AOI22_X1 U8825 ( .A1(n7669), .A2(\adder_stage2[6][12] ), .B1(n8105), .B2(
        n7668), .ZN(n7670) );
  INV_X1 U8826 ( .A(n7670), .ZN(n9791) );
  FA_X1 U8827 ( .A(n3447), .B(n3466), .CI(n7671), .CO(n7672), .S(n3511) );
  INV_X1 U8828 ( .A(n7672), .ZN(n7673) );
  AOI22_X1 U8829 ( .A1(n7673), .A2(n8334), .B1(n7855), .B2(
        \adder_stage1[6][20] ), .ZN(n7674) );
  INV_X1 U8830 ( .A(n7674), .ZN(n10054) );
  FA_X1 U8831 ( .A(\adder_stage1[4][15] ), .B(\adder_stage1[5][15] ), .CI(
        n7675), .CO(n7990), .S(n5407) );
  NAND2_X1 U8832 ( .A1(n7676), .A2(n7819), .ZN(n7678) );
  NAND2_X1 U8833 ( .A1(n7928), .A2(\adder_stage2[2][16] ), .ZN(n7677) );
  NAND2_X1 U8834 ( .A1(n7678), .A2(n7677), .ZN(n9854) );
  AND2_X1 U8835 ( .A1(n7679), .A2(n7683), .ZN(n7680) );
  NAND2_X1 U8836 ( .A1(n8270), .A2(n7680), .ZN(n7686) );
  INV_X1 U8837 ( .A(n7681), .ZN(n7682) );
  AOI21_X1 U8838 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n7685) );
  NAND2_X1 U8839 ( .A1(n7686), .A2(n7685), .ZN(n7688) );
  XOR2_X1 U8840 ( .A(\adder_stage3[1][20] ), .B(\adder_stage3[0][20] ), .Z(
        n7687) );
  XOR2_X1 U8841 ( .A(n7688), .B(n7687), .Z(n7689) );
  NAND2_X1 U8842 ( .A1(n7689), .A2(n6875), .ZN(n7691) );
  NAND2_X1 U8843 ( .A1(n8313), .A2(\adder_stage4[0][20] ), .ZN(n7690) );
  NAND2_X1 U8844 ( .A1(n7691), .A2(n7690), .ZN(n9667) );
  FA_X1 U8845 ( .A(\x_mult_f[16][14] ), .B(\x_mult_f[17][14] ), .CI(n7692), 
        .CO(n8123), .S(n5229) );
  NAND2_X1 U8846 ( .A1(n7693), .A2(n8078), .ZN(n7695) );
  NAND2_X1 U8847 ( .A1(n8319), .A2(\adder_stage1[8][15] ), .ZN(n7694) );
  NAND2_X1 U8848 ( .A1(n7695), .A2(n7694), .ZN(n10021) );
  FA_X1 U8849 ( .A(n3461), .B(n8795), .CI(n7696), .CO(n7501), .S(n7697) );
  NAND2_X1 U8850 ( .A1(n7697), .A2(n7862), .ZN(n7700) );
  NAND2_X1 U8851 ( .A1(n7698), .A2(\adder_stage1[9][15] ), .ZN(n7699) );
  NAND2_X1 U8852 ( .A1(n7700), .A2(n7699), .ZN(n10004) );
  FA_X1 U8853 ( .A(n3462), .B(n8793), .CI(n7701), .CO(n4665), .S(n7703) );
  AND2_X1 U8854 ( .A1(n8313), .A2(\adder_stage1[5][15] ), .ZN(n7702) );
  AOI21_X1 U8855 ( .B1(n7703), .B2(n8314), .A(n7702), .ZN(n8863) );
  FA_X1 U8856 ( .A(\x_mult_f[28][14] ), .B(\x_mult_f[29][14] ), .CI(n7704), 
        .CO(n8034), .S(n6280) );
  NAND2_X1 U8857 ( .A1(n7705), .A2(n8235), .ZN(n7707) );
  NAND2_X1 U8858 ( .A1(n8434), .A2(\adder_stage1[14][15] ), .ZN(n7706) );
  NAND2_X1 U8859 ( .A1(n7707), .A2(n7706), .ZN(n9920) );
  AND2_X1 U8860 ( .A1(n7708), .A2(n7710), .ZN(n8062) );
  OR2_X1 U8861 ( .A1(\adder_stage3[2][19] ), .A2(\adder_stage3[3][19] ), .ZN(
        n8064) );
  AND2_X1 U8862 ( .A1(n8062), .A2(n8064), .ZN(n7709) );
  NAND2_X1 U8863 ( .A1(n8137), .A2(n7709), .ZN(n7716) );
  INV_X1 U8864 ( .A(n7710), .ZN(n7712) );
  OAI21_X1 U8865 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n8061) );
  NAND2_X1 U8866 ( .A1(\adder_stage3[2][19] ), .A2(\adder_stage3[3][19] ), 
        .ZN(n8063) );
  INV_X1 U8867 ( .A(n8063), .ZN(n7714) );
  AOI21_X1 U8868 ( .B1(n8061), .B2(n8064), .A(n7714), .ZN(n7715) );
  NAND2_X1 U8869 ( .A1(n7716), .A2(n7715), .ZN(n7718) );
  XOR2_X1 U8870 ( .A(\adder_stage3[3][20] ), .B(\adder_stage3[2][20] ), .Z(
        n7717) );
  XOR2_X1 U8871 ( .A(n7718), .B(n7717), .Z(n7719) );
  NAND2_X1 U8872 ( .A1(n7719), .A2(n4311), .ZN(n7721) );
  NAND2_X1 U8873 ( .A1(n8398), .A2(\adder_stage4[1][20] ), .ZN(n7720) );
  NAND2_X1 U8874 ( .A1(n7721), .A2(n7720), .ZN(n9646) );
  FA_X1 U8875 ( .A(\x_mult_f[2][14] ), .B(\x_mult_f[3][14] ), .CI(n7722), .CO(
        n7961), .S(n5517) );
  INV_X1 U8876 ( .A(n7723), .ZN(n7724) );
  NAND2_X1 U8877 ( .A1(n7724), .A2(n7962), .ZN(n7726) );
  NAND2_X1 U8878 ( .A1(n8319), .A2(\adder_stage1[1][20] ), .ZN(n7725) );
  NAND2_X1 U8879 ( .A1(n7726), .A2(n7725), .ZN(n10136) );
  FA_X1 U8880 ( .A(\x_mult_f[0][14] ), .B(\x_mult_f[1][14] ), .CI(n7727), .CO(
        n8026), .S(n6071) );
  NAND2_X1 U8881 ( .A1(n7728), .A2(n7627), .ZN(n7730) );
  NAND2_X1 U8882 ( .A1(n7928), .A2(\adder_stage1[0][15] ), .ZN(n7729) );
  NAND2_X1 U8883 ( .A1(n7730), .A2(n7729), .ZN(n10154) );
  FA_X1 U8884 ( .A(\x_mult_f[22][14] ), .B(\x_mult_f[23][14] ), .CI(n7731), 
        .CO(n8012), .S(n5160) );
  NAND2_X1 U8885 ( .A1(n7732), .A2(n8078), .ZN(n7734) );
  NAND2_X1 U8886 ( .A1(n7622), .A2(\adder_stage1[11][15] ), .ZN(n7733) );
  NAND2_X1 U8887 ( .A1(n7734), .A2(n7733), .ZN(n9971) );
  AND2_X1 U8888 ( .A1(n8248), .A2(n7738), .ZN(n8418) );
  NOR2_X1 U8889 ( .A1(\adder_stage2[2][18] ), .A2(\adder_stage2[3][18] ), .ZN(
        n7740) );
  INV_X1 U8890 ( .A(n7740), .ZN(n8423) );
  AND2_X1 U8891 ( .A1(n8418), .A2(n8423), .ZN(n8412) );
  OR2_X1 U8892 ( .A1(\adder_stage2[2][19] ), .A2(\adder_stage2[3][19] ), .ZN(
        n8414) );
  AND2_X1 U8893 ( .A1(n8412), .A2(n8414), .ZN(n7735) );
  NAND2_X1 U8894 ( .A1(n8419), .A2(n7735), .ZN(n7743) );
  INV_X1 U8895 ( .A(n7736), .ZN(n7737) );
  AOI21_X1 U8896 ( .B1(n7739), .B2(n7738), .A(n7737), .ZN(n8420) );
  NAND2_X1 U8897 ( .A1(\adder_stage2[2][18] ), .A2(\adder_stage2[3][18] ), 
        .ZN(n8422) );
  OAI21_X1 U8898 ( .B1(n8420), .B2(n7740), .A(n8422), .ZN(n8411) );
  NAND2_X1 U8899 ( .A1(\adder_stage2[2][19] ), .A2(\adder_stage2[3][19] ), 
        .ZN(n8413) );
  INV_X1 U8900 ( .A(n8413), .ZN(n7741) );
  AOI21_X1 U8901 ( .B1(n8411), .B2(n8414), .A(n7741), .ZN(n7742) );
  NAND2_X1 U8902 ( .A1(n7743), .A2(n7742), .ZN(n7745) );
  XOR2_X1 U8903 ( .A(\adder_stage2[3][20] ), .B(\adder_stage2[2][20] ), .Z(
        n7744) );
  XOR2_X1 U8904 ( .A(n7745), .B(n7744), .Z(n7746) );
  NAND2_X1 U8905 ( .A1(n7746), .A2(n7862), .ZN(n7748) );
  NAND2_X1 U8906 ( .A1(n7952), .A2(\adder_stage3[1][20] ), .ZN(n7747) );
  NAND2_X1 U8907 ( .A1(n7748), .A2(n7747), .ZN(n9730) );
  FA_X1 U8908 ( .A(\x_mult_f[8][14] ), .B(\x_mult_f[9][14] ), .CI(n7749), .CO(
        n7808), .S(n6058) );
  NAND2_X1 U8909 ( .A1(n7750), .A2(n6636), .ZN(n7752) );
  NAND2_X1 U8910 ( .A1(n7959), .A2(\adder_stage1[4][15] ), .ZN(n7751) );
  NAND2_X1 U8911 ( .A1(n7752), .A2(n7751), .ZN(n10088) );
  AND2_X1 U8912 ( .A1(n7753), .A2(n7757), .ZN(n7754) );
  NAND2_X1 U8913 ( .A1(n8263), .A2(n7754), .ZN(n7760) );
  INV_X1 U8914 ( .A(n7755), .ZN(n7756) );
  AOI21_X1 U8915 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7759) );
  NAND2_X1 U8916 ( .A1(n7760), .A2(n7759), .ZN(n7762) );
  XOR2_X1 U8917 ( .A(\adder_stage2[7][20] ), .B(\adder_stage2[6][20] ), .Z(
        n7761) );
  XOR2_X1 U8918 ( .A(n7762), .B(n7761), .Z(n7763) );
  NAND2_X1 U8919 ( .A1(n7763), .A2(n8281), .ZN(n7765) );
  NAND2_X1 U8920 ( .A1(n7525), .A2(\adder_stage3[3][20] ), .ZN(n7764) );
  NAND2_X1 U8921 ( .A1(n7765), .A2(n7764), .ZN(n9688) );
  FA_X1 U8922 ( .A(\x_mult_f[26][14] ), .B(\x_mult_f[27][14] ), .CI(n7766), 
        .CO(n7817), .S(n4860) );
  NAND2_X1 U8923 ( .A1(n7767), .A2(n7819), .ZN(n7769) );
  NAND2_X1 U8924 ( .A1(n6273), .A2(\adder_stage1[13][15] ), .ZN(n7768) );
  NAND2_X1 U8925 ( .A1(n7769), .A2(n7768), .ZN(n9937) );
  FA_X1 U8926 ( .A(\x_mult_f[14][14] ), .B(\x_mult_f[15][14] ), .CI(n7770), 
        .CO(n7853), .S(n6889) );
  NAND2_X1 U8927 ( .A1(n7771), .A2(n8294), .ZN(n7773) );
  NAND2_X1 U8928 ( .A1(n7855), .A2(\adder_stage1[7][15] ), .ZN(n7772) );
  NAND2_X1 U8929 ( .A1(n7773), .A2(n7772), .ZN(n10038) );
  FA_X1 U8930 ( .A(\adder_stage1[8][15] ), .B(\adder_stage1[9][15] ), .CI(
        n7774), .CO(n7796), .S(n5385) );
  NAND2_X1 U8931 ( .A1(n7775), .A2(n8314), .ZN(n7777) );
  NAND2_X1 U8932 ( .A1(n8309), .A2(\adder_stage2[4][16] ), .ZN(n7776) );
  NAND2_X1 U8933 ( .A1(n7777), .A2(n7776), .ZN(n9820) );
  FA_X1 U8934 ( .A(\x_mult_f[20][14] ), .B(\x_mult_f[21][14] ), .CI(n7778), 
        .CO(n7930), .S(n5155) );
  INV_X1 U8935 ( .A(n7779), .ZN(n7780) );
  NAND2_X1 U8936 ( .A1(n7780), .A2(n6307), .ZN(n7782) );
  NAND2_X1 U8937 ( .A1(n8328), .A2(\adder_stage1[10][20] ), .ZN(n7781) );
  NAND2_X1 U8938 ( .A1(n7782), .A2(n7781), .ZN(n9987) );
  AND2_X1 U8939 ( .A1(n7783), .A2(n7787), .ZN(n7784) );
  NAND2_X1 U8940 ( .A1(n8256), .A2(n7784), .ZN(n7790) );
  INV_X1 U8941 ( .A(n7785), .ZN(n7786) );
  AOI21_X1 U8942 ( .B1(n7788), .B2(n7787), .A(n7786), .ZN(n7789) );
  NAND2_X1 U8943 ( .A1(n7790), .A2(n7789), .ZN(n7792) );
  XOR2_X1 U8944 ( .A(\adder_stage2[5][20] ), .B(\adder_stage2[4][20] ), .Z(
        n7791) );
  XOR2_X1 U8945 ( .A(n7792), .B(n7791), .Z(n7793) );
  NAND2_X1 U8946 ( .A1(n7793), .A2(n8311), .ZN(n7795) );
  NAND2_X1 U8947 ( .A1(n8306), .A2(\adder_stage3[2][20] ), .ZN(n7794) );
  NAND2_X1 U8948 ( .A1(n7795), .A2(n7794), .ZN(n9709) );
  OR2_X1 U8949 ( .A1(n7978), .A2(n8846), .ZN(n7799) );
  FA_X1 U8950 ( .A(n3463), .B(n8803), .CI(n7796), .CO(n7797), .S(n7775) );
  INV_X1 U8951 ( .A(n7797), .ZN(n7798) );
  NAND2_X1 U8952 ( .A1(n7798), .A2(n6279), .ZN(n7980) );
  NAND2_X1 U8953 ( .A1(n7799), .A2(n7980), .ZN(n1972) );
  FA_X1 U8954 ( .A(\adder_stage1[6][15] ), .B(\adder_stage1[7][15] ), .CI(
        n7800), .CO(n7974), .S(n5436) );
  AOI22_X1 U8955 ( .A1(n7801), .A2(n8332), .B1(n8434), .B2(
        \adder_stage2[3][16] ), .ZN(n7802) );
  INV_X1 U8956 ( .A(n7802), .ZN(n9837) );
  OR2_X1 U8957 ( .A1(\x_mult_f[22][0] ), .A2(\x_mult_f[23][0] ), .ZN(n7804) );
  AND2_X1 U8958 ( .A1(n7804), .A2(n7803), .ZN(n7805) );
  AOI22_X1 U8959 ( .A1(n7556), .A2(\adder_stage1[11][0] ), .B1(n8265), .B2(
        n7805), .ZN(n7806) );
  INV_X1 U8960 ( .A(n7806), .ZN(n9986) );
  AOI22_X1 U8961 ( .A1(n7959), .A2(\x_mult_f[31][0] ), .B1(n8175), .B2(
        \x_mult_f_int[31][0] ), .ZN(n7807) );
  INV_X1 U8962 ( .A(n7807), .ZN(n9389) );
  FA_X1 U8963 ( .A(n8791), .B(n8792), .CI(n7808), .CO(n7809), .S(n7750) );
  INV_X1 U8964 ( .A(n7809), .ZN(n7810) );
  AOI22_X1 U8965 ( .A1(n7810), .A2(n4257), .B1(n8427), .B2(
        \adder_stage1[4][20] ), .ZN(n7811) );
  INV_X1 U8966 ( .A(n7811), .ZN(n10087) );
  AOI22_X1 U8967 ( .A1(n7815), .A2(n8294), .B1(n8434), .B2(
        \adder_stage2[7][16] ), .ZN(n7816) );
  INV_X1 U8968 ( .A(n7816), .ZN(n9770) );
  FA_X1 U8969 ( .A(n3448), .B(n3467), .CI(n7817), .CO(n7818), .S(n7767) );
  INV_X1 U8970 ( .A(n7818), .ZN(n7820) );
  AOI22_X1 U8971 ( .A1(n7820), .A2(n7819), .B1(n8434), .B2(
        \adder_stage1[13][20] ), .ZN(n7821) );
  INV_X1 U8972 ( .A(n7821), .ZN(n9936) );
  FA_X1 U8973 ( .A(\x_mult_f[6][14] ), .B(\x_mult_f[7][14] ), .CI(n7822), .CO(
        n8038), .S(n5469) );
  INV_X1 U8974 ( .A(n7823), .ZN(n7824) );
  AOI22_X1 U8975 ( .A1(n7824), .A2(n6875), .B1(n8296), .B2(
        \adder_stage1[3][20] ), .ZN(n7825) );
  INV_X1 U8976 ( .A(n7825), .ZN(n10104) );
  AOI22_X1 U8977 ( .A1(\x_mult_f_int[5][13] ), .A2(n7862), .B1(n8336), .B2(
        \x_mult_f[5][13] ), .ZN(n7826) );
  INV_X1 U8978 ( .A(n7826), .ZN(n8979) );
  AOI22_X1 U8979 ( .A1(\x_mult_f_int[14][14] ), .A2(n8334), .B1(n8336), .B2(
        \x_mult_f[14][14] ), .ZN(n7827) );
  INV_X1 U8980 ( .A(n7827), .ZN(n9096) );
  AOI22_X1 U8981 ( .A1(\x_mult_f_int[0][14] ), .A2(n8294), .B1(n8427), .B2(
        \x_mult_f[0][14] ), .ZN(n7828) );
  INV_X1 U8982 ( .A(n7828), .ZN(n8914) );
  AOI22_X1 U8983 ( .A1(\x_mult_f_int[30][13] ), .A2(n7962), .B1(n7669), .B2(
        \x_mult_f[30][13] ), .ZN(n7829) );
  INV_X1 U8984 ( .A(n7829), .ZN(n9302) );
  AOI22_X1 U8985 ( .A1(\x_mult_f_int[4][13] ), .A2(n7819), .B1(n8338), .B2(
        \x_mult_f[4][13] ), .ZN(n7830) );
  INV_X1 U8986 ( .A(n7830), .ZN(n8971) );
  AOI22_X1 U8987 ( .A1(\x_mult_f_int[0][12] ), .A2(n7627), .B1(n8409), .B2(
        \x_mult_f[0][12] ), .ZN(n7831) );
  INV_X1 U8988 ( .A(n7831), .ZN(n8916) );
  AOI22_X1 U8989 ( .A1(\x_mult_f_int[14][12] ), .A2(n8334), .B1(n8309), .B2(
        \x_mult_f[14][12] ), .ZN(n7832) );
  INV_X1 U8990 ( .A(n7832), .ZN(n9098) );
  AOI22_X1 U8991 ( .A1(\x_mult_f_int[0][13] ), .A2(n5175), .B1(n8336), .B2(
        \x_mult_f[0][13] ), .ZN(n7833) );
  INV_X1 U8992 ( .A(n7833), .ZN(n8915) );
  FA_X1 U8993 ( .A(n3449), .B(n3468), .CI(n7834), .CO(n7328), .S(n7835) );
  AOI22_X1 U8994 ( .A1(n7835), .A2(n7862), .B1(n8428), .B2(
        \adder_stage1[15][15] ), .ZN(n8854) );
  AOI22_X1 U8995 ( .A1(\x_mult_f_int[27][12] ), .A2(n7819), .B1(n8336), .B2(
        \x_mult_f[27][12] ), .ZN(n7836) );
  INV_X1 U8996 ( .A(n7836), .ZN(n9261) );
  AOI22_X1 U8997 ( .A1(\x_mult_f_int[27][13] ), .A2(n8281), .B1(n7864), .B2(
        \x_mult_f[27][13] ), .ZN(n7837) );
  INV_X1 U8998 ( .A(n7837), .ZN(n9260) );
  AOI22_X1 U8999 ( .A1(\x_mult_f_int[2][14] ), .A2(n7450), .B1(n7698), .B2(
        \x_mult_f[2][14] ), .ZN(n7838) );
  INV_X1 U9000 ( .A(n7838), .ZN(n8942) );
  AOI22_X1 U9001 ( .A1(\x_mult_f_int[4][12] ), .A2(n8314), .B1(n8338), .B2(
        \x_mult_f[4][12] ), .ZN(n7839) );
  INV_X1 U9002 ( .A(n7839), .ZN(n8972) );
  AOI22_X1 U9003 ( .A1(\x_mult_f_int[10][12] ), .A2(n8311), .B1(n8336), .B2(
        \x_mult_f[10][12] ), .ZN(n7840) );
  INV_X1 U9004 ( .A(n7840), .ZN(n9043) );
  AOI22_X1 U9005 ( .A1(\x_mult_f_int[14][13] ), .A2(n8334), .B1(n7698), .B2(
        \x_mult_f[14][13] ), .ZN(n7841) );
  INV_X1 U9006 ( .A(n7841), .ZN(n9097) );
  AOI22_X1 U9007 ( .A1(\x_mult_f_int[16][13] ), .A2(n8301), .B1(n8409), .B2(
        \x_mult_f[16][13] ), .ZN(n7842) );
  INV_X1 U9008 ( .A(n7842), .ZN(n9125) );
  AOI22_X1 U9009 ( .A1(\x_mult_f_int[26][12] ), .A2(n8117), .B1(n8401), .B2(
        \x_mult_f[26][12] ), .ZN(n7843) );
  INV_X1 U9010 ( .A(n7843), .ZN(n9247) );
  AOI22_X1 U9011 ( .A1(\x_mult_f_int[30][12] ), .A2(n7507), .B1(n8434), .B2(
        \x_mult_f[30][12] ), .ZN(n7844) );
  INV_X1 U9012 ( .A(n7844), .ZN(n9303) );
  AOI22_X1 U9013 ( .A1(\x_mult_f_int[23][12] ), .A2(n8216), .B1(n8330), .B2(
        \x_mult_f[23][12] ), .ZN(n7845) );
  INV_X1 U9014 ( .A(n7845), .ZN(n9213) );
  AOI22_X1 U9015 ( .A1(\x_mult_f_int[25][12] ), .A2(n8332), .B1(n8176), .B2(
        \x_mult_f[25][12] ), .ZN(n7846) );
  INV_X1 U9016 ( .A(n7846), .ZN(n9233) );
  AOI22_X1 U9017 ( .A1(\x_mult_f_int[22][12] ), .A2(n6636), .B1(n8328), .B2(
        \x_mult_f[22][12] ), .ZN(n7847) );
  INV_X1 U9018 ( .A(n7847), .ZN(n9199) );
  AOI22_X1 U9019 ( .A1(\x_mult_f_int[22][13] ), .A2(n6636), .B1(n8328), .B2(
        \x_mult_f[22][13] ), .ZN(n7848) );
  INV_X1 U9020 ( .A(n7848), .ZN(n9198) );
  AOI22_X1 U9021 ( .A1(\x_mult_f_int[19][12] ), .A2(n5175), .B1(n7855), .B2(
        \x_mult_f[19][12] ), .ZN(n7849) );
  INV_X1 U9022 ( .A(n7849), .ZN(n9157) );
  AOI22_X1 U9023 ( .A1(\x_mult_f_int[3][13] ), .A2(n8301), .B1(n8428), .B2(
        \x_mult_f[3][13] ), .ZN(n7850) );
  INV_X1 U9024 ( .A(n7850), .ZN(n8957) );
  AOI22_X1 U9025 ( .A1(\x_mult_f_int[28][14] ), .A2(n7819), .B1(n8338), .B2(
        \x_mult_f[28][14] ), .ZN(n7851) );
  INV_X1 U9026 ( .A(n7851), .ZN(n9273) );
  AOI22_X1 U9027 ( .A1(\x_mult_f_int[20][14] ), .A2(n8292), .B1(n8323), .B2(
        \x_mult_f[20][14] ), .ZN(n7852) );
  INV_X1 U9028 ( .A(n7852), .ZN(n9169) );
  FA_X1 U9029 ( .A(n3450), .B(n3469), .CI(n7853), .CO(n7854), .S(n7771) );
  INV_X1 U9030 ( .A(n7854), .ZN(n7856) );
  AOI22_X1 U9031 ( .A1(n7856), .A2(n8294), .B1(n7855), .B2(
        \adder_stage1[7][20] ), .ZN(n7857) );
  INV_X1 U9032 ( .A(n7857), .ZN(n10037) );
  AOI22_X1 U9033 ( .A1(\x_mult_f_int[6][13] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[6][13] ), .ZN(n7858) );
  INV_X1 U9034 ( .A(n7858), .ZN(n8986) );
  AOI22_X1 U9035 ( .A1(\x_mult_f_int[9][13] ), .A2(n5707), .B1(n8309), .B2(
        \x_mult_f[9][13] ), .ZN(n7859) );
  INV_X1 U9036 ( .A(n7859), .ZN(n9028) );
  AOI22_X1 U9037 ( .A1(\x_mult_f_int[10][14] ), .A2(n8311), .B1(n7864), .B2(
        \x_mult_f[10][14] ), .ZN(n7860) );
  INV_X1 U9038 ( .A(n7860), .ZN(n9041) );
  AOI22_X1 U9039 ( .A1(\x_mult_f_int[21][13] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][13] ), .ZN(n7861) );
  INV_X1 U9040 ( .A(n7861), .ZN(n9184) );
  AOI22_X1 U9041 ( .A1(\x_mult_f_int[24][13] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[24][13] ), .ZN(n8855) );
  AOI22_X1 U9042 ( .A1(\x_mult_f_int[29][12] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][12] ), .ZN(n7863) );
  INV_X1 U9043 ( .A(n7863), .ZN(n9289) );
  AOI22_X1 U9044 ( .A1(\x_mult_f_int[5][14] ), .A2(n7862), .B1(n7864), .B2(
        \x_mult_f[5][14] ), .ZN(n8856) );
  AOI22_X1 U9045 ( .A1(\x_mult_f_int[30][14] ), .A2(n6875), .B1(n8323), .B2(
        \x_mult_f[30][14] ), .ZN(n7865) );
  INV_X1 U9046 ( .A(n7865), .ZN(n9301) );
  AOI22_X1 U9047 ( .A1(\x_mult_f_int[1][14] ), .A2(n8298), .B1(n8398), .B2(
        \x_mult_f[1][14] ), .ZN(n7866) );
  INV_X1 U9048 ( .A(n7866), .ZN(n8928) );
  AOI22_X1 U9049 ( .A1(\x_mult_f_int[2][12] ), .A2(n8301), .B1(n8340), .B2(
        \x_mult_f[2][12] ), .ZN(n7867) );
  INV_X1 U9050 ( .A(n7867), .ZN(n8944) );
  AOI22_X1 U9051 ( .A1(\x_mult_f_int[1][13] ), .A2(n8298), .B1(n8401), .B2(
        \x_mult_f[1][13] ), .ZN(n7868) );
  INV_X1 U9052 ( .A(n7868), .ZN(n8929) );
  AOI22_X1 U9053 ( .A1(\x_mult_f_int[22][14] ), .A2(n6636), .B1(n8328), .B2(
        \x_mult_f[22][14] ), .ZN(n7869) );
  INV_X1 U9054 ( .A(n7869), .ZN(n9197) );
  AOI22_X1 U9055 ( .A1(\x_mult_f_int[3][14] ), .A2(n8301), .B1(n8428), .B2(
        \x_mult_f[3][14] ), .ZN(n7870) );
  INV_X1 U9056 ( .A(n7870), .ZN(n8956) );
  AOI22_X1 U9057 ( .A1(\x_mult_f_int[13][13] ), .A2(n7862), .B1(n8296), .B2(
        \x_mult_f[13][13] ), .ZN(n7871) );
  INV_X1 U9058 ( .A(n7871), .ZN(n9083) );
  AOI22_X1 U9059 ( .A1(\x_mult_f_int[11][13] ), .A2(n8314), .B1(n8323), .B2(
        \x_mult_f[11][13] ), .ZN(n7872) );
  INV_X1 U9060 ( .A(n7872), .ZN(n9055) );
  AOI22_X1 U9061 ( .A1(\x_mult_f_int[19][13] ), .A2(n5175), .B1(n8434), .B2(
        \x_mult_f[19][13] ), .ZN(n7873) );
  INV_X1 U9062 ( .A(n7873), .ZN(n9156) );
  AOI22_X1 U9063 ( .A1(\x_mult_f_int[7][14] ), .A2(n8216), .B1(n8306), .B2(
        \x_mult_f[7][14] ), .ZN(n7874) );
  INV_X1 U9064 ( .A(n7874), .ZN(n8999) );
  AOI22_X1 U9065 ( .A1(\x_mult_f_int[11][14] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][14] ), .ZN(n7875) );
  INV_X1 U9066 ( .A(n7875), .ZN(n9054) );
  AOI22_X1 U9067 ( .A1(\x_mult_f_int[18][14] ), .A2(n5175), .B1(n8319), .B2(
        \x_mult_f[18][14] ), .ZN(n7876) );
  INV_X1 U9068 ( .A(n7876), .ZN(n9141) );
  AOI22_X1 U9069 ( .A1(\x_mult_f_int[23][14] ), .A2(n8265), .B1(n8330), .B2(
        \x_mult_f[23][14] ), .ZN(n7877) );
  INV_X1 U9070 ( .A(n7877), .ZN(n9211) );
  AOI22_X1 U9071 ( .A1(\x_mult_f_int[12][13] ), .A2(n8311), .B1(n8434), .B2(
        \x_mult_f[12][13] ), .ZN(n7878) );
  INV_X1 U9072 ( .A(n7878), .ZN(n9069) );
  AOI22_X1 U9073 ( .A1(\x_mult_f_int[26][13] ), .A2(n6609), .B1(n8409), .B2(
        \x_mult_f[26][13] ), .ZN(n7879) );
  INV_X1 U9074 ( .A(n7879), .ZN(n9246) );
  AOI22_X1 U9075 ( .A1(\x_mult_f_int[15][13] ), .A2(n6279), .B1(n8434), .B2(
        \x_mult_f[15][13] ), .ZN(n7880) );
  INV_X1 U9076 ( .A(n7880), .ZN(n9111) );
  AOI22_X1 U9077 ( .A1(\x_mult_f_int[23][13] ), .A2(n8167), .B1(n8330), .B2(
        \x_mult_f[23][13] ), .ZN(n7881) );
  INV_X1 U9078 ( .A(n7881), .ZN(n9212) );
  AOI22_X1 U9079 ( .A1(\x_mult_f_int[6][14] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[6][14] ), .ZN(n7882) );
  INV_X1 U9080 ( .A(n7882), .ZN(n8985) );
  AOI22_X1 U9081 ( .A1(\x_mult_f_int[13][14] ), .A2(n7570), .B1(n8296), .B2(
        \x_mult_f[13][14] ), .ZN(n7883) );
  INV_X1 U9082 ( .A(n7883), .ZN(n9082) );
  FA_X1 U9083 ( .A(\adder_stage1[0][15] ), .B(\adder_stage1[1][15] ), .CI(
        n7884), .CO(n7985), .S(n7316) );
  AOI22_X1 U9084 ( .A1(n7885), .A2(n4840), .B1(n8306), .B2(
        \adder_stage2[0][16] ), .ZN(n7886) );
  INV_X1 U9085 ( .A(n7886), .ZN(n9888) );
  AOI22_X1 U9086 ( .A1(\x_mult_f_int[12][14] ), .A2(n4645), .B1(n8409), .B2(
        \x_mult_f[12][14] ), .ZN(n7887) );
  INV_X1 U9087 ( .A(n7887), .ZN(n9068) );
  AOI22_X1 U9088 ( .A1(\x_mult_f_int[19][14] ), .A2(n5175), .B1(n8427), .B2(
        \x_mult_f[19][14] ), .ZN(n7888) );
  INV_X1 U9089 ( .A(n7888), .ZN(n9155) );
  AOI22_X1 U9090 ( .A1(\x_mult_f_int[26][14] ), .A2(n8251), .B1(n8398), .B2(
        \x_mult_f[26][14] ), .ZN(n7889) );
  INV_X1 U9091 ( .A(n7889), .ZN(n9245) );
  AOI22_X1 U9092 ( .A1(\x_mult_f_int[2][13] ), .A2(n5707), .B1(n8340), .B2(
        \x_mult_f[2][13] ), .ZN(n7890) );
  INV_X1 U9093 ( .A(n7890), .ZN(n8943) );
  AOI22_X1 U9094 ( .A1(\x_mult_f_int[10][13] ), .A2(n8311), .B1(n8336), .B2(
        \x_mult_f[10][13] ), .ZN(n7891) );
  INV_X1 U9095 ( .A(n7891), .ZN(n9042) );
  AOI22_X1 U9096 ( .A1(\x_mult_f_int[25][13] ), .A2(n8332), .B1(n8434), .B2(
        \x_mult_f[25][13] ), .ZN(n7892) );
  INV_X1 U9097 ( .A(n7892), .ZN(n9232) );
  AOI22_X1 U9098 ( .A1(\x_mult_f_int[29][13] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][13] ), .ZN(n7893) );
  INV_X1 U9099 ( .A(n7893), .ZN(n9288) );
  AOI22_X1 U9100 ( .A1(\x_mult_f_int[16][12] ), .A2(n7819), .B1(n7928), .B2(
        \x_mult_f[16][12] ), .ZN(n8857) );
  AOI22_X1 U9101 ( .A1(\x_mult_f_int[24][12] ), .A2(n8167), .B1(n8427), .B2(
        \x_mult_f[24][12] ), .ZN(n7894) );
  INV_X1 U9102 ( .A(n7894), .ZN(n9224) );
  AOI22_X1 U9103 ( .A1(\x_mult_f_int[1][12] ), .A2(n8298), .B1(n8398), .B2(
        \x_mult_f[1][12] ), .ZN(n7895) );
  INV_X1 U9104 ( .A(n7895), .ZN(n8930) );
  AOI22_X1 U9105 ( .A1(\x_mult_f_int[5][12] ), .A2(n7862), .B1(n8401), .B2(
        \x_mult_f[5][12] ), .ZN(n8858) );
  AOI22_X1 U9106 ( .A1(\x_mult_f_int[9][12] ), .A2(n8301), .B1(n8309), .B2(
        \x_mult_f[9][12] ), .ZN(n7896) );
  INV_X1 U9107 ( .A(n7896), .ZN(n9029) );
  AOI22_X1 U9108 ( .A1(\x_mult_f_int[17][13] ), .A2(n8292), .B1(n7614), .B2(
        \x_mult_f[17][13] ), .ZN(n8859) );
  AOI22_X1 U9109 ( .A1(\x_mult_f_int[6][12] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[6][12] ), .ZN(n7897) );
  INV_X1 U9110 ( .A(n7897), .ZN(n8987) );
  AOI22_X1 U9111 ( .A1(\x_mult_f_int[13][12] ), .A2(n7155), .B1(n8328), .B2(
        \x_mult_f[13][12] ), .ZN(n7898) );
  INV_X1 U9112 ( .A(n7898), .ZN(n9084) );
  AOI22_X1 U9113 ( .A1(\x_mult_f_int[21][12] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][12] ), .ZN(n7899) );
  INV_X1 U9114 ( .A(n7899), .ZN(n9185) );
  AOI22_X1 U9115 ( .A1(\x_mult_f_int[4][14] ), .A2(n8117), .B1(n8338), .B2(
        \x_mult_f[4][14] ), .ZN(n7900) );
  INV_X1 U9116 ( .A(n7900), .ZN(n8970) );
  AOI22_X1 U9117 ( .A1(\x_mult_f_int[31][12] ), .A2(n8304), .B1(n8296), .B2(
        \x_mult_f[31][12] ), .ZN(n7901) );
  INV_X1 U9118 ( .A(n7901), .ZN(n9317) );
  FA_X1 U9119 ( .A(\adder_stage1[12][15] ), .B(\adder_stage1[13][15] ), .CI(
        n7902), .CO(n7981), .S(n6974) );
  AOI22_X1 U9120 ( .A1(n7903), .A2(n8311), .B1(n8338), .B2(
        \adder_stage2[6][16] ), .ZN(n7904) );
  INV_X1 U9121 ( .A(n7904), .ZN(n9787) );
  AOI22_X1 U9122 ( .A1(\x_mult_f_int[17][12] ), .A2(n6626), .B1(n7041), .B2(
        \x_mult_f[17][12] ), .ZN(n8860) );
  AOI22_X1 U9123 ( .A1(\x_mult_f_int[17][14] ), .A2(n6307), .B1(n7525), .B2(
        \x_mult_f[17][14] ), .ZN(n8861) );
  AOI22_X1 U9124 ( .A1(\x_mult_f_int[24][14] ), .A2(n8311), .B1(n8427), .B2(
        \x_mult_f[24][14] ), .ZN(n8862) );
  FA_X1 U9125 ( .A(\x_mult_f[12][14] ), .B(\x_mult_f[13][14] ), .CI(n7905), 
        .CO(n7671), .S(n7906) );
  AOI22_X1 U9126 ( .A1(n7906), .A2(n8334), .B1(n8319), .B2(
        \adder_stage1[6][14] ), .ZN(n7907) );
  INV_X1 U9127 ( .A(n7907), .ZN(n10056) );
  AOI22_X1 U9128 ( .A1(\x_mult_f_int[25][14] ), .A2(n8332), .B1(n8330), .B2(
        \x_mult_f[25][14] ), .ZN(n7908) );
  INV_X1 U9129 ( .A(n7908), .ZN(n9231) );
  AOI22_X1 U9130 ( .A1(\x_mult_f_int[15][14] ), .A2(n8235), .B1(n8309), .B2(
        \x_mult_f[15][14] ), .ZN(n7909) );
  INV_X1 U9131 ( .A(n7909), .ZN(n9110) );
  OAI21_X1 U9132 ( .B1(n7912), .B2(n7911), .A(n7910), .ZN(n7917) );
  INV_X1 U9133 ( .A(n7913), .ZN(n7915) );
  NAND2_X1 U9134 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  XNOR2_X1 U9135 ( .A(n7917), .B(n7916), .ZN(n7918) );
  AOI22_X1 U9136 ( .A1(n7920), .A2(\adder_stage1[9][12] ), .B1(n7919), .B2(
        n7918), .ZN(n7921) );
  INV_X1 U9137 ( .A(n7921), .ZN(n10007) );
  NAND2_X1 U9138 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  XNOR2_X1 U9139 ( .A(n3425), .B(n7924), .ZN(n7926) );
  AOI22_X1 U9140 ( .A1(n7928), .A2(\adder_stage1[14][12] ), .B1(n7927), .B2(
        n7926), .ZN(n7929) );
  INV_X1 U9141 ( .A(n7929), .ZN(n9923) );
  FA_X1 U9142 ( .A(n8796), .B(n3470), .CI(n7930), .CO(n7779), .S(n7931) );
  AOI22_X1 U9143 ( .A1(n7931), .A2(n6307), .B1(n8328), .B2(
        \adder_stage1[10][15] ), .ZN(n7932) );
  INV_X1 U9144 ( .A(n7932), .ZN(n9988) );
  INV_X1 U9145 ( .A(n7933), .ZN(n7939) );
  OAI21_X1 U9146 ( .B1(n7936), .B2(n7935), .A(n7934), .ZN(n7937) );
  AOI21_X1 U9147 ( .B1(n7939), .B2(n3419), .A(n7937), .ZN(n7943) );
  NAND2_X1 U9148 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  XOR2_X1 U9149 ( .A(n7943), .B(n7942), .Z(n7944) );
  AOI22_X1 U9150 ( .A1(n8057), .A2(\adder_stage1[1][11] ), .B1(n8054), .B2(
        n7944), .ZN(n7945) );
  INV_X1 U9151 ( .A(n7945), .ZN(n10141) );
  AOI22_X1 U9152 ( .A1(\x_mult_f_int[21][14] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][14] ), .ZN(n7946) );
  INV_X1 U9153 ( .A(n7946), .ZN(n9183) );
  NAND2_X1 U9154 ( .A1(n7948), .A2(n7947), .ZN(n7949) );
  XNOR2_X1 U9155 ( .A(n7950), .B(n7949), .ZN(n7951) );
  AOI22_X1 U9156 ( .A1(n7952), .A2(\adder_stage1[14][4] ), .B1(n8301), .B2(
        n7951), .ZN(n7953) );
  INV_X1 U9157 ( .A(n7953), .ZN(n9931) );
  NAND2_X1 U9158 ( .A1(n7955), .A2(n7954), .ZN(n7956) );
  XNOR2_X1 U9159 ( .A(n3411), .B(n7956), .ZN(n7958) );
  AOI22_X1 U9160 ( .A1(n7959), .A2(\adder_stage1[15][12] ), .B1(n8294), .B2(
        n7958), .ZN(n7960) );
  INV_X1 U9161 ( .A(n7960), .ZN(n9906) );
  FA_X1 U9162 ( .A(n8789), .B(n3471), .CI(n7961), .CO(n7723), .S(n7963) );
  AOI22_X1 U9163 ( .A1(n7963), .A2(n7962), .B1(n8428), .B2(
        \adder_stage1[1][15] ), .ZN(n7964) );
  INV_X1 U9164 ( .A(n7964), .ZN(n10137) );
  AOI22_X1 U9165 ( .A1(\x_mult_f_int[31][13] ), .A2(n8265), .B1(n8434), .B2(
        \x_mult_f[31][13] ), .ZN(n7965) );
  INV_X1 U9166 ( .A(n7965), .ZN(n9316) );
  NAND2_X1 U9167 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  XNOR2_X1 U9168 ( .A(n7969), .B(n7968), .ZN(n7970) );
  AOI22_X1 U9169 ( .A1(n7972), .A2(\adder_stage1[2][12] ), .B1(n7971), .B2(
        n7970), .ZN(n7973) );
  INV_X1 U9170 ( .A(n7973), .ZN(n10123) );
  FA_X1 U9171 ( .A(n3451), .B(n3472), .CI(n7974), .CO(n7975), .S(n7801) );
  INV_X1 U9172 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U9173 ( .A1(n7976), .A2(n6279), .ZN(n7977) );
  OAI21_X1 U9174 ( .B1(n7978), .B2(n8850), .A(n7977), .ZN(n1993) );
  OAI21_X1 U9175 ( .B1(n7978), .B2(n8816), .A(n7977), .ZN(n1996) );
  OAI21_X1 U9176 ( .B1(n7978), .B2(n8817), .A(n7977), .ZN(n1995) );
  OAI21_X1 U9177 ( .B1(n7978), .B2(n8818), .A(n7977), .ZN(n1994) );
  OAI21_X1 U9178 ( .B1(n8000), .B2(n8828), .A(n7980), .ZN(n1975) );
  OAI21_X1 U9179 ( .B1(n8000), .B2(n8829), .A(n7980), .ZN(n1974) );
  OAI21_X1 U9180 ( .B1(n7978), .B2(n8830), .A(n7980), .ZN(n1973) );
  FA_X1 U9181 ( .A(n3452), .B(n3473), .CI(n7981), .CO(n7982), .S(n7903) );
  INV_X1 U9182 ( .A(n7982), .ZN(n7983) );
  NAND2_X1 U9183 ( .A1(n7983), .A2(n6279), .ZN(n7984) );
  OAI21_X1 U9184 ( .B1(n8000), .B2(n8847), .A(n7984), .ZN(n1930) );
  OAI21_X1 U9185 ( .B1(n7978), .B2(n8831), .A(n7984), .ZN(n1933) );
  OAI21_X1 U9186 ( .B1(n8000), .B2(n8832), .A(n7984), .ZN(n1932) );
  OAI21_X1 U9187 ( .B1(n7978), .B2(n8833), .A(n7984), .ZN(n1931) );
  FA_X1 U9188 ( .A(n8799), .B(n3481), .CI(n7985), .CO(n7986), .S(n7885) );
  INV_X1 U9189 ( .A(n7986), .ZN(n7987) );
  NAND2_X1 U9190 ( .A1(n7987), .A2(n6279), .ZN(n7988) );
  OAI21_X1 U9191 ( .B1(n7978), .B2(n8834), .A(n7988), .ZN(n2059) );
  OAI21_X1 U9192 ( .B1(n8000), .B2(n8835), .A(n7988), .ZN(n2058) );
  OAI21_X1 U9193 ( .B1(n7978), .B2(n8836), .A(n7988), .ZN(n2057) );
  OAI21_X1 U9194 ( .B1(n8000), .B2(n8848), .A(n7988), .ZN(n2056) );
  FA_X1 U9195 ( .A(n8801), .B(n8802), .CI(n7990), .CO(n7991), .S(n7676) );
  INV_X1 U9196 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U9197 ( .A1(n7992), .A2(n6279), .ZN(n7993) );
  OAI21_X1 U9198 ( .B1(n7978), .B2(n8849), .A(n7993), .ZN(n2014) );
  OAI21_X1 U9199 ( .B1(n8000), .B2(n8837), .A(n7993), .ZN(n2017) );
  OAI21_X1 U9200 ( .B1(n7978), .B2(n8838), .A(n7993), .ZN(n2016) );
  OAI21_X1 U9201 ( .B1(n8000), .B2(n8839), .A(n7993), .ZN(n2015) );
  FA_X1 U9202 ( .A(\adder_stage1[10][15] ), .B(\adder_stage1[11][15] ), .CI(
        n7994), .CO(n8133), .S(n7161) );
  OAI211_X1 U9203 ( .C1(n7998), .C2(n7997), .A(n6279), .B(n7996), .ZN(n7995)
         );
  OAI21_X1 U9204 ( .B1(n8000), .B2(n8819), .A(n7995), .ZN(n1954) );
  OAI21_X1 U9205 ( .B1(n8000), .B2(n8820), .A(n7995), .ZN(n1953) );
  OAI211_X1 U9206 ( .C1(n7998), .C2(n7997), .A(n6279), .B(n7996), .ZN(n7999)
         );
  OAI21_X1 U9207 ( .B1(n8000), .B2(n8821), .A(n7999), .ZN(n1952) );
  OAI21_X1 U9208 ( .B1(n8000), .B2(n8851), .A(n7999), .ZN(n1951) );
  FA_X1 U9209 ( .A(n3453), .B(n3474), .CI(n8001), .CO(n8002), .S(n7815) );
  INV_X1 U9210 ( .A(n8002), .ZN(n8003) );
  NAND2_X1 U9211 ( .A1(n8003), .A2(n6279), .ZN(n8005) );
  OAI21_X1 U9212 ( .B1(n7978), .B2(n8852), .A(n8005), .ZN(n1909) );
  OAI21_X1 U9213 ( .B1(n8000), .B2(n8822), .A(n8005), .ZN(n1912) );
  OAI21_X1 U9214 ( .B1(n7978), .B2(n8823), .A(n8005), .ZN(n1911) );
  OAI21_X1 U9215 ( .B1(n8000), .B2(n8824), .A(n8005), .ZN(n1910) );
  INV_X1 U9216 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U9217 ( .A1(n8010), .A2(n6279), .ZN(n8011) );
  OAI21_X1 U9218 ( .B1(n8000), .B2(n8825), .A(n8011), .ZN(n2038) );
  OAI21_X1 U9219 ( .B1(n7978), .B2(n8826), .A(n8011), .ZN(n2037) );
  OAI21_X1 U9220 ( .B1(n7978), .B2(n8827), .A(n3442), .ZN(n2036) );
  OAI21_X1 U9221 ( .B1(n8000), .B2(n8853), .A(n3442), .ZN(n2035) );
  FA_X1 U9222 ( .A(n3454), .B(n3475), .CI(n8012), .CO(n8013), .S(n7732) );
  INV_X1 U9223 ( .A(n8013), .ZN(n8014) );
  AOI22_X1 U9224 ( .A1(n8014), .A2(n7627), .B1(n8309), .B2(
        \adder_stage1[11][20] ), .ZN(n8015) );
  INV_X1 U9225 ( .A(n8015), .ZN(n9970) );
  AOI21_X1 U9226 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8022) );
  NAND2_X1 U9227 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  XOR2_X1 U9228 ( .A(n8022), .B(n8021), .Z(n8023) );
  AOI22_X1 U9229 ( .A1(n7920), .A2(\adder_stage1[8][9] ), .B1(n8024), .B2(
        n8023), .ZN(n8025) );
  INV_X1 U9230 ( .A(n8025), .ZN(n10027) );
  FA_X1 U9231 ( .A(n8788), .B(n3476), .CI(n8026), .CO(n8027), .S(n7728) );
  INV_X1 U9232 ( .A(n8027), .ZN(n8028) );
  AOI22_X1 U9233 ( .A1(n8028), .A2(n7919), .B1(n8176), .B2(
        \adder_stage1[0][20] ), .ZN(n8029) );
  INV_X1 U9234 ( .A(n8029), .ZN(n10153) );
  FA_X1 U9235 ( .A(\x_mult_f[24][14] ), .B(\x_mult_f[25][14] ), .CI(n8030), 
        .CO(n8041), .S(n6457) );
  INV_X1 U9236 ( .A(n8031), .ZN(n8032) );
  AOI22_X1 U9237 ( .A1(n8032), .A2(n7862), .B1(n8336), .B2(
        \adder_stage1[12][20] ), .ZN(n8033) );
  INV_X1 U9238 ( .A(n8033), .ZN(n9953) );
  FA_X1 U9239 ( .A(n8798), .B(n3477), .CI(n8034), .CO(n8035), .S(n7705) );
  INV_X1 U9240 ( .A(n8035), .ZN(n8036) );
  AOI22_X1 U9241 ( .A1(n8036), .A2(n8298), .B1(n8434), .B2(
        \adder_stage1[14][20] ), .ZN(n8037) );
  INV_X1 U9242 ( .A(n8037), .ZN(n9919) );
  FA_X1 U9243 ( .A(n3455), .B(n3478), .CI(n8038), .CO(n7823), .S(n8039) );
  AOI22_X1 U9244 ( .A1(n8039), .A2(n7971), .B1(n8296), .B2(
        \adder_stage1[3][15] ), .ZN(n8040) );
  INV_X1 U9245 ( .A(n8040), .ZN(n10105) );
  FA_X1 U9246 ( .A(n8797), .B(n3479), .CI(n8041), .CO(n8031), .S(n8042) );
  AOI22_X1 U9247 ( .A1(n8042), .A2(n6279), .B1(n8409), .B2(
        \adder_stage1[12][15] ), .ZN(n8043) );
  INV_X1 U9248 ( .A(n8043), .ZN(n9954) );
  FA_X1 U9249 ( .A(\x_mult_f[4][14] ), .B(\x_mult_f[5][14] ), .CI(n8044), .CO(
        n8399), .S(n7322) );
  AOI21_X1 U9250 ( .B1(n8047), .B2(n7862), .A(n8046), .ZN(n8048) );
  INV_X1 U9251 ( .A(n8048), .ZN(n10121) );
  NAND2_X1 U9252 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  XNOR2_X1 U9253 ( .A(n8052), .B(n8051), .ZN(n8053) );
  AOI22_X1 U9254 ( .A1(n8057), .A2(\adder_stage1[1][12] ), .B1(n8054), .B2(
        n8053), .ZN(n8055) );
  INV_X1 U9255 ( .A(n8055), .ZN(n10140) );
  AOI22_X1 U9256 ( .A1(n8057), .A2(\x_mult_f[9][0] ), .B1(n8087), .B2(
        \x_mult_f_int[9][0] ), .ZN(n8056) );
  INV_X1 U9257 ( .A(n8056), .ZN(n9345) );
  AOI22_X1 U9258 ( .A1(n8057), .A2(\x_mult_f[9][1] ), .B1(n8087), .B2(
        \x_mult_f_int[9][1] ), .ZN(n8058) );
  INV_X1 U9259 ( .A(n8058), .ZN(n9344) );
  AOI22_X1 U9260 ( .A1(\x_mult_f_int[8][14] ), .A2(n8294), .B1(n8323), .B2(
        \x_mult_f[8][14] ), .ZN(n8059) );
  INV_X1 U9261 ( .A(n8059), .ZN(n9013) );
  AOI22_X1 U9262 ( .A1(\x_mult_f_int[27][14] ), .A2(n8153), .B1(n8336), .B2(
        \x_mult_f[27][14] ), .ZN(n8060) );
  INV_X1 U9263 ( .A(n8060), .ZN(n9259) );
  AOI21_X1 U9264 ( .B1(n8137), .B2(n8062), .A(n8061), .ZN(n8066) );
  NAND2_X1 U9265 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  XOR2_X1 U9266 ( .A(n8066), .B(n8065), .Z(n8067) );
  AOI22_X1 U9267 ( .A1(n8067), .A2(n5175), .B1(n8401), .B2(
        \adder_stage4[1][19] ), .ZN(n8068) );
  INV_X1 U9268 ( .A(n8068), .ZN(n9647) );
  NAND2_X1 U9269 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U9270 ( .A1(n8072), .A2(n8071), .ZN(n8076) );
  NAND2_X1 U9271 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  XNOR2_X1 U9272 ( .A(n8076), .B(n8075), .ZN(n8077) );
  AOI22_X1 U9273 ( .A1(n7972), .A2(\adder_stage1[5][12] ), .B1(n8078), .B2(
        n8077), .ZN(n8079) );
  INV_X1 U9274 ( .A(n8079), .ZN(n10074) );
  OAI21_X1 U9275 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n8084) );
  XOR2_X1 U9276 ( .A(\adder_stage2[1][20] ), .B(\adder_stage2[0][20] ), .Z(
        n8083) );
  XOR2_X1 U9277 ( .A(n8084), .B(n8083), .Z(n8085) );
  AOI22_X1 U9278 ( .A1(n8085), .A2(n8298), .B1(n8328), .B2(
        \adder_stage3[0][20] ), .ZN(n8086) );
  INV_X1 U9279 ( .A(n8086), .ZN(n9749) );
  AOI22_X1 U9280 ( .A1(n8088), .A2(\x_mult_f[9][5] ), .B1(n8087), .B2(
        \x_mult_f_int[9][5] ), .ZN(n8089) );
  INV_X1 U9281 ( .A(n8089), .ZN(n9036) );
  OAI21_X1 U9282 ( .B1(n8202), .B2(n8091), .A(n8090), .ZN(n8095) );
  NAND2_X1 U9283 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  XNOR2_X1 U9284 ( .A(n8095), .B(n8094), .ZN(n8096) );
  AOI22_X1 U9285 ( .A1(n8097), .A2(\adder_stage2[4][14] ), .B1(n8209), .B2(
        n8096), .ZN(n8098) );
  INV_X1 U9286 ( .A(n8098), .ZN(n9822) );
  INV_X1 U9287 ( .A(n8099), .ZN(n8101) );
  NAND2_X1 U9288 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  XOR2_X1 U9289 ( .A(n8103), .B(n8102), .Z(n8104) );
  AOI22_X1 U9290 ( .A1(n8273), .A2(\adder_stage3[3][8] ), .B1(n8105), .B2(
        n8104), .ZN(n8106) );
  INV_X1 U9291 ( .A(n8106), .ZN(n9700) );
  INV_X1 U9292 ( .A(n8107), .ZN(n8108) );
  AOI21_X1 U9293 ( .B1(n8110), .B2(n8109), .A(n8108), .ZN(n8115) );
  INV_X1 U9294 ( .A(n8111), .ZN(n8113) );
  NAND2_X1 U9295 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  XOR2_X1 U9296 ( .A(n8115), .B(n8114), .Z(n8116) );
  AOI22_X1 U9297 ( .A1(n8118), .A2(\adder_stage2[2][5] ), .B1(n8117), .B2(
        n8116), .ZN(n8119) );
  INV_X1 U9298 ( .A(n8119), .ZN(n9865) );
  AOI22_X1 U9299 ( .A1(\x_mult_f_int[29][14] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][14] ), .ZN(n8120) );
  INV_X1 U9300 ( .A(n8120), .ZN(n9287) );
  AOI22_X1 U9301 ( .A1(\x_mult_f_int[31][14] ), .A2(n8105), .B1(n8428), .B2(
        \x_mult_f[31][14] ), .ZN(n8121) );
  INV_X1 U9302 ( .A(n8121), .ZN(n9315) );
  AOI22_X1 U9303 ( .A1(\x_mult_f_int[16][14] ), .A2(n6279), .B1(n8313), .B2(
        \x_mult_f[16][14] ), .ZN(n8122) );
  INV_X1 U9304 ( .A(n8122), .ZN(n9124) );
  FA_X1 U9305 ( .A(n3464), .B(n8794), .CI(n8123), .CO(n8124), .S(n7693) );
  INV_X1 U9306 ( .A(n8124), .ZN(n8125) );
  AOI22_X1 U9307 ( .A1(n8125), .A2(n8298), .B1(n8319), .B2(
        \adder_stage1[8][20] ), .ZN(n8126) );
  INV_X1 U9308 ( .A(n8126), .ZN(n10020) );
  FA_X1 U9309 ( .A(\x_mult_f[30][14] ), .B(\x_mult_f[31][14] ), .CI(n8127), 
        .CO(n7834), .S(n8128) );
  AOI22_X1 U9310 ( .A1(n8128), .A2(n7862), .B1(n8434), .B2(
        \adder_stage1[15][14] ), .ZN(n8864) );
  FA_X1 U9311 ( .A(n8800), .B(n3480), .CI(n8129), .CO(n8009), .S(n8130) );
  AOI22_X1 U9312 ( .A1(n8130), .A2(n8298), .B1(n8118), .B2(
        \adder_stage2[1][16] ), .ZN(n8131) );
  INV_X1 U9313 ( .A(n8131), .ZN(n9871) );
  AOI22_X1 U9314 ( .A1(n8134), .A2(n8314), .B1(n8296), .B2(
        \adder_stage2[5][16] ), .ZN(n8865) );
  AOI21_X1 U9315 ( .B1(n8137), .B2(n8136), .A(n8135), .ZN(n8141) );
  NAND2_X1 U9316 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  XOR2_X1 U9317 ( .A(n8141), .B(n8140), .Z(n8142) );
  AOI22_X1 U9318 ( .A1(n8142), .A2(n8294), .B1(n8409), .B2(
        \adder_stage4[1][17] ), .ZN(n8143) );
  INV_X1 U9319 ( .A(n8143), .ZN(n9649) );
  NAND2_X1 U9320 ( .A1(n8145), .A2(n8144), .ZN(n8147) );
  NAND2_X1 U9321 ( .A1(n8147), .A2(n8146), .ZN(n8151) );
  NAND2_X1 U9322 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  XNOR2_X1 U9323 ( .A(n8151), .B(n8150), .ZN(n8152) );
  AOI22_X1 U9324 ( .A1(n8336), .A2(\adder_stage1[7][12] ), .B1(n8153), .B2(
        n8152), .ZN(n8154) );
  INV_X1 U9325 ( .A(n8154), .ZN(n10041) );
  INV_X1 U9326 ( .A(n8155), .ZN(n8157) );
  NAND2_X1 U9327 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  XOR2_X1 U9328 ( .A(n8159), .B(n8158), .Z(n8160) );
  AOI22_X1 U9329 ( .A1(n7928), .A2(\adder_stage1[10][2] ), .B1(n8292), .B2(
        n8160), .ZN(n8161) );
  INV_X1 U9330 ( .A(n8161), .ZN(n10000) );
  NAND2_X1 U9331 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  XNOR2_X1 U9332 ( .A(n8165), .B(n8164), .ZN(n8166) );
  AOI22_X1 U9333 ( .A1(n8168), .A2(\adder_stage1[11][4] ), .B1(n8167), .B2(
        n8166), .ZN(n8169) );
  INV_X1 U9334 ( .A(n8169), .ZN(n9982) );
  NAND2_X1 U9335 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  XNOR2_X1 U9336 ( .A(n8173), .B(n8172), .ZN(n8174) );
  AOI22_X1 U9337 ( .A1(n8176), .A2(\adder_stage1[12][12] ), .B1(n8175), .B2(
        n8174), .ZN(n8177) );
  INV_X1 U9338 ( .A(n8177), .ZN(n9957) );
  NAND2_X1 U9339 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  XNOR2_X1 U9340 ( .A(n8181), .B(n8180), .ZN(n8182) );
  AOI22_X1 U9341 ( .A1(n7041), .A2(\adder_stage1[13][12] ), .B1(n7962), .B2(
        n8182), .ZN(n8183) );
  INV_X1 U9342 ( .A(n8183), .ZN(n9940) );
  NAND2_X1 U9343 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  XNOR2_X1 U9344 ( .A(n8187), .B(n8186), .ZN(n8188) );
  AOI22_X1 U9345 ( .A1(n8245), .A2(\adder_stage2[1][12] ), .B1(n8189), .B2(
        n8188), .ZN(n8190) );
  INV_X1 U9346 ( .A(n8190), .ZN(n9875) );
  OAI21_X1 U9347 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8197) );
  NAND2_X1 U9348 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  XNOR2_X1 U9349 ( .A(n8197), .B(n8196), .ZN(n8198) );
  AOI22_X1 U9350 ( .A1(n7622), .A2(\adder_stage2[3][14] ), .B1(n6875), .B2(
        n8198), .ZN(n8199) );
  INV_X1 U9351 ( .A(n8199), .ZN(n9839) );
  OAI21_X1 U9352 ( .B1(n8202), .B2(n8201), .A(n8200), .ZN(n8203) );
  INV_X1 U9353 ( .A(n8203), .ZN(n8207) );
  NAND2_X1 U9354 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  XOR2_X1 U9355 ( .A(n8207), .B(n8206), .Z(n8208) );
  AOI22_X1 U9356 ( .A1(n8313), .A2(\adder_stage2[4][13] ), .B1(n8209), .B2(
        n8208), .ZN(n8210) );
  INV_X1 U9357 ( .A(n8210), .ZN(n9823) );
  NAND2_X1 U9358 ( .A1(n8212), .A2(n8211), .ZN(n8213) );
  XNOR2_X1 U9359 ( .A(n8214), .B(n8213), .ZN(n8215) );
  AOI22_X1 U9360 ( .A1(n8097), .A2(\adder_stage2[5][14] ), .B1(n8216), .B2(
        n8215), .ZN(n8217) );
  INV_X1 U9361 ( .A(n8217), .ZN(n9805) );
  NAND2_X1 U9362 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  XNOR2_X1 U9363 ( .A(n8222), .B(n8221), .ZN(n8223) );
  AOI22_X1 U9364 ( .A1(n7698), .A2(\adder_stage2[7][14] ), .B1(n8258), .B2(
        n8223), .ZN(n8224) );
  INV_X1 U9365 ( .A(n8224), .ZN(n9772) );
  INV_X1 U9366 ( .A(n8225), .ZN(n8226) );
  AOI21_X1 U9367 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8233) );
  INV_X1 U9368 ( .A(n8229), .ZN(n8231) );
  NAND2_X1 U9369 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  XOR2_X1 U9370 ( .A(n8233), .B(n8232), .Z(n8234) );
  AOI22_X1 U9371 ( .A1(n8428), .A2(\adder_stage3[0][5] ), .B1(n8235), .B2(
        n8234), .ZN(n8236) );
  INV_X1 U9372 ( .A(n8236), .ZN(n9764) );
  OAI21_X1 U9373 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8243) );
  NAND2_X1 U9374 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  XNOR2_X1 U9375 ( .A(n8243), .B(n8242), .ZN(n8244) );
  AOI22_X1 U9376 ( .A1(n8245), .A2(\adder_stage3[0][16] ), .B1(n7971), .B2(
        n8244), .ZN(n8246) );
  INV_X1 U9377 ( .A(n8246), .ZN(n9753) );
  NAND2_X1 U9378 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  XNOR2_X1 U9379 ( .A(n8419), .B(n8249), .ZN(n8250) );
  AOI22_X1 U9380 ( .A1(n7855), .A2(\adder_stage3[1][16] ), .B1(n8251), .B2(
        n8250), .ZN(n8252) );
  INV_X1 U9381 ( .A(n8252), .ZN(n9732) );
  NAND2_X1 U9382 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  XNOR2_X1 U9383 ( .A(n8256), .B(n8255), .ZN(n8257) );
  AOI22_X1 U9384 ( .A1(n7622), .A2(\adder_stage3[2][16] ), .B1(n8258), .B2(
        n8257), .ZN(n8259) );
  INV_X1 U9385 ( .A(n8259), .ZN(n9713) );
  NAND2_X1 U9386 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  XNOR2_X1 U9387 ( .A(n8263), .B(n8262), .ZN(n8264) );
  AOI22_X1 U9388 ( .A1(n8273), .A2(\adder_stage3[3][16] ), .B1(n8265), .B2(
        n8264), .ZN(n8266) );
  INV_X1 U9389 ( .A(n8266), .ZN(n9692) );
  NAND2_X1 U9390 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  XNOR2_X1 U9391 ( .A(n8270), .B(n8269), .ZN(n8271) );
  AOI22_X1 U9392 ( .A1(n8273), .A2(\adder_stage4[0][16] ), .B1(n8272), .B2(
        n8271), .ZN(n8274) );
  INV_X1 U9393 ( .A(n8274), .ZN(n9671) );
  INV_X1 U9394 ( .A(n8275), .ZN(n8277) );
  NAND2_X1 U9395 ( .A1(n8277), .A2(n8276), .ZN(n8279) );
  XOR2_X1 U9396 ( .A(n8279), .B(n8278), .Z(n8280) );
  AOI22_X1 U9397 ( .A1(n8273), .A2(\adder_stage4[1][1] ), .B1(n8281), .B2(
        n8280), .ZN(n8282) );
  INV_X1 U9398 ( .A(n8282), .ZN(n9665) );
  OAI21_X1 U9399 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8290) );
  INV_X1 U9400 ( .A(n8286), .ZN(n8288) );
  NAND2_X1 U9401 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  XNOR2_X1 U9402 ( .A(n8290), .B(n8289), .ZN(n8291) );
  AOI22_X1 U9403 ( .A1(n8306), .A2(\adder_stage4[1][7] ), .B1(n8292), .B2(
        n8291), .ZN(n8293) );
  INV_X1 U9404 ( .A(n8293), .ZN(n9659) );
  AOI22_X1 U9405 ( .A1(\x_mult_f_int[0][15] ), .A2(n8294), .B1(n8427), .B2(
        \x_mult_f[0][15] ), .ZN(n8295) );
  INV_X1 U9406 ( .A(n8295), .ZN(n8913) );
  AOI22_X1 U9407 ( .A1(\x_mult_f_int[13][15] ), .A2(n8272), .B1(n8296), .B2(
        \x_mult_f[13][15] ), .ZN(n8297) );
  INV_X1 U9408 ( .A(n8297), .ZN(n9081) );
  AOI22_X1 U9409 ( .A1(\x_mult_f_int[1][15] ), .A2(n8298), .B1(n8409), .B2(
        \x_mult_f[1][15] ), .ZN(n8299) );
  INV_X1 U9410 ( .A(n8299), .ZN(n8927) );
  AOI22_X1 U9411 ( .A1(\x_mult_f_int[2][15] ), .A2(n8054), .B1(n7864), .B2(
        \x_mult_f[2][15] ), .ZN(n8300) );
  INV_X1 U9412 ( .A(n8300), .ZN(n8941) );
  AOI22_X1 U9413 ( .A1(\x_mult_f_int[3][15] ), .A2(n8301), .B1(n8319), .B2(
        \x_mult_f[3][15] ), .ZN(n8302) );
  INV_X1 U9414 ( .A(n8302), .ZN(n8955) );
  AOI22_X1 U9415 ( .A1(\x_mult_f_int[4][15] ), .A2(n7862), .B1(n8338), .B2(
        \x_mult_f[4][15] ), .ZN(n8303) );
  INV_X1 U9416 ( .A(n8303), .ZN(n8969) );
  AOI22_X1 U9417 ( .A1(\x_mult_f_int[5][15] ), .A2(n7862), .B1(n8338), .B2(
        \x_mult_f[5][15] ), .ZN(n8866) );
  AOI22_X1 U9418 ( .A1(\x_mult_f_int[6][15] ), .A2(n8304), .B1(n8427), .B2(
        \x_mult_f[6][15] ), .ZN(n8305) );
  INV_X1 U9419 ( .A(n8305), .ZN(n8984) );
  AOI22_X1 U9420 ( .A1(\x_mult_f_int[7][15] ), .A2(n8314), .B1(n8306), .B2(
        \x_mult_f[7][15] ), .ZN(n8307) );
  INV_X1 U9421 ( .A(n8307), .ZN(n8998) );
  AOI22_X1 U9422 ( .A1(\x_mult_f_int[8][15] ), .A2(n7927), .B1(n8323), .B2(
        \x_mult_f[8][15] ), .ZN(n8308) );
  INV_X1 U9423 ( .A(n8308), .ZN(n9012) );
  AOI22_X1 U9424 ( .A1(\x_mult_f_int[9][15] ), .A2(n5175), .B1(n8309), .B2(
        \x_mult_f[9][15] ), .ZN(n8310) );
  INV_X1 U9425 ( .A(n8310), .ZN(n9026) );
  AOI22_X1 U9426 ( .A1(\x_mult_f_int[10][15] ), .A2(n8311), .B1(n8306), .B2(
        \x_mult_f[10][15] ), .ZN(n8312) );
  INV_X1 U9427 ( .A(n8312), .ZN(n9040) );
  AOI22_X1 U9428 ( .A1(\x_mult_f_int[11][15] ), .A2(n8314), .B1(n8313), .B2(
        \x_mult_f[11][15] ), .ZN(n8867) );
  AOI22_X1 U9429 ( .A1(\x_mult_f_int[12][15] ), .A2(n8301), .B1(n8336), .B2(
        \x_mult_f[12][15] ), .ZN(n8315) );
  INV_X1 U9430 ( .A(n8315), .ZN(n9067) );
  AOI22_X1 U9431 ( .A1(\x_mult_f_int[14][15] ), .A2(n8334), .B1(n8340), .B2(
        \x_mult_f[14][15] ), .ZN(n8316) );
  INV_X1 U9432 ( .A(n8316), .ZN(n9095) );
  AOI22_X1 U9433 ( .A1(\x_mult_f_int[15][15] ), .A2(n7862), .B1(n8340), .B2(
        \x_mult_f[15][15] ), .ZN(n8317) );
  INV_X1 U9434 ( .A(n8317), .ZN(n9109) );
  AOI22_X1 U9435 ( .A1(\x_mult_f_int[16][15] ), .A2(n7507), .B1(n8409), .B2(
        \x_mult_f[16][15] ), .ZN(n8318) );
  INV_X1 U9436 ( .A(n8318), .ZN(n9123) );
  AOI22_X1 U9437 ( .A1(\x_mult_f_int[17][15] ), .A2(n8332), .B1(n6273), .B2(
        \x_mult_f[17][15] ), .ZN(n8868) );
  AOI22_X1 U9438 ( .A1(\x_mult_f_int[18][15] ), .A2(n6636), .B1(n8319), .B2(
        \x_mult_f[18][15] ), .ZN(n8320) );
  INV_X1 U9439 ( .A(n8320), .ZN(n9140) );
  AOI22_X1 U9440 ( .A1(\x_mult_f_int[19][15] ), .A2(n5175), .B1(n7855), .B2(
        \x_mult_f[19][15] ), .ZN(n8322) );
  INV_X1 U9441 ( .A(n8322), .ZN(n9154) );
  AOI22_X1 U9442 ( .A1(\x_mult_f_int[20][15] ), .A2(n6626), .B1(n8323), .B2(
        \x_mult_f[20][15] ), .ZN(n8324) );
  INV_X1 U9443 ( .A(n8324), .ZN(n9168) );
  AOI22_X1 U9444 ( .A1(\x_mult_f_int[21][15] ), .A2(n6307), .B1(n8325), .B2(
        \x_mult_f[21][15] ), .ZN(n8327) );
  INV_X1 U9445 ( .A(n8327), .ZN(n9182) );
  AOI22_X1 U9446 ( .A1(\x_mult_f_int[22][15] ), .A2(n8281), .B1(n8328), .B2(
        \x_mult_f[22][15] ), .ZN(n8329) );
  INV_X1 U9447 ( .A(n8329), .ZN(n9196) );
  AOI22_X1 U9448 ( .A1(\x_mult_f_int[23][15] ), .A2(n8105), .B1(n8330), .B2(
        \x_mult_f[23][15] ), .ZN(n8331) );
  INV_X1 U9449 ( .A(n8331), .ZN(n9210) );
  AOI22_X1 U9450 ( .A1(\x_mult_f_int[24][15] ), .A2(n8311), .B1(n8427), .B2(
        \x_mult_f[24][15] ), .ZN(n8869) );
  AOI22_X1 U9451 ( .A1(\x_mult_f_int[25][15] ), .A2(n8332), .B1(n8401), .B2(
        \x_mult_f[25][15] ), .ZN(n8333) );
  INV_X1 U9452 ( .A(n8333), .ZN(n9230) );
  AOI22_X1 U9453 ( .A1(\x_mult_f_int[26][15] ), .A2(n8334), .B1(n8401), .B2(
        \x_mult_f[26][15] ), .ZN(n8335) );
  INV_X1 U9454 ( .A(n8335), .ZN(n9244) );
  AOI22_X1 U9455 ( .A1(\x_mult_f_int[27][15] ), .A2(n5981), .B1(n8336), .B2(
        \x_mult_f[27][15] ), .ZN(n8337) );
  INV_X1 U9456 ( .A(n8337), .ZN(n9258) );
  AOI22_X1 U9457 ( .A1(\x_mult_f_int[28][15] ), .A2(n8175), .B1(n8338), .B2(
        \x_mult_f[28][15] ), .ZN(n8339) );
  INV_X1 U9458 ( .A(n8339), .ZN(n9272) );
  AOI22_X1 U9459 ( .A1(\x_mult_f_int[29][15] ), .A2(n8298), .B1(n8340), .B2(
        \x_mult_f[29][15] ), .ZN(n8341) );
  INV_X1 U9460 ( .A(n8341), .ZN(n9286) );
  AOI22_X1 U9461 ( .A1(\x_mult_f_int[30][15] ), .A2(n8298), .B1(n8434), .B2(
        \x_mult_f[30][15] ), .ZN(n8343) );
  INV_X1 U9462 ( .A(n8343), .ZN(n9300) );
  AOI22_X1 U9463 ( .A1(\x_mult_f_int[31][15] ), .A2(n7819), .B1(n8428), .B2(
        \x_mult_f[31][15] ), .ZN(n8344) );
  INV_X1 U9464 ( .A(n8344), .ZN(n9314) );
  INV_X1 U9465 ( .A(n8345), .ZN(n8351) );
  INV_X1 U9466 ( .A(n8392), .ZN(n8346) );
  OAI21_X1 U9467 ( .B1(n8348), .B2(n8347), .A(n8346), .ZN(n8376) );
  NAND2_X1 U9468 ( .A1(n8376), .A2(n8394), .ZN(n8381) );
  NOR2_X1 U9469 ( .A1(n8349), .A2(n8352), .ZN(n8350) );
  AOI211_X1 U9470 ( .C1(n8351), .C2(n3650), .A(n8381), .B(n8350), .ZN(n8353)
         );
  NAND3_X1 U9471 ( .A1(\ctrl_inst/pline_cntr [0]), .A2(
        \ctrl_inst/pline_cntr [1]), .A3(n8355), .ZN(n8359) );
  NOR2_X1 U9472 ( .A1(\ctrl_inst/pline_cntr [2]), .A2(n8359), .ZN(n8362) );
  AOI21_X1 U9473 ( .B1(n8365), .B2(n8352), .A(n8362), .ZN(n8358) );
  NAND2_X1 U9474 ( .A1(n8355), .A2(n8810), .ZN(n8366) );
  INV_X1 U9475 ( .A(n8353), .ZN(n8783) );
  NAND2_X1 U9476 ( .A1(n8366), .A2(n8783), .ZN(n8354) );
  AOI21_X1 U9477 ( .B1(\ctrl_inst/pline_cntr [0]), .B2(n8365), .A(n8354), .ZN(
        n8785) );
  NAND2_X1 U9478 ( .A1(n8355), .A2(n8840), .ZN(n8356) );
  OAI211_X1 U9479 ( .C1(n8373), .C2(n8840), .A(n8785), .B(n8356), .ZN(n8361)
         );
  NAND2_X1 U9480 ( .A1(n8361), .A2(\ctrl_inst/pline_cntr [2]), .ZN(n8357) );
  OAI21_X1 U9481 ( .B1(n8367), .B2(n8358), .A(n8357), .ZN(n3119) );
  INV_X1 U9482 ( .A(n8359), .ZN(n8360) );
  NAND3_X1 U9483 ( .A1(n8841), .A2(\ctrl_inst/pline_cntr [2]), .A3(n8360), 
        .ZN(n8364) );
  AOI211_X1 U9484 ( .C1(\ctrl_inst/pline_cntr [2]), .C2(n8365), .A(n8362), .B(
        n8361), .ZN(n8363) );
  OAI22_X1 U9485 ( .A1(n8367), .A2(n8364), .B1(n8363), .B2(n8841), .ZN(n3118)
         );
  NAND3_X1 U9486 ( .A1(n8365), .A2(n8810), .A3(n8371), .ZN(n8780) );
  NAND2_X1 U9487 ( .A1(n8780), .A2(n8366), .ZN(n8368) );
  MUX2_X1 U9488 ( .A(n8368), .B(\ctrl_inst/pline_cntr [0]), .S(n8367), .Z(
        n3121) );
  INV_X1 U9489 ( .A(n8369), .ZN(n8370) );
  OAI33_X1 U9490 ( .A1(n8373), .A2(n8372), .A3(n8371), .B1(n8844), .B2(n8370), 
        .B3(reset), .ZN(n3390) );
  MUX2_X1 U9491 ( .A(n8375), .B(n8374), .S(\ctrl_inst/xmem_tracker [0]), .Z(
        n3383) );
  INV_X1 U9492 ( .A(n8376), .ZN(n8377) );
  NOR3_X1 U9493 ( .A1(n8379), .A2(n8378), .A3(n8377), .ZN(n8380) );
  NOR2_X1 U9494 ( .A1(n8380), .A2(reset), .ZN(n8387) );
  NOR2_X1 U9495 ( .A1(n8382), .A2(n8381), .ZN(n8385) );
  OR2_X1 U9496 ( .A1(n3666), .A2(n8383), .ZN(n8393) );
  NAND3_X1 U9497 ( .A1(n8385), .A2(n8384), .A3(n8393), .ZN(n8386) );
  MUX2_X1 U9498 ( .A(\ctrl_inst/s_ready_fsm ), .B(n8387), .S(n8386), .Z(n3385)
         );
  INV_X4 U9499 ( .A(n8388), .ZN(n8389) );
  MUX2_X1 U9500 ( .A(s_data_in_x[0]), .B(\xmem_data[31][0] ), .S(n8389), .Z(
        n3370) );
  INV_X4 U9501 ( .A(n8388), .ZN(n8390) );
  MUX2_X1 U9502 ( .A(\xmem_data[31][0] ), .B(\xmem_data[30][0] ), .S(n8390), 
        .Z(n10410) );
  MUX2_X1 U9503 ( .A(\xmem_data[30][0] ), .B(\xmem_data[29][0] ), .S(n8389), 
        .Z(n10402) );
  MUX2_X1 U9504 ( .A(\xmem_data[29][0] ), .B(\xmem_data[28][0] ), .S(n8391), 
        .Z(n10394) );
  MUX2_X1 U9505 ( .A(\xmem_data[28][0] ), .B(\xmem_data[27][0] ), .S(n8391), 
        .Z(n10386) );
  MUX2_X1 U9506 ( .A(\xmem_data[27][0] ), .B(\xmem_data[26][0] ), .S(n8391), 
        .Z(n10378) );
  MUX2_X1 U9507 ( .A(\xmem_data[26][0] ), .B(\xmem_data[25][0] ), .S(n8390), 
        .Z(n10245) );
  MUX2_X1 U9508 ( .A(\xmem_data[25][0] ), .B(\xmem_data[24][0] ), .S(n8389), 
        .Z(n10244) );
  MUX2_X1 U9509 ( .A(\xmem_data[24][0] ), .B(\xmem_data[23][0] ), .S(n8390), 
        .Z(n10243) );
  MUX2_X1 U9510 ( .A(\xmem_data[23][0] ), .B(\xmem_data[22][0] ), .S(n8391), 
        .Z(n10242) );
  MUX2_X1 U9511 ( .A(\xmem_data[22][0] ), .B(\xmem_data[21][0] ), .S(n8389), 
        .Z(n10241) );
  MUX2_X1 U9512 ( .A(\xmem_data[21][0] ), .B(\xmem_data[20][0] ), .S(n8391), 
        .Z(n10240) );
  MUX2_X1 U9513 ( .A(\xmem_data[20][0] ), .B(\xmem_data[19][0] ), .S(n8389), 
        .Z(n10239) );
  MUX2_X1 U9514 ( .A(\xmem_data[19][0] ), .B(\xmem_data[18][0] ), .S(n8390), 
        .Z(n10238) );
  MUX2_X1 U9515 ( .A(\xmem_data[18][0] ), .B(\xmem_data[17][0] ), .S(n8390), 
        .Z(n10237) );
  MUX2_X1 U9516 ( .A(\xmem_data[17][0] ), .B(\xmem_data[16][0] ), .S(n8389), 
        .Z(n10236) );
  MUX2_X1 U9517 ( .A(\xmem_data[16][0] ), .B(\xmem_data[15][0] ), .S(n8391), 
        .Z(n10235) );
  MUX2_X1 U9518 ( .A(\xmem_data[15][0] ), .B(\xmem_data[14][0] ), .S(n8391), 
        .Z(n10234) );
  MUX2_X1 U9519 ( .A(\xmem_data[14][0] ), .B(\xmem_data[13][0] ), .S(n8389), 
        .Z(n10233) );
  MUX2_X1 U9520 ( .A(\xmem_data[13][0] ), .B(\xmem_data[12][0] ), .S(n8389), 
        .Z(n10232) );
  MUX2_X1 U9521 ( .A(\xmem_data[12][0] ), .B(\xmem_data[11][0] ), .S(n8390), 
        .Z(n10231) );
  MUX2_X1 U9522 ( .A(\xmem_data[11][0] ), .B(\xmem_data[10][0] ), .S(n8391), 
        .Z(n10230) );
  MUX2_X1 U9523 ( .A(\xmem_data[10][0] ), .B(\xmem_data[9][0] ), .S(n8389), 
        .Z(n10229) );
  MUX2_X1 U9524 ( .A(\xmem_data[9][0] ), .B(\xmem_data[8][0] ), .S(n8390), .Z(
        n10228) );
  MUX2_X1 U9525 ( .A(\xmem_data[8][0] ), .B(\xmem_data[7][0] ), .S(n8389), .Z(
        n10227) );
  MUX2_X1 U9526 ( .A(\xmem_data[7][0] ), .B(\xmem_data[6][0] ), .S(n8390), .Z(
        n10226) );
  MUX2_X1 U9527 ( .A(\xmem_data[6][0] ), .B(\xmem_data[5][0] ), .S(n8391), .Z(
        n10225) );
  MUX2_X1 U9528 ( .A(\xmem_data[5][0] ), .B(\xmem_data[4][0] ), .S(n8390), .Z(
        n10224) );
  MUX2_X1 U9529 ( .A(\xmem_data[4][0] ), .B(\xmem_data[3][0] ), .S(n8390), .Z(
        n10223) );
  MUX2_X1 U9530 ( .A(\xmem_data[3][0] ), .B(\xmem_data[2][0] ), .S(n8391), .Z(
        n10222) );
  MUX2_X1 U9531 ( .A(\xmem_data[2][0] ), .B(\xmem_data[1][0] ), .S(n8391), .Z(
        n10221) );
  MUX2_X1 U9532 ( .A(\xmem_data[1][0] ), .B(\xmem_data[0][0] ), .S(n8389), .Z(
        n10220) );
  MUX2_X1 U9533 ( .A(s_data_in_x[1]), .B(\xmem_data[31][1] ), .S(n8389), .Z(
        n3371) );
  MUX2_X1 U9534 ( .A(\xmem_data[31][1] ), .B(\xmem_data[30][1] ), .S(n8389), 
        .Z(n10411) );
  MUX2_X1 U9535 ( .A(\xmem_data[30][1] ), .B(\xmem_data[29][1] ), .S(n8390), 
        .Z(n10403) );
  MUX2_X1 U9536 ( .A(\xmem_data[29][1] ), .B(\xmem_data[28][1] ), .S(n8390), 
        .Z(n10395) );
  MUX2_X1 U9537 ( .A(\xmem_data[28][1] ), .B(\xmem_data[27][1] ), .S(n8389), 
        .Z(n10387) );
  MUX2_X1 U9538 ( .A(\xmem_data[27][1] ), .B(\xmem_data[26][1] ), .S(n8390), 
        .Z(n10379) );
  MUX2_X1 U9539 ( .A(\xmem_data[26][1] ), .B(\xmem_data[25][1] ), .S(n8389), 
        .Z(n10271) );
  MUX2_X1 U9540 ( .A(\xmem_data[25][1] ), .B(\xmem_data[24][1] ), .S(n8391), 
        .Z(n10270) );
  MUX2_X1 U9541 ( .A(\xmem_data[24][1] ), .B(\xmem_data[23][1] ), .S(n8391), 
        .Z(n10269) );
  MUX2_X1 U9542 ( .A(\xmem_data[23][1] ), .B(\xmem_data[22][1] ), .S(n8391), 
        .Z(n10268) );
  MUX2_X1 U9543 ( .A(\xmem_data[22][1] ), .B(\xmem_data[21][1] ), .S(n8389), 
        .Z(n10267) );
  MUX2_X1 U9544 ( .A(\xmem_data[21][1] ), .B(\xmem_data[20][1] ), .S(n8391), 
        .Z(n10266) );
  MUX2_X1 U9545 ( .A(\xmem_data[20][1] ), .B(\xmem_data[19][1] ), .S(n8389), 
        .Z(n10265) );
  MUX2_X1 U9546 ( .A(\xmem_data[19][1] ), .B(\xmem_data[18][1] ), .S(n8389), 
        .Z(n10264) );
  MUX2_X1 U9547 ( .A(\xmem_data[18][1] ), .B(\xmem_data[17][1] ), .S(n8390), 
        .Z(n10263) );
  MUX2_X1 U9548 ( .A(\xmem_data[17][1] ), .B(\xmem_data[16][1] ), .S(n8389), 
        .Z(n10262) );
  MUX2_X1 U9549 ( .A(\xmem_data[16][1] ), .B(\xmem_data[15][1] ), .S(n8389), 
        .Z(n10261) );
  MUX2_X1 U9550 ( .A(\xmem_data[15][1] ), .B(\xmem_data[14][1] ), .S(n8390), 
        .Z(n10260) );
  MUX2_X1 U9551 ( .A(\xmem_data[14][1] ), .B(\xmem_data[13][1] ), .S(n8389), 
        .Z(n10259) );
  MUX2_X1 U9552 ( .A(\xmem_data[13][1] ), .B(\xmem_data[12][1] ), .S(n8389), 
        .Z(n10258) );
  MUX2_X1 U9553 ( .A(\xmem_data[12][1] ), .B(\xmem_data[11][1] ), .S(n8391), 
        .Z(n10257) );
  MUX2_X1 U9554 ( .A(\xmem_data[11][1] ), .B(\xmem_data[10][1] ), .S(n8390), 
        .Z(n10256) );
  MUX2_X1 U9555 ( .A(\xmem_data[10][1] ), .B(\xmem_data[9][1] ), .S(n8391), 
        .Z(n10255) );
  MUX2_X1 U9556 ( .A(\xmem_data[9][1] ), .B(\xmem_data[8][1] ), .S(n8390), .Z(
        n10254) );
  MUX2_X1 U9557 ( .A(\xmem_data[8][1] ), .B(\xmem_data[7][1] ), .S(n8390), .Z(
        n10253) );
  MUX2_X1 U9558 ( .A(\xmem_data[7][1] ), .B(\xmem_data[6][1] ), .S(n8389), .Z(
        n10252) );
  MUX2_X1 U9559 ( .A(\xmem_data[6][1] ), .B(\xmem_data[5][1] ), .S(n8391), .Z(
        n10251) );
  MUX2_X1 U9560 ( .A(\xmem_data[5][1] ), .B(\xmem_data[4][1] ), .S(n8390), .Z(
        n10250) );
  MUX2_X1 U9561 ( .A(\xmem_data[4][1] ), .B(\xmem_data[3][1] ), .S(n8389), .Z(
        n10249) );
  MUX2_X1 U9562 ( .A(\xmem_data[3][1] ), .B(\xmem_data[2][1] ), .S(n8390), .Z(
        n10248) );
  MUX2_X1 U9563 ( .A(\xmem_data[2][1] ), .B(\xmem_data[1][1] ), .S(n8390), .Z(
        n10247) );
  MUX2_X1 U9564 ( .A(\xmem_data[1][1] ), .B(\xmem_data[0][1] ), .S(n8390), .Z(
        n10246) );
  MUX2_X1 U9565 ( .A(s_data_in_x[2]), .B(\xmem_data[31][2] ), .S(n8389), .Z(
        n3372) );
  MUX2_X1 U9566 ( .A(\xmem_data[31][2] ), .B(\xmem_data[30][2] ), .S(n8389), 
        .Z(n10412) );
  MUX2_X1 U9567 ( .A(\xmem_data[30][2] ), .B(\xmem_data[29][2] ), .S(n8390), 
        .Z(n10404) );
  MUX2_X1 U9568 ( .A(\xmem_data[29][2] ), .B(\xmem_data[28][2] ), .S(n8390), 
        .Z(n10396) );
  MUX2_X1 U9569 ( .A(\xmem_data[28][2] ), .B(\xmem_data[27][2] ), .S(n8391), 
        .Z(n10388) );
  MUX2_X1 U9570 ( .A(\xmem_data[27][2] ), .B(\xmem_data[26][2] ), .S(n8389), 
        .Z(n10380) );
  MUX2_X1 U9571 ( .A(\xmem_data[26][2] ), .B(\xmem_data[25][2] ), .S(n8390), 
        .Z(n10297) );
  MUX2_X1 U9572 ( .A(\xmem_data[25][2] ), .B(\xmem_data[24][2] ), .S(n8391), 
        .Z(n10296) );
  MUX2_X1 U9573 ( .A(\xmem_data[24][2] ), .B(\xmem_data[23][2] ), .S(n8389), 
        .Z(n10295) );
  MUX2_X1 U9574 ( .A(\xmem_data[23][2] ), .B(\xmem_data[22][2] ), .S(n8391), 
        .Z(n10294) );
  MUX2_X1 U9575 ( .A(\xmem_data[22][2] ), .B(\xmem_data[21][2] ), .S(n8391), 
        .Z(n10293) );
  MUX2_X1 U9576 ( .A(\xmem_data[21][2] ), .B(\xmem_data[20][2] ), .S(n8389), 
        .Z(n10292) );
  MUX2_X1 U9577 ( .A(\xmem_data[20][2] ), .B(\xmem_data[19][2] ), .S(n8391), 
        .Z(n10291) );
  MUX2_X1 U9578 ( .A(\xmem_data[19][2] ), .B(\xmem_data[18][2] ), .S(n8390), 
        .Z(n10290) );
  MUX2_X1 U9579 ( .A(\xmem_data[18][2] ), .B(\xmem_data[17][2] ), .S(n8390), 
        .Z(n10289) );
  MUX2_X1 U9580 ( .A(\xmem_data[17][2] ), .B(\xmem_data[16][2] ), .S(n8389), 
        .Z(n10288) );
  MUX2_X1 U9581 ( .A(\xmem_data[16][2] ), .B(\xmem_data[15][2] ), .S(n8389), 
        .Z(n10287) );
  MUX2_X1 U9582 ( .A(\xmem_data[15][2] ), .B(\xmem_data[14][2] ), .S(n8389), 
        .Z(n10286) );
  MUX2_X1 U9583 ( .A(\xmem_data[14][2] ), .B(\xmem_data[13][2] ), .S(n8389), 
        .Z(n10285) );
  MUX2_X1 U9584 ( .A(\xmem_data[13][2] ), .B(\xmem_data[12][2] ), .S(n8390), 
        .Z(n10284) );
  MUX2_X1 U9585 ( .A(\xmem_data[12][2] ), .B(\xmem_data[11][2] ), .S(n8390), 
        .Z(n10283) );
  MUX2_X1 U9586 ( .A(\xmem_data[11][2] ), .B(\xmem_data[10][2] ), .S(n8390), 
        .Z(n10282) );
  MUX2_X1 U9587 ( .A(\xmem_data[10][2] ), .B(\xmem_data[9][2] ), .S(n8391), 
        .Z(n10281) );
  MUX2_X1 U9588 ( .A(\xmem_data[9][2] ), .B(\xmem_data[8][2] ), .S(n8391), .Z(
        n10280) );
  MUX2_X1 U9589 ( .A(\xmem_data[8][2] ), .B(\xmem_data[7][2] ), .S(n8391), .Z(
        n10279) );
  MUX2_X1 U9590 ( .A(\xmem_data[7][2] ), .B(\xmem_data[6][2] ), .S(n8389), .Z(
        n10278) );
  MUX2_X1 U9591 ( .A(\xmem_data[6][2] ), .B(\xmem_data[5][2] ), .S(n8390), .Z(
        n10277) );
  MUX2_X1 U9592 ( .A(\xmem_data[5][2] ), .B(\xmem_data[4][2] ), .S(n8390), .Z(
        n10276) );
  MUX2_X1 U9593 ( .A(\xmem_data[4][2] ), .B(\xmem_data[3][2] ), .S(n8390), .Z(
        n10275) );
  MUX2_X1 U9594 ( .A(\xmem_data[3][2] ), .B(\xmem_data[2][2] ), .S(n8391), .Z(
        n10274) );
  MUX2_X1 U9595 ( .A(\xmem_data[2][2] ), .B(\xmem_data[1][2] ), .S(n8389), .Z(
        n10273) );
  MUX2_X1 U9596 ( .A(\xmem_data[1][2] ), .B(\xmem_data[0][2] ), .S(n8390), .Z(
        n10272) );
  MUX2_X1 U9597 ( .A(s_data_in_x[3]), .B(\xmem_data[31][3] ), .S(n8391), .Z(
        n3373) );
  MUX2_X1 U9598 ( .A(\xmem_data[31][3] ), .B(\xmem_data[30][3] ), .S(n8389), 
        .Z(n10413) );
  MUX2_X1 U9599 ( .A(\xmem_data[30][3] ), .B(\xmem_data[29][3] ), .S(n8391), 
        .Z(n10405) );
  MUX2_X1 U9600 ( .A(\xmem_data[29][3] ), .B(\xmem_data[28][3] ), .S(n8391), 
        .Z(n10397) );
  MUX2_X1 U9601 ( .A(\xmem_data[28][3] ), .B(\xmem_data[27][3] ), .S(n8390), 
        .Z(n10389) );
  MUX2_X1 U9602 ( .A(\xmem_data[27][3] ), .B(\xmem_data[26][3] ), .S(n8391), 
        .Z(n10381) );
  MUX2_X1 U9603 ( .A(\xmem_data[26][3] ), .B(\xmem_data[25][3] ), .S(n8390), 
        .Z(n10323) );
  MUX2_X1 U9604 ( .A(\xmem_data[25][3] ), .B(\xmem_data[24][3] ), .S(n8389), 
        .Z(n10322) );
  MUX2_X1 U9605 ( .A(\xmem_data[24][3] ), .B(\xmem_data[23][3] ), .S(n8391), 
        .Z(n10321) );
  MUX2_X1 U9606 ( .A(\xmem_data[23][3] ), .B(\xmem_data[22][3] ), .S(n8391), 
        .Z(n10320) );
  MUX2_X1 U9607 ( .A(\xmem_data[22][3] ), .B(\xmem_data[21][3] ), .S(n8390), 
        .Z(n10319) );
  MUX2_X1 U9608 ( .A(\xmem_data[21][3] ), .B(\xmem_data[20][3] ), .S(n8389), 
        .Z(n10318) );
  MUX2_X1 U9609 ( .A(\xmem_data[20][3] ), .B(\xmem_data[19][3] ), .S(n8391), 
        .Z(n10317) );
  MUX2_X1 U9610 ( .A(\xmem_data[19][3] ), .B(\xmem_data[18][3] ), .S(n8390), 
        .Z(n10316) );
  MUX2_X1 U9611 ( .A(\xmem_data[18][3] ), .B(\xmem_data[17][3] ), .S(n8389), 
        .Z(n10315) );
  MUX2_X1 U9612 ( .A(\xmem_data[17][3] ), .B(\xmem_data[16][3] ), .S(n8391), 
        .Z(n10314) );
  MUX2_X1 U9613 ( .A(\xmem_data[16][3] ), .B(\xmem_data[15][3] ), .S(n8390), 
        .Z(n10313) );
  MUX2_X1 U9614 ( .A(\xmem_data[15][3] ), .B(\xmem_data[14][3] ), .S(n8391), 
        .Z(n10312) );
  MUX2_X1 U9615 ( .A(\xmem_data[14][3] ), .B(\xmem_data[13][3] ), .S(n8389), 
        .Z(n10311) );
  MUX2_X1 U9616 ( .A(\xmem_data[13][3] ), .B(\xmem_data[12][3] ), .S(n8389), 
        .Z(n10310) );
  MUX2_X1 U9617 ( .A(\xmem_data[12][3] ), .B(\xmem_data[11][3] ), .S(n8389), 
        .Z(n10309) );
  MUX2_X1 U9618 ( .A(\xmem_data[11][3] ), .B(\xmem_data[10][3] ), .S(n8391), 
        .Z(n10308) );
  MUX2_X1 U9619 ( .A(\xmem_data[10][3] ), .B(\xmem_data[9][3] ), .S(n8391), 
        .Z(n10307) );
  MUX2_X1 U9620 ( .A(\xmem_data[9][3] ), .B(\xmem_data[8][3] ), .S(n8390), .Z(
        n10306) );
  MUX2_X1 U9621 ( .A(\xmem_data[8][3] ), .B(\xmem_data[7][3] ), .S(n8389), .Z(
        n10305) );
  MUX2_X1 U9622 ( .A(\xmem_data[7][3] ), .B(\xmem_data[6][3] ), .S(n8390), .Z(
        n10304) );
  MUX2_X1 U9623 ( .A(\xmem_data[6][3] ), .B(\xmem_data[5][3] ), .S(n8391), .Z(
        n10303) );
  MUX2_X1 U9624 ( .A(\xmem_data[5][3] ), .B(\xmem_data[4][3] ), .S(n8390), .Z(
        n10302) );
  MUX2_X1 U9625 ( .A(\xmem_data[4][3] ), .B(\xmem_data[3][3] ), .S(n8391), .Z(
        n10301) );
  MUX2_X1 U9626 ( .A(\xmem_data[3][3] ), .B(\xmem_data[2][3] ), .S(n8390), .Z(
        n10300) );
  MUX2_X1 U9627 ( .A(\xmem_data[2][3] ), .B(\xmem_data[1][3] ), .S(n8391), .Z(
        n10299) );
  MUX2_X1 U9628 ( .A(\xmem_data[1][3] ), .B(\xmem_data[0][3] ), .S(n8390), .Z(
        n10298) );
  MUX2_X1 U9629 ( .A(s_data_in_x[4]), .B(\xmem_data[31][4] ), .S(n8391), .Z(
        n3374) );
  MUX2_X1 U9630 ( .A(\xmem_data[31][4] ), .B(\xmem_data[30][4] ), .S(n8391), 
        .Z(n10414) );
  MUX2_X1 U9631 ( .A(\xmem_data[30][4] ), .B(\xmem_data[29][4] ), .S(n8390), 
        .Z(n10406) );
  MUX2_X1 U9632 ( .A(\xmem_data[29][4] ), .B(\xmem_data[28][4] ), .S(n8391), 
        .Z(n10398) );
  MUX2_X1 U9633 ( .A(\xmem_data[28][4] ), .B(\xmem_data[27][4] ), .S(n8389), 
        .Z(n10390) );
  MUX2_X1 U9634 ( .A(\xmem_data[27][4] ), .B(\xmem_data[26][4] ), .S(n8391), 
        .Z(n10382) );
  MUX2_X1 U9635 ( .A(\xmem_data[26][4] ), .B(\xmem_data[25][4] ), .S(n8389), 
        .Z(n10349) );
  MUX2_X1 U9636 ( .A(\xmem_data[25][4] ), .B(\xmem_data[24][4] ), .S(n8390), 
        .Z(n10348) );
  MUX2_X1 U9637 ( .A(\xmem_data[24][4] ), .B(\xmem_data[23][4] ), .S(n8391), 
        .Z(n10347) );
  MUX2_X1 U9638 ( .A(\xmem_data[23][4] ), .B(\xmem_data[22][4] ), .S(n8389), 
        .Z(n10346) );
  MUX2_X1 U9639 ( .A(\xmem_data[22][4] ), .B(\xmem_data[21][4] ), .S(n8391), 
        .Z(n10345) );
  MUX2_X1 U9640 ( .A(\xmem_data[21][4] ), .B(\xmem_data[20][4] ), .S(n8390), 
        .Z(n10344) );
  MUX2_X1 U9641 ( .A(\xmem_data[20][4] ), .B(\xmem_data[19][4] ), .S(n8391), 
        .Z(n10343) );
  MUX2_X1 U9642 ( .A(\xmem_data[19][4] ), .B(\xmem_data[18][4] ), .S(n8389), 
        .Z(n10342) );
  MUX2_X1 U9643 ( .A(\xmem_data[18][4] ), .B(\xmem_data[17][4] ), .S(n8391), 
        .Z(n10341) );
  MUX2_X1 U9644 ( .A(\xmem_data[17][4] ), .B(\xmem_data[16][4] ), .S(n8390), 
        .Z(n10340) );
  MUX2_X1 U9645 ( .A(\xmem_data[16][4] ), .B(\xmem_data[15][4] ), .S(n8390), 
        .Z(n10339) );
  MUX2_X1 U9646 ( .A(\xmem_data[15][4] ), .B(\xmem_data[14][4] ), .S(n8389), 
        .Z(n10338) );
  MUX2_X1 U9647 ( .A(\xmem_data[14][4] ), .B(\xmem_data[13][4] ), .S(n8390), 
        .Z(n10337) );
  MUX2_X1 U9648 ( .A(\xmem_data[13][4] ), .B(\xmem_data[12][4] ), .S(n8389), 
        .Z(n10336) );
  MUX2_X1 U9649 ( .A(\xmem_data[12][4] ), .B(\xmem_data[11][4] ), .S(n8390), 
        .Z(n10335) );
  MUX2_X1 U9650 ( .A(\xmem_data[11][4] ), .B(\xmem_data[10][4] ), .S(n8391), 
        .Z(n10334) );
  MUX2_X1 U9651 ( .A(\xmem_data[10][4] ), .B(\xmem_data[9][4] ), .S(n8390), 
        .Z(n10333) );
  MUX2_X1 U9652 ( .A(\xmem_data[9][4] ), .B(\xmem_data[8][4] ), .S(n8389), .Z(
        n10332) );
  MUX2_X1 U9653 ( .A(\xmem_data[8][4] ), .B(\xmem_data[7][4] ), .S(n8391), .Z(
        n10331) );
  MUX2_X1 U9654 ( .A(\xmem_data[7][4] ), .B(\xmem_data[6][4] ), .S(n8389), .Z(
        n10330) );
  MUX2_X1 U9655 ( .A(\xmem_data[6][4] ), .B(\xmem_data[5][4] ), .S(n8389), .Z(
        n10329) );
  MUX2_X1 U9656 ( .A(\xmem_data[5][4] ), .B(\xmem_data[4][4] ), .S(n8390), .Z(
        n10328) );
  MUX2_X1 U9657 ( .A(\xmem_data[4][4] ), .B(\xmem_data[3][4] ), .S(n8390), .Z(
        n10327) );
  MUX2_X1 U9658 ( .A(\xmem_data[3][4] ), .B(\xmem_data[2][4] ), .S(n8391), .Z(
        n10326) );
  MUX2_X1 U9659 ( .A(\xmem_data[2][4] ), .B(\xmem_data[1][4] ), .S(n8390), .Z(
        n10325) );
  MUX2_X1 U9660 ( .A(\xmem_data[1][4] ), .B(\xmem_data[0][4] ), .S(n8389), .Z(
        n10324) );
  MUX2_X1 U9661 ( .A(s_data_in_x[5]), .B(\xmem_data[31][5] ), .S(n8389), .Z(
        n3375) );
  MUX2_X1 U9662 ( .A(\xmem_data[31][5] ), .B(\xmem_data[30][5] ), .S(n8390), 
        .Z(n10415) );
  MUX2_X1 U9663 ( .A(\xmem_data[30][5] ), .B(\xmem_data[29][5] ), .S(n8391), 
        .Z(n10407) );
  MUX2_X1 U9664 ( .A(\xmem_data[29][5] ), .B(\xmem_data[28][5] ), .S(n8391), 
        .Z(n10399) );
  MUX2_X1 U9665 ( .A(\xmem_data[28][5] ), .B(\xmem_data[27][5] ), .S(n8391), 
        .Z(n10391) );
  MUX2_X1 U9666 ( .A(\xmem_data[27][5] ), .B(\xmem_data[26][5] ), .S(n8389), 
        .Z(n10383) );
  MUX2_X1 U9667 ( .A(\xmem_data[26][5] ), .B(\xmem_data[25][5] ), .S(n8390), 
        .Z(n10375) );
  MUX2_X1 U9668 ( .A(\xmem_data[25][5] ), .B(\xmem_data[24][5] ), .S(n8390), 
        .Z(n10374) );
  MUX2_X1 U9669 ( .A(\xmem_data[24][5] ), .B(\xmem_data[23][5] ), .S(n8389), 
        .Z(n10373) );
  MUX2_X1 U9670 ( .A(\xmem_data[23][5] ), .B(\xmem_data[22][5] ), .S(n8390), 
        .Z(n10372) );
  MUX2_X1 U9671 ( .A(\xmem_data[22][5] ), .B(\xmem_data[21][5] ), .S(n8389), 
        .Z(n10371) );
  MUX2_X1 U9672 ( .A(\xmem_data[21][5] ), .B(\xmem_data[20][5] ), .S(n8390), 
        .Z(n10370) );
  MUX2_X1 U9673 ( .A(\xmem_data[20][5] ), .B(\xmem_data[19][5] ), .S(n8389), 
        .Z(n10369) );
  MUX2_X1 U9674 ( .A(\xmem_data[19][5] ), .B(\xmem_data[18][5] ), .S(n8391), 
        .Z(n10368) );
  MUX2_X1 U9675 ( .A(\xmem_data[18][5] ), .B(\xmem_data[17][5] ), .S(n8391), 
        .Z(n10367) );
  MUX2_X1 U9676 ( .A(\xmem_data[17][5] ), .B(\xmem_data[16][5] ), .S(n8391), 
        .Z(n10366) );
  MUX2_X1 U9677 ( .A(\xmem_data[16][5] ), .B(\xmem_data[15][5] ), .S(n8391), 
        .Z(n10365) );
  MUX2_X1 U9678 ( .A(\xmem_data[15][5] ), .B(\xmem_data[14][5] ), .S(n8390), 
        .Z(n10364) );
  MUX2_X1 U9679 ( .A(\xmem_data[14][5] ), .B(\xmem_data[13][5] ), .S(n8391), 
        .Z(n10363) );
  MUX2_X1 U9680 ( .A(\xmem_data[13][5] ), .B(\xmem_data[12][5] ), .S(n8389), 
        .Z(n10362) );
  MUX2_X1 U9681 ( .A(\xmem_data[12][5] ), .B(\xmem_data[11][5] ), .S(n8390), 
        .Z(n10361) );
  MUX2_X1 U9682 ( .A(\xmem_data[11][5] ), .B(\xmem_data[10][5] ), .S(n8389), 
        .Z(n10360) );
  MUX2_X1 U9683 ( .A(\xmem_data[10][5] ), .B(\xmem_data[9][5] ), .S(n8389), 
        .Z(n10359) );
  MUX2_X1 U9684 ( .A(\xmem_data[9][5] ), .B(\xmem_data[8][5] ), .S(n8391), .Z(
        n10358) );
  MUX2_X1 U9685 ( .A(\xmem_data[8][5] ), .B(\xmem_data[7][5] ), .S(n8391), .Z(
        n10357) );
  MUX2_X1 U9686 ( .A(\xmem_data[7][5] ), .B(\xmem_data[6][5] ), .S(n8389), .Z(
        n10356) );
  MUX2_X1 U9687 ( .A(\xmem_data[6][5] ), .B(\xmem_data[5][5] ), .S(n8391), .Z(
        n10355) );
  MUX2_X1 U9688 ( .A(\xmem_data[5][5] ), .B(\xmem_data[4][5] ), .S(n8389), .Z(
        n10354) );
  MUX2_X1 U9689 ( .A(\xmem_data[4][5] ), .B(\xmem_data[3][5] ), .S(n8391), .Z(
        n10353) );
  MUX2_X1 U9690 ( .A(\xmem_data[3][5] ), .B(\xmem_data[2][5] ), .S(n8390), .Z(
        n10352) );
  MUX2_X1 U9691 ( .A(\xmem_data[2][5] ), .B(\xmem_data[1][5] ), .S(n8389), .Z(
        n10351) );
  MUX2_X1 U9692 ( .A(\xmem_data[1][5] ), .B(\xmem_data[0][5] ), .S(n8390), .Z(
        n10350) );
  MUX2_X1 U9693 ( .A(s_data_in_x[6]), .B(\xmem_data[31][6] ), .S(n8389), .Z(
        n3376) );
  MUX2_X1 U9694 ( .A(\xmem_data[31][6] ), .B(\xmem_data[30][6] ), .S(n8389), 
        .Z(n10416) );
  MUX2_X1 U9695 ( .A(\xmem_data[30][6] ), .B(\xmem_data[29][6] ), .S(n8390), 
        .Z(n10408) );
  MUX2_X1 U9696 ( .A(\xmem_data[29][6] ), .B(\xmem_data[28][6] ), .S(n8391), 
        .Z(n10400) );
  MUX2_X1 U9697 ( .A(\xmem_data[28][6] ), .B(\xmem_data[27][6] ), .S(n8390), 
        .Z(n10392) );
  MUX2_X1 U9698 ( .A(\xmem_data[27][6] ), .B(\xmem_data[26][6] ), .S(n8391), 
        .Z(n10384) );
  MUX2_X1 U9699 ( .A(\xmem_data[26][6] ), .B(\xmem_data[25][6] ), .S(n8391), 
        .Z(n10376) );
  MUX2_X1 U9700 ( .A(\xmem_data[25][6] ), .B(\xmem_data[24][6] ), .S(n8390), 
        .Z(n10194) );
  MUX2_X1 U9701 ( .A(\xmem_data[24][6] ), .B(\xmem_data[23][6] ), .S(n8391), 
        .Z(n10193) );
  MUX2_X1 U9702 ( .A(\xmem_data[23][6] ), .B(\xmem_data[22][6] ), .S(n8390), 
        .Z(n10192) );
  MUX2_X1 U9703 ( .A(\xmem_data[22][6] ), .B(\xmem_data[21][6] ), .S(n8389), 
        .Z(n10191) );
  MUX2_X1 U9704 ( .A(\xmem_data[21][6] ), .B(\xmem_data[20][6] ), .S(n8389), 
        .Z(n10190) );
  MUX2_X1 U9705 ( .A(\xmem_data[20][6] ), .B(\xmem_data[19][6] ), .S(n8389), 
        .Z(n10189) );
  MUX2_X1 U9706 ( .A(\xmem_data[19][6] ), .B(\xmem_data[18][6] ), .S(n8390), 
        .Z(n10188) );
  MUX2_X1 U9707 ( .A(\xmem_data[18][6] ), .B(\xmem_data[17][6] ), .S(n8390), 
        .Z(n10187) );
  MUX2_X1 U9708 ( .A(\xmem_data[17][6] ), .B(\xmem_data[16][6] ), .S(n8391), 
        .Z(n10186) );
  MUX2_X1 U9709 ( .A(\xmem_data[16][6] ), .B(\xmem_data[15][6] ), .S(n8391), 
        .Z(n10185) );
  MUX2_X1 U9710 ( .A(\xmem_data[15][6] ), .B(\xmem_data[14][6] ), .S(n8390), 
        .Z(n10184) );
  MUX2_X1 U9711 ( .A(\xmem_data[14][6] ), .B(\xmem_data[13][6] ), .S(n8390), 
        .Z(n10183) );
  MUX2_X1 U9712 ( .A(\xmem_data[13][6] ), .B(\xmem_data[12][6] ), .S(n8391), 
        .Z(n10182) );
  MUX2_X1 U9713 ( .A(\xmem_data[12][6] ), .B(\xmem_data[11][6] ), .S(n8391), 
        .Z(n10181) );
  MUX2_X1 U9714 ( .A(\xmem_data[11][6] ), .B(\xmem_data[10][6] ), .S(n8389), 
        .Z(n10180) );
  MUX2_X1 U9715 ( .A(\xmem_data[10][6] ), .B(\xmem_data[9][6] ), .S(n8390), 
        .Z(n10179) );
  MUX2_X1 U9716 ( .A(\xmem_data[9][6] ), .B(\xmem_data[8][6] ), .S(n8389), .Z(
        n10178) );
  MUX2_X1 U9717 ( .A(\xmem_data[8][6] ), .B(\xmem_data[7][6] ), .S(n8389), .Z(
        n10177) );
  MUX2_X1 U9718 ( .A(\xmem_data[7][6] ), .B(\xmem_data[6][6] ), .S(n8389), .Z(
        n10176) );
  MUX2_X1 U9719 ( .A(\xmem_data[6][6] ), .B(\xmem_data[5][6] ), .S(n8389), .Z(
        n10175) );
  MUX2_X1 U9720 ( .A(\xmem_data[5][6] ), .B(\xmem_data[4][6] ), .S(n8390), .Z(
        n10174) );
  MUX2_X1 U9721 ( .A(\xmem_data[4][6] ), .B(\xmem_data[3][6] ), .S(n8389), .Z(
        n10173) );
  MUX2_X1 U9722 ( .A(\xmem_data[3][6] ), .B(\xmem_data[2][6] ), .S(n8389), .Z(
        n10172) );
  MUX2_X1 U9723 ( .A(\xmem_data[2][6] ), .B(\xmem_data[1][6] ), .S(n8391), .Z(
        n10171) );
  MUX2_X1 U9724 ( .A(\xmem_data[1][6] ), .B(\xmem_data[0][6] ), .S(n8391), .Z(
        n10170) );
  MUX2_X1 U9725 ( .A(s_data_in_x[7]), .B(\xmem_data[31][7] ), .S(n8390), .Z(
        n3377) );
  MUX2_X1 U9726 ( .A(\xmem_data[31][7] ), .B(\xmem_data[30][7] ), .S(n8389), 
        .Z(n10417) );
  MUX2_X1 U9727 ( .A(\xmem_data[30][7] ), .B(\xmem_data[29][7] ), .S(n8389), 
        .Z(n10409) );
  MUX2_X1 U9728 ( .A(\xmem_data[29][7] ), .B(\xmem_data[28][7] ), .S(n8389), 
        .Z(n10401) );
  MUX2_X1 U9729 ( .A(\xmem_data[28][7] ), .B(\xmem_data[27][7] ), .S(n8390), 
        .Z(n10393) );
  MUX2_X1 U9730 ( .A(\xmem_data[27][7] ), .B(\xmem_data[26][7] ), .S(n8391), 
        .Z(n10385) );
  MUX2_X1 U9731 ( .A(\xmem_data[26][7] ), .B(\xmem_data[25][7] ), .S(n8389), 
        .Z(n10377) );
  MUX2_X1 U9732 ( .A(\xmem_data[25][7] ), .B(\xmem_data[24][7] ), .S(n8390), 
        .Z(n10219) );
  MUX2_X1 U9733 ( .A(\xmem_data[24][7] ), .B(\xmem_data[23][7] ), .S(n8390), 
        .Z(n10218) );
  MUX2_X1 U9734 ( .A(\xmem_data[23][7] ), .B(\xmem_data[22][7] ), .S(n8390), 
        .Z(n10217) );
  MUX2_X1 U9735 ( .A(\xmem_data[22][7] ), .B(\xmem_data[21][7] ), .S(n8391), 
        .Z(n10216) );
  MUX2_X1 U9736 ( .A(\xmem_data[21][7] ), .B(\xmem_data[20][7] ), .S(n8391), 
        .Z(n10215) );
  MUX2_X1 U9737 ( .A(\xmem_data[20][7] ), .B(\xmem_data[19][7] ), .S(n8389), 
        .Z(n10214) );
  MUX2_X1 U9738 ( .A(\xmem_data[19][7] ), .B(\xmem_data[18][7] ), .S(n8389), 
        .Z(n10213) );
  MUX2_X1 U9739 ( .A(\xmem_data[18][7] ), .B(\xmem_data[17][7] ), .S(n8390), 
        .Z(n10212) );
  MUX2_X1 U9740 ( .A(\xmem_data[17][7] ), .B(\xmem_data[16][7] ), .S(n8391), 
        .Z(n10211) );
  MUX2_X1 U9741 ( .A(\xmem_data[16][7] ), .B(\xmem_data[15][7] ), .S(n8389), 
        .Z(n10210) );
  MUX2_X1 U9742 ( .A(\xmem_data[15][7] ), .B(\xmem_data[14][7] ), .S(n8390), 
        .Z(n10209) );
  MUX2_X1 U9743 ( .A(\xmem_data[14][7] ), .B(\xmem_data[13][7] ), .S(n8391), 
        .Z(n10208) );
  MUX2_X1 U9744 ( .A(\xmem_data[13][7] ), .B(\xmem_data[12][7] ), .S(n8391), 
        .Z(n10207) );
  MUX2_X1 U9745 ( .A(\xmem_data[12][7] ), .B(\xmem_data[11][7] ), .S(n8389), 
        .Z(n10206) );
  MUX2_X1 U9746 ( .A(\xmem_data[11][7] ), .B(\xmem_data[10][7] ), .S(n8390), 
        .Z(n10205) );
  MUX2_X1 U9747 ( .A(\xmem_data[10][7] ), .B(\xmem_data[9][7] ), .S(n8390), 
        .Z(n10204) );
  MUX2_X1 U9748 ( .A(\xmem_data[9][7] ), .B(\xmem_data[8][7] ), .S(n8391), .Z(
        n10203) );
  MUX2_X1 U9749 ( .A(\xmem_data[8][7] ), .B(\xmem_data[7][7] ), .S(n8391), .Z(
        n10202) );
  MUX2_X1 U9750 ( .A(\xmem_data[7][7] ), .B(\xmem_data[6][7] ), .S(n8391), .Z(
        n10201) );
  MUX2_X1 U9751 ( .A(\xmem_data[6][7] ), .B(\xmem_data[5][7] ), .S(n8389), .Z(
        n10200) );
  MUX2_X1 U9752 ( .A(\xmem_data[5][7] ), .B(\xmem_data[4][7] ), .S(n8391), .Z(
        n10199) );
  MUX2_X1 U9753 ( .A(\xmem_data[4][7] ), .B(\xmem_data[3][7] ), .S(n8390), .Z(
        n10198) );
  MUX2_X1 U9754 ( .A(\xmem_data[3][7] ), .B(\xmem_data[2][7] ), .S(n8391), .Z(
        n10197) );
  MUX2_X1 U9755 ( .A(\xmem_data[2][7] ), .B(\xmem_data[1][7] ), .S(n8389), .Z(
        n10196) );
  MUX2_X1 U9756 ( .A(\xmem_data[1][7] ), .B(\xmem_data[0][7] ), .S(n8390), .Z(
        n10195) );
  NOR2_X1 U9757 ( .A1(n8392), .A2(reset), .ZN(n8397) );
  NAND3_X1 U9758 ( .A1(n8395), .A2(n8394), .A3(n8393), .ZN(n8396) );
  MUX2_X1 U9759 ( .A(xmem_full), .B(n8397), .S(n8396), .Z(n3391) );
  AOI22_X1 U9760 ( .A1(\x_mult_f_int[4][9] ), .A2(n7862), .B1(n6877), .B2(
        \x_mult_f[4][9] ), .ZN(n8872) );
  AOI22_X1 U9761 ( .A1(\x_mult_f_int[4][8] ), .A2(n7862), .B1(n8088), .B2(
        \x_mult_f[4][8] ), .ZN(n8873) );
  AOI22_X1 U9762 ( .A1(\x_mult_f_int[4][7] ), .A2(n7862), .B1(n8245), .B2(
        \x_mult_f[4][7] ), .ZN(n8874) );
  AOI22_X1 U9763 ( .A1(\x_mult_f_int[4][6] ), .A2(n7862), .B1(n8428), .B2(
        \x_mult_f[4][6] ), .ZN(n8875) );
  AOI22_X1 U9764 ( .A1(\x_mult_f_int[5][11] ), .A2(n7862), .B1(n8401), .B2(
        \x_mult_f[5][11] ), .ZN(n8876) );
  AOI22_X1 U9765 ( .A1(\x_mult_f_int[5][10] ), .A2(n7862), .B1(n8401), .B2(
        \x_mult_f[5][10] ), .ZN(n8877) );
  AOI22_X1 U9766 ( .A1(\x_mult_f_int[5][9] ), .A2(n7862), .B1(n8409), .B2(
        \x_mult_f[5][9] ), .ZN(n8878) );
  AOI22_X1 U9767 ( .A1(\x_mult_f_int[5][8] ), .A2(n7862), .B1(n8398), .B2(
        \x_mult_f[5][8] ), .ZN(n8879) );
  AOI22_X1 U9768 ( .A1(\x_mult_f_int[5][7] ), .A2(n7862), .B1(n8401), .B2(
        \x_mult_f[5][7] ), .ZN(n8880) );
  AOI22_X1 U9769 ( .A1(\x_mult_f_int[5][6] ), .A2(n8258), .B1(n8398), .B2(
        \x_mult_f[5][6] ), .ZN(n8881) );
  FA_X1 U9770 ( .A(n3465), .B(n8790), .CI(n8399), .CO(n8400), .S(n8047) );
  INV_X1 U9771 ( .A(n8400), .ZN(n8402) );
  AOI22_X1 U9772 ( .A1(n8402), .A2(n8078), .B1(n8401), .B2(
        \adder_stage1[2][20] ), .ZN(n8882) );
  INV_X1 U9773 ( .A(n8404), .ZN(n8406) );
  NAND2_X1 U9774 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  XOR2_X1 U9775 ( .A(n8408), .B(n8407), .Z(n8410) );
  AOI22_X1 U9776 ( .A1(n8410), .A2(n8117), .B1(n8409), .B2(
        \adder_stage1[2][13] ), .ZN(n8883) );
  AOI21_X1 U9777 ( .B1(n8419), .B2(n8412), .A(n8411), .ZN(n8416) );
  NAND2_X1 U9778 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  XOR2_X1 U9779 ( .A(n8416), .B(n8415), .Z(n8417) );
  AOI22_X1 U9780 ( .A1(n8417), .A2(n8334), .B1(n7959), .B2(
        \adder_stage3[1][19] ), .ZN(n8884) );
  NAND2_X1 U9781 ( .A1(n8419), .A2(n8418), .ZN(n8421) );
  NAND2_X1 U9782 ( .A1(n8421), .A2(n8420), .ZN(n8425) );
  NAND2_X1 U9783 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  XNOR2_X1 U9784 ( .A(n8425), .B(n8424), .ZN(n8426) );
  AOI22_X1 U9785 ( .A1(n8426), .A2(n8078), .B1(n7959), .B2(
        \adder_stage3[1][18] ), .ZN(n8885) );
  AOI22_X1 U9786 ( .A1(\x_mult_f_int[16][11] ), .A2(n8117), .B1(n7959), .B2(
        \x_mult_f[16][11] ), .ZN(n8886) );
  AOI22_X1 U9787 ( .A1(\x_mult_f_int[16][10] ), .A2(n8251), .B1(n7928), .B2(
        \x_mult_f[16][10] ), .ZN(n8887) );
  AOI22_X1 U9788 ( .A1(\x_mult_f_int[16][9] ), .A2(n8272), .B1(n6273), .B2(
        \x_mult_f[16][9] ), .ZN(n8888) );
  AOI22_X1 U9789 ( .A1(\x_mult_f_int[16][8] ), .A2(n7570), .B1(n7525), .B2(
        \x_mult_f[16][8] ), .ZN(n8889) );
  AOI22_X1 U9790 ( .A1(\x_mult_f_int[16][7] ), .A2(n7155), .B1(n7920), .B2(
        \x_mult_f[16][7] ), .ZN(n8890) );
  AOI22_X1 U9791 ( .A1(\x_mult_f_int[16][6] ), .A2(n6609), .B1(n6273), .B2(
        \x_mult_f[16][6] ), .ZN(n8891) );
  AOI22_X1 U9792 ( .A1(\x_mult_f_int[24][11] ), .A2(n4894), .B1(n8427), .B2(
        \x_mult_f[24][11] ), .ZN(n8893) );
  AOI22_X1 U9793 ( .A1(\x_mult_f_int[24][10] ), .A2(n8334), .B1(n8427), .B2(
        \x_mult_f[24][10] ), .ZN(n8894) );
  AOI22_X1 U9794 ( .A1(\x_mult_f_int[24][9] ), .A2(n8311), .B1(n8427), .B2(
        \x_mult_f[24][9] ), .ZN(n8895) );
  AOI22_X1 U9795 ( .A1(\x_mult_f_int[24][8] ), .A2(n6875), .B1(n6854), .B2(
        \x_mult_f[24][8] ), .ZN(n8896) );
  AOI22_X1 U9796 ( .A1(\x_mult_f_int[24][7] ), .A2(n7507), .B1(n6273), .B2(
        \x_mult_f[24][7] ), .ZN(n8897) );
  AOI22_X1 U9797 ( .A1(\x_mult_f_int[31][7] ), .A2(n8251), .B1(n7920), .B2(
        \x_mult_f[31][7] ), .ZN(n8898) );
  AOI22_X1 U9798 ( .A1(\x_mult_f_int[31][6] ), .A2(n8272), .B1(n8428), .B2(
        \x_mult_f[31][6] ), .ZN(n8899) );
  INV_X1 U9799 ( .A(n8429), .ZN(n8431) );
  NAND2_X1 U9800 ( .A1(n8431), .A2(n8430), .ZN(n8432) );
  XOR2_X1 U9801 ( .A(n8433), .B(n8432), .Z(n8435) );
  AOI22_X1 U9802 ( .A1(n8435), .A2(n5175), .B1(n8434), .B2(
        \adder_stage1[15][13] ), .ZN(n8900) );
  NAND3_X1 U9803 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .A3(fmem_addr[2]), 
        .ZN(n8766) );
  NAND2_X1 U9804 ( .A1(n8771), .A2(fmem_addr[4]), .ZN(n8515) );
  OAI22_X1 U9805 ( .A1(n3444), .A2(s_data_in_f[7]), .B1(\fmem_data[31][7] ), 
        .B2(n8779), .ZN(n8436) );
  INV_X1 U9806 ( .A(n8436), .ZN(n9390) );
  OAI22_X1 U9807 ( .A1(n3444), .A2(s_data_in_f[6]), .B1(\fmem_data[31][6] ), 
        .B2(n8779), .ZN(n8437) );
  INV_X1 U9808 ( .A(n8437), .ZN(n9391) );
  OAI22_X1 U9809 ( .A1(n3444), .A2(s_data_in_f[5]), .B1(\fmem_data[31][5] ), 
        .B2(n8779), .ZN(n8438) );
  INV_X1 U9810 ( .A(n8438), .ZN(n9392) );
  OAI22_X1 U9811 ( .A1(n3444), .A2(s_data_in_f[4]), .B1(\fmem_data[31][4] ), 
        .B2(n8779), .ZN(n8439) );
  INV_X1 U9812 ( .A(n8439), .ZN(n9393) );
  OAI22_X1 U9813 ( .A1(n3444), .A2(s_data_in_f[3]), .B1(\fmem_data[31][3] ), 
        .B2(n8779), .ZN(n8440) );
  INV_X1 U9814 ( .A(n8440), .ZN(n9394) );
  OAI22_X1 U9815 ( .A1(n3444), .A2(s_data_in_f[2]), .B1(\fmem_data[31][2] ), 
        .B2(n8779), .ZN(n8441) );
  INV_X1 U9816 ( .A(n8441), .ZN(n9395) );
  OAI22_X1 U9817 ( .A1(n3444), .A2(s_data_in_f[1]), .B1(\fmem_data[31][1] ), 
        .B2(n8779), .ZN(n8442) );
  INV_X1 U9818 ( .A(n8442), .ZN(n9396) );
  OAI22_X1 U9819 ( .A1(n3444), .A2(s_data_in_f[0]), .B1(\fmem_data[31][0] ), 
        .B2(n8779), .ZN(n8443) );
  INV_X1 U9820 ( .A(n8443), .ZN(n9397) );
  NAND3_X1 U9821 ( .A1(fmem_addr[1]), .A2(fmem_addr[2]), .A3(n8805), .ZN(n8688) );
  OAI22_X1 U9822 ( .A1(n8452), .A2(s_data_in_f[7]), .B1(\fmem_data[30][7] ), 
        .B2(n8451), .ZN(n8444) );
  INV_X1 U9823 ( .A(n8444), .ZN(n9398) );
  OAI22_X1 U9824 ( .A1(n8452), .A2(s_data_in_f[6]), .B1(\fmem_data[30][6] ), 
        .B2(n8451), .ZN(n8445) );
  INV_X1 U9825 ( .A(n8445), .ZN(n9399) );
  OAI22_X1 U9826 ( .A1(n8452), .A2(s_data_in_f[5]), .B1(\fmem_data[30][5] ), 
        .B2(n8451), .ZN(n8446) );
  INV_X1 U9827 ( .A(n8446), .ZN(n9400) );
  OAI22_X1 U9828 ( .A1(n8452), .A2(s_data_in_f[4]), .B1(\fmem_data[30][4] ), 
        .B2(n8451), .ZN(n8447) );
  INV_X1 U9829 ( .A(n8447), .ZN(n9401) );
  OAI22_X1 U9830 ( .A1(n8452), .A2(s_data_in_f[3]), .B1(\fmem_data[30][3] ), 
        .B2(n8451), .ZN(n8448) );
  INV_X1 U9831 ( .A(n8448), .ZN(n9402) );
  OAI22_X1 U9832 ( .A1(n8452), .A2(s_data_in_f[2]), .B1(\fmem_data[30][2] ), 
        .B2(n8451), .ZN(n8449) );
  INV_X1 U9833 ( .A(n8449), .ZN(n9403) );
  OAI22_X1 U9834 ( .A1(n8452), .A2(s_data_in_f[1]), .B1(\fmem_data[30][1] ), 
        .B2(n8451), .ZN(n8450) );
  INV_X1 U9835 ( .A(n8450), .ZN(n9404) );
  OAI22_X1 U9836 ( .A1(n8452), .A2(s_data_in_f[0]), .B1(\fmem_data[30][0] ), 
        .B2(n8451), .ZN(n8453) );
  INV_X1 U9837 ( .A(n8453), .ZN(n9405) );
  NAND3_X1 U9838 ( .A1(fmem_addr[0]), .A2(fmem_addr[2]), .A3(n8808), .ZN(n8699) );
  OAI22_X1 U9839 ( .A1(n8462), .A2(s_data_in_f[7]), .B1(\fmem_data[29][7] ), 
        .B2(n8461), .ZN(n8454) );
  INV_X1 U9840 ( .A(n8454), .ZN(n9406) );
  OAI22_X1 U9841 ( .A1(n8462), .A2(s_data_in_f[6]), .B1(\fmem_data[29][6] ), 
        .B2(n8461), .ZN(n8455) );
  INV_X1 U9842 ( .A(n8455), .ZN(n9407) );
  OAI22_X1 U9843 ( .A1(n8462), .A2(s_data_in_f[5]), .B1(\fmem_data[29][5] ), 
        .B2(n8461), .ZN(n8456) );
  INV_X1 U9844 ( .A(n8456), .ZN(n9408) );
  OAI22_X1 U9845 ( .A1(n8462), .A2(s_data_in_f[4]), .B1(\fmem_data[29][4] ), 
        .B2(n8461), .ZN(n8457) );
  INV_X1 U9846 ( .A(n8457), .ZN(n9409) );
  OAI22_X1 U9847 ( .A1(n8462), .A2(s_data_in_f[3]), .B1(\fmem_data[29][3] ), 
        .B2(n8461), .ZN(n8458) );
  INV_X1 U9848 ( .A(n8458), .ZN(n9410) );
  OAI22_X1 U9849 ( .A1(n8462), .A2(s_data_in_f[2]), .B1(\fmem_data[29][2] ), 
        .B2(n8461), .ZN(n8459) );
  INV_X1 U9850 ( .A(n8459), .ZN(n9411) );
  OAI22_X1 U9851 ( .A1(n8462), .A2(s_data_in_f[1]), .B1(\fmem_data[29][1] ), 
        .B2(n8461), .ZN(n8460) );
  INV_X1 U9852 ( .A(n8460), .ZN(n9412) );
  OAI22_X1 U9853 ( .A1(n8462), .A2(s_data_in_f[0]), .B1(\fmem_data[29][0] ), 
        .B2(n8461), .ZN(n8463) );
  INV_X1 U9854 ( .A(n8463), .ZN(n9413) );
  NAND3_X1 U9855 ( .A1(fmem_addr[2]), .A2(n8805), .A3(n8808), .ZN(n8710) );
  OAI22_X1 U9856 ( .A1(n8472), .A2(s_data_in_f[7]), .B1(\fmem_data[28][7] ), 
        .B2(n8471), .ZN(n8464) );
  INV_X1 U9857 ( .A(n8464), .ZN(n9414) );
  OAI22_X1 U9858 ( .A1(n8472), .A2(s_data_in_f[6]), .B1(\fmem_data[28][6] ), 
        .B2(n8471), .ZN(n8465) );
  INV_X1 U9859 ( .A(n8465), .ZN(n9415) );
  OAI22_X1 U9860 ( .A1(n8472), .A2(s_data_in_f[5]), .B1(\fmem_data[28][5] ), 
        .B2(n8471), .ZN(n8466) );
  INV_X1 U9861 ( .A(n8466), .ZN(n9416) );
  OAI22_X1 U9862 ( .A1(n8472), .A2(s_data_in_f[4]), .B1(\fmem_data[28][4] ), 
        .B2(n8471), .ZN(n8467) );
  INV_X1 U9863 ( .A(n8467), .ZN(n9417) );
  OAI22_X1 U9864 ( .A1(n8472), .A2(s_data_in_f[3]), .B1(\fmem_data[28][3] ), 
        .B2(n8471), .ZN(n8468) );
  INV_X1 U9865 ( .A(n8468), .ZN(n9418) );
  OAI22_X1 U9866 ( .A1(n8472), .A2(s_data_in_f[2]), .B1(\fmem_data[28][2] ), 
        .B2(n8471), .ZN(n8469) );
  INV_X1 U9867 ( .A(n8469), .ZN(n9419) );
  OAI22_X1 U9868 ( .A1(n8472), .A2(s_data_in_f[1]), .B1(\fmem_data[28][1] ), 
        .B2(n8471), .ZN(n8470) );
  INV_X1 U9869 ( .A(n8470), .ZN(n9420) );
  OAI22_X1 U9870 ( .A1(n8472), .A2(s_data_in_f[0]), .B1(\fmem_data[28][0] ), 
        .B2(n8471), .ZN(n8473) );
  INV_X1 U9871 ( .A(n8473), .ZN(n9421) );
  NAND3_X1 U9872 ( .A1(fmem_addr[1]), .A2(fmem_addr[0]), .A3(n8804), .ZN(n8775) );
  OAI22_X1 U9873 ( .A1(n8482), .A2(s_data_in_f[7]), .B1(\fmem_data[27][7] ), 
        .B2(n8481), .ZN(n8474) );
  INV_X1 U9874 ( .A(n8474), .ZN(n9422) );
  OAI22_X1 U9875 ( .A1(n8482), .A2(s_data_in_f[6]), .B1(\fmem_data[27][6] ), 
        .B2(n8481), .ZN(n8475) );
  INV_X1 U9876 ( .A(n8475), .ZN(n9423) );
  OAI22_X1 U9877 ( .A1(n8482), .A2(s_data_in_f[5]), .B1(\fmem_data[27][5] ), 
        .B2(n8481), .ZN(n8476) );
  INV_X1 U9878 ( .A(n8476), .ZN(n9424) );
  OAI22_X1 U9879 ( .A1(n8482), .A2(s_data_in_f[4]), .B1(\fmem_data[27][4] ), 
        .B2(n8481), .ZN(n8477) );
  INV_X1 U9880 ( .A(n8477), .ZN(n9425) );
  OAI22_X1 U9881 ( .A1(n8482), .A2(s_data_in_f[3]), .B1(\fmem_data[27][3] ), 
        .B2(n8481), .ZN(n8478) );
  INV_X1 U9882 ( .A(n8478), .ZN(n9426) );
  OAI22_X1 U9883 ( .A1(n8482), .A2(s_data_in_f[2]), .B1(\fmem_data[27][2] ), 
        .B2(n8481), .ZN(n8479) );
  INV_X1 U9884 ( .A(n8479), .ZN(n9427) );
  OAI22_X1 U9885 ( .A1(n8482), .A2(s_data_in_f[1]), .B1(\fmem_data[27][1] ), 
        .B2(n8481), .ZN(n8480) );
  INV_X1 U9886 ( .A(n8480), .ZN(n9428) );
  OAI22_X1 U9887 ( .A1(n8482), .A2(s_data_in_f[0]), .B1(\fmem_data[27][0] ), 
        .B2(n8481), .ZN(n8483) );
  INV_X1 U9888 ( .A(n8483), .ZN(n9429) );
  NAND3_X1 U9889 ( .A1(fmem_addr[1]), .A2(n8805), .A3(n8804), .ZN(n8731) );
  OAI22_X1 U9890 ( .A1(n8492), .A2(s_data_in_f[7]), .B1(\fmem_data[26][7] ), 
        .B2(n8491), .ZN(n8484) );
  INV_X1 U9891 ( .A(n8484), .ZN(n9430) );
  OAI22_X1 U9892 ( .A1(n8492), .A2(s_data_in_f[6]), .B1(\fmem_data[26][6] ), 
        .B2(n8491), .ZN(n8485) );
  INV_X1 U9893 ( .A(n8485), .ZN(n9431) );
  OAI22_X1 U9894 ( .A1(n8492), .A2(s_data_in_f[5]), .B1(\fmem_data[26][5] ), 
        .B2(n8491), .ZN(n8486) );
  INV_X1 U9895 ( .A(n8486), .ZN(n9432) );
  OAI22_X1 U9896 ( .A1(n8492), .A2(s_data_in_f[4]), .B1(\fmem_data[26][4] ), 
        .B2(n8491), .ZN(n8487) );
  INV_X1 U9897 ( .A(n8487), .ZN(n9433) );
  OAI22_X1 U9898 ( .A1(n8492), .A2(s_data_in_f[3]), .B1(\fmem_data[26][3] ), 
        .B2(n8491), .ZN(n8488) );
  INV_X1 U9899 ( .A(n8488), .ZN(n9434) );
  OAI22_X1 U9900 ( .A1(n8492), .A2(s_data_in_f[2]), .B1(\fmem_data[26][2] ), 
        .B2(n8491), .ZN(n8489) );
  INV_X1 U9901 ( .A(n8489), .ZN(n9435) );
  OAI22_X1 U9902 ( .A1(n8492), .A2(s_data_in_f[1]), .B1(\fmem_data[26][1] ), 
        .B2(n8491), .ZN(n8490) );
  INV_X1 U9903 ( .A(n8490), .ZN(n9436) );
  OAI22_X1 U9904 ( .A1(n8492), .A2(s_data_in_f[0]), .B1(\fmem_data[26][0] ), 
        .B2(n8491), .ZN(n8493) );
  INV_X1 U9905 ( .A(n8493), .ZN(n9437) );
  NAND3_X1 U9906 ( .A1(fmem_addr[0]), .A2(n8808), .A3(n8804), .ZN(n8742) );
  OAI22_X1 U9907 ( .A1(n8502), .A2(s_data_in_f[7]), .B1(\fmem_data[25][7] ), 
        .B2(n8501), .ZN(n8494) );
  INV_X1 U9908 ( .A(n8494), .ZN(n9438) );
  OAI22_X1 U9909 ( .A1(n8502), .A2(s_data_in_f[6]), .B1(\fmem_data[25][6] ), 
        .B2(n8501), .ZN(n8495) );
  INV_X1 U9910 ( .A(n8495), .ZN(n9439) );
  OAI22_X1 U9911 ( .A1(n8502), .A2(s_data_in_f[5]), .B1(\fmem_data[25][5] ), 
        .B2(n8501), .ZN(n8496) );
  INV_X1 U9912 ( .A(n8496), .ZN(n9440) );
  OAI22_X1 U9913 ( .A1(n8502), .A2(s_data_in_f[4]), .B1(\fmem_data[25][4] ), 
        .B2(n8501), .ZN(n8497) );
  INV_X1 U9914 ( .A(n8497), .ZN(n9441) );
  OAI22_X1 U9915 ( .A1(n8502), .A2(s_data_in_f[3]), .B1(\fmem_data[25][3] ), 
        .B2(n8501), .ZN(n8498) );
  INV_X1 U9916 ( .A(n8498), .ZN(n9442) );
  OAI22_X1 U9917 ( .A1(n8502), .A2(s_data_in_f[2]), .B1(\fmem_data[25][2] ), 
        .B2(n8501), .ZN(n8499) );
  INV_X1 U9918 ( .A(n8499), .ZN(n9443) );
  OAI22_X1 U9919 ( .A1(n8502), .A2(s_data_in_f[1]), .B1(\fmem_data[25][1] ), 
        .B2(n8501), .ZN(n8500) );
  INV_X1 U9920 ( .A(n8500), .ZN(n9444) );
  OAI22_X1 U9921 ( .A1(n8502), .A2(s_data_in_f[0]), .B1(\fmem_data[25][0] ), 
        .B2(n8501), .ZN(n8503) );
  INV_X1 U9922 ( .A(n8503), .ZN(n9445) );
  NAND3_X1 U9923 ( .A1(n8805), .A2(n8808), .A3(n8804), .ZN(n8754) );
  OAI22_X1 U9924 ( .A1(n8513), .A2(s_data_in_f[7]), .B1(\fmem_data[24][7] ), 
        .B2(n8512), .ZN(n8505) );
  INV_X1 U9925 ( .A(n8505), .ZN(n9446) );
  OAI22_X1 U9926 ( .A1(n8513), .A2(s_data_in_f[6]), .B1(\fmem_data[24][6] ), 
        .B2(n8512), .ZN(n8506) );
  INV_X1 U9927 ( .A(n8506), .ZN(n9447) );
  OAI22_X1 U9928 ( .A1(n8513), .A2(s_data_in_f[5]), .B1(\fmem_data[24][5] ), 
        .B2(n8512), .ZN(n8507) );
  INV_X1 U9929 ( .A(n8507), .ZN(n9448) );
  OAI22_X1 U9930 ( .A1(n8513), .A2(s_data_in_f[4]), .B1(\fmem_data[24][4] ), 
        .B2(n8512), .ZN(n8508) );
  INV_X1 U9931 ( .A(n8508), .ZN(n9449) );
  OAI22_X1 U9932 ( .A1(n8513), .A2(s_data_in_f[3]), .B1(\fmem_data[24][3] ), 
        .B2(n8512), .ZN(n8509) );
  INV_X1 U9933 ( .A(n8509), .ZN(n9450) );
  OAI22_X1 U9934 ( .A1(n8513), .A2(s_data_in_f[2]), .B1(\fmem_data[24][2] ), 
        .B2(n8512), .ZN(n8510) );
  INV_X1 U9935 ( .A(n8510), .ZN(n9451) );
  OAI22_X1 U9936 ( .A1(n8513), .A2(s_data_in_f[1]), .B1(\fmem_data[24][1] ), 
        .B2(n8512), .ZN(n8511) );
  INV_X1 U9937 ( .A(n8511), .ZN(n9452) );
  OAI22_X1 U9938 ( .A1(n8513), .A2(s_data_in_f[0]), .B1(\fmem_data[24][0] ), 
        .B2(n8512), .ZN(n8514) );
  INV_X1 U9939 ( .A(n8514), .ZN(n9453) );
  OAI22_X1 U9940 ( .A1(n8524), .A2(s_data_in_f[7]), .B1(\fmem_data[23][7] ), 
        .B2(n8523), .ZN(n8516) );
  INV_X1 U9941 ( .A(n8516), .ZN(n9454) );
  OAI22_X1 U9942 ( .A1(n8524), .A2(s_data_in_f[6]), .B1(\fmem_data[23][6] ), 
        .B2(n8523), .ZN(n8517) );
  INV_X1 U9943 ( .A(n8517), .ZN(n9455) );
  OAI22_X1 U9944 ( .A1(n8524), .A2(s_data_in_f[5]), .B1(\fmem_data[23][5] ), 
        .B2(n8523), .ZN(n8518) );
  INV_X1 U9945 ( .A(n8518), .ZN(n9456) );
  OAI22_X1 U9946 ( .A1(n8524), .A2(s_data_in_f[4]), .B1(\fmem_data[23][4] ), 
        .B2(n8523), .ZN(n8519) );
  INV_X1 U9947 ( .A(n8519), .ZN(n9457) );
  OAI22_X1 U9948 ( .A1(n8524), .A2(s_data_in_f[3]), .B1(\fmem_data[23][3] ), 
        .B2(n8523), .ZN(n8520) );
  INV_X1 U9949 ( .A(n8520), .ZN(n9458) );
  OAI22_X1 U9950 ( .A1(n8524), .A2(s_data_in_f[2]), .B1(\fmem_data[23][2] ), 
        .B2(n8523), .ZN(n8521) );
  INV_X1 U9951 ( .A(n8521), .ZN(n9459) );
  OAI22_X1 U9952 ( .A1(n8524), .A2(s_data_in_f[1]), .B1(\fmem_data[23][1] ), 
        .B2(n8523), .ZN(n8522) );
  INV_X1 U9953 ( .A(n8522), .ZN(n9460) );
  OAI22_X1 U9954 ( .A1(n8524), .A2(s_data_in_f[0]), .B1(\fmem_data[23][0] ), 
        .B2(n8523), .ZN(n8525) );
  INV_X1 U9955 ( .A(n8525), .ZN(n9461) );
  OAI22_X1 U9956 ( .A1(n8534), .A2(s_data_in_f[7]), .B1(\fmem_data[22][7] ), 
        .B2(n8533), .ZN(n8526) );
  INV_X1 U9957 ( .A(n8526), .ZN(n9462) );
  OAI22_X1 U9958 ( .A1(n8534), .A2(s_data_in_f[6]), .B1(\fmem_data[22][6] ), 
        .B2(n8533), .ZN(n8527) );
  INV_X1 U9959 ( .A(n8527), .ZN(n9463) );
  OAI22_X1 U9960 ( .A1(n8534), .A2(s_data_in_f[5]), .B1(\fmem_data[22][5] ), 
        .B2(n8533), .ZN(n8528) );
  INV_X1 U9961 ( .A(n8528), .ZN(n9464) );
  OAI22_X1 U9962 ( .A1(n8534), .A2(s_data_in_f[4]), .B1(\fmem_data[22][4] ), 
        .B2(n8533), .ZN(n8529) );
  INV_X1 U9963 ( .A(n8529), .ZN(n9465) );
  OAI22_X1 U9964 ( .A1(n8534), .A2(s_data_in_f[3]), .B1(\fmem_data[22][3] ), 
        .B2(n8533), .ZN(n8530) );
  INV_X1 U9965 ( .A(n8530), .ZN(n9466) );
  OAI22_X1 U9966 ( .A1(n8534), .A2(s_data_in_f[2]), .B1(\fmem_data[22][2] ), 
        .B2(n8533), .ZN(n8531) );
  INV_X1 U9967 ( .A(n8531), .ZN(n9467) );
  OAI22_X1 U9968 ( .A1(n8534), .A2(s_data_in_f[1]), .B1(\fmem_data[22][1] ), 
        .B2(n8533), .ZN(n8532) );
  INV_X1 U9969 ( .A(n8532), .ZN(n9468) );
  OAI22_X1 U9970 ( .A1(n8534), .A2(s_data_in_f[0]), .B1(\fmem_data[22][0] ), 
        .B2(n8533), .ZN(n8535) );
  INV_X1 U9971 ( .A(n8535), .ZN(n9469) );
  OAI22_X1 U9972 ( .A1(n8544), .A2(s_data_in_f[7]), .B1(\fmem_data[21][7] ), 
        .B2(n8543), .ZN(n8536) );
  INV_X1 U9973 ( .A(n8536), .ZN(n9470) );
  OAI22_X1 U9974 ( .A1(n8544), .A2(s_data_in_f[6]), .B1(\fmem_data[21][6] ), 
        .B2(n8543), .ZN(n8537) );
  INV_X1 U9975 ( .A(n8537), .ZN(n9471) );
  OAI22_X1 U9976 ( .A1(n8544), .A2(s_data_in_f[5]), .B1(\fmem_data[21][5] ), 
        .B2(n8543), .ZN(n8538) );
  INV_X1 U9977 ( .A(n8538), .ZN(n9472) );
  OAI22_X1 U9978 ( .A1(n8544), .A2(s_data_in_f[4]), .B1(\fmem_data[21][4] ), 
        .B2(n8543), .ZN(n8539) );
  INV_X1 U9979 ( .A(n8539), .ZN(n9473) );
  OAI22_X1 U9980 ( .A1(n8544), .A2(s_data_in_f[3]), .B1(\fmem_data[21][3] ), 
        .B2(n8543), .ZN(n8540) );
  INV_X1 U9981 ( .A(n8540), .ZN(n9474) );
  OAI22_X1 U9982 ( .A1(n8544), .A2(s_data_in_f[2]), .B1(\fmem_data[21][2] ), 
        .B2(n8543), .ZN(n8541) );
  INV_X1 U9983 ( .A(n8541), .ZN(n9475) );
  OAI22_X1 U9984 ( .A1(n8544), .A2(s_data_in_f[1]), .B1(\fmem_data[21][1] ), 
        .B2(n8543), .ZN(n8542) );
  INV_X1 U9985 ( .A(n8542), .ZN(n9476) );
  OAI22_X1 U9986 ( .A1(n8544), .A2(s_data_in_f[0]), .B1(\fmem_data[21][0] ), 
        .B2(n8543), .ZN(n8545) );
  INV_X1 U9987 ( .A(n8545), .ZN(n9477) );
  OAI22_X1 U9988 ( .A1(n8554), .A2(s_data_in_f[7]), .B1(\fmem_data[20][7] ), 
        .B2(n8553), .ZN(n8546) );
  INV_X1 U9989 ( .A(n8546), .ZN(n9478) );
  OAI22_X1 U9990 ( .A1(n8554), .A2(s_data_in_f[6]), .B1(\fmem_data[20][6] ), 
        .B2(n8553), .ZN(n8547) );
  INV_X1 U9991 ( .A(n8547), .ZN(n9479) );
  OAI22_X1 U9992 ( .A1(n8554), .A2(s_data_in_f[5]), .B1(\fmem_data[20][5] ), 
        .B2(n8553), .ZN(n8548) );
  INV_X1 U9993 ( .A(n8548), .ZN(n9480) );
  OAI22_X1 U9994 ( .A1(n8554), .A2(s_data_in_f[4]), .B1(\fmem_data[20][4] ), 
        .B2(n8553), .ZN(n8549) );
  INV_X1 U9995 ( .A(n8549), .ZN(n9481) );
  OAI22_X1 U9996 ( .A1(n8554), .A2(s_data_in_f[3]), .B1(\fmem_data[20][3] ), 
        .B2(n8553), .ZN(n8550) );
  INV_X1 U9997 ( .A(n8550), .ZN(n9482) );
  OAI22_X1 U9998 ( .A1(n8554), .A2(s_data_in_f[2]), .B1(\fmem_data[20][2] ), 
        .B2(n8553), .ZN(n8551) );
  INV_X1 U9999 ( .A(n8551), .ZN(n9483) );
  OAI22_X1 U10000 ( .A1(n8554), .A2(s_data_in_f[1]), .B1(\fmem_data[20][1] ), 
        .B2(n8553), .ZN(n8552) );
  INV_X1 U10001 ( .A(n8552), .ZN(n9484) );
  OAI22_X1 U10002 ( .A1(n8554), .A2(s_data_in_f[0]), .B1(\fmem_data[20][0] ), 
        .B2(n8553), .ZN(n8555) );
  INV_X1 U10003 ( .A(n8555), .ZN(n9485) );
  OAI22_X1 U10004 ( .A1(n8564), .A2(s_data_in_f[7]), .B1(\fmem_data[19][7] ), 
        .B2(n8563), .ZN(n8556) );
  INV_X1 U10005 ( .A(n8556), .ZN(n9486) );
  OAI22_X1 U10006 ( .A1(n8564), .A2(s_data_in_f[6]), .B1(\fmem_data[19][6] ), 
        .B2(n8563), .ZN(n8557) );
  INV_X1 U10007 ( .A(n8557), .ZN(n9487) );
  OAI22_X1 U10008 ( .A1(n8564), .A2(s_data_in_f[5]), .B1(\fmem_data[19][5] ), 
        .B2(n8563), .ZN(n8558) );
  INV_X1 U10009 ( .A(n8558), .ZN(n9488) );
  OAI22_X1 U10010 ( .A1(n8564), .A2(s_data_in_f[4]), .B1(\fmem_data[19][4] ), 
        .B2(n8563), .ZN(n8559) );
  INV_X1 U10011 ( .A(n8559), .ZN(n9489) );
  OAI22_X1 U10012 ( .A1(n8564), .A2(s_data_in_f[3]), .B1(\fmem_data[19][3] ), 
        .B2(n8563), .ZN(n8560) );
  INV_X1 U10013 ( .A(n8560), .ZN(n9490) );
  OAI22_X1 U10014 ( .A1(n8564), .A2(s_data_in_f[2]), .B1(\fmem_data[19][2] ), 
        .B2(n8563), .ZN(n8561) );
  INV_X1 U10015 ( .A(n8561), .ZN(n9491) );
  OAI22_X1 U10016 ( .A1(n8564), .A2(s_data_in_f[1]), .B1(\fmem_data[19][1] ), 
        .B2(n8563), .ZN(n8562) );
  INV_X1 U10017 ( .A(n8562), .ZN(n9492) );
  OAI22_X1 U10018 ( .A1(n8564), .A2(s_data_in_f[0]), .B1(\fmem_data[19][0] ), 
        .B2(n8563), .ZN(n8565) );
  INV_X1 U10019 ( .A(n8565), .ZN(n9493) );
  OAI22_X1 U10020 ( .A1(n8574), .A2(s_data_in_f[7]), .B1(\fmem_data[18][7] ), 
        .B2(n8573), .ZN(n8566) );
  INV_X1 U10021 ( .A(n8566), .ZN(n9494) );
  OAI22_X1 U10022 ( .A1(n8574), .A2(s_data_in_f[6]), .B1(\fmem_data[18][6] ), 
        .B2(n8573), .ZN(n8567) );
  INV_X1 U10023 ( .A(n8567), .ZN(n9495) );
  OAI22_X1 U10024 ( .A1(n8574), .A2(s_data_in_f[5]), .B1(\fmem_data[18][5] ), 
        .B2(n8573), .ZN(n8568) );
  INV_X1 U10025 ( .A(n8568), .ZN(n9496) );
  OAI22_X1 U10026 ( .A1(n8574), .A2(s_data_in_f[4]), .B1(\fmem_data[18][4] ), 
        .B2(n8573), .ZN(n8569) );
  INV_X1 U10027 ( .A(n8569), .ZN(n9497) );
  OAI22_X1 U10028 ( .A1(n8574), .A2(s_data_in_f[3]), .B1(\fmem_data[18][3] ), 
        .B2(n8573), .ZN(n8570) );
  INV_X1 U10029 ( .A(n8570), .ZN(n9498) );
  OAI22_X1 U10030 ( .A1(n8574), .A2(s_data_in_f[2]), .B1(\fmem_data[18][2] ), 
        .B2(n8573), .ZN(n8571) );
  INV_X1 U10031 ( .A(n8571), .ZN(n9499) );
  OAI22_X1 U10032 ( .A1(n8574), .A2(s_data_in_f[1]), .B1(\fmem_data[18][1] ), 
        .B2(n8573), .ZN(n8572) );
  INV_X1 U10033 ( .A(n8572), .ZN(n9500) );
  OAI22_X1 U10034 ( .A1(n8574), .A2(s_data_in_f[0]), .B1(\fmem_data[18][0] ), 
        .B2(n8573), .ZN(n8575) );
  INV_X1 U10035 ( .A(n8575), .ZN(n9501) );
  OAI22_X1 U10036 ( .A1(n8584), .A2(s_data_in_f[7]), .B1(\fmem_data[17][7] ), 
        .B2(n8583), .ZN(n8576) );
  INV_X1 U10037 ( .A(n8576), .ZN(n9502) );
  OAI22_X1 U10038 ( .A1(n8584), .A2(s_data_in_f[6]), .B1(\fmem_data[17][6] ), 
        .B2(n8583), .ZN(n8577) );
  INV_X1 U10039 ( .A(n8577), .ZN(n9503) );
  OAI22_X1 U10040 ( .A1(n8584), .A2(s_data_in_f[5]), .B1(\fmem_data[17][5] ), 
        .B2(n8583), .ZN(n8578) );
  INV_X1 U10041 ( .A(n8578), .ZN(n9504) );
  OAI22_X1 U10042 ( .A1(n8584), .A2(s_data_in_f[4]), .B1(\fmem_data[17][4] ), 
        .B2(n8583), .ZN(n8579) );
  INV_X1 U10043 ( .A(n8579), .ZN(n9505) );
  OAI22_X1 U10044 ( .A1(n8584), .A2(s_data_in_f[3]), .B1(\fmem_data[17][3] ), 
        .B2(n8583), .ZN(n8580) );
  INV_X1 U10045 ( .A(n8580), .ZN(n9506) );
  OAI22_X1 U10046 ( .A1(n8584), .A2(s_data_in_f[2]), .B1(\fmem_data[17][2] ), 
        .B2(n8583), .ZN(n8581) );
  INV_X1 U10047 ( .A(n8581), .ZN(n9507) );
  OAI22_X1 U10048 ( .A1(n8584), .A2(s_data_in_f[1]), .B1(\fmem_data[17][1] ), 
        .B2(n8583), .ZN(n8582) );
  INV_X1 U10049 ( .A(n8582), .ZN(n9508) );
  OAI22_X1 U10050 ( .A1(n8584), .A2(s_data_in_f[0]), .B1(\fmem_data[17][0] ), 
        .B2(n8583), .ZN(n8585) );
  INV_X1 U10051 ( .A(n8585), .ZN(n9509) );
  OAI22_X1 U10052 ( .A1(n8595), .A2(s_data_in_f[7]), .B1(\fmem_data[16][7] ), 
        .B2(n8594), .ZN(n8587) );
  INV_X1 U10053 ( .A(n8587), .ZN(n9510) );
  OAI22_X1 U10054 ( .A1(n8595), .A2(s_data_in_f[6]), .B1(\fmem_data[16][6] ), 
        .B2(n8594), .ZN(n8588) );
  INV_X1 U10055 ( .A(n8588), .ZN(n9511) );
  OAI22_X1 U10056 ( .A1(n8595), .A2(s_data_in_f[5]), .B1(\fmem_data[16][5] ), 
        .B2(n8594), .ZN(n8589) );
  INV_X1 U10057 ( .A(n8589), .ZN(n9512) );
  OAI22_X1 U10058 ( .A1(n8595), .A2(s_data_in_f[4]), .B1(\fmem_data[16][4] ), 
        .B2(n8594), .ZN(n8590) );
  INV_X1 U10059 ( .A(n8590), .ZN(n9513) );
  OAI22_X1 U10060 ( .A1(n8595), .A2(s_data_in_f[3]), .B1(\fmem_data[16][3] ), 
        .B2(n8594), .ZN(n8591) );
  INV_X1 U10061 ( .A(n8591), .ZN(n9514) );
  OAI22_X1 U10062 ( .A1(n8595), .A2(s_data_in_f[2]), .B1(\fmem_data[16][2] ), 
        .B2(n8594), .ZN(n8592) );
  INV_X1 U10063 ( .A(n8592), .ZN(n9515) );
  OAI22_X1 U10064 ( .A1(n8595), .A2(s_data_in_f[1]), .B1(\fmem_data[16][1] ), 
        .B2(n8594), .ZN(n8593) );
  INV_X1 U10065 ( .A(n8593), .ZN(n9516) );
  OAI22_X1 U10066 ( .A1(n8595), .A2(s_data_in_f[0]), .B1(\fmem_data[16][0] ), 
        .B2(n8594), .ZN(n8596) );
  INV_X1 U10067 ( .A(n8596), .ZN(n9517) );
  NOR2_X1 U10068 ( .A1(fmem_addr[4]), .A2(n8772), .ZN(n8677) );
  OAI22_X1 U10069 ( .A1(n8768), .A2(s_data_in_f[7]), .B1(\fmem_data[15][7] ), 
        .B2(n8604), .ZN(n8597) );
  INV_X1 U10070 ( .A(n8597), .ZN(n9518) );
  OAI22_X1 U10071 ( .A1(n8768), .A2(s_data_in_f[6]), .B1(\fmem_data[15][6] ), 
        .B2(n8604), .ZN(n8598) );
  INV_X1 U10072 ( .A(n8598), .ZN(n9519) );
  OAI22_X1 U10073 ( .A1(n8768), .A2(s_data_in_f[5]), .B1(\fmem_data[15][5] ), 
        .B2(n8604), .ZN(n8599) );
  INV_X1 U10074 ( .A(n8599), .ZN(n9520) );
  OAI22_X1 U10075 ( .A1(n8768), .A2(s_data_in_f[4]), .B1(\fmem_data[15][4] ), 
        .B2(n8604), .ZN(n8600) );
  INV_X1 U10076 ( .A(n8600), .ZN(n9521) );
  OAI22_X1 U10077 ( .A1(n8768), .A2(s_data_in_f[3]), .B1(\fmem_data[15][3] ), 
        .B2(n8604), .ZN(n8601) );
  INV_X1 U10078 ( .A(n8601), .ZN(n9522) );
  OAI22_X1 U10079 ( .A1(n8768), .A2(s_data_in_f[2]), .B1(\fmem_data[15][2] ), 
        .B2(n8604), .ZN(n8602) );
  INV_X1 U10080 ( .A(n8602), .ZN(n9523) );
  OAI22_X1 U10081 ( .A1(n8768), .A2(s_data_in_f[1]), .B1(\fmem_data[15][1] ), 
        .B2(n8604), .ZN(n8603) );
  INV_X1 U10082 ( .A(n8603), .ZN(n9524) );
  OAI22_X1 U10083 ( .A1(n8768), .A2(s_data_in_f[0]), .B1(\fmem_data[15][0] ), 
        .B2(n8604), .ZN(n8605) );
  INV_X1 U10084 ( .A(n8605), .ZN(n9525) );
  OAI22_X1 U10085 ( .A1(n8614), .A2(s_data_in_f[7]), .B1(\fmem_data[14][7] ), 
        .B2(n8613), .ZN(n8606) );
  INV_X1 U10086 ( .A(n8606), .ZN(n9526) );
  OAI22_X1 U10087 ( .A1(n8614), .A2(s_data_in_f[6]), .B1(\fmem_data[14][6] ), 
        .B2(n8613), .ZN(n8607) );
  INV_X1 U10088 ( .A(n8607), .ZN(n9527) );
  OAI22_X1 U10089 ( .A1(n8614), .A2(s_data_in_f[5]), .B1(\fmem_data[14][5] ), 
        .B2(n8613), .ZN(n8608) );
  INV_X1 U10090 ( .A(n8608), .ZN(n9528) );
  OAI22_X1 U10091 ( .A1(n8614), .A2(s_data_in_f[4]), .B1(\fmem_data[14][4] ), 
        .B2(n8613), .ZN(n8609) );
  INV_X1 U10092 ( .A(n8609), .ZN(n9529) );
  OAI22_X1 U10093 ( .A1(n8614), .A2(s_data_in_f[3]), .B1(\fmem_data[14][3] ), 
        .B2(n8613), .ZN(n8610) );
  INV_X1 U10094 ( .A(n8610), .ZN(n9530) );
  OAI22_X1 U10095 ( .A1(n8614), .A2(s_data_in_f[2]), .B1(\fmem_data[14][2] ), 
        .B2(n8613), .ZN(n8611) );
  INV_X1 U10096 ( .A(n8611), .ZN(n9531) );
  OAI22_X1 U10097 ( .A1(n8614), .A2(s_data_in_f[1]), .B1(\fmem_data[14][1] ), 
        .B2(n8613), .ZN(n8612) );
  INV_X1 U10098 ( .A(n8612), .ZN(n9532) );
  OAI22_X1 U10099 ( .A1(n8614), .A2(s_data_in_f[0]), .B1(\fmem_data[14][0] ), 
        .B2(n8613), .ZN(n8615) );
  INV_X1 U10100 ( .A(n8615), .ZN(n9533) );
  OAI22_X1 U10101 ( .A1(n8624), .A2(s_data_in_f[7]), .B1(\fmem_data[13][7] ), 
        .B2(n8623), .ZN(n8616) );
  INV_X1 U10102 ( .A(n8616), .ZN(n9534) );
  OAI22_X1 U10103 ( .A1(n8624), .A2(s_data_in_f[6]), .B1(\fmem_data[13][6] ), 
        .B2(n8623), .ZN(n8617) );
  INV_X1 U10104 ( .A(n8617), .ZN(n9535) );
  OAI22_X1 U10105 ( .A1(n8624), .A2(s_data_in_f[5]), .B1(\fmem_data[13][5] ), 
        .B2(n8623), .ZN(n8618) );
  INV_X1 U10106 ( .A(n8618), .ZN(n9536) );
  OAI22_X1 U10107 ( .A1(n8624), .A2(s_data_in_f[4]), .B1(\fmem_data[13][4] ), 
        .B2(n8623), .ZN(n8619) );
  INV_X1 U10108 ( .A(n8619), .ZN(n9537) );
  OAI22_X1 U10109 ( .A1(n8624), .A2(s_data_in_f[3]), .B1(\fmem_data[13][3] ), 
        .B2(n8623), .ZN(n8620) );
  INV_X1 U10110 ( .A(n8620), .ZN(n9538) );
  OAI22_X1 U10111 ( .A1(n8624), .A2(s_data_in_f[2]), .B1(\fmem_data[13][2] ), 
        .B2(n8623), .ZN(n8621) );
  INV_X1 U10112 ( .A(n8621), .ZN(n9539) );
  OAI22_X1 U10113 ( .A1(n8624), .A2(s_data_in_f[1]), .B1(\fmem_data[13][1] ), 
        .B2(n8623), .ZN(n8622) );
  INV_X1 U10114 ( .A(n8622), .ZN(n9540) );
  OAI22_X1 U10115 ( .A1(n8624), .A2(s_data_in_f[0]), .B1(\fmem_data[13][0] ), 
        .B2(n8623), .ZN(n8625) );
  INV_X1 U10116 ( .A(n8625), .ZN(n9541) );
  OAI22_X1 U10117 ( .A1(n8634), .A2(s_data_in_f[7]), .B1(\fmem_data[12][7] ), 
        .B2(n8633), .ZN(n8626) );
  INV_X1 U10118 ( .A(n8626), .ZN(n9542) );
  OAI22_X1 U10119 ( .A1(n8634), .A2(s_data_in_f[6]), .B1(\fmem_data[12][6] ), 
        .B2(n8633), .ZN(n8627) );
  INV_X1 U10120 ( .A(n8627), .ZN(n9543) );
  OAI22_X1 U10121 ( .A1(n8634), .A2(s_data_in_f[5]), .B1(\fmem_data[12][5] ), 
        .B2(n8633), .ZN(n8628) );
  INV_X1 U10122 ( .A(n8628), .ZN(n9544) );
  OAI22_X1 U10123 ( .A1(n8634), .A2(s_data_in_f[4]), .B1(\fmem_data[12][4] ), 
        .B2(n8633), .ZN(n8629) );
  INV_X1 U10124 ( .A(n8629), .ZN(n9545) );
  OAI22_X1 U10125 ( .A1(n8634), .A2(s_data_in_f[3]), .B1(\fmem_data[12][3] ), 
        .B2(n8633), .ZN(n8630) );
  INV_X1 U10126 ( .A(n8630), .ZN(n9546) );
  OAI22_X1 U10127 ( .A1(n8634), .A2(s_data_in_f[2]), .B1(\fmem_data[12][2] ), 
        .B2(n8633), .ZN(n8631) );
  INV_X1 U10128 ( .A(n8631), .ZN(n9547) );
  OAI22_X1 U10129 ( .A1(n8634), .A2(s_data_in_f[1]), .B1(\fmem_data[12][1] ), 
        .B2(n8633), .ZN(n8632) );
  INV_X1 U10130 ( .A(n8632), .ZN(n9548) );
  OAI22_X1 U10131 ( .A1(n8634), .A2(s_data_in_f[0]), .B1(\fmem_data[12][0] ), 
        .B2(n8633), .ZN(n8635) );
  INV_X1 U10132 ( .A(n8635), .ZN(n9549) );
  OAI22_X1 U10133 ( .A1(n8644), .A2(s_data_in_f[7]), .B1(\fmem_data[11][7] ), 
        .B2(n8643), .ZN(n8636) );
  INV_X1 U10134 ( .A(n8636), .ZN(n9550) );
  OAI22_X1 U10135 ( .A1(n8644), .A2(s_data_in_f[6]), .B1(\fmem_data[11][6] ), 
        .B2(n8643), .ZN(n8637) );
  INV_X1 U10136 ( .A(n8637), .ZN(n9551) );
  OAI22_X1 U10137 ( .A1(n8644), .A2(s_data_in_f[5]), .B1(\fmem_data[11][5] ), 
        .B2(n8643), .ZN(n8638) );
  INV_X1 U10138 ( .A(n8638), .ZN(n9552) );
  OAI22_X1 U10139 ( .A1(n8644), .A2(s_data_in_f[4]), .B1(\fmem_data[11][4] ), 
        .B2(n8643), .ZN(n8639) );
  INV_X1 U10140 ( .A(n8639), .ZN(n9553) );
  OAI22_X1 U10141 ( .A1(n8644), .A2(s_data_in_f[3]), .B1(\fmem_data[11][3] ), 
        .B2(n8643), .ZN(n8640) );
  INV_X1 U10142 ( .A(n8640), .ZN(n9554) );
  OAI22_X1 U10143 ( .A1(n8644), .A2(s_data_in_f[2]), .B1(\fmem_data[11][2] ), 
        .B2(n8643), .ZN(n8641) );
  INV_X1 U10144 ( .A(n8641), .ZN(n9555) );
  OAI22_X1 U10145 ( .A1(n8644), .A2(s_data_in_f[1]), .B1(\fmem_data[11][1] ), 
        .B2(n8643), .ZN(n8642) );
  INV_X1 U10146 ( .A(n8642), .ZN(n9556) );
  OAI22_X1 U10147 ( .A1(n8644), .A2(s_data_in_f[0]), .B1(\fmem_data[11][0] ), 
        .B2(n8643), .ZN(n8645) );
  INV_X1 U10148 ( .A(n8645), .ZN(n9557) );
  OAI22_X1 U10149 ( .A1(n8654), .A2(s_data_in_f[7]), .B1(\fmem_data[10][7] ), 
        .B2(n8653), .ZN(n8646) );
  INV_X1 U10150 ( .A(n8646), .ZN(n9558) );
  OAI22_X1 U10151 ( .A1(n8654), .A2(s_data_in_f[6]), .B1(\fmem_data[10][6] ), 
        .B2(n8653), .ZN(n8647) );
  INV_X1 U10152 ( .A(n8647), .ZN(n9559) );
  OAI22_X1 U10153 ( .A1(n8654), .A2(s_data_in_f[5]), .B1(\fmem_data[10][5] ), 
        .B2(n8653), .ZN(n8648) );
  INV_X1 U10154 ( .A(n8648), .ZN(n9560) );
  OAI22_X1 U10155 ( .A1(n8654), .A2(s_data_in_f[4]), .B1(\fmem_data[10][4] ), 
        .B2(n8653), .ZN(n8649) );
  INV_X1 U10156 ( .A(n8649), .ZN(n9561) );
  OAI22_X1 U10157 ( .A1(n8654), .A2(s_data_in_f[3]), .B1(\fmem_data[10][3] ), 
        .B2(n8653), .ZN(n8650) );
  INV_X1 U10158 ( .A(n8650), .ZN(n9562) );
  OAI22_X1 U10159 ( .A1(n8654), .A2(s_data_in_f[2]), .B1(\fmem_data[10][2] ), 
        .B2(n8653), .ZN(n8651) );
  INV_X1 U10160 ( .A(n8651), .ZN(n9563) );
  OAI22_X1 U10161 ( .A1(n8654), .A2(s_data_in_f[1]), .B1(\fmem_data[10][1] ), 
        .B2(n8653), .ZN(n8652) );
  INV_X1 U10162 ( .A(n8652), .ZN(n9564) );
  OAI22_X1 U10163 ( .A1(n8654), .A2(s_data_in_f[0]), .B1(\fmem_data[10][0] ), 
        .B2(n8653), .ZN(n8655) );
  INV_X1 U10164 ( .A(n8655), .ZN(n9565) );
  OAI22_X1 U10165 ( .A1(n8664), .A2(s_data_in_f[7]), .B1(\fmem_data[9][7] ), 
        .B2(n8663), .ZN(n8656) );
  INV_X1 U10166 ( .A(n8656), .ZN(n9566) );
  OAI22_X1 U10167 ( .A1(n8664), .A2(s_data_in_f[6]), .B1(\fmem_data[9][6] ), 
        .B2(n8663), .ZN(n8657) );
  INV_X1 U10168 ( .A(n8657), .ZN(n9567) );
  OAI22_X1 U10169 ( .A1(n8664), .A2(s_data_in_f[5]), .B1(\fmem_data[9][5] ), 
        .B2(n8663), .ZN(n8658) );
  INV_X1 U10170 ( .A(n8658), .ZN(n9568) );
  OAI22_X1 U10171 ( .A1(n8664), .A2(s_data_in_f[4]), .B1(\fmem_data[9][4] ), 
        .B2(n8663), .ZN(n8659) );
  INV_X1 U10172 ( .A(n8659), .ZN(n9569) );
  OAI22_X1 U10173 ( .A1(n8664), .A2(s_data_in_f[3]), .B1(\fmem_data[9][3] ), 
        .B2(n8663), .ZN(n8660) );
  INV_X1 U10174 ( .A(n8660), .ZN(n9570) );
  OAI22_X1 U10175 ( .A1(n8664), .A2(s_data_in_f[2]), .B1(\fmem_data[9][2] ), 
        .B2(n8663), .ZN(n8661) );
  INV_X1 U10176 ( .A(n8661), .ZN(n9571) );
  OAI22_X1 U10177 ( .A1(n8664), .A2(s_data_in_f[1]), .B1(\fmem_data[9][1] ), 
        .B2(n8663), .ZN(n8662) );
  INV_X1 U10178 ( .A(n8662), .ZN(n9572) );
  OAI22_X1 U10179 ( .A1(n8664), .A2(s_data_in_f[0]), .B1(\fmem_data[9][0] ), 
        .B2(n8663), .ZN(n8665) );
  INV_X1 U10180 ( .A(n8665), .ZN(n9573) );
  OAI22_X1 U10181 ( .A1(n8675), .A2(s_data_in_f[7]), .B1(\fmem_data[8][7] ), 
        .B2(n8674), .ZN(n8667) );
  INV_X1 U10182 ( .A(n8667), .ZN(n9574) );
  OAI22_X1 U10183 ( .A1(n8675), .A2(s_data_in_f[6]), .B1(\fmem_data[8][6] ), 
        .B2(n8674), .ZN(n8668) );
  INV_X1 U10184 ( .A(n8668), .ZN(n9575) );
  OAI22_X1 U10185 ( .A1(n8675), .A2(s_data_in_f[5]), .B1(\fmem_data[8][5] ), 
        .B2(n8674), .ZN(n8669) );
  INV_X1 U10186 ( .A(n8669), .ZN(n9576) );
  OAI22_X1 U10187 ( .A1(n8675), .A2(s_data_in_f[4]), .B1(\fmem_data[8][4] ), 
        .B2(n8674), .ZN(n8670) );
  INV_X1 U10188 ( .A(n8670), .ZN(n9577) );
  OAI22_X1 U10189 ( .A1(n8675), .A2(s_data_in_f[3]), .B1(\fmem_data[8][3] ), 
        .B2(n8674), .ZN(n8671) );
  INV_X1 U10190 ( .A(n8671), .ZN(n9578) );
  OAI22_X1 U10191 ( .A1(n8675), .A2(s_data_in_f[2]), .B1(\fmem_data[8][2] ), 
        .B2(n8674), .ZN(n8672) );
  INV_X1 U10192 ( .A(n8672), .ZN(n9579) );
  OAI22_X1 U10193 ( .A1(n8675), .A2(s_data_in_f[1]), .B1(\fmem_data[8][1] ), 
        .B2(n8674), .ZN(n8673) );
  INV_X1 U10194 ( .A(n8673), .ZN(n9580) );
  OAI22_X1 U10195 ( .A1(n8675), .A2(s_data_in_f[0]), .B1(\fmem_data[8][0] ), 
        .B2(n8674), .ZN(n8676) );
  INV_X1 U10196 ( .A(n8676), .ZN(n9581) );
  OAI22_X1 U10197 ( .A1(n8686), .A2(s_data_in_f[7]), .B1(\fmem_data[7][7] ), 
        .B2(n8685), .ZN(n8678) );
  INV_X1 U10198 ( .A(n8678), .ZN(n9582) );
  OAI22_X1 U10199 ( .A1(n8686), .A2(s_data_in_f[6]), .B1(\fmem_data[7][6] ), 
        .B2(n8685), .ZN(n8679) );
  INV_X1 U10200 ( .A(n8679), .ZN(n9583) );
  OAI22_X1 U10201 ( .A1(n8686), .A2(s_data_in_f[5]), .B1(\fmem_data[7][5] ), 
        .B2(n8685), .ZN(n8680) );
  INV_X1 U10202 ( .A(n8680), .ZN(n9584) );
  OAI22_X1 U10203 ( .A1(n8686), .A2(s_data_in_f[4]), .B1(\fmem_data[7][4] ), 
        .B2(n8685), .ZN(n8681) );
  INV_X1 U10204 ( .A(n8681), .ZN(n9585) );
  OAI22_X1 U10205 ( .A1(n8686), .A2(s_data_in_f[3]), .B1(\fmem_data[7][3] ), 
        .B2(n8685), .ZN(n8682) );
  INV_X1 U10206 ( .A(n8682), .ZN(n9586) );
  OAI22_X1 U10207 ( .A1(n8686), .A2(s_data_in_f[2]), .B1(\fmem_data[7][2] ), 
        .B2(n8685), .ZN(n8683) );
  INV_X1 U10208 ( .A(n8683), .ZN(n9587) );
  OAI22_X1 U10209 ( .A1(n8686), .A2(s_data_in_f[1]), .B1(\fmem_data[7][1] ), 
        .B2(n8685), .ZN(n8684) );
  INV_X1 U10210 ( .A(n8684), .ZN(n9588) );
  OAI22_X1 U10211 ( .A1(n8686), .A2(s_data_in_f[0]), .B1(\fmem_data[7][0] ), 
        .B2(n8685), .ZN(n8687) );
  INV_X1 U10212 ( .A(n8687), .ZN(n9589) );
  OAI22_X1 U10213 ( .A1(n8697), .A2(s_data_in_f[7]), .B1(\fmem_data[6][7] ), 
        .B2(n8696), .ZN(n8689) );
  INV_X1 U10214 ( .A(n8689), .ZN(n9590) );
  OAI22_X1 U10215 ( .A1(n8697), .A2(s_data_in_f[6]), .B1(\fmem_data[6][6] ), 
        .B2(n8696), .ZN(n8690) );
  INV_X1 U10216 ( .A(n8690), .ZN(n9591) );
  OAI22_X1 U10217 ( .A1(n8697), .A2(s_data_in_f[5]), .B1(\fmem_data[6][5] ), 
        .B2(n8696), .ZN(n8691) );
  INV_X1 U10218 ( .A(n8691), .ZN(n9592) );
  OAI22_X1 U10219 ( .A1(n8697), .A2(s_data_in_f[4]), .B1(\fmem_data[6][4] ), 
        .B2(n8696), .ZN(n8692) );
  INV_X1 U10220 ( .A(n8692), .ZN(n9593) );
  OAI22_X1 U10221 ( .A1(n8697), .A2(s_data_in_f[3]), .B1(\fmem_data[6][3] ), 
        .B2(n8696), .ZN(n8693) );
  INV_X1 U10222 ( .A(n8693), .ZN(n9594) );
  OAI22_X1 U10223 ( .A1(n8697), .A2(s_data_in_f[2]), .B1(\fmem_data[6][2] ), 
        .B2(n8696), .ZN(n8694) );
  INV_X1 U10224 ( .A(n8694), .ZN(n9595) );
  OAI22_X1 U10225 ( .A1(n8697), .A2(s_data_in_f[1]), .B1(\fmem_data[6][1] ), 
        .B2(n8696), .ZN(n8695) );
  INV_X1 U10226 ( .A(n8695), .ZN(n9596) );
  OAI22_X1 U10227 ( .A1(n8697), .A2(s_data_in_f[0]), .B1(\fmem_data[6][0] ), 
        .B2(n8696), .ZN(n8698) );
  INV_X1 U10228 ( .A(n8698), .ZN(n9597) );
  OAI22_X1 U10229 ( .A1(n8708), .A2(s_data_in_f[7]), .B1(\fmem_data[5][7] ), 
        .B2(n8707), .ZN(n8700) );
  INV_X1 U10230 ( .A(n8700), .ZN(n9598) );
  OAI22_X1 U10231 ( .A1(n8708), .A2(s_data_in_f[6]), .B1(\fmem_data[5][6] ), 
        .B2(n8707), .ZN(n8701) );
  INV_X1 U10232 ( .A(n8701), .ZN(n9599) );
  OAI22_X1 U10233 ( .A1(n8708), .A2(s_data_in_f[5]), .B1(\fmem_data[5][5] ), 
        .B2(n8707), .ZN(n8702) );
  INV_X1 U10234 ( .A(n8702), .ZN(n9600) );
  OAI22_X1 U10235 ( .A1(n8708), .A2(s_data_in_f[4]), .B1(\fmem_data[5][4] ), 
        .B2(n8707), .ZN(n8703) );
  INV_X1 U10236 ( .A(n8703), .ZN(n9601) );
  OAI22_X1 U10237 ( .A1(n8708), .A2(s_data_in_f[3]), .B1(\fmem_data[5][3] ), 
        .B2(n8707), .ZN(n8704) );
  INV_X1 U10238 ( .A(n8704), .ZN(n9602) );
  OAI22_X1 U10239 ( .A1(n8708), .A2(s_data_in_f[2]), .B1(\fmem_data[5][2] ), 
        .B2(n8707), .ZN(n8705) );
  INV_X1 U10240 ( .A(n8705), .ZN(n9603) );
  OAI22_X1 U10241 ( .A1(n8708), .A2(s_data_in_f[1]), .B1(\fmem_data[5][1] ), 
        .B2(n8707), .ZN(n8706) );
  INV_X1 U10242 ( .A(n8706), .ZN(n9604) );
  OAI22_X1 U10243 ( .A1(n8708), .A2(s_data_in_f[0]), .B1(\fmem_data[5][0] ), 
        .B2(n8707), .ZN(n8709) );
  INV_X1 U10244 ( .A(n8709), .ZN(n9605) );
  OAI22_X1 U10245 ( .A1(n8719), .A2(s_data_in_f[7]), .B1(\fmem_data[4][7] ), 
        .B2(n8718), .ZN(n8711) );
  INV_X1 U10246 ( .A(n8711), .ZN(n9606) );
  OAI22_X1 U10247 ( .A1(n8719), .A2(s_data_in_f[6]), .B1(\fmem_data[4][6] ), 
        .B2(n8718), .ZN(n8712) );
  INV_X1 U10248 ( .A(n8712), .ZN(n9607) );
  OAI22_X1 U10249 ( .A1(n8719), .A2(s_data_in_f[5]), .B1(\fmem_data[4][5] ), 
        .B2(n8718), .ZN(n8713) );
  INV_X1 U10250 ( .A(n8713), .ZN(n9608) );
  OAI22_X1 U10251 ( .A1(n8719), .A2(s_data_in_f[4]), .B1(\fmem_data[4][4] ), 
        .B2(n8718), .ZN(n8714) );
  INV_X1 U10252 ( .A(n8714), .ZN(n9609) );
  OAI22_X1 U10253 ( .A1(n8719), .A2(s_data_in_f[3]), .B1(\fmem_data[4][3] ), 
        .B2(n8718), .ZN(n8715) );
  INV_X1 U10254 ( .A(n8715), .ZN(n9610) );
  OAI22_X1 U10255 ( .A1(n8719), .A2(s_data_in_f[2]), .B1(\fmem_data[4][2] ), 
        .B2(n8718), .ZN(n8716) );
  INV_X1 U10256 ( .A(n8716), .ZN(n9611) );
  OAI22_X1 U10257 ( .A1(n8719), .A2(s_data_in_f[1]), .B1(\fmem_data[4][1] ), 
        .B2(n8718), .ZN(n8717) );
  INV_X1 U10258 ( .A(n8717), .ZN(n9612) );
  OAI22_X1 U10259 ( .A1(n8719), .A2(s_data_in_f[0]), .B1(\fmem_data[4][0] ), 
        .B2(n8718), .ZN(n8720) );
  INV_X1 U10260 ( .A(n8720), .ZN(n9613) );
  OAI22_X1 U10261 ( .A1(n8729), .A2(s_data_in_f[7]), .B1(\fmem_data[3][7] ), 
        .B2(n8728), .ZN(n8721) );
  INV_X1 U10262 ( .A(n8721), .ZN(n9614) );
  OAI22_X1 U10263 ( .A1(n8729), .A2(s_data_in_f[6]), .B1(\fmem_data[3][6] ), 
        .B2(n8728), .ZN(n8722) );
  INV_X1 U10264 ( .A(n8722), .ZN(n9615) );
  OAI22_X1 U10265 ( .A1(n8729), .A2(s_data_in_f[5]), .B1(\fmem_data[3][5] ), 
        .B2(n8728), .ZN(n8723) );
  INV_X1 U10266 ( .A(n8723), .ZN(n9616) );
  OAI22_X1 U10267 ( .A1(n8729), .A2(s_data_in_f[4]), .B1(\fmem_data[3][4] ), 
        .B2(n8728), .ZN(n8724) );
  INV_X1 U10268 ( .A(n8724), .ZN(n9617) );
  OAI22_X1 U10269 ( .A1(n8729), .A2(s_data_in_f[3]), .B1(\fmem_data[3][3] ), 
        .B2(n8728), .ZN(n8725) );
  INV_X1 U10270 ( .A(n8725), .ZN(n9618) );
  OAI22_X1 U10271 ( .A1(n8729), .A2(s_data_in_f[2]), .B1(\fmem_data[3][2] ), 
        .B2(n8728), .ZN(n8726) );
  INV_X1 U10272 ( .A(n8726), .ZN(n9619) );
  OAI22_X1 U10273 ( .A1(n8729), .A2(s_data_in_f[1]), .B1(\fmem_data[3][1] ), 
        .B2(n8728), .ZN(n8727) );
  INV_X1 U10274 ( .A(n8727), .ZN(n9620) );
  OAI22_X1 U10275 ( .A1(n8729), .A2(s_data_in_f[0]), .B1(\fmem_data[3][0] ), 
        .B2(n8728), .ZN(n8730) );
  INV_X1 U10276 ( .A(n8730), .ZN(n9621) );
  OAI22_X1 U10277 ( .A1(n8740), .A2(s_data_in_f[7]), .B1(\fmem_data[2][7] ), 
        .B2(n8739), .ZN(n8732) );
  INV_X1 U10278 ( .A(n8732), .ZN(n9622) );
  OAI22_X1 U10279 ( .A1(n8740), .A2(s_data_in_f[6]), .B1(\fmem_data[2][6] ), 
        .B2(n8739), .ZN(n8733) );
  INV_X1 U10280 ( .A(n8733), .ZN(n9623) );
  OAI22_X1 U10281 ( .A1(n8740), .A2(s_data_in_f[5]), .B1(\fmem_data[2][5] ), 
        .B2(n8739), .ZN(n8734) );
  INV_X1 U10282 ( .A(n8734), .ZN(n9624) );
  OAI22_X1 U10283 ( .A1(n8740), .A2(s_data_in_f[4]), .B1(\fmem_data[2][4] ), 
        .B2(n8739), .ZN(n8735) );
  INV_X1 U10284 ( .A(n8735), .ZN(n9625) );
  OAI22_X1 U10285 ( .A1(n8740), .A2(s_data_in_f[3]), .B1(\fmem_data[2][3] ), 
        .B2(n8739), .ZN(n8736) );
  INV_X1 U10286 ( .A(n8736), .ZN(n9626) );
  OAI22_X1 U10287 ( .A1(n8740), .A2(s_data_in_f[2]), .B1(\fmem_data[2][2] ), 
        .B2(n8739), .ZN(n8737) );
  INV_X1 U10288 ( .A(n8737), .ZN(n9627) );
  OAI22_X1 U10289 ( .A1(n8740), .A2(s_data_in_f[1]), .B1(\fmem_data[2][1] ), 
        .B2(n8739), .ZN(n8738) );
  INV_X1 U10290 ( .A(n8738), .ZN(n9628) );
  OAI22_X1 U10291 ( .A1(n8740), .A2(s_data_in_f[0]), .B1(\fmem_data[2][0] ), 
        .B2(n8739), .ZN(n8741) );
  INV_X1 U10292 ( .A(n8741), .ZN(n9629) );
  OAI22_X1 U10293 ( .A1(n8751), .A2(s_data_in_f[7]), .B1(\fmem_data[1][7] ), 
        .B2(n8750), .ZN(n8743) );
  INV_X1 U10294 ( .A(n8743), .ZN(n9630) );
  OAI22_X1 U10295 ( .A1(n8751), .A2(s_data_in_f[6]), .B1(\fmem_data[1][6] ), 
        .B2(n8750), .ZN(n8744) );
  INV_X1 U10296 ( .A(n8744), .ZN(n9631) );
  OAI22_X1 U10297 ( .A1(n8751), .A2(s_data_in_f[5]), .B1(\fmem_data[1][5] ), 
        .B2(n8750), .ZN(n8745) );
  INV_X1 U10298 ( .A(n8745), .ZN(n9632) );
  OAI22_X1 U10299 ( .A1(n8751), .A2(s_data_in_f[4]), .B1(\fmem_data[1][4] ), 
        .B2(n8750), .ZN(n8746) );
  INV_X1 U10300 ( .A(n8746), .ZN(n9633) );
  OAI22_X1 U10301 ( .A1(n8751), .A2(s_data_in_f[3]), .B1(\fmem_data[1][3] ), 
        .B2(n8750), .ZN(n8747) );
  INV_X1 U10302 ( .A(n8747), .ZN(n9634) );
  OAI22_X1 U10303 ( .A1(n8751), .A2(s_data_in_f[2]), .B1(\fmem_data[1][2] ), 
        .B2(n8750), .ZN(n8748) );
  INV_X1 U10304 ( .A(n8748), .ZN(n9635) );
  OAI22_X1 U10305 ( .A1(n8751), .A2(s_data_in_f[1]), .B1(\fmem_data[1][1] ), 
        .B2(n8750), .ZN(n8749) );
  INV_X1 U10306 ( .A(n8749), .ZN(n9636) );
  OAI22_X1 U10307 ( .A1(n8751), .A2(s_data_in_f[0]), .B1(\fmem_data[1][0] ), 
        .B2(n8750), .ZN(n8752) );
  INV_X1 U10308 ( .A(n8752), .ZN(n9637) );
  OAI22_X1 U10309 ( .A1(n8763), .A2(s_data_in_f[7]), .B1(\fmem_data[0][7] ), 
        .B2(n8762), .ZN(n8755) );
  INV_X1 U10310 ( .A(n8755), .ZN(n9638) );
  OAI22_X1 U10311 ( .A1(n8763), .A2(s_data_in_f[6]), .B1(\fmem_data[0][6] ), 
        .B2(n8762), .ZN(n8756) );
  INV_X1 U10312 ( .A(n8756), .ZN(n9639) );
  OAI22_X1 U10313 ( .A1(n8763), .A2(s_data_in_f[5]), .B1(\fmem_data[0][5] ), 
        .B2(n8762), .ZN(n8757) );
  INV_X1 U10314 ( .A(n8757), .ZN(n9640) );
  OAI22_X1 U10315 ( .A1(n8763), .A2(s_data_in_f[4]), .B1(\fmem_data[0][4] ), 
        .B2(n8762), .ZN(n8758) );
  INV_X1 U10316 ( .A(n8758), .ZN(n9641) );
  OAI22_X1 U10317 ( .A1(n8763), .A2(s_data_in_f[3]), .B1(\fmem_data[0][3] ), 
        .B2(n8762), .ZN(n8759) );
  INV_X1 U10318 ( .A(n8759), .ZN(n9642) );
  OAI22_X1 U10319 ( .A1(n8763), .A2(s_data_in_f[2]), .B1(\fmem_data[0][2] ), 
        .B2(n8762), .ZN(n8760) );
  INV_X1 U10320 ( .A(n8760), .ZN(n9643) );
  OAI22_X1 U10321 ( .A1(n8763), .A2(s_data_in_f[1]), .B1(\fmem_data[0][1] ), 
        .B2(n8762), .ZN(n8761) );
  INV_X1 U10322 ( .A(n8761), .ZN(n9644) );
  OAI22_X1 U10323 ( .A1(n8763), .A2(s_data_in_f[0]), .B1(\fmem_data[0][0] ), 
        .B2(n8762), .ZN(n8764) );
  INV_X1 U10324 ( .A(n8764), .ZN(n9645) );
  NAND2_X1 U10325 ( .A1(n8778), .A2(n3444), .ZN(n8769) );
  AOI21_X1 U10326 ( .B1(n8845), .B2(n8768), .A(n8769), .ZN(n3397) );
  INV_X1 U10327 ( .A(n8769), .ZN(n8765) );
  NAND2_X1 U10328 ( .A1(n8771), .A2(n8765), .ZN(n8776) );
  OAI22_X1 U10329 ( .A1(n8766), .A2(n8776), .B1(n8809), .B2(n8769), .ZN(n8767)
         );
  AND2_X1 U10330 ( .A1(n8768), .A2(n8767), .ZN(n3396) );
  OAI33_X1 U10331 ( .A1(n8771), .A2(n8805), .A3(n8770), .B1(n8772), .B2(n8769), 
        .B3(fmem_addr[0]), .ZN(n3395) );
  NAND2_X1 U10332 ( .A1(fmem_addr[0]), .A2(n8771), .ZN(n8774) );
  NAND2_X1 U10333 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n8773) );
  OAI21_X1 U10334 ( .B1(n8773), .B2(n8772), .A(n8778), .ZN(n8777) );
  AOI21_X1 U10335 ( .B1(n8808), .B2(n8774), .A(n8777), .ZN(n3394) );
  OAI22_X1 U10336 ( .A1(n8804), .A2(n8777), .B1(n8776), .B2(n8775), .ZN(n3393)
         );
  OAI21_X1 U10337 ( .B1(n8779), .B2(n8811), .A(n8778), .ZN(n3392) );
  OAI21_X1 U10338 ( .B1(n8781), .B2(n8810), .A(n8780), .ZN(n8782) );
  NAND2_X1 U10339 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  AOI22_X1 U10340 ( .A1(\ctrl_inst/pline_cntr [1]), .A2(n8785), .B1(n8784), 
        .B2(n8840), .ZN(n3120) );
endmodule

