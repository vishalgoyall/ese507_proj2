
module conv_8_4 ( clk, reset, s_valid_x, s_valid_f, m_ready_y, s_data_in_x, 
        s_data_in_f, s_ready_f, s_ready_x, m_valid_y, m_data_out_y );
  input [7:0] s_data_in_x;
  input [7:0] s_data_in_f;
  output [17:0] m_data_out_y;
  input clk, reset, s_valid_x, s_valid_f, m_ready_y;
  output s_ready_f, s_ready_x, m_valid_y;
  wire   conv_done, conv_pre_start, N6, \xmem_inst/N20 , \xmem_inst/N19 ,
         \xmem_inst/N18 , \xmem_inst/N17 , \xmem_inst/N16 , \xmem_inst/N15 ,
         \xmem_inst/N14 , \xmem_inst/N13 , \xmem_inst/mem[7][7] ,
         \xmem_inst/mem[7][6] , \xmem_inst/mem[7][5] , \xmem_inst/mem[7][4] ,
         \xmem_inst/mem[7][3] , \xmem_inst/mem[7][2] , \xmem_inst/mem[7][1] ,
         \xmem_inst/mem[7][0] , \xmem_inst/mem[6][7] , \xmem_inst/mem[6][6] ,
         \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] , \xmem_inst/mem[6][3] ,
         \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] , \xmem_inst/mem[6][0] ,
         \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] , \xmem_inst/mem[5][5] ,
         \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] , \xmem_inst/mem[5][2] ,
         \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] , \xmem_inst/mem[4][7] ,
         \xmem_inst/mem[4][6] , \xmem_inst/mem[4][5] , \xmem_inst/mem[4][4] ,
         \xmem_inst/mem[4][3] , \xmem_inst/mem[4][2] , \xmem_inst/mem[4][1] ,
         \xmem_inst/mem[4][0] , \xmem_inst/mem[3][7] , \xmem_inst/mem[3][6] ,
         \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] , \xmem_inst/mem[3][3] ,
         \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] , \xmem_inst/mem[3][0] ,
         \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] , \xmem_inst/mem[2][5] ,
         \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] , \xmem_inst/mem[2][2] ,
         \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] , \xmem_inst/mem[1][7] ,
         \xmem_inst/mem[1][6] , \xmem_inst/mem[1][5] , \xmem_inst/mem[1][4] ,
         \xmem_inst/mem[1][3] , \xmem_inst/mem[1][2] , \xmem_inst/mem[1][1] ,
         \xmem_inst/mem[1][0] , \xmem_inst/mem[0][7] , \xmem_inst/mem[0][6] ,
         \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] , \xmem_inst/mem[0][3] ,
         \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] , \xmem_inst/mem[0][0] ,
         \fmem_inst/N13 , \fmem_inst/N11 , \fmem_inst/mem[1][7] ,
         \fmem_inst/mem[1][6] , \fmem_inst/mem[1][5] , \fmem_inst/mem[1][4] ,
         \fmem_inst/mem[1][3] , \fmem_inst/mem[1][2] , \fmem_inst/mem[1][1] ,
         \fmem_inst/mem[1][0] , \fmem_inst/mem[0][7] , \fmem_inst/mem[0][6] ,
         \fmem_inst/mem[0][5] , \fmem_inst/mem[0][4] , \fmem_inst/mem[0][3] ,
         \fmem_inst/mem[0][2] , \fmem_inst/mem[0][1] , \fmem_inst/mem[0][0] ,
         \ctrl_conv_output_inst/N71 , \ctrl_conv_output_inst/N68 ,
         \ctrl_conv_output_inst/m_pre_valid_int ,
         \ctrl_conv_output_inst/conv_start_accum ,
         \ctrl_conv_output_inst/m_pre_valid , n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, \DP_OP_61J1_122_4588/n326 , n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074;
  wire   [2:0] xmem_addr;
  wire   [7:0] xmem_data;
  wire   [1:0] fmem_addr;
  wire   [7:0] fmem_data;
  wire   [2:0] \ctrl_conv_output_inst/cnt_conv ;

  DFF_X1 \xmem_inst/data_out_reg[1]  ( .D(\xmem_inst/N19 ), .CK(clk), .Q(
        xmem_data[1]), .QN(n1030) );
  DFF_X1 \xmem_inst/data_out_reg[2]  ( .D(\xmem_inst/N18 ), .CK(clk), .Q(
        xmem_data[2]), .QN(n1029) );
  DFF_X1 \fmem_inst/data_out_reg[2]  ( .D(\fmem_inst/N13 ), .CK(clk), .Q(
        fmem_data[2]), .QN(n1032) );
  DFF_X1 \fmem_inst/data_out_reg[4]  ( .D(\fmem_inst/N11 ), .CK(clk), .Q(
        fmem_data[4]), .QN(n1034) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n344), .CK(clk), .Q(
        xmem_addr[2]), .QN(n1059) );
  DFF_X1 \ctrl_conv_output_inst/conv_start_accum_reg  ( .D(
        \ctrl_conv_output_inst/N68 ), .CK(clk), .Q(
        \ctrl_conv_output_inst/conv_start_accum ), .QN(n1073) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[1]  ( .D(n380), .CK(clk), .Q(
        fmem_addr[1]), .QN(n1064) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_int_reg  ( .D(n388), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid_int ), .QN(n1060) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[0]  ( .D(n381), .CK(clk), .Q(
        fmem_addr[0]), .QN(n1048) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_reg  ( .D(n384), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid ), .QN(n1074) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[0]  ( .D(n386), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [0]), .QN(n1061) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n346), .CK(clk), .Q(
        xmem_addr[0]), .QN(n1062) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[1]  ( .D(n385), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [1]), .QN(n1049) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[2]  ( .D(n387), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [2]), .QN(n1063) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n345), .CK(clk), .Q(
        xmem_addr[1]), .QN(n1050) );
  DFF_X1 \fmem_inst/mem_reg[2][0]  ( .D(n363), .CK(clk), .QN(n1065) );
  DFF_X1 \fmem_inst/mem_reg[2][1]  ( .D(n362), .CK(clk), .QN(n1066) );
  DFF_X1 \fmem_inst/mem_reg[2][2]  ( .D(n361), .CK(clk), .QN(n1067) );
  DFF_X1 \fmem_inst/mem_reg[2][3]  ( .D(n360), .CK(clk), .QN(n1068) );
  DFF_X1 \fmem_inst/mem_reg[2][4]  ( .D(n359), .CK(clk), .QN(n1069) );
  DFF_X1 \fmem_inst/mem_reg[2][5]  ( .D(n358), .CK(clk), .QN(n1070) );
  DFF_X1 \fmem_inst/mem_reg[2][6]  ( .D(n357), .CK(clk), .QN(n1071) );
  DFF_X1 \fmem_inst/mem_reg[2][7]  ( .D(n356), .CK(clk), .QN(n1072) );
  DFF_X1 \fmem_inst/mem_reg[3][0]  ( .D(n355), .CK(clk), .QN(n1051) );
  DFF_X1 \fmem_inst/mem_reg[3][1]  ( .D(n354), .CK(clk), .QN(n1052) );
  DFF_X1 \fmem_inst/mem_reg[3][2]  ( .D(n353), .CK(clk), .QN(n1053) );
  DFF_X1 \fmem_inst/mem_reg[3][3]  ( .D(n352), .CK(clk), .QN(n1054) );
  DFF_X1 \fmem_inst/mem_reg[3][4]  ( .D(n351), .CK(clk), .QN(n1055) );
  DFF_X1 \fmem_inst/mem_reg[3][5]  ( .D(n350), .CK(clk), .QN(n1056) );
  DFF_X1 \fmem_inst/mem_reg[3][6]  ( .D(n349), .CK(clk), .QN(n1057) );
  DFF_X1 \fmem_inst/mem_reg[3][7]  ( .D(n348), .CK(clk), .QN(n1058) );
  DFF_X1 \accum_out_reg[16]  ( .D(n262), .CK(clk), .Q(m_data_out_y[16]), .QN(
        n397) );
  DFF_X1 \fmem_inst/data_out_reg[7]  ( .D(n411), .CK(clk), .Q(n1043), .QN(
        fmem_data[7]) );
  DFF_X1 \fmem_inst/data_out_reg[5]  ( .D(n410), .CK(clk), .Q(n1031), .QN(
        fmem_data[5]) );
  DFF_X1 \fmem_inst/data_out_reg[6]  ( .D(n409), .CK(clk), .Q(n1045), .QN(
        fmem_data[6]) );
  DFF_X1 \fmem_inst/data_out_reg[3]  ( .D(n408), .CK(clk), .Q(n1035), .QN(
        fmem_data[3]) );
  DFF_X1 \fmem_inst/data_out_reg[0]  ( .D(n407), .CK(clk), .Q(n1042), .QN(
        fmem_data[0]) );
  DFF_X1 \fmem_inst/data_out_reg[1]  ( .D(n406), .CK(clk), .Q(n1033), .QN(
        \DP_OP_61J1_122_4588/n326 ) );
  DFF_X1 \accum_out_reg[15]  ( .D(n263), .CK(clk), .Q(m_data_out_y[15]), .QN(
        n1038) );
  DFF_X1 \accum_out_reg[17]  ( .D(n279), .CK(clk), .Q(m_data_out_y[17]), .QN(
        n1037) );
  DFF_X1 \accum_out_reg[13]  ( .D(n265), .CK(clk), .Q(m_data_out_y[13]), .QN(
        n1039) );
  DFF_X1 conv_pre_start_reg ( .D(N6), .CK(clk), .Q(conv_pre_start) );
  DFF_X1 \ctrl_conv_output_inst/conv_done_reg  ( .D(
        \ctrl_conv_output_inst/N71 ), .CK(clk), .Q(conv_done) );
  DFF_X1 \xmem_inst/data_out_reg[7]  ( .D(\xmem_inst/N13 ), .CK(clk), .Q(
        xmem_data[7]) );
  DFF_X1 \xmem_inst/data_out_reg[6]  ( .D(\xmem_inst/N14 ), .CK(clk), .Q(
        xmem_data[6]) );
  DFF_X1 \xmem_inst/data_out_reg[5]  ( .D(\xmem_inst/N15 ), .CK(clk), .Q(
        xmem_data[5]) );
  DFF_X1 \xmem_inst/data_out_reg[4]  ( .D(\xmem_inst/N16 ), .CK(clk), .Q(
        xmem_data[4]) );
  DFF_X1 \xmem_inst/data_out_reg[3]  ( .D(\xmem_inst/N17 ), .CK(clk), .Q(
        xmem_data[3]) );
  DFF_X1 \xmem_inst/data_out_reg[0]  ( .D(\xmem_inst/N20 ), .CK(clk), .Q(
        xmem_data[0]) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n383), .CK(clk), .Q(
        m_valid_y) );
  DFF_X1 \fmem_inst/mem_reg[0][7]  ( .D(n372), .CK(clk), .Q(
        \fmem_inst/mem[0][7] ) );
  DFF_X1 \fmem_inst/mem_reg[0][6]  ( .D(n373), .CK(clk), .Q(
        \fmem_inst/mem[0][6] ) );
  DFF_X1 \fmem_inst/mem_reg[0][5]  ( .D(n374), .CK(clk), .Q(
        \fmem_inst/mem[0][5] ) );
  DFF_X1 \fmem_inst/mem_reg[0][4]  ( .D(n375), .CK(clk), .Q(
        \fmem_inst/mem[0][4] ) );
  DFF_X1 \fmem_inst/mem_reg[0][3]  ( .D(n376), .CK(clk), .Q(
        \fmem_inst/mem[0][3] ) );
  DFF_X1 \fmem_inst/mem_reg[0][2]  ( .D(n377), .CK(clk), .Q(
        \fmem_inst/mem[0][2] ) );
  DFF_X1 \fmem_inst/mem_reg[0][1]  ( .D(n378), .CK(clk), .Q(
        \fmem_inst/mem[0][1] ) );
  DFF_X1 \fmem_inst/mem_reg[0][0]  ( .D(n379), .CK(clk), .Q(
        \fmem_inst/mem[0][0] ) );
  DFF_X1 \accum_out_reg[0]  ( .D(n278), .CK(clk), .Q(m_data_out_y[0]) );
  DFF_X1 \fmem_inst/mem_reg[1][7]  ( .D(n364), .CK(clk), .Q(
        \fmem_inst/mem[1][7] ) );
  DFF_X1 \fmem_inst/mem_reg[1][6]  ( .D(n365), .CK(clk), .Q(
        \fmem_inst/mem[1][6] ) );
  DFF_X1 \fmem_inst/mem_reg[1][5]  ( .D(n366), .CK(clk), .Q(
        \fmem_inst/mem[1][5] ) );
  DFF_X1 \fmem_inst/mem_reg[1][4]  ( .D(n367), .CK(clk), .Q(
        \fmem_inst/mem[1][4] ) );
  DFF_X1 \fmem_inst/mem_reg[1][3]  ( .D(n368), .CK(clk), .Q(
        \fmem_inst/mem[1][3] ) );
  DFF_X1 \fmem_inst/mem_reg[1][2]  ( .D(n369), .CK(clk), .Q(
        \fmem_inst/mem[1][2] ) );
  DFF_X1 \fmem_inst/mem_reg[1][1]  ( .D(n370), .CK(clk), .Q(
        \fmem_inst/mem[1][1] ) );
  DFF_X1 \fmem_inst/mem_reg[1][0]  ( .D(n371), .CK(clk), .Q(
        \fmem_inst/mem[1][0] ) );
  DFF_X1 \ctrl_fmem_write_inst/s_ready_reg  ( .D(n382), .CK(clk), .Q(s_ready_f) );
  DFF_X1 \accum_out_reg[1]  ( .D(n277), .CK(clk), .Q(m_data_out_y[1]), .QN(
        n1044) );
  DFF_X1 \accum_out_reg[2]  ( .D(n276), .CK(clk), .Q(m_data_out_y[2]) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n288), .CK(clk), .Q(
        \xmem_inst/mem[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n289), .CK(clk), .Q(
        \xmem_inst/mem[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n290), .CK(clk), .Q(
        \xmem_inst/mem[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n291), .CK(clk), .Q(
        \xmem_inst/mem[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n292), .CK(clk), .Q(
        \xmem_inst/mem[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n293), .CK(clk), .Q(
        \xmem_inst/mem[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n294), .CK(clk), .Q(
        \xmem_inst/mem[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n295), .CK(clk), .Q(
        \xmem_inst/mem[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n296), .CK(clk), .Q(
        \xmem_inst/mem[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n297), .CK(clk), .Q(
        \xmem_inst/mem[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n298), .CK(clk), .Q(
        \xmem_inst/mem[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n299), .CK(clk), .Q(
        \xmem_inst/mem[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n300), .CK(clk), .Q(
        \xmem_inst/mem[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n301), .CK(clk), .Q(
        \xmem_inst/mem[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n302), .CK(clk), .Q(
        \xmem_inst/mem[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n303), .CK(clk), .Q(
        \xmem_inst/mem[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n304), .CK(clk), .Q(
        \xmem_inst/mem[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n305), .CK(clk), .Q(
        \xmem_inst/mem[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n306), .CK(clk), .Q(
        \xmem_inst/mem[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n307), .CK(clk), .Q(
        \xmem_inst/mem[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n308), .CK(clk), .Q(
        \xmem_inst/mem[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n309), .CK(clk), .Q(
        \xmem_inst/mem[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n310), .CK(clk), .Q(
        \xmem_inst/mem[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n311), .CK(clk), .Q(
        \xmem_inst/mem[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n312), .CK(clk), .Q(
        \xmem_inst/mem[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n313), .CK(clk), .Q(
        \xmem_inst/mem[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n314), .CK(clk), .Q(
        \xmem_inst/mem[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n315), .CK(clk), .Q(
        \xmem_inst/mem[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n316), .CK(clk), .Q(
        \xmem_inst/mem[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n317), .CK(clk), .Q(
        \xmem_inst/mem[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n318), .CK(clk), .Q(
        \xmem_inst/mem[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n319), .CK(clk), .Q(
        \xmem_inst/mem[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n320), .CK(clk), .Q(
        \xmem_inst/mem[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n321), .CK(clk), .Q(
        \xmem_inst/mem[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n322), .CK(clk), .Q(
        \xmem_inst/mem[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n323), .CK(clk), .Q(
        \xmem_inst/mem[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n324), .CK(clk), .Q(
        \xmem_inst/mem[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n325), .CK(clk), .Q(
        \xmem_inst/mem[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n326), .CK(clk), .Q(
        \xmem_inst/mem[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n327), .CK(clk), .Q(
        \xmem_inst/mem[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n328), .CK(clk), .Q(
        \xmem_inst/mem[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n329), .CK(clk), .Q(
        \xmem_inst/mem[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n330), .CK(clk), .Q(
        \xmem_inst/mem[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n331), .CK(clk), .Q(
        \xmem_inst/mem[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n332), .CK(clk), .Q(
        \xmem_inst/mem[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n333), .CK(clk), .Q(
        \xmem_inst/mem[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n334), .CK(clk), .Q(
        \xmem_inst/mem[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n335), .CK(clk), .Q(
        \xmem_inst/mem[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n336), .CK(clk), .Q(
        \xmem_inst/mem[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n337), .CK(clk), .Q(
        \xmem_inst/mem[0][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n338), .CK(clk), .Q(
        \xmem_inst/mem[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n339), .CK(clk), .Q(
        \xmem_inst/mem[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n340), .CK(clk), .Q(
        \xmem_inst/mem[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n341), .CK(clk), .Q(
        \xmem_inst/mem[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n342), .CK(clk), .Q(
        \xmem_inst/mem[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n343), .CK(clk), .Q(
        \xmem_inst/mem[0][0] ) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n347), .CK(clk), .Q(s_ready_x) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n280), .CK(clk), .Q(
        \xmem_inst/mem[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n281), .CK(clk), .Q(
        \xmem_inst/mem[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n282), .CK(clk), .Q(
        \xmem_inst/mem[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n283), .CK(clk), .Q(
        \xmem_inst/mem[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n284), .CK(clk), .Q(
        \xmem_inst/mem[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n285), .CK(clk), .Q(
        \xmem_inst/mem[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n286), .CK(clk), .Q(
        \xmem_inst/mem[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n287), .CK(clk), .Q(
        \xmem_inst/mem[7][0] ) );
  DFF_X1 \accum_out_reg[3]  ( .D(n275), .CK(clk), .Q(m_data_out_y[3]) );
  DFF_X1 \accum_out_reg[4]  ( .D(n274), .CK(clk), .Q(m_data_out_y[4]), .QN(
        n1036) );
  DFF_X1 \accum_out_reg[5]  ( .D(n273), .CK(clk), .Q(m_data_out_y[5]) );
  DFF_X1 \accum_out_reg[6]  ( .D(n272), .CK(clk), .Q(m_data_out_y[6]) );
  DFF_X1 \accum_out_reg[8]  ( .D(n270), .CK(clk), .Q(m_data_out_y[8]) );
  DFF_X1 \accum_out_reg[7]  ( .D(n271), .CK(clk), .Q(m_data_out_y[7]), .QN(
        n1046) );
  DFF_X1 \accum_out_reg[10]  ( .D(n268), .CK(clk), .Q(m_data_out_y[10]) );
  DFF_X1 \accum_out_reg[9]  ( .D(n269), .CK(clk), .Q(m_data_out_y[9]), .QN(
        n1041) );
  DFF_X1 \accum_out_reg[11]  ( .D(n267), .CK(clk), .Q(m_data_out_y[11]), .QN(
        n1040) );
  DFF_X1 \accum_out_reg[12]  ( .D(n266), .CK(clk), .Q(m_data_out_y[12]), .QN(
        n1047) );
  DFFRS_X1 \accum_out_reg[14]  ( .D(n264), .CK(clk), .RN(1'b1), .SN(1'b1), .Q(
        m_data_out_y[14]) );
  BUF_X1 U410 ( .A(\DP_OP_61J1_122_4588/n326 ), .Z(n488) );
  OAI21_X1 U411 ( .B1(n860), .B2(n599), .A(n631), .ZN(n656) );
  CLKBUF_X1 U412 ( .A(n576), .Z(n391) );
  INV_X1 U413 ( .A(n534), .ZN(n535) );
  INV_X1 U414 ( .A(n566), .ZN(n562) );
  NAND2_X1 U415 ( .A1(n460), .A2(n1036), .ZN(n461) );
  BUF_X1 U416 ( .A(\DP_OP_61J1_122_4588/n326 ), .Z(n470) );
  CLKBUF_X1 U417 ( .A(n1043), .Z(n392) );
  BUF_X1 U418 ( .A(fmem_data[3]), .Z(n393) );
  INV_X1 U419 ( .A(n466), .ZN(n607) );
  BUF_X1 U420 ( .A(n607), .Z(n661) );
  NAND2_X1 U421 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U422 ( .A1(n624), .A2(n623), .ZN(n649) );
  CLKBUF_X1 U423 ( .A(n647), .Z(n593) );
  NAND2_X1 U424 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U425 ( .A1(n465), .A2(n464), .ZN(n513) );
  NAND2_X1 U426 ( .A1(n462), .A2(n461), .ZN(n465) );
  CLKBUF_X1 U427 ( .A(n652), .Z(n639) );
  CLKBUF_X1 U428 ( .A(n822), .Z(n836) );
  INV_X1 U429 ( .A(n492), .ZN(n389) );
  OAI21_X1 U430 ( .B1(n479), .B2(n478), .A(n839), .ZN(n390) );
  OR2_X1 U431 ( .A1(fmem_data[0]), .A2(n1033), .ZN(n542) );
  BUF_X1 U432 ( .A(n656), .Z(n394) );
  XNOR2_X1 U433 ( .A(fmem_data[5]), .B(fmem_data[6]), .ZN(n395) );
  XNOR2_X1 U434 ( .A(n1032), .B(fmem_data[3]), .ZN(n447) );
  XNOR2_X1 U435 ( .A(\DP_OP_61J1_122_4588/n326 ), .B(fmem_data[2]), .ZN(n446)
         );
  OR2_X1 U436 ( .A1(n898), .A2(n798), .ZN(n396) );
  NOR3_X2 U437 ( .A1(n1073), .A2(m_valid_y), .A3(reset), .ZN(n871) );
  OR2_X1 U438 ( .A1(n741), .A2(n740), .ZN(n398) );
  NAND2_X1 U439 ( .A1(n632), .A2(n631), .ZN(n399) );
  NAND2_X1 U440 ( .A1(n699), .A2(n701), .ZN(n400) );
  NAND2_X1 U441 ( .A1(n725), .A2(n709), .ZN(n401) );
  NAND2_X1 U442 ( .A1(n714), .A2(n727), .ZN(n402) );
  NAND2_X1 U443 ( .A1(n640), .A2(n639), .ZN(n403) );
  NAND2_X1 U444 ( .A1(n733), .A2(n732), .ZN(n404) );
  NAND2_X1 U445 ( .A1(n625), .A2(n651), .ZN(n405) );
  AND2_X1 U446 ( .A1(n414), .A2(n413), .ZN(n406) );
  AND2_X1 U447 ( .A1(n417), .A2(n416), .ZN(n407) );
  AND2_X1 U448 ( .A1(n420), .A2(n419), .ZN(n408) );
  AND2_X1 U449 ( .A1(n423), .A2(n422), .ZN(n409) );
  AND2_X1 U450 ( .A1(n426), .A2(n425), .ZN(n410) );
  AND2_X1 U451 ( .A1(n429), .A2(n428), .ZN(n411) );
  NAND2_X1 U453 ( .A1(n1048), .A2(fmem_addr[1]), .ZN(n886) );
  NAND2_X1 U454 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n888) );
  OAI22_X1 U455 ( .A1(n886), .A2(n1066), .B1(n888), .B2(n1052), .ZN(n412) );
  INV_X1 U456 ( .A(n412), .ZN(n414) );
  NAND2_X1 U457 ( .A1(n1048), .A2(n1064), .ZN(n798) );
  INV_X1 U458 ( .A(n798), .ZN(n749) );
  NOR2_X1 U459 ( .A1(fmem_addr[1]), .A2(n1048), .ZN(n899) );
  AOI22_X1 U460 ( .A1(n749), .A2(\fmem_inst/mem[0][1] ), .B1(n899), .B2(
        \fmem_inst/mem[1][1] ), .ZN(n413) );
  OAI22_X1 U461 ( .A1(n886), .A2(n1065), .B1(n888), .B2(n1051), .ZN(n415) );
  INV_X1 U462 ( .A(n415), .ZN(n417) );
  AOI22_X1 U463 ( .A1(n749), .A2(\fmem_inst/mem[0][0] ), .B1(n899), .B2(
        \fmem_inst/mem[1][0] ), .ZN(n416) );
  OAI22_X1 U464 ( .A1(n886), .A2(n1068), .B1(n888), .B2(n1054), .ZN(n418) );
  INV_X1 U465 ( .A(n418), .ZN(n420) );
  AOI22_X1 U466 ( .A1(n749), .A2(\fmem_inst/mem[0][3] ), .B1(n899), .B2(
        \fmem_inst/mem[1][3] ), .ZN(n419) );
  OAI22_X1 U467 ( .A1(n886), .A2(n1071), .B1(n888), .B2(n1057), .ZN(n421) );
  INV_X1 U468 ( .A(n421), .ZN(n423) );
  AOI22_X1 U469 ( .A1(n749), .A2(\fmem_inst/mem[0][6] ), .B1(n899), .B2(
        \fmem_inst/mem[1][6] ), .ZN(n422) );
  OAI22_X1 U470 ( .A1(n886), .A2(n1070), .B1(n888), .B2(n1056), .ZN(n424) );
  INV_X1 U471 ( .A(n424), .ZN(n426) );
  AOI22_X1 U472 ( .A1(n749), .A2(\fmem_inst/mem[0][5] ), .B1(n899), .B2(
        \fmem_inst/mem[1][5] ), .ZN(n425) );
  OAI22_X1 U473 ( .A1(n886), .A2(n1072), .B1(n888), .B2(n1058), .ZN(n427) );
  INV_X1 U474 ( .A(n427), .ZN(n429) );
  AOI22_X1 U475 ( .A1(n749), .A2(\fmem_inst/mem[0][7] ), .B1(n899), .B2(
        \fmem_inst/mem[1][7] ), .ZN(n428) );
  INV_X1 U476 ( .A(n446), .ZN(n448) );
  AND2_X1 U477 ( .A1(xmem_data[0]), .A2(n448), .ZN(n443) );
  XNOR2_X1 U478 ( .A(n488), .B(xmem_data[1]), .ZN(n430) );
  XNOR2_X1 U479 ( .A(n488), .B(xmem_data[2]), .ZN(n441) );
  OAI22_X1 U480 ( .A1(n542), .A2(n430), .B1(n441), .B2(n1042), .ZN(n442) );
  OAI22_X1 U481 ( .A1(n430), .A2(n1042), .B1(n542), .B2(xmem_data[0]), .ZN(
        n431) );
  AND2_X1 U482 ( .A1(n431), .A2(m_data_out_y[1]), .ZN(n435) );
  OR2_X1 U483 ( .A1(n436), .A2(n435), .ZN(n816) );
  XNOR2_X1 U484 ( .A(n431), .B(n1044), .ZN(n434) );
  OR2_X1 U485 ( .A1(xmem_data[0]), .A2(n1033), .ZN(n432) );
  NAND2_X1 U486 ( .A1(n432), .A2(n542), .ZN(n433) );
  NOR2_X1 U487 ( .A1(n434), .A2(n433), .ZN(n807) );
  AND2_X1 U488 ( .A1(xmem_data[0]), .A2(fmem_data[0]), .ZN(n755) );
  NAND2_X1 U489 ( .A1(n755), .A2(m_data_out_y[0]), .ZN(n810) );
  NAND2_X1 U490 ( .A1(n434), .A2(n433), .ZN(n808) );
  OAI21_X1 U491 ( .B1(n807), .B2(n810), .A(n808), .ZN(n817) );
  NAND2_X1 U492 ( .A1(n436), .A2(n435), .ZN(n815) );
  INV_X1 U493 ( .A(n815), .ZN(n437) );
  AOI21_X1 U494 ( .B1(n816), .B2(n817), .A(n437), .ZN(n830) );
  NAND2_X1 U495 ( .A1(n447), .A2(n446), .ZN(n583) );
  BUF_X2 U496 ( .A(fmem_data[3]), .Z(n532) );
  INV_X1 U497 ( .A(n393), .ZN(n439) );
  OR2_X1 U498 ( .A1(xmem_data[0]), .A2(n439), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n1032), .B(n1033), .ZN(n468) );
  BUF_X2 U500 ( .A(n468), .Z(n584) );
  OAI22_X1 U501 ( .A1(n533), .A2(n439), .B1(n438), .B2(n584), .ZN(n455) );
  XNOR2_X1 U502 ( .A(n393), .B(xmem_data[0]), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n532), .B(xmem_data[1]), .ZN(n450) );
  OAI22_X1 U504 ( .A1(n533), .A2(n440), .B1(n584), .B2(n450), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n488), .B(xmem_data[3]), .ZN(n451) );
  OAI22_X1 U506 ( .A1(n542), .A2(n441), .B1(n451), .B2(n1042), .ZN(n445) );
  FA_X1 U507 ( .A(n443), .B(m_data_out_y[2]), .CI(n442), .CO(n826), .S(n436)
         );
  NOR2_X1 U508 ( .A1(n827), .A2(n826), .ZN(n444) );
  NAND2_X1 U509 ( .A1(n827), .A2(n826), .ZN(n828) );
  OAI21_X1 U510 ( .B1(n830), .B2(n444), .A(n828), .ZN(n822) );
  HA_X1 U511 ( .A(n445), .B(m_data_out_y[3]), .CO(n477), .S(n453) );
  NAND2_X1 U512 ( .A1(n447), .A2(n446), .ZN(n533) );
  INV_X1 U513 ( .A(n448), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n393), .B(xmem_data[2]), .ZN(n469) );
  OAI22_X1 U515 ( .A1(n533), .A2(n450), .B1(n449), .B2(n469), .ZN(n476) );
  XNOR2_X1 U516 ( .A(n488), .B(xmem_data[4]), .ZN(n471) );
  OAI22_X1 U517 ( .A1(n542), .A2(n451), .B1(n471), .B2(n1042), .ZN(n462) );
  XNOR2_X1 U518 ( .A(fmem_data[4]), .B(n1035), .ZN(n466) );
  AND2_X1 U519 ( .A1(xmem_data[0]), .A2(n466), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(m_data_out_y[4]), .ZN(n452) );
  XNOR2_X1 U521 ( .A(n462), .B(n452), .ZN(n475) );
  INV_X1 U522 ( .A(n459), .ZN(n457) );
  FA_X1 U523 ( .A(n455), .B(n454), .CI(n453), .CO(n458), .S(n827) );
  INV_X1 U524 ( .A(n458), .ZN(n456) );
  NAND2_X1 U525 ( .A1(n457), .A2(n456), .ZN(n835) );
  NAND2_X1 U526 ( .A1(n459), .A2(n458), .ZN(n821) );
  INV_X1 U527 ( .A(n821), .ZN(n834) );
  AOI21_X1 U528 ( .B1(n822), .B2(n835), .A(n834), .ZN(n479) );
  INV_X1 U529 ( .A(n463), .ZN(n460) );
  NAND2_X1 U530 ( .A1(n463), .A2(m_data_out_y[4]), .ZN(n464) );
  XOR2_X1 U531 ( .A(fmem_data[5]), .B(fmem_data[4]), .Z(n472) );
  XNOR2_X1 U532 ( .A(n1034), .B(n1035), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n472), .A2(n484), .ZN(n540) );
  INV_X1 U534 ( .A(n1031), .ZN(n606) );
  XNOR2_X1 U535 ( .A(n606), .B(xmem_data[0]), .ZN(n467) );
  BUF_X2 U536 ( .A(fmem_data[5]), .Z(n538) );
  XNOR2_X1 U537 ( .A(n538), .B(xmem_data[1]), .ZN(n480) );
  OAI22_X1 U538 ( .A1(n540), .A2(n467), .B1(n607), .B2(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n532), .B(xmem_data[3]), .ZN(n481) );
  OAI22_X1 U540 ( .A1(n583), .A2(n469), .B1(n584), .B2(n481), .ZN(n501) );
  XNOR2_X1 U541 ( .A(n470), .B(xmem_data[5]), .ZN(n494) );
  OAI22_X1 U542 ( .A1(n542), .A2(n471), .B1(n494), .B2(n1042), .ZN(n500) );
  NAND2_X1 U543 ( .A1(n472), .A2(n484), .ZN(n662) );
  INV_X1 U544 ( .A(n538), .ZN(n474) );
  OR2_X1 U545 ( .A1(xmem_data[0]), .A2(n474), .ZN(n473) );
  OAI22_X1 U546 ( .A1(n662), .A2(n474), .B1(n473), .B2(n607), .ZN(n499) );
  FA_X1 U547 ( .A(n477), .B(n476), .CI(n475), .CO(n837), .S(n459) );
  NOR2_X1 U548 ( .A1(n838), .A2(n837), .ZN(n478) );
  NAND2_X1 U549 ( .A1(n838), .A2(n837), .ZN(n839) );
  OAI21_X1 U550 ( .B1(n479), .B2(n478), .A(n839), .ZN(n845) );
  XNOR2_X1 U551 ( .A(n538), .B(xmem_data[2]), .ZN(n485) );
  OAI22_X1 U552 ( .A1(n662), .A2(n480), .B1(n661), .B2(n485), .ZN(n498) );
  XNOR2_X1 U553 ( .A(n532), .B(xmem_data[4]), .ZN(n483) );
  OAI22_X1 U554 ( .A1(n583), .A2(n481), .B1(n483), .B2(n584), .ZN(n497) );
  HA_X1 U555 ( .A(n482), .B(m_data_out_y[5]), .CO(n496), .S(n512) );
  XNOR2_X1 U556 ( .A(fmem_data[3]), .B(xmem_data[5]), .ZN(n537) );
  OAI22_X1 U557 ( .A1(n533), .A2(n483), .B1(n537), .B2(n468), .ZN(n521) );
  XNOR2_X1 U558 ( .A(n538), .B(xmem_data[3]), .ZN(n539) );
  OAI22_X1 U559 ( .A1(n540), .A2(n485), .B1(n539), .B2(n484), .ZN(n520) );
  XNOR2_X1 U560 ( .A(n1045), .B(fmem_data[7]), .ZN(n522) );
  XNOR2_X1 U561 ( .A(fmem_data[5]), .B(fmem_data[6]), .ZN(n523) );
  NAND2_X1 U562 ( .A1(n522), .A2(n523), .ZN(n687) );
  INV_X1 U563 ( .A(n1043), .ZN(n604) );
  XNOR2_X1 U564 ( .A(n604), .B(xmem_data[0]), .ZN(n487) );
  XNOR2_X1 U565 ( .A(fmem_data[6]), .B(n1031), .ZN(n492) );
  INV_X1 U566 ( .A(n492), .ZN(n689) );
  XNOR2_X1 U567 ( .A(n392), .B(n1030), .ZN(n486) );
  OAI22_X1 U568 ( .A1(n687), .A2(n487), .B1(n689), .B2(n486), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n567), .B(n566), .ZN(n495) );
  XNOR2_X1 U570 ( .A(n470), .B(xmem_data[6]), .ZN(n493) );
  XNOR2_X1 U571 ( .A(n488), .B(xmem_data[7]), .ZN(n541) );
  OAI22_X1 U572 ( .A1(n542), .A2(n493), .B1(n541), .B2(n1042), .ZN(n549) );
  OR2_X1 U573 ( .A1(xmem_data[0]), .A2(n1043), .ZN(n489) );
  OR2_X1 U574 ( .A1(n489), .A2(n395), .ZN(n491) );
  NAND3_X1 U575 ( .A1(n522), .A2(n395), .A3(n604), .ZN(n490) );
  NAND2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n528) );
  XNOR2_X1 U577 ( .A(n528), .B(n1046), .ZN(n548) );
  AND2_X1 U578 ( .A1(n492), .A2(xmem_data[0]), .ZN(n503) );
  OAI22_X1 U579 ( .A1(n542), .A2(n494), .B1(n493), .B2(n1042), .ZN(n502) );
  XNOR2_X1 U580 ( .A(n495), .B(n564), .ZN(n517) );
  FA_X1 U581 ( .A(n498), .B(n497), .CI(n496), .CO(n567), .S(n510) );
  FA_X1 U582 ( .A(n501), .B(n500), .CI(n499), .CO(n508), .S(n511) );
  FA_X1 U583 ( .A(n503), .B(m_data_out_y[6]), .CI(n502), .CO(n547), .S(n507)
         );
  OR2_X1 U584 ( .A1(n508), .A2(n507), .ZN(n504) );
  NAND2_X1 U585 ( .A1(n510), .A2(n504), .ZN(n506) );
  NAND2_X1 U586 ( .A1(n508), .A2(n507), .ZN(n505) );
  NAND2_X1 U587 ( .A1(n506), .A2(n505), .ZN(n516) );
  NOR2_X1 U588 ( .A1(n517), .A2(n516), .ZN(n853) );
  XNOR2_X1 U589 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U590 ( .A(n510), .B(n509), .ZN(n515) );
  FA_X1 U591 ( .A(n513), .B(n512), .CI(n511), .CO(n514), .S(n838) );
  NOR2_X1 U592 ( .A1(n515), .A2(n514), .ZN(n851) );
  NOR2_X1 U593 ( .A1(n853), .A2(n851), .ZN(n719) );
  NOR2_X1 U594 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U595 ( .A1(n515), .A2(n514), .ZN(n850) );
  NAND2_X1 U596 ( .A1(n517), .A2(n516), .ZN(n854) );
  OAI21_X1 U597 ( .B1(n518), .B2(n850), .A(n854), .ZN(n718) );
  AOI21_X1 U598 ( .B1(n845), .B2(n719), .A(n718), .ZN(n657) );
  INV_X1 U599 ( .A(n657), .ZN(n863) );
  FA_X1 U600 ( .A(n520), .B(n521), .CI(n519), .CO(n558), .S(n566) );
  AND2_X1 U601 ( .A1(n523), .A2(n522), .ZN(n525) );
  XOR2_X1 U602 ( .A(n1043), .B(n1030), .Z(n524) );
  NAND2_X1 U603 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U604 ( .A(fmem_data[7]), .B(n1029), .ZN(n534) );
  NAND2_X1 U605 ( .A1(n534), .A2(n492), .ZN(n526) );
  NAND2_X1 U606 ( .A1(n527), .A2(n526), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n545), .B(m_data_out_y[8]), .ZN(n556) );
  AND2_X1 U608 ( .A1(n528), .A2(m_data_out_y[7]), .ZN(n555) );
  OR2_X1 U609 ( .A1(n556), .A2(n555), .ZN(n529) );
  NAND2_X1 U610 ( .A1(n558), .A2(n529), .ZN(n531) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n530) );
  NAND2_X1 U612 ( .A1(n531), .A2(n530), .ZN(n592) );
  XNOR2_X1 U613 ( .A(n393), .B(xmem_data[6]), .ZN(n536) );
  XNOR2_X1 U614 ( .A(n532), .B(xmem_data[7]), .ZN(n582) );
  OAI22_X1 U615 ( .A1(n533), .A2(n536), .B1(n584), .B2(n582), .ZN(n581) );
  XNOR2_X1 U616 ( .A(n604), .B(xmem_data[3]), .ZN(n578) );
  OAI22_X1 U617 ( .A1(n687), .A2(n535), .B1(n689), .B2(n578), .ZN(n580) );
  OAI22_X1 U618 ( .A1(n583), .A2(n537), .B1(n584), .B2(n536), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n538), .B(xmem_data[4]), .ZN(n544) );
  OAI22_X1 U620 ( .A1(n540), .A2(n539), .B1(n607), .B2(n544), .ZN(n551) );
  AOI21_X1 U621 ( .B1(n542), .B2(n1042), .A(n541), .ZN(n543) );
  INV_X1 U622 ( .A(n543), .ZN(n550) );
  XNOR2_X1 U623 ( .A(n606), .B(xmem_data[5]), .ZN(n587) );
  OAI22_X1 U624 ( .A1(n662), .A2(n544), .B1(n607), .B2(n587), .ZN(n576) );
  OR2_X1 U625 ( .A1(n545), .A2(m_data_out_y[8]), .ZN(n577) );
  XNOR2_X1 U626 ( .A(n576), .B(n577), .ZN(n546) );
  XNOR2_X1 U627 ( .A(n575), .B(n546), .ZN(n590) );
  FA_X1 U628 ( .A(n549), .B(n548), .CI(n547), .CO(n570), .S(n564) );
  INV_X1 U629 ( .A(n570), .ZN(n554) );
  FA_X1 U630 ( .A(n552), .B(n551), .CI(n550), .CO(n575), .S(n571) );
  INV_X1 U631 ( .A(n571), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n554), .A2(n553), .ZN(n559) );
  XNOR2_X1 U633 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U634 ( .A(n558), .B(n557), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n559), .A2(n572), .ZN(n561) );
  NAND2_X1 U636 ( .A1(n570), .A2(n571), .ZN(n560) );
  NAND2_X1 U637 ( .A1(n561), .A2(n560), .ZN(n597) );
  NOR2_X1 U638 ( .A1(n598), .A2(n597), .ZN(n645) );
  BUF_X1 U639 ( .A(n645), .Z(n636) );
  INV_X1 U640 ( .A(n567), .ZN(n563) );
  NAND2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n569), .A2(n568), .ZN(n595) );
  XNOR2_X1 U644 ( .A(n571), .B(n570), .ZN(n573) );
  XNOR2_X1 U645 ( .A(n573), .B(n572), .ZN(n596) );
  NOR2_X1 U646 ( .A1(n595), .A2(n596), .ZN(n644) );
  OR2_X1 U647 ( .A1(n636), .A2(n644), .ZN(n594) );
  OR2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n619) );
  NAND2_X1 U650 ( .A1(n577), .A2(n391), .ZN(n618) );
  NAND2_X1 U651 ( .A1(n619), .A2(n618), .ZN(n579) );
  INV_X1 U652 ( .A(n1043), .ZN(n671) );
  XNOR2_X1 U653 ( .A(n671), .B(xmem_data[4]), .ZN(n605) );
  OAI22_X1 U654 ( .A1(n687), .A2(n578), .B1(n689), .B2(n605), .ZN(n609) );
  XNOR2_X1 U655 ( .A(n579), .B(n621), .ZN(n589) );
  FA_X1 U656 ( .A(n581), .B(n1041), .CI(n580), .CO(n612), .S(n591) );
  AOI21_X1 U657 ( .B1(n584), .B2(n583), .A(n582), .ZN(n585) );
  INV_X1 U658 ( .A(n585), .ZN(n613) );
  XNOR2_X1 U659 ( .A(n606), .B(xmem_data[6]), .ZN(n608) );
  OR2_X1 U660 ( .A1(n607), .A2(n608), .ZN(n586) );
  OAI21_X1 U661 ( .B1(n662), .B2(n587), .A(n586), .ZN(n614) );
  XNOR2_X1 U662 ( .A(n613), .B(n614), .ZN(n588) );
  XNOR2_X1 U663 ( .A(n612), .B(n588), .ZN(n620) );
  XNOR2_X1 U664 ( .A(n589), .B(n620), .ZN(n601) );
  FA_X1 U665 ( .A(n592), .B(n591), .CI(n590), .CO(n600), .S(n598) );
  NOR2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n647) );
  INV_X1 U667 ( .A(n593), .ZN(n640) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n860) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n631) );
  INV_X1 U672 ( .A(n394), .ZN(n637) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n652) );
  OAI21_X1 U674 ( .B1(n637), .B2(n593), .A(n639), .ZN(n602) );
  AOI21_X1 U675 ( .B1(n863), .B2(n603), .A(n602), .ZN(n626) );
  XNOR2_X1 U676 ( .A(n604), .B(xmem_data[5]), .ZN(n664) );
  OAI22_X1 U677 ( .A1(n687), .A2(n605), .B1(n689), .B2(n664), .ZN(n659) );
  XNOR2_X1 U678 ( .A(n606), .B(xmem_data[7]), .ZN(n660) );
  OAI22_X1 U679 ( .A1(n662), .A2(n608), .B1(n607), .B2(n660), .ZN(n658) );
  FA_X1 U680 ( .A(m_data_out_y[9]), .B(m_data_out_y[10]), .CI(n609), .CO(n667), 
        .S(n621) );
  XNOR2_X1 U681 ( .A(n668), .B(n667), .ZN(n617) );
  INV_X1 U682 ( .A(n614), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n610), .A2(n585), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n666) );
  XNOR2_X1 U687 ( .A(n617), .B(n666), .ZN(n650) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n622) );
  OAI21_X1 U689 ( .B1(n622), .B2(n621), .A(n620), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U691 ( .A1(n650), .A2(n649), .ZN(n646) );
  INV_X1 U692 ( .A(n646), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U694 ( .A(n626), .B(n405), .ZN(n629) );
  INV_X1 U695 ( .A(reset), .ZN(n877) );
  NAND2_X1 U696 ( .A1(m_valid_y), .A2(n877), .ZN(n627) );
  NOR2_X1 U697 ( .A1(m_ready_y), .A2(n627), .ZN(n752) );
  AND2_X1 U698 ( .A1(n752), .A2(\ctrl_conv_output_inst/conv_start_accum ), 
        .ZN(n870) );
  NAND2_X1 U699 ( .A1(n870), .A2(m_data_out_y[11]), .ZN(n628) );
  OAI21_X1 U700 ( .B1(n629), .B2(n695), .A(n628), .ZN(n267) );
  INV_X1 U701 ( .A(n644), .ZN(n861) );
  INV_X1 U702 ( .A(n860), .ZN(n630) );
  AOI21_X1 U703 ( .B1(n863), .B2(n861), .A(n630), .ZN(n633) );
  INV_X1 U704 ( .A(n636), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n633), .B(n399), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n870), .A2(m_data_out_y[9]), .ZN(n634) );
  OAI21_X1 U707 ( .B1(n635), .B2(n695), .A(n634), .ZN(n269) );
  NOR2_X1 U708 ( .A1(n636), .A2(n644), .ZN(n638) );
  AOI21_X1 U709 ( .B1(n863), .B2(n638), .A(n394), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(n403), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n870), .A2(m_data_out_y[10]), .ZN(n642) );
  OAI21_X1 U712 ( .B1(n643), .B2(n695), .A(n642), .ZN(n268) );
  NOR2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n648), .A2(n655), .ZN(n722) );
  NOR2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n653) );
  OAI21_X1 U717 ( .B1(n653), .B2(n652), .A(n651), .ZN(n654) );
  AOI21_X1 U718 ( .B1(n656), .B2(n655), .A(n654), .ZN(n720) );
  OAI21_X1 U719 ( .B1(n722), .B2(n657), .A(n720), .ZN(n713) );
  FA_X1 U720 ( .A(n659), .B(n1040), .CI(n658), .CO(n679), .S(n668) );
  AOI21_X1 U721 ( .B1(n662), .B2(n661), .A(n660), .ZN(n663) );
  INV_X1 U722 ( .A(n663), .ZN(n678) );
  XNOR2_X1 U723 ( .A(n671), .B(xmem_data[6]), .ZN(n672) );
  OAI22_X1 U724 ( .A1(n389), .A2(n672), .B1(n687), .B2(n664), .ZN(n674) );
  XNOR2_X1 U725 ( .A(m_data_out_y[11]), .B(m_data_out_y[12]), .ZN(n665) );
  XNOR2_X1 U726 ( .A(n674), .B(n665), .ZN(n677) );
  OAI21_X1 U727 ( .B1(n668), .B2(n667), .A(n666), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n670), .A2(n669), .ZN(n680) );
  NOR2_X1 U729 ( .A1(n681), .A2(n680), .ZN(n737) );
  XNOR2_X1 U730 ( .A(n671), .B(xmem_data[7]), .ZN(n688) );
  OAI22_X1 U731 ( .A1(n687), .A2(n672), .B1(n389), .B2(n688), .ZN(n686) );
  NAND2_X1 U732 ( .A1(n1040), .A2(n1047), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n676) );
  NAND2_X1 U734 ( .A1(m_data_out_y[11]), .A2(m_data_out_y[12]), .ZN(n675) );
  NAND2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n685) );
  FA_X1 U736 ( .A(n679), .B(n678), .CI(n677), .CO(n682), .S(n681) );
  NOR2_X1 U737 ( .A1(n683), .A2(n682), .ZN(n741) );
  OR2_X1 U738 ( .A1(n737), .A2(n741), .ZN(n698) );
  INV_X1 U739 ( .A(n698), .ZN(n684) );
  NAND2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n866) );
  NAND2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n739) );
  OAI21_X1 U742 ( .B1(n866), .B2(n741), .A(n739), .ZN(n700) );
  AOI21_X1 U743 ( .B1(n713), .B2(n684), .A(n700), .ZN(n693) );
  FA_X1 U744 ( .A(n686), .B(n1039), .CI(n685), .CO(n692), .S(n683) );
  AOI21_X1 U745 ( .B1(n389), .B2(n687), .A(n688), .ZN(n690) );
  INV_X1 U746 ( .A(n690), .ZN(n703) );
  NOR2_X1 U747 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U748 ( .A(n697), .ZN(n699) );
  NAND2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n701) );
  XNOR2_X1 U750 ( .A(n693), .B(n400), .ZN(n696) );
  INV_X1 U751 ( .A(n871), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n870), .A2(m_data_out_y[14]), .ZN(n694) );
  OAI21_X1 U753 ( .B1(n696), .B2(n695), .A(n694), .ZN(n264) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n708) );
  NAND2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n726) );
  AOI21_X1 U757 ( .B1(n713), .B2(n708), .A(n726), .ZN(n705) );
  FA_X1 U758 ( .A(m_data_out_y[13]), .B(m_data_out_y[14]), .CI(n703), .CO(n704), .S(n691) );
  OR2_X1 U759 ( .A1(n704), .A2(n1038), .ZN(n725) );
  NAND2_X1 U760 ( .A1(n704), .A2(n1038), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n705), .B(n401), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n870), .A2(m_data_out_y[15]), .ZN(n706) );
  OAI21_X1 U763 ( .B1(n707), .B2(n695), .A(n706), .ZN(n263) );
  NAND2_X1 U764 ( .A1(n708), .A2(n725), .ZN(n723) );
  INV_X1 U765 ( .A(n723), .ZN(n712) );
  INV_X1 U766 ( .A(n709), .ZN(n724) );
  AOI21_X1 U767 ( .B1(n726), .B2(n725), .A(n724), .ZN(n710) );
  INV_X1 U768 ( .A(n710), .ZN(n711) );
  AOI21_X1 U769 ( .B1(n713), .B2(n712), .A(n711), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n397), .A2(m_data_out_y[15]), .ZN(n728) );
  INV_X1 U771 ( .A(n728), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n397), .A2(m_data_out_y[15]), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n715), .B(n402), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n870), .A2(m_data_out_y[16]), .ZN(n716) );
  OAI21_X1 U775 ( .B1(n717), .B2(n695), .A(n716), .ZN(n262) );
  AOI21_X1 U776 ( .B1(n390), .B2(n719), .A(n718), .ZN(n721) );
  OAI21_X1 U777 ( .B1(n722), .B2(n721), .A(n720), .ZN(n869) );
  NOR2_X1 U778 ( .A1(n723), .A2(n728), .ZN(n731) );
  AOI21_X1 U779 ( .B1(n726), .B2(n725), .A(n724), .ZN(n729) );
  OAI21_X1 U780 ( .B1(n729), .B2(n728), .A(n727), .ZN(n730) );
  AOI21_X1 U781 ( .B1(n869), .B2(n731), .A(n730), .ZN(n734) );
  OR2_X1 U782 ( .A1(n1037), .A2(m_data_out_y[16]), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n1037), .A2(m_data_out_y[16]), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n734), .B(n404), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n870), .A2(m_data_out_y[17]), .ZN(n735) );
  OAI21_X1 U786 ( .B1(n736), .B2(n695), .A(n735), .ZN(n279) );
  INV_X1 U787 ( .A(n737), .ZN(n867) );
  INV_X1 U788 ( .A(n866), .ZN(n738) );
  AOI21_X1 U789 ( .B1(n869), .B2(n867), .A(n738), .ZN(n742) );
  INV_X1 U790 ( .A(n739), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n742), .B(n398), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n870), .A2(m_data_out_y[13]), .ZN(n743) );
  OAI21_X1 U793 ( .B1(n744), .B2(n695), .A(n743), .ZN(n265) );
  OAI22_X1 U794 ( .A1(n886), .A2(n1067), .B1(n888), .B2(n1053), .ZN(n745) );
  INV_X1 U795 ( .A(n745), .ZN(n747) );
  AOI22_X1 U796 ( .A1(n749), .A2(\fmem_inst/mem[0][2] ), .B1(n899), .B2(
        \fmem_inst/mem[1][2] ), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n747), .A2(n746), .ZN(\fmem_inst/N13 ) );
  OAI22_X1 U798 ( .A1(n886), .A2(n1069), .B1(n888), .B2(n1055), .ZN(n748) );
  INV_X1 U799 ( .A(n748), .ZN(n751) );
  AOI22_X1 U800 ( .A1(n749), .A2(\fmem_inst/mem[0][4] ), .B1(n899), .B2(
        \fmem_inst/mem[1][4] ), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(\fmem_inst/N11 ) );
  NAND2_X1 U802 ( .A1(m_valid_y), .A2(m_ready_y), .ZN(n879) );
  NOR2_X1 U803 ( .A1(s_ready_x), .A2(s_ready_f), .ZN(n878) );
  NAND2_X1 U804 ( .A1(n878), .A2(conv_pre_start), .ZN(n880) );
  INV_X1 U805 ( .A(n880), .ZN(n891) );
  NAND2_X1 U806 ( .A1(n879), .A2(n891), .ZN(n892) );
  NOR2_X1 U807 ( .A1(reset), .A2(n892), .ZN(\ctrl_conv_output_inst/N68 ) );
  INV_X1 U808 ( .A(\ctrl_conv_output_inst/N68 ), .ZN(n754) );
  INV_X1 U809 ( .A(n752), .ZN(n753) );
  OAI21_X1 U810 ( .B1(n754), .B2(n1060), .A(n753), .ZN(n383) );
  OR2_X1 U811 ( .A1(n755), .A2(m_data_out_y[0]), .ZN(n756) );
  AND2_X1 U812 ( .A1(n756), .A2(n810), .ZN(n757) );
  AOI22_X1 U813 ( .A1(n870), .A2(m_data_out_y[0]), .B1(n871), .B2(n757), .ZN(
        n758) );
  INV_X1 U814 ( .A(n758), .ZN(n278) );
  NAND2_X1 U815 ( .A1(xmem_addr[0]), .A2(xmem_addr[1]), .ZN(n973) );
  NOR2_X1 U816 ( .A1(n1059), .A2(n973), .ZN(n934) );
  NAND2_X1 U817 ( .A1(xmem_addr[1]), .A2(n1062), .ZN(n1007) );
  NOR2_X1 U818 ( .A1(xmem_addr[2]), .A2(n1007), .ZN(n787) );
  AOI22_X1 U819 ( .A1(n934), .A2(\xmem_inst/mem[7][6] ), .B1(n787), .B2(
        \xmem_inst/mem[2][6] ), .ZN(n762) );
  NAND2_X1 U820 ( .A1(xmem_addr[0]), .A2(n1050), .ZN(n995) );
  NOR2_X1 U821 ( .A1(xmem_addr[2]), .A2(n995), .ZN(n789) );
  NAND2_X1 U822 ( .A1(n1062), .A2(n1050), .ZN(n984) );
  NOR2_X1 U823 ( .A1(xmem_addr[2]), .A2(n984), .ZN(n788) );
  AOI22_X1 U824 ( .A1(n789), .A2(\xmem_inst/mem[1][6] ), .B1(n788), .B2(
        \xmem_inst/mem[0][6] ), .ZN(n761) );
  NOR2_X1 U825 ( .A1(n1059), .A2(n984), .ZN(n791) );
  NOR2_X1 U826 ( .A1(n1007), .A2(n1059), .ZN(n790) );
  AOI22_X1 U827 ( .A1(n791), .A2(\xmem_inst/mem[4][6] ), .B1(n790), .B2(
        \xmem_inst/mem[6][6] ), .ZN(n760) );
  NOR2_X1 U828 ( .A1(n995), .A2(n1059), .ZN(n793) );
  NOR2_X1 U829 ( .A1(xmem_addr[2]), .A2(n973), .ZN(n792) );
  AOI22_X1 U830 ( .A1(n793), .A2(\xmem_inst/mem[5][6] ), .B1(n792), .B2(
        \xmem_inst/mem[3][6] ), .ZN(n759) );
  NAND4_X1 U831 ( .A1(n762), .A2(n761), .A3(n760), .A4(n759), .ZN(
        \xmem_inst/N14 ) );
  AOI22_X1 U832 ( .A1(n934), .A2(\xmem_inst/mem[7][4] ), .B1(n787), .B2(
        \xmem_inst/mem[2][4] ), .ZN(n766) );
  AOI22_X1 U833 ( .A1(n789), .A2(\xmem_inst/mem[1][4] ), .B1(n788), .B2(
        \xmem_inst/mem[0][4] ), .ZN(n765) );
  AOI22_X1 U834 ( .A1(n791), .A2(\xmem_inst/mem[4][4] ), .B1(n790), .B2(
        \xmem_inst/mem[6][4] ), .ZN(n764) );
  AOI22_X1 U835 ( .A1(n793), .A2(\xmem_inst/mem[5][4] ), .B1(n792), .B2(
        \xmem_inst/mem[3][4] ), .ZN(n763) );
  NAND4_X1 U836 ( .A1(n766), .A2(n765), .A3(n764), .A4(n763), .ZN(
        \xmem_inst/N16 ) );
  AOI22_X1 U837 ( .A1(n934), .A2(\xmem_inst/mem[7][1] ), .B1(n787), .B2(
        \xmem_inst/mem[2][1] ), .ZN(n770) );
  AOI22_X1 U838 ( .A1(n789), .A2(\xmem_inst/mem[1][1] ), .B1(n788), .B2(
        \xmem_inst/mem[0][1] ), .ZN(n769) );
  AOI22_X1 U839 ( .A1(n791), .A2(\xmem_inst/mem[4][1] ), .B1(n790), .B2(
        \xmem_inst/mem[6][1] ), .ZN(n768) );
  AOI22_X1 U840 ( .A1(n793), .A2(\xmem_inst/mem[5][1] ), .B1(n792), .B2(
        \xmem_inst/mem[3][1] ), .ZN(n767) );
  NAND4_X1 U841 ( .A1(n770), .A2(n769), .A3(n768), .A4(n767), .ZN(
        \xmem_inst/N19 ) );
  AOI22_X1 U842 ( .A1(n934), .A2(\xmem_inst/mem[7][7] ), .B1(n787), .B2(
        \xmem_inst/mem[2][7] ), .ZN(n774) );
  AOI22_X1 U843 ( .A1(n789), .A2(\xmem_inst/mem[1][7] ), .B1(n788), .B2(
        \xmem_inst/mem[0][7] ), .ZN(n773) );
  AOI22_X1 U844 ( .A1(n791), .A2(\xmem_inst/mem[4][7] ), .B1(n790), .B2(
        \xmem_inst/mem[6][7] ), .ZN(n772) );
  AOI22_X1 U845 ( .A1(n793), .A2(\xmem_inst/mem[5][7] ), .B1(n792), .B2(
        \xmem_inst/mem[3][7] ), .ZN(n771) );
  NAND4_X1 U846 ( .A1(n774), .A2(n773), .A3(n772), .A4(n771), .ZN(
        \xmem_inst/N13 ) );
  AOI22_X1 U847 ( .A1(n934), .A2(\xmem_inst/mem[7][3] ), .B1(n787), .B2(
        \xmem_inst/mem[2][3] ), .ZN(n778) );
  AOI22_X1 U848 ( .A1(n789), .A2(\xmem_inst/mem[1][3] ), .B1(n788), .B2(
        \xmem_inst/mem[0][3] ), .ZN(n777) );
  AOI22_X1 U849 ( .A1(n791), .A2(\xmem_inst/mem[4][3] ), .B1(n790), .B2(
        \xmem_inst/mem[6][3] ), .ZN(n776) );
  AOI22_X1 U850 ( .A1(n793), .A2(\xmem_inst/mem[5][3] ), .B1(n792), .B2(
        \xmem_inst/mem[3][3] ), .ZN(n775) );
  NAND4_X1 U851 ( .A1(n778), .A2(n777), .A3(n776), .A4(n775), .ZN(
        \xmem_inst/N17 ) );
  AOI22_X1 U852 ( .A1(n934), .A2(\xmem_inst/mem[7][5] ), .B1(n787), .B2(
        \xmem_inst/mem[2][5] ), .ZN(n782) );
  AOI22_X1 U853 ( .A1(n789), .A2(\xmem_inst/mem[1][5] ), .B1(n788), .B2(
        \xmem_inst/mem[0][5] ), .ZN(n781) );
  AOI22_X1 U854 ( .A1(n791), .A2(\xmem_inst/mem[4][5] ), .B1(n790), .B2(
        \xmem_inst/mem[6][5] ), .ZN(n780) );
  AOI22_X1 U855 ( .A1(n793), .A2(\xmem_inst/mem[5][5] ), .B1(n792), .B2(
        \xmem_inst/mem[3][5] ), .ZN(n779) );
  NAND4_X1 U856 ( .A1(n782), .A2(n781), .A3(n780), .A4(n779), .ZN(
        \xmem_inst/N15 ) );
  AOI22_X1 U857 ( .A1(n934), .A2(\xmem_inst/mem[7][2] ), .B1(n787), .B2(
        \xmem_inst/mem[2][2] ), .ZN(n786) );
  AOI22_X1 U858 ( .A1(n789), .A2(\xmem_inst/mem[1][2] ), .B1(n788), .B2(
        \xmem_inst/mem[0][2] ), .ZN(n785) );
  AOI22_X1 U859 ( .A1(n791), .A2(\xmem_inst/mem[4][2] ), .B1(n790), .B2(
        \xmem_inst/mem[6][2] ), .ZN(n784) );
  AOI22_X1 U860 ( .A1(n793), .A2(\xmem_inst/mem[5][2] ), .B1(n792), .B2(
        \xmem_inst/mem[3][2] ), .ZN(n783) );
  NAND4_X1 U861 ( .A1(n786), .A2(n785), .A3(n784), .A4(n783), .ZN(
        \xmem_inst/N18 ) );
  AOI22_X1 U862 ( .A1(n934), .A2(\xmem_inst/mem[7][0] ), .B1(n787), .B2(
        \xmem_inst/mem[2][0] ), .ZN(n797) );
  AOI22_X1 U863 ( .A1(n789), .A2(\xmem_inst/mem[1][0] ), .B1(n788), .B2(
        \xmem_inst/mem[0][0] ), .ZN(n796) );
  AOI22_X1 U864 ( .A1(n791), .A2(\xmem_inst/mem[4][0] ), .B1(n790), .B2(
        \xmem_inst/mem[6][0] ), .ZN(n795) );
  AOI22_X1 U865 ( .A1(n793), .A2(\xmem_inst/mem[5][0] ), .B1(n792), .B2(
        \xmem_inst/mem[3][0] ), .ZN(n794) );
  NAND4_X1 U866 ( .A1(n797), .A2(n796), .A3(n795), .A4(n794), .ZN(
        \xmem_inst/N20 ) );
  INV_X1 U867 ( .A(s_data_in_f[3]), .ZN(n917) );
  NAND2_X1 U868 ( .A1(s_ready_f), .A2(s_valid_f), .ZN(n898) );
  NAND2_X1 U869 ( .A1(n396), .A2(\fmem_inst/mem[0][3] ), .ZN(n799) );
  OAI21_X1 U870 ( .B1(n917), .B2(n396), .A(n799), .ZN(n376) );
  INV_X1 U871 ( .A(s_data_in_f[5]), .ZN(n919) );
  NAND2_X1 U872 ( .A1(n396), .A2(\fmem_inst/mem[0][5] ), .ZN(n800) );
  OAI21_X1 U873 ( .B1(n919), .B2(n396), .A(n800), .ZN(n374) );
  INV_X1 U874 ( .A(s_data_in_f[6]), .ZN(n920) );
  NAND2_X1 U875 ( .A1(n396), .A2(\fmem_inst/mem[0][6] ), .ZN(n801) );
  OAI21_X1 U876 ( .B1(n920), .B2(n396), .A(n801), .ZN(n373) );
  INV_X1 U877 ( .A(s_data_in_f[7]), .ZN(n922) );
  NAND2_X1 U878 ( .A1(n396), .A2(\fmem_inst/mem[0][7] ), .ZN(n802) );
  OAI21_X1 U879 ( .B1(n922), .B2(n396), .A(n802), .ZN(n372) );
  INV_X1 U880 ( .A(s_data_in_f[2]), .ZN(n916) );
  NAND2_X1 U881 ( .A1(n396), .A2(\fmem_inst/mem[0][2] ), .ZN(n803) );
  OAI21_X1 U882 ( .B1(n916), .B2(n396), .A(n803), .ZN(n377) );
  INV_X1 U883 ( .A(s_data_in_f[0]), .ZN(n914) );
  NAND2_X1 U884 ( .A1(n396), .A2(\fmem_inst/mem[0][0] ), .ZN(n804) );
  OAI21_X1 U885 ( .B1(n914), .B2(n396), .A(n804), .ZN(n379) );
  INV_X1 U886 ( .A(s_data_in_f[1]), .ZN(n915) );
  NAND2_X1 U887 ( .A1(n396), .A2(\fmem_inst/mem[0][1] ), .ZN(n805) );
  OAI21_X1 U888 ( .B1(n915), .B2(n396), .A(n805), .ZN(n378) );
  INV_X1 U889 ( .A(s_data_in_f[4]), .ZN(n918) );
  NAND2_X1 U890 ( .A1(n396), .A2(\fmem_inst/mem[0][4] ), .ZN(n806) );
  OAI21_X1 U891 ( .B1(n918), .B2(n396), .A(n806), .ZN(n375) );
  INV_X1 U892 ( .A(n807), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n812) );
  INV_X1 U894 ( .A(n810), .ZN(n811) );
  XNOR2_X1 U895 ( .A(n812), .B(n811), .ZN(n813) );
  AOI22_X1 U896 ( .A1(n813), .A2(n871), .B1(n870), .B2(m_data_out_y[1]), .ZN(
        n814) );
  INV_X1 U897 ( .A(n814), .ZN(n277) );
  NAND2_X1 U898 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U899 ( .A(n818), .B(n817), .ZN(n819) );
  AOI22_X1 U900 ( .A1(n819), .A2(n871), .B1(n870), .B2(m_data_out_y[2]), .ZN(
        n820) );
  INV_X1 U901 ( .A(n820), .ZN(n276) );
  NAND2_X1 U902 ( .A1(n835), .A2(n821), .ZN(n823) );
  XNOR2_X1 U903 ( .A(n823), .B(n836), .ZN(n824) );
  AOI22_X1 U904 ( .A1(n824), .A2(n871), .B1(n870), .B2(m_data_out_y[4]), .ZN(
        n825) );
  INV_X1 U905 ( .A(n825), .ZN(n274) );
  OR2_X1 U906 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U907 ( .A1(n829), .A2(n828), .ZN(n831) );
  XOR2_X1 U908 ( .A(n831), .B(n830), .Z(n832) );
  AOI22_X1 U909 ( .A1(n832), .A2(n871), .B1(n870), .B2(m_data_out_y[3]), .ZN(
        n833) );
  INV_X1 U910 ( .A(n833), .ZN(n275) );
  AOI21_X1 U911 ( .B1(n836), .B2(n835), .A(n834), .ZN(n842) );
  OR2_X1 U912 ( .A1(n838), .A2(n837), .ZN(n840) );
  NAND2_X1 U913 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U914 ( .A(n842), .B(n841), .Z(n843) );
  AOI22_X1 U915 ( .A1(n843), .A2(n871), .B1(n870), .B2(m_data_out_y[5]), .ZN(
        n844) );
  INV_X1 U916 ( .A(n844), .ZN(n273) );
  INV_X1 U917 ( .A(n390), .ZN(n852) );
  INV_X1 U918 ( .A(n851), .ZN(n846) );
  NAND2_X1 U919 ( .A1(n846), .A2(n850), .ZN(n847) );
  XOR2_X1 U920 ( .A(n852), .B(n847), .Z(n848) );
  AOI22_X1 U921 ( .A1(n848), .A2(n871), .B1(n870), .B2(m_data_out_y[6]), .ZN(
        n849) );
  INV_X1 U922 ( .A(n849), .ZN(n272) );
  OAI21_X1 U923 ( .B1(n852), .B2(n851), .A(n850), .ZN(n857) );
  INV_X1 U924 ( .A(n853), .ZN(n855) );
  NAND2_X1 U925 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U926 ( .A(n857), .B(n856), .ZN(n858) );
  AOI22_X1 U927 ( .A1(n858), .A2(n871), .B1(n870), .B2(m_data_out_y[7]), .ZN(
        n859) );
  INV_X1 U928 ( .A(n859), .ZN(n271) );
  NAND2_X1 U929 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U930 ( .A(n863), .B(n862), .ZN(n864) );
  AOI22_X1 U931 ( .A1(n864), .A2(n871), .B1(n870), .B2(m_data_out_y[8]), .ZN(
        n865) );
  INV_X1 U932 ( .A(n865), .ZN(n270) );
  NAND2_X1 U933 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U934 ( .A(n869), .B(n868), .ZN(n872) );
  AOI22_X1 U935 ( .A1(n872), .A2(n871), .B1(n870), .B2(m_data_out_y[12]), .ZN(
        n873) );
  INV_X1 U936 ( .A(n873), .ZN(n266) );
  NOR2_X1 U937 ( .A1(reset), .A2(conv_done), .ZN(n927) );
  NAND3_X1 U938 ( .A1(n1060), .A2(\ctrl_conv_output_inst/m_pre_valid ), .A3(
        n927), .ZN(n884) );
  NAND2_X1 U939 ( .A1(n1060), .A2(\ctrl_conv_output_inst/m_pre_valid ), .ZN(
        n882) );
  OAI21_X1 U940 ( .B1(n1061), .B2(n882), .A(n927), .ZN(n885) );
  OAI21_X1 U941 ( .B1(n884), .B2(\ctrl_conv_output_inst/cnt_conv [1]), .A(n885), .ZN(n874) );
  INV_X1 U942 ( .A(n874), .ZN(n876) );
  OR3_X1 U943 ( .A1(n1061), .A2(n1049), .A3(n884), .ZN(n875) );
  AOI22_X1 U944 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(n876), .B1(
        n875), .B2(n1063), .ZN(n387) );
  NAND2_X1 U945 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n1049), .ZN(
        n883) );
  NOR4_X1 U946 ( .A1(reset), .A2(n879), .A3(n1063), .A4(n883), .ZN(
        \ctrl_conv_output_inst/N71 ) );
  AND2_X1 U947 ( .A1(n878), .A2(n877), .ZN(N6) );
  INV_X1 U948 ( .A(n879), .ZN(n890) );
  OR2_X1 U949 ( .A1(n880), .A2(n888), .ZN(n881) );
  AOI221_X1 U950 ( .B1(n890), .B2(\ctrl_conv_output_inst/m_pre_valid_int ), 
        .C1(n881), .C2(n1060), .A(reset), .ZN(n388) );
  AOI21_X1 U951 ( .B1(n1061), .B2(n882), .A(n885), .ZN(n386) );
  OAI22_X1 U952 ( .A1(n1049), .A2(n885), .B1(n884), .B2(n883), .ZN(n385) );
  INV_X1 U953 ( .A(n886), .ZN(n910) );
  NAND2_X1 U954 ( .A1(n891), .A2(n910), .ZN(n887) );
  AOI221_X1 U955 ( .B1(n890), .B2(\ctrl_conv_output_inst/m_pre_valid ), .C1(
        n887), .C2(n1074), .A(reset), .ZN(n384) );
  NOR2_X1 U956 ( .A1(n898), .A2(n888), .ZN(n923) );
  INV_X1 U957 ( .A(n923), .ZN(n921) );
  INV_X1 U958 ( .A(n927), .ZN(n930) );
  AOI21_X1 U959 ( .B1(n921), .B2(s_ready_f), .A(n930), .ZN(n889) );
  INV_X1 U960 ( .A(n889), .ZN(n382) );
  NAND2_X1 U961 ( .A1(n891), .A2(n890), .ZN(n931) );
  NAND2_X1 U962 ( .A1(n927), .A2(n931), .ZN(n929) );
  INV_X1 U963 ( .A(n929), .ZN(n893) );
  OR2_X1 U964 ( .A1(n892), .A2(\ctrl_conv_output_inst/m_pre_valid ), .ZN(n925)
         );
  NAND3_X1 U965 ( .A1(n893), .A2(n925), .A3(n898), .ZN(n895) );
  NAND2_X1 U966 ( .A1(n925), .A2(n898), .ZN(n894) );
  NAND2_X1 U967 ( .A1(n927), .A2(n894), .ZN(n896) );
  AOI22_X1 U968 ( .A1(fmem_addr[0]), .A2(n895), .B1(n896), .B2(n1048), .ZN(
        n381) );
  NOR2_X1 U969 ( .A1(n899), .A2(n910), .ZN(n897) );
  OAI22_X1 U970 ( .A1(n897), .A2(n896), .B1(n895), .B2(n1064), .ZN(n380) );
  INV_X1 U971 ( .A(n898), .ZN(n911) );
  NAND2_X1 U972 ( .A1(n911), .A2(n899), .ZN(n908) );
  INV_X1 U973 ( .A(n908), .ZN(n907) );
  OAI22_X1 U974 ( .A1(n908), .A2(s_data_in_f[0]), .B1(\fmem_inst/mem[1][0] ), 
        .B2(n907), .ZN(n900) );
  INV_X1 U975 ( .A(n900), .ZN(n371) );
  OAI22_X1 U976 ( .A1(n908), .A2(s_data_in_f[1]), .B1(\fmem_inst/mem[1][1] ), 
        .B2(n907), .ZN(n901) );
  INV_X1 U977 ( .A(n901), .ZN(n370) );
  OAI22_X1 U978 ( .A1(n908), .A2(s_data_in_f[2]), .B1(\fmem_inst/mem[1][2] ), 
        .B2(n907), .ZN(n902) );
  INV_X1 U979 ( .A(n902), .ZN(n369) );
  OAI22_X1 U980 ( .A1(n908), .A2(s_data_in_f[3]), .B1(\fmem_inst/mem[1][3] ), 
        .B2(n907), .ZN(n903) );
  INV_X1 U981 ( .A(n903), .ZN(n368) );
  OAI22_X1 U982 ( .A1(n908), .A2(s_data_in_f[4]), .B1(\fmem_inst/mem[1][4] ), 
        .B2(n907), .ZN(n904) );
  INV_X1 U983 ( .A(n904), .ZN(n367) );
  OAI22_X1 U984 ( .A1(n908), .A2(s_data_in_f[5]), .B1(\fmem_inst/mem[1][5] ), 
        .B2(n907), .ZN(n905) );
  INV_X1 U985 ( .A(n905), .ZN(n366) );
  OAI22_X1 U986 ( .A1(n908), .A2(s_data_in_f[6]), .B1(\fmem_inst/mem[1][6] ), 
        .B2(n907), .ZN(n906) );
  INV_X1 U987 ( .A(n906), .ZN(n365) );
  OAI22_X1 U988 ( .A1(n908), .A2(s_data_in_f[7]), .B1(\fmem_inst/mem[1][7] ), 
        .B2(n907), .ZN(n909) );
  INV_X1 U989 ( .A(n909), .ZN(n364) );
  NAND2_X1 U990 ( .A1(n911), .A2(n910), .ZN(n912) );
  INV_X1 U991 ( .A(n912), .ZN(n913) );
  AOI22_X1 U992 ( .A1(n913), .A2(n914), .B1(n1065), .B2(n912), .ZN(n363) );
  AOI22_X1 U993 ( .A1(n913), .A2(n915), .B1(n1066), .B2(n912), .ZN(n362) );
  AOI22_X1 U994 ( .A1(n913), .A2(n916), .B1(n1067), .B2(n912), .ZN(n361) );
  AOI22_X1 U995 ( .A1(n913), .A2(n917), .B1(n1068), .B2(n912), .ZN(n360) );
  AOI22_X1 U996 ( .A1(n913), .A2(n918), .B1(n1069), .B2(n912), .ZN(n359) );
  AOI22_X1 U997 ( .A1(n913), .A2(n919), .B1(n1070), .B2(n912), .ZN(n358) );
  AOI22_X1 U998 ( .A1(n913), .A2(n920), .B1(n1071), .B2(n912), .ZN(n357) );
  AOI22_X1 U999 ( .A1(n913), .A2(n922), .B1(n1072), .B2(n912), .ZN(n356) );
  AOI22_X1 U1000 ( .A1(n923), .A2(n914), .B1(n1051), .B2(n921), .ZN(n355) );
  AOI22_X1 U1001 ( .A1(n923), .A2(n915), .B1(n1052), .B2(n921), .ZN(n354) );
  AOI22_X1 U1002 ( .A1(n923), .A2(n916), .B1(n1053), .B2(n921), .ZN(n353) );
  AOI22_X1 U1003 ( .A1(n923), .A2(n917), .B1(n1054), .B2(n921), .ZN(n352) );
  AOI22_X1 U1004 ( .A1(n923), .A2(n918), .B1(n1055), .B2(n921), .ZN(n351) );
  AOI22_X1 U1005 ( .A1(n923), .A2(n919), .B1(n1056), .B2(n921), .ZN(n350) );
  AOI22_X1 U1006 ( .A1(n923), .A2(n920), .B1(n1057), .B2(n921), .ZN(n349) );
  AOI22_X1 U1007 ( .A1(n923), .A2(n922), .B1(n1058), .B2(n921), .ZN(n348) );
  NAND2_X1 U1008 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n926) );
  INV_X1 U1009 ( .A(n926), .ZN(n941) );
  NAND2_X1 U1010 ( .A1(n941), .A2(xmem_addr[2]), .ZN(n1006) );
  NOR2_X1 U1011 ( .A1(n973), .A2(n1006), .ZN(n1025) );
  INV_X1 U1012 ( .A(n1025), .ZN(n1026) );
  AOI21_X1 U1013 ( .B1(n1026), .B2(s_ready_x), .A(n930), .ZN(n924) );
  INV_X1 U1014 ( .A(n924), .ZN(n347) );
  NAND2_X1 U1015 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1016 ( .A1(n927), .A2(n928), .ZN(n940) );
  NOR2_X1 U1017 ( .A1(n929), .A2(n928), .ZN(n937) );
  NOR2_X1 U1018 ( .A1(n931), .A2(n930), .ZN(n936) );
  AOI22_X1 U1019 ( .A1(xmem_addr[0]), .A2(n937), .B1(n936), .B2(
        \ctrl_conv_output_inst/cnt_conv [0]), .ZN(n932) );
  OAI21_X1 U1020 ( .B1(xmem_addr[0]), .B2(n940), .A(n932), .ZN(n346) );
  AOI22_X1 U1021 ( .A1(n937), .A2(xmem_addr[1]), .B1(n936), .B2(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n933) );
  OAI221_X1 U1022 ( .B1(n940), .B2(n1007), .C1(n940), .C2(n995), .A(n933), 
        .ZN(n345) );
  AOI21_X1 U1023 ( .B1(n1059), .B2(n973), .A(n934), .ZN(n935) );
  INV_X1 U1024 ( .A(n935), .ZN(n939) );
  AOI22_X1 U1025 ( .A1(n937), .A2(xmem_addr[2]), .B1(n936), .B2(
        \ctrl_conv_output_inst/cnt_conv [2]), .ZN(n938) );
  OAI21_X1 U1026 ( .B1(n940), .B2(n939), .A(n938), .ZN(n344) );
  NAND2_X1 U1027 ( .A1(n941), .A2(n1059), .ZN(n972) );
  NOR2_X1 U1028 ( .A1(n984), .A2(n972), .ZN(n949) );
  INV_X1 U1029 ( .A(n949), .ZN(n950) );
  OAI22_X1 U1030 ( .A1(n950), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[0][0] ), 
        .B2(n949), .ZN(n942) );
  INV_X1 U1031 ( .A(n942), .ZN(n343) );
  OAI22_X1 U1032 ( .A1(n950), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[0][1] ), 
        .B2(n949), .ZN(n943) );
  INV_X1 U1033 ( .A(n943), .ZN(n342) );
  OAI22_X1 U1034 ( .A1(n950), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[0][2] ), 
        .B2(n949), .ZN(n944) );
  INV_X1 U1035 ( .A(n944), .ZN(n341) );
  OAI22_X1 U1036 ( .A1(n950), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[0][3] ), 
        .B2(n949), .ZN(n945) );
  INV_X1 U1037 ( .A(n945), .ZN(n340) );
  OAI22_X1 U1038 ( .A1(n950), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[0][4] ), 
        .B2(n949), .ZN(n946) );
  INV_X1 U1039 ( .A(n946), .ZN(n339) );
  OAI22_X1 U1040 ( .A1(n950), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[0][5] ), 
        .B2(n949), .ZN(n947) );
  INV_X1 U1041 ( .A(n947), .ZN(n338) );
  OAI22_X1 U1042 ( .A1(n950), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[0][6] ), 
        .B2(n949), .ZN(n948) );
  INV_X1 U1043 ( .A(n948), .ZN(n337) );
  OAI22_X1 U1044 ( .A1(n950), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[0][7] ), 
        .B2(n949), .ZN(n951) );
  INV_X1 U1045 ( .A(n951), .ZN(n336) );
  NOR2_X1 U1046 ( .A1(n995), .A2(n972), .ZN(n959) );
  INV_X1 U1047 ( .A(n959), .ZN(n960) );
  OAI22_X1 U1048 ( .A1(n960), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[1][0] ), 
        .B2(n959), .ZN(n952) );
  INV_X1 U1049 ( .A(n952), .ZN(n335) );
  OAI22_X1 U1050 ( .A1(n960), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[1][1] ), 
        .B2(n959), .ZN(n953) );
  INV_X1 U1051 ( .A(n953), .ZN(n334) );
  OAI22_X1 U1052 ( .A1(n960), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[1][2] ), 
        .B2(n959), .ZN(n954) );
  INV_X1 U1053 ( .A(n954), .ZN(n333) );
  OAI22_X1 U1054 ( .A1(n960), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[1][3] ), 
        .B2(n959), .ZN(n955) );
  INV_X1 U1055 ( .A(n955), .ZN(n332) );
  OAI22_X1 U1056 ( .A1(n960), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[1][4] ), 
        .B2(n959), .ZN(n956) );
  INV_X1 U1057 ( .A(n956), .ZN(n331) );
  OAI22_X1 U1058 ( .A1(n960), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[1][5] ), 
        .B2(n959), .ZN(n957) );
  INV_X1 U1059 ( .A(n957), .ZN(n330) );
  OAI22_X1 U1060 ( .A1(n960), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[1][6] ), 
        .B2(n959), .ZN(n958) );
  INV_X1 U1061 ( .A(n958), .ZN(n329) );
  OAI22_X1 U1062 ( .A1(n960), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[1][7] ), 
        .B2(n959), .ZN(n961) );
  INV_X1 U1063 ( .A(n961), .ZN(n328) );
  NOR2_X1 U1064 ( .A1(n1007), .A2(n972), .ZN(n969) );
  INV_X1 U1065 ( .A(n969), .ZN(n970) );
  OAI22_X1 U1066 ( .A1(n970), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[2][0] ), 
        .B2(n969), .ZN(n962) );
  INV_X1 U1067 ( .A(n962), .ZN(n327) );
  OAI22_X1 U1068 ( .A1(n970), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[2][1] ), 
        .B2(n969), .ZN(n963) );
  INV_X1 U1069 ( .A(n963), .ZN(n326) );
  OAI22_X1 U1070 ( .A1(n970), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[2][2] ), 
        .B2(n969), .ZN(n964) );
  INV_X1 U1071 ( .A(n964), .ZN(n325) );
  OAI22_X1 U1072 ( .A1(n970), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[2][3] ), 
        .B2(n969), .ZN(n965) );
  INV_X1 U1073 ( .A(n965), .ZN(n324) );
  OAI22_X1 U1074 ( .A1(n970), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[2][4] ), 
        .B2(n969), .ZN(n966) );
  INV_X1 U1075 ( .A(n966), .ZN(n323) );
  OAI22_X1 U1076 ( .A1(n970), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[2][5] ), 
        .B2(n969), .ZN(n967) );
  INV_X1 U1077 ( .A(n967), .ZN(n322) );
  OAI22_X1 U1078 ( .A1(n970), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[2][6] ), 
        .B2(n969), .ZN(n968) );
  INV_X1 U1079 ( .A(n968), .ZN(n321) );
  OAI22_X1 U1080 ( .A1(n970), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[2][7] ), 
        .B2(n969), .ZN(n971) );
  INV_X1 U1081 ( .A(n971), .ZN(n320) );
  NOR2_X1 U1082 ( .A1(n973), .A2(n972), .ZN(n981) );
  INV_X1 U1083 ( .A(n981), .ZN(n982) );
  OAI22_X1 U1084 ( .A1(n982), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[3][0] ), 
        .B2(n981), .ZN(n974) );
  INV_X1 U1085 ( .A(n974), .ZN(n319) );
  OAI22_X1 U1086 ( .A1(n982), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[3][1] ), 
        .B2(n981), .ZN(n975) );
  INV_X1 U1087 ( .A(n975), .ZN(n318) );
  OAI22_X1 U1088 ( .A1(n982), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[3][2] ), 
        .B2(n981), .ZN(n976) );
  INV_X1 U1089 ( .A(n976), .ZN(n317) );
  OAI22_X1 U1090 ( .A1(n982), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[3][3] ), 
        .B2(n981), .ZN(n977) );
  INV_X1 U1091 ( .A(n977), .ZN(n316) );
  OAI22_X1 U1092 ( .A1(n982), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[3][4] ), 
        .B2(n981), .ZN(n978) );
  INV_X1 U1093 ( .A(n978), .ZN(n315) );
  OAI22_X1 U1094 ( .A1(n982), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[3][5] ), 
        .B2(n981), .ZN(n979) );
  INV_X1 U1095 ( .A(n979), .ZN(n314) );
  OAI22_X1 U1096 ( .A1(n982), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[3][6] ), 
        .B2(n981), .ZN(n980) );
  INV_X1 U1097 ( .A(n980), .ZN(n313) );
  OAI22_X1 U1098 ( .A1(n982), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[3][7] ), 
        .B2(n981), .ZN(n983) );
  INV_X1 U1099 ( .A(n983), .ZN(n312) );
  NOR2_X1 U1100 ( .A1(n984), .A2(n1006), .ZN(n992) );
  INV_X1 U1101 ( .A(n992), .ZN(n993) );
  OAI22_X1 U1102 ( .A1(n993), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[4][0] ), 
        .B2(n992), .ZN(n985) );
  INV_X1 U1103 ( .A(n985), .ZN(n311) );
  OAI22_X1 U1104 ( .A1(n993), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[4][1] ), 
        .B2(n992), .ZN(n986) );
  INV_X1 U1105 ( .A(n986), .ZN(n310) );
  OAI22_X1 U1106 ( .A1(n993), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[4][2] ), 
        .B2(n992), .ZN(n987) );
  INV_X1 U1107 ( .A(n987), .ZN(n309) );
  OAI22_X1 U1108 ( .A1(n993), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[4][3] ), 
        .B2(n992), .ZN(n988) );
  INV_X1 U1109 ( .A(n988), .ZN(n308) );
  OAI22_X1 U1110 ( .A1(n993), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[4][4] ), 
        .B2(n992), .ZN(n989) );
  INV_X1 U1111 ( .A(n989), .ZN(n307) );
  OAI22_X1 U1112 ( .A1(n993), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[4][5] ), 
        .B2(n992), .ZN(n990) );
  INV_X1 U1113 ( .A(n990), .ZN(n306) );
  OAI22_X1 U1114 ( .A1(n993), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[4][6] ), 
        .B2(n992), .ZN(n991) );
  INV_X1 U1115 ( .A(n991), .ZN(n305) );
  OAI22_X1 U1116 ( .A1(n993), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[4][7] ), 
        .B2(n992), .ZN(n994) );
  INV_X1 U1117 ( .A(n994), .ZN(n304) );
  NOR2_X1 U1118 ( .A1(n995), .A2(n1006), .ZN(n1003) );
  INV_X1 U1119 ( .A(n1003), .ZN(n1004) );
  OAI22_X1 U1120 ( .A1(n1004), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[5][0] ), 
        .B2(n1003), .ZN(n996) );
  INV_X1 U1121 ( .A(n996), .ZN(n303) );
  OAI22_X1 U1122 ( .A1(n1004), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[5][1] ), 
        .B2(n1003), .ZN(n997) );
  INV_X1 U1123 ( .A(n997), .ZN(n302) );
  OAI22_X1 U1124 ( .A1(n1004), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[5][2] ), 
        .B2(n1003), .ZN(n998) );
  INV_X1 U1125 ( .A(n998), .ZN(n301) );
  OAI22_X1 U1126 ( .A1(n1004), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[5][3] ), 
        .B2(n1003), .ZN(n999) );
  INV_X1 U1127 ( .A(n999), .ZN(n300) );
  OAI22_X1 U1128 ( .A1(n1004), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[5][4] ), 
        .B2(n1003), .ZN(n1000) );
  INV_X1 U1129 ( .A(n1000), .ZN(n299) );
  OAI22_X1 U1130 ( .A1(n1004), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[5][5] ), 
        .B2(n1003), .ZN(n1001) );
  INV_X1 U1131 ( .A(n1001), .ZN(n298) );
  OAI22_X1 U1132 ( .A1(n1004), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[5][6] ), 
        .B2(n1003), .ZN(n1002) );
  INV_X1 U1133 ( .A(n1002), .ZN(n297) );
  OAI22_X1 U1134 ( .A1(n1004), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[5][7] ), 
        .B2(n1003), .ZN(n1005) );
  INV_X1 U1135 ( .A(n1005), .ZN(n296) );
  NOR2_X1 U1136 ( .A1(n1007), .A2(n1006), .ZN(n1015) );
  INV_X1 U1137 ( .A(n1015), .ZN(n1016) );
  OAI22_X1 U1138 ( .A1(n1016), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[6][0] ), 
        .B2(n1015), .ZN(n1008) );
  INV_X1 U1139 ( .A(n1008), .ZN(n295) );
  OAI22_X1 U1140 ( .A1(n1016), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[6][1] ), 
        .B2(n1015), .ZN(n1009) );
  INV_X1 U1141 ( .A(n1009), .ZN(n294) );
  OAI22_X1 U1142 ( .A1(n1016), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[6][2] ), 
        .B2(n1015), .ZN(n1010) );
  INV_X1 U1143 ( .A(n1010), .ZN(n293) );
  OAI22_X1 U1144 ( .A1(n1016), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[6][3] ), 
        .B2(n1015), .ZN(n1011) );
  INV_X1 U1145 ( .A(n1011), .ZN(n292) );
  OAI22_X1 U1146 ( .A1(n1016), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[6][4] ), 
        .B2(n1015), .ZN(n1012) );
  INV_X1 U1147 ( .A(n1012), .ZN(n291) );
  OAI22_X1 U1148 ( .A1(n1016), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[6][5] ), 
        .B2(n1015), .ZN(n1013) );
  INV_X1 U1149 ( .A(n1013), .ZN(n290) );
  OAI22_X1 U1150 ( .A1(n1016), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[6][6] ), 
        .B2(n1015), .ZN(n1014) );
  INV_X1 U1151 ( .A(n1014), .ZN(n289) );
  OAI22_X1 U1152 ( .A1(n1016), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[6][7] ), 
        .B2(n1015), .ZN(n1017) );
  INV_X1 U1153 ( .A(n1017), .ZN(n288) );
  OAI22_X1 U1154 ( .A1(n1026), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[7][0] ), 
        .B2(n1025), .ZN(n1018) );
  INV_X1 U1155 ( .A(n1018), .ZN(n287) );
  OAI22_X1 U1156 ( .A1(n1026), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[7][1] ), 
        .B2(n1025), .ZN(n1019) );
  INV_X1 U1157 ( .A(n1019), .ZN(n286) );
  OAI22_X1 U1158 ( .A1(n1026), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[7][2] ), 
        .B2(n1025), .ZN(n1020) );
  INV_X1 U1159 ( .A(n1020), .ZN(n285) );
  OAI22_X1 U1160 ( .A1(n1026), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[7][3] ), 
        .B2(n1025), .ZN(n1021) );
  INV_X1 U1161 ( .A(n1021), .ZN(n284) );
  OAI22_X1 U1162 ( .A1(n1026), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[7][4] ), 
        .B2(n1025), .ZN(n1022) );
  INV_X1 U1163 ( .A(n1022), .ZN(n283) );
  OAI22_X1 U1164 ( .A1(n1026), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[7][5] ), 
        .B2(n1025), .ZN(n1023) );
  INV_X1 U1165 ( .A(n1023), .ZN(n282) );
  OAI22_X1 U1166 ( .A1(n1026), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[7][6] ), 
        .B2(n1025), .ZN(n1024) );
  INV_X1 U1167 ( .A(n1024), .ZN(n281) );
  OAI22_X1 U1168 ( .A1(n1026), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[7][7] ), 
        .B2(n1025), .ZN(n1027) );
  INV_X1 U1169 ( .A(n1027), .ZN(n280) );
endmodule

