
module conv_128_32_DW_mult_pipe_J1_0 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n356, n358,
         n360, n362, n364, n366, n368, n370, n372, n374, n376, n378, n380,
         n382, n384, n386, n388, n390, n392, n394, n396, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n408, n410, n412, n414, n416,
         n418, n420, n422, n424, n426, n428, n430, n432, n434, n436, n438,
         n440, n442, n444, n446, n448, n450, n452, n454, n456, n458, n460,
         n462, n464, n466, n468, n470, n472, n474, n476, n478, n480, n482,
         n484, n486, n488, n490, n492, n494, n496, n498, n500, n502, n504,
         n506, n508, n510, n512, n514, n516, n517, n519, n520, n522, n523,
         n525, n526, n528, n529, n531, n533, n535, n537, n539, n541, n543,
         n545, n547, n549, n551, n552, n553;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n404), .SE(n514), .CK(clk), .Q(n552), 
        .QN(n39) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n404), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n36) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n404), .SE(n506), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n329) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n404), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n404), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n26) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n404), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n404), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n35) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n405), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n32) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n406), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n404), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n31) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n404), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n34) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n404), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n33) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n404), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n404), .SE(n480), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n404), .SE(n478), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n404), .SE(n476), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n404), .SE(n474), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n404), .SE(n472), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n406), .SE(n470), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n404), .SE(n468), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n405), .SE(n466), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n404), .SE(n464), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n404), .SE(n462), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n404), .SE(n460), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n404), .SE(n458), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n404), .SE(n456), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n404), .SE(n454), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n404), .SE(n452), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n406), .SE(n450), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n406), .SE(n448), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n406), .SE(n446), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n406), .SE(n444), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n406), .SE(n442), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n406), .SE(n440), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n406), .SE(n438), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n406), .SE(n436), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n406), .SE(n434), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n406), .SE(n432), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n406), .SE(n430), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n405), .SE(n428), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n405), .SE(n426), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n405), .SE(n424), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n405), .SE(n422), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n405), .SE(n420), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n405), .SE(n418), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n405), .SE(n416), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n405), .SE(n414), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n405), .SE(n412), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n405), .SE(n410), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n405), .SE(n408), .CK(clk), .Q(
        product[0]) );
  SDFF_X2 clk_r_REG51_S1 ( .D(1'b0), .SI(n404), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n330) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n404), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n553), .SE(n396), .CK(
        clk), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n553), .SE(n394), .CK(
        clk), .QN(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n553), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n553), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n553), .SE(n388), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n553), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n348), .QN(n37) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2_IP  ( .D(1'b1), .SI(n553), .SE(n384), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n553), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n553), .SE(n380), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n553), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n553), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n343), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n553), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n342), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n553), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n553), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n340), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n553), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n339), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2  ( .D(n553), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n553), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n337), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n553), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n336), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n553), .SE(n360), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n553), .SE(n358), .CK(
        clk), .QN(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n553), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n553), .SE(n354), .CK(
        clk), .QN(n332) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n404), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n331) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n404), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n27) );
  INV_X1 U2 ( .A(n331), .ZN(n25) );
  INV_X1 U3 ( .A(n112), .ZN(n247) );
  BUF_X1 U4 ( .A(n404), .Z(n405) );
  INV_X2 U5 ( .A(n553), .ZN(n404) );
  BUF_X1 U6 ( .A(n49), .Z(n50) );
  INV_X1 U7 ( .A(n20), .ZN(n23) );
  INV_X1 U8 ( .A(n20), .ZN(n22) );
  INV_X1 U9 ( .A(n20), .ZN(n21) );
  NAND2_X1 U10 ( .A1(n15), .A2(n14), .ZN(n238) );
  INV_X1 U11 ( .A(n112), .ZN(n188) );
  NAND2_X1 U12 ( .A1(n239), .A2(n16), .ZN(n15) );
  BUF_X1 U13 ( .A(n404), .Z(n406) );
  NAND2_X1 U14 ( .A1(n240), .A2(n38), .ZN(n14) );
  OR2_X1 U15 ( .A1(n240), .A2(n38), .ZN(n16) );
  INV_X1 U16 ( .A(rst_n), .ZN(n553) );
  INV_X1 U17 ( .A(n46), .ZN(n146) );
  NAND2_X1 U18 ( .A1(\mult_x_1/n313 ), .A2(n26), .ZN(n209) );
  AND2_X1 U19 ( .A1(n552), .A2(\mult_x_1/n281 ), .ZN(n113) );
  NAND2_X1 U20 ( .A1(n8), .A2(n7), .ZN(n366) );
  NAND2_X1 U21 ( .A1(n112), .A2(n338), .ZN(n7) );
  NAND2_X1 U22 ( .A1(n9), .A2(n188), .ZN(n8) );
  NAND2_X1 U23 ( .A1(n175), .A2(n174), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n11), .A2(n10), .ZN(n390) );
  NAND2_X1 U25 ( .A1(n20), .A2(n350), .ZN(n10) );
  NAND2_X1 U26 ( .A1(n12), .A2(n247), .ZN(n11) );
  XNOR2_X1 U27 ( .A(n13), .B(n239), .ZN(n12) );
  XNOR2_X1 U28 ( .A(n240), .B(n38), .ZN(n13) );
  XNOR2_X1 U29 ( .A(n102), .B(n101), .ZN(n224) );
  XNOR2_X1 U30 ( .A(n100), .B(n99), .ZN(n101) );
  INV_X1 U31 ( .A(en), .ZN(n20) );
  XNOR2_X1 U32 ( .A(n220), .B(n219), .ZN(n222) );
  NAND2_X1 U33 ( .A1(n228), .A2(n227), .ZN(n229) );
  NAND2_X1 U34 ( .A1(n226), .A2(n225), .ZN(n227) );
  OAI21_X1 U35 ( .B1(n225), .B2(n226), .A(n224), .ZN(n228) );
  XNOR2_X1 U36 ( .A(n103), .B(n224), .ZN(n104) );
  INV_X1 U37 ( .A(n27), .ZN(n17) );
  INV_X1 U38 ( .A(\mult_x_1/n312 ), .ZN(n18) );
  XNOR2_X1 U39 ( .A(n329), .B(n330), .ZN(n19) );
  NAND2_X2 U40 ( .A1(n43), .A2(n19), .ZN(n136) );
  XNOR2_X1 U41 ( .A(n222), .B(n221), .ZN(n223) );
  XNOR2_X1 U42 ( .A(n226), .B(n225), .ZN(n103) );
  INV_X1 U43 ( .A(n28), .ZN(n24) );
  AND2_X1 U44 ( .A1(n231), .A2(n230), .ZN(n38) );
  XOR2_X1 U45 ( .A(n231), .B(n230), .Z(n40) );
  INV_X1 U46 ( .A(en), .ZN(n112) );
  OR2_X1 U47 ( .A1(n188), .A2(n37), .ZN(n41) );
  AND2_X1 U48 ( .A1(n57), .A2(n56), .ZN(n42) );
  XOR2_X1 U49 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n43) );
  XNOR2_X1 U50 ( .A(n329), .B(n330), .ZN(n44) );
  XNOR2_X1 U51 ( .A(n25), .B(\mult_x_1/n281 ), .ZN(n54) );
  XNOR2_X1 U52 ( .A(n113), .B(n25), .ZN(n66) );
  INV_X1 U53 ( .A(n44), .ZN(n45) );
  OAI22_X1 U54 ( .A1(n136), .A2(n54), .B1(n66), .B2(n44), .ZN(n116) );
  INV_X1 U55 ( .A(n116), .ZN(n64) );
  XNOR2_X1 U56 ( .A(n36), .B(n17), .ZN(n75) );
  XNOR2_X1 U57 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n74) );
  NAND2_X1 U58 ( .A1(n75), .A2(n74), .ZN(n145) );
  XNOR2_X1 U59 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n47) );
  INV_X1 U60 ( .A(n74), .ZN(n46) );
  XNOR2_X1 U61 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n65) );
  OAI22_X1 U62 ( .A1(n145), .A2(n47), .B1(n146), .B2(n65), .ZN(n63) );
  NAND2_X1 U63 ( .A1(n39), .A2(\mult_x_1/n310 ), .ZN(n148) );
  NOR2_X1 U64 ( .A1(n30), .A2(n148), .ZN(n62) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n53) );
  OAI22_X1 U66 ( .A1(n145), .A2(n53), .B1(n146), .B2(n47), .ZN(n98) );
  XOR2_X1 U67 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n48) );
  XNOR2_X1 U68 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n49) );
  NAND2_X2 U69 ( .A1(n48), .A2(n49), .ZN(n205) );
  XNOR2_X1 U70 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n81) );
  XNOR2_X1 U71 ( .A(n113), .B(\mult_x_1/n312 ), .ZN(n51) );
  OAI22_X1 U72 ( .A1(n205), .A2(n81), .B1(n51), .B2(n50), .ZN(n97) );
  AOI21_X1 U73 ( .B1(n50), .B2(n205), .A(n51), .ZN(n52) );
  INV_X1 U74 ( .A(n52), .ZN(n96) );
  XNOR2_X1 U75 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n76) );
  OAI22_X1 U76 ( .A1(n145), .A2(n76), .B1(n146), .B2(n53), .ZN(n234) );
  XNOR2_X1 U77 ( .A(n25), .B(\mult_x_1/n283 ), .ZN(n79) );
  XNOR2_X1 U78 ( .A(n25), .B(\mult_x_1/n282 ), .ZN(n55) );
  OAI22_X1 U79 ( .A1(n136), .A2(n79), .B1(n44), .B2(n55), .ZN(n233) );
  INV_X1 U80 ( .A(n97), .ZN(n232) );
  INV_X1 U81 ( .A(n102), .ZN(n59) );
  NOR2_X1 U82 ( .A1(n31), .A2(n148), .ZN(n100) );
  INV_X1 U83 ( .A(n100), .ZN(n57) );
  OAI22_X1 U84 ( .A1(n136), .A2(n55), .B1(n44), .B2(n54), .ZN(n99) );
  INV_X1 U85 ( .A(n99), .ZN(n56) );
  NAND2_X1 U86 ( .A1(n99), .A2(n100), .ZN(n58) );
  OAI21_X1 U87 ( .B1(n59), .B2(n42), .A(n58), .ZN(n221) );
  OAI21_X1 U88 ( .B1(n220), .B2(n219), .A(n221), .ZN(n61) );
  NAND2_X1 U89 ( .A1(n220), .A2(n219), .ZN(n60) );
  NAND2_X1 U90 ( .A1(n61), .A2(n60), .ZN(n193) );
  INV_X1 U91 ( .A(n193), .ZN(n69) );
  FA_X1 U92 ( .A(n64), .B(n63), .CI(n62), .CO(n120), .S(n220) );
  NOR2_X1 U93 ( .A1(n32), .A2(n148), .ZN(n119) );
  XNOR2_X1 U94 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n114) );
  OAI22_X1 U95 ( .A1(n145), .A2(n65), .B1(n146), .B2(n114), .ZN(n117) );
  AOI21_X1 U96 ( .B1(n44), .B2(n136), .A(n66), .ZN(n67) );
  INV_X1 U97 ( .A(n67), .ZN(n115) );
  INV_X1 U98 ( .A(n194), .ZN(n68) );
  NAND2_X1 U99 ( .A1(n69), .A2(n68), .ZN(n70) );
  NAND2_X1 U100 ( .A1(n70), .A2(n247), .ZN(n72) );
  NAND2_X1 U101 ( .A1(n20), .A2(n344), .ZN(n71) );
  NAND2_X1 U102 ( .A1(n72), .A2(n71), .ZN(n378) );
  XNOR2_X1 U103 ( .A(n113), .B(n24), .ZN(n86) );
  AOI21_X1 U104 ( .B1(n209), .B2(n26), .A(n86), .ZN(n73) );
  INV_X1 U105 ( .A(n73), .ZN(n95) );
  NAND2_X1 U106 ( .A1(n75), .A2(n74), .ZN(n85) );
  XNOR2_X1 U107 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n83) );
  OAI22_X1 U108 ( .A1(n85), .A2(n83), .B1(n146), .B2(n76), .ZN(n94) );
  NOR2_X1 U109 ( .A1(n33), .A2(n148), .ZN(n93) );
  XNOR2_X1 U110 ( .A(n25), .B(\mult_x_1/n285 ), .ZN(n127) );
  XNOR2_X1 U111 ( .A(n25), .B(\mult_x_1/n284 ), .ZN(n80) );
  OAI22_X1 U112 ( .A1(n136), .A2(n127), .B1(n44), .B2(n80), .ZN(n169) );
  XNOR2_X1 U113 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n130) );
  XNOR2_X1 U114 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n82) );
  OAI22_X1 U115 ( .A1(n205), .A2(n130), .B1(n50), .B2(n82), .ZN(n168) );
  OR2_X1 U116 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n77) );
  OAI22_X1 U117 ( .A1(n85), .A2(n27), .B1(n77), .B2(n146), .ZN(n126) );
  XNOR2_X1 U118 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n78) );
  XNOR2_X1 U119 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n84) );
  OAI22_X1 U120 ( .A1(n85), .A2(n78), .B1(n146), .B2(n84), .ZN(n125) );
  OAI22_X1 U121 ( .A1(n136), .A2(n80), .B1(n44), .B2(n79), .ZN(n92) );
  OAI22_X1 U122 ( .A1(n205), .A2(n82), .B1(n50), .B2(n81), .ZN(n91) );
  XNOR2_X1 U123 ( .A(n92), .B(n91), .ZN(n231) );
  OAI22_X1 U124 ( .A1(n85), .A2(n84), .B1(n146), .B2(n83), .ZN(n163) );
  XNOR2_X1 U125 ( .A(n24), .B(\mult_x_1/n281 ), .ZN(n128) );
  OAI22_X1 U126 ( .A1(n209), .A2(n128), .B1(n86), .B2(n26), .ZN(n162) );
  INV_X1 U127 ( .A(n148), .ZN(n87) );
  AND2_X1 U128 ( .A1(\mult_x_1/n288 ), .A2(n87), .ZN(n161) );
  NAND2_X1 U129 ( .A1(n88), .A2(n247), .ZN(n90) );
  NAND2_X1 U130 ( .A1(n112), .A2(n352), .ZN(n89) );
  NAND2_X1 U131 ( .A1(n90), .A2(n89), .ZN(n394) );
  OR2_X1 U132 ( .A1(n92), .A2(n91), .ZN(n237) );
  NOR2_X1 U133 ( .A1(n34), .A2(n148), .ZN(n236) );
  FA_X1 U134 ( .A(n95), .B(n94), .CI(n93), .CO(n235), .S(n242) );
  FA_X1 U135 ( .A(n98), .B(n97), .CI(n96), .CO(n219), .S(n225) );
  NAND2_X1 U136 ( .A1(n104), .A2(n247), .ZN(n105) );
  NAND2_X1 U137 ( .A1(n105), .A2(n41), .ZN(n386) );
  XNOR2_X1 U160 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n109) );
  XNOR2_X1 U161 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n124) );
  OAI22_X1 U162 ( .A1(n205), .A2(n109), .B1(n50), .B2(n124), .ZN(n184) );
  XNOR2_X1 U163 ( .A(n24), .B(\mult_x_1/n284 ), .ZN(n108) );
  XNOR2_X1 U164 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n122) );
  OAI22_X1 U165 ( .A1(n209), .A2(n108), .B1(n122), .B2(n26), .ZN(n183) );
  OR2_X1 U166 ( .A1(\mult_x_1/n288 ), .A2(n331), .ZN(n106) );
  OAI22_X1 U167 ( .A1(n136), .A2(n331), .B1(n106), .B2(n44), .ZN(n133) );
  XNOR2_X1 U168 ( .A(n25), .B(\mult_x_1/n288 ), .ZN(n107) );
  XNOR2_X1 U169 ( .A(n25), .B(\mult_x_1/n287 ), .ZN(n135) );
  OAI22_X1 U170 ( .A1(n136), .A2(n107), .B1(n44), .B2(n135), .ZN(n132) );
  XNOR2_X1 U171 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n201) );
  OAI22_X1 U172 ( .A1(n209), .A2(n201), .B1(n108), .B2(n26), .ZN(n198) );
  AND2_X1 U173 ( .A1(\mult_x_1/n288 ), .A2(n45), .ZN(n197) );
  XNOR2_X1 U174 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n199) );
  OAI22_X1 U175 ( .A1(n205), .A2(n199), .B1(n50), .B2(n109), .ZN(n196) );
  NOR2_X1 U176 ( .A1(n191), .A2(n190), .ZN(n111) );
  NAND2_X1 U177 ( .A1(n112), .A2(n332), .ZN(n110) );
  OAI21_X1 U178 ( .B1(n112), .B2(n111), .A(n110), .ZN(n354) );
  NOR2_X1 U179 ( .A1(n35), .A2(n148), .ZN(n143) );
  XNOR2_X1 U180 ( .A(n113), .B(\mult_x_1/n310 ), .ZN(n144) );
  OAI22_X1 U181 ( .A1(n145), .A2(n114), .B1(n144), .B2(n146), .ZN(n152) );
  INV_X1 U182 ( .A(n152), .ZN(n142) );
  FA_X1 U183 ( .A(n117), .B(n116), .CI(n115), .CO(n141), .S(n118) );
  FA_X1 U184 ( .A(n120), .B(n119), .CI(n118), .CO(n158), .S(n194) );
  OR2_X1 U185 ( .A1(n159), .A2(n158), .ZN(n121) );
  MUX2_X1 U186 ( .A(n333), .B(n121), .S(n188), .Z(n356) );
  XNOR2_X1 U187 ( .A(n24), .B(\mult_x_1/n282 ), .ZN(n129) );
  OAI22_X1 U188 ( .A1(n209), .A2(n122), .B1(n129), .B2(n26), .ZN(n139) );
  INV_X1 U189 ( .A(n146), .ZN(n123) );
  AND2_X1 U190 ( .A1(\mult_x_1/n288 ), .A2(n123), .ZN(n138) );
  XNOR2_X1 U191 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n131) );
  OAI22_X1 U192 ( .A1(n205), .A2(n124), .B1(n50), .B2(n131), .ZN(n137) );
  HA_X1 U193 ( .A(n126), .B(n125), .CO(n167), .S(n171) );
  XNOR2_X1 U194 ( .A(n25), .B(\mult_x_1/n286 ), .ZN(n134) );
  OAI22_X1 U195 ( .A1(n136), .A2(n134), .B1(n44), .B2(n127), .ZN(n166) );
  OAI22_X1 U196 ( .A1(n209), .A2(n129), .B1(n128), .B2(n26), .ZN(n165) );
  OAI22_X1 U197 ( .A1(n205), .A2(n131), .B1(n50), .B2(n130), .ZN(n164) );
  HA_X1 U198 ( .A(n133), .B(n132), .CO(n181), .S(n182) );
  OAI22_X1 U199 ( .A1(n136), .A2(n135), .B1(n44), .B2(n134), .ZN(n180) );
  FA_X1 U200 ( .A(n139), .B(n138), .CI(n137), .CO(n172), .S(n179) );
  OR2_X1 U201 ( .A1(n177), .A2(n176), .ZN(n140) );
  MUX2_X1 U202 ( .A(n334), .B(n140), .S(n188), .Z(n358) );
  FA_X1 U203 ( .A(n143), .B(n142), .CI(n141), .CO(n154), .S(n159) );
  AOI21_X1 U204 ( .B1(n146), .B2(n145), .A(n144), .ZN(n147) );
  INV_X1 U205 ( .A(n147), .ZN(n150) );
  NOR2_X1 U206 ( .A1(n29), .A2(n148), .ZN(n149) );
  XOR2_X1 U207 ( .A(n150), .B(n149), .Z(n151) );
  XOR2_X1 U208 ( .A(n152), .B(n151), .Z(n153) );
  OR2_X1 U209 ( .A1(n154), .A2(n153), .ZN(n156) );
  NAND2_X1 U210 ( .A1(n154), .A2(n153), .ZN(n155) );
  NAND2_X1 U211 ( .A1(n156), .A2(n155), .ZN(n157) );
  MUX2_X1 U212 ( .A(n335), .B(n157), .S(n188), .Z(n360) );
  NAND2_X1 U213 ( .A1(n159), .A2(n158), .ZN(n160) );
  MUX2_X1 U214 ( .A(n336), .B(n160), .S(n188), .Z(n362) );
  FA_X1 U215 ( .A(n163), .B(n162), .CI(n161), .CO(n230), .S(n246) );
  FA_X1 U216 ( .A(n166), .B(n165), .CI(n164), .CO(n245), .S(n170) );
  FA_X1 U217 ( .A(n169), .B(n168), .CI(n167), .CO(n241), .S(n244) );
  FA_X1 U218 ( .A(n172), .B(n171), .CI(n170), .CO(n174), .S(n177) );
  NOR2_X1 U219 ( .A1(n175), .A2(n174), .ZN(n173) );
  MUX2_X1 U220 ( .A(n337), .B(n173), .S(n188), .Z(n364) );
  NAND2_X1 U221 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2_X1 U222 ( .A(n339), .B(n178), .S(n188), .Z(n368) );
  FA_X1 U223 ( .A(n181), .B(n180), .CI(n179), .CO(n176), .S(n187) );
  FA_X1 U224 ( .A(n184), .B(n183), .CI(n182), .CO(n186), .S(n191) );
  NOR2_X1 U225 ( .A1(n187), .A2(n186), .ZN(n185) );
  MUX2_X1 U226 ( .A(n340), .B(n185), .S(n188), .Z(n370) );
  NAND2_X1 U227 ( .A1(n187), .A2(n186), .ZN(n189) );
  MUX2_X1 U228 ( .A(n341), .B(n189), .S(n188), .Z(n372) );
  NAND2_X1 U229 ( .A1(n191), .A2(n190), .ZN(n192) );
  MUX2_X1 U230 ( .A(n342), .B(n192), .S(n247), .Z(n374) );
  NAND2_X1 U231 ( .A1(n194), .A2(n193), .ZN(n195) );
  MUX2_X1 U232 ( .A(n343), .B(n195), .S(n247), .Z(n376) );
  FA_X1 U233 ( .A(n198), .B(n197), .CI(n196), .CO(n190), .S(n217) );
  XNOR2_X1 U234 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n200) );
  OAI22_X1 U235 ( .A1(n205), .A2(n200), .B1(n50), .B2(n199), .ZN(n203) );
  XNOR2_X1 U236 ( .A(n24), .B(\mult_x_1/n286 ), .ZN(n206) );
  OAI22_X1 U237 ( .A1(n209), .A2(n206), .B1(n201), .B2(n26), .ZN(n202) );
  NOR2_X1 U238 ( .A1(n217), .A2(n216), .ZN(n265) );
  HA_X1 U239 ( .A(n203), .B(n202), .CO(n216), .S(n214) );
  OR2_X1 U240 ( .A1(\mult_x_1/n288 ), .A2(n18), .ZN(n204) );
  OAI22_X1 U241 ( .A1(n205), .A2(n18), .B1(n204), .B2(n50), .ZN(n213) );
  OR2_X1 U242 ( .A1(n214), .A2(n213), .ZN(n261) );
  XNOR2_X1 U243 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n208) );
  OAI22_X1 U244 ( .A1(n209), .A2(n208), .B1(n206), .B2(n26), .ZN(n212) );
  INV_X1 U245 ( .A(n50), .ZN(n207) );
  AND2_X1 U246 ( .A1(\mult_x_1/n288 ), .A2(n207), .ZN(n211) );
  NOR2_X1 U247 ( .A1(n212), .A2(n211), .ZN(n254) );
  OAI22_X1 U248 ( .A1(n209), .A2(\mult_x_1/n288 ), .B1(n208), .B2(n26), .ZN(
        n251) );
  OR2_X1 U249 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n210) );
  NAND2_X1 U250 ( .A1(n210), .A2(n209), .ZN(n250) );
  NAND2_X1 U251 ( .A1(n251), .A2(n250), .ZN(n257) );
  NAND2_X1 U252 ( .A1(n212), .A2(n211), .ZN(n255) );
  OAI21_X1 U253 ( .B1(n254), .B2(n257), .A(n255), .ZN(n262) );
  NAND2_X1 U254 ( .A1(n214), .A2(n213), .ZN(n260) );
  INV_X1 U255 ( .A(n260), .ZN(n215) );
  AOI21_X1 U256 ( .B1(n261), .B2(n262), .A(n215), .ZN(n268) );
  NAND2_X1 U257 ( .A1(n217), .A2(n216), .ZN(n266) );
  OAI21_X1 U258 ( .B1(n265), .B2(n268), .A(n266), .ZN(n218) );
  MUX2_X1 U259 ( .A(n345), .B(n218), .S(n247), .Z(n380) );
  MUX2_X1 U260 ( .A(n346), .B(n223), .S(n247), .Z(n382) );
  MUX2_X1 U261 ( .A(n347), .B(n229), .S(n247), .Z(n384) );
  FA_X1 U262 ( .A(n234), .B(n233), .CI(n232), .CO(n102), .S(n240) );
  FA_X1 U263 ( .A(n237), .B(n236), .CI(n235), .CO(n226), .S(n239) );
  MUX2_X1 U264 ( .A(n349), .B(n238), .S(n247), .Z(n388) );
  FA_X1 U265 ( .A(n242), .B(n241), .CI(n40), .CO(n243), .S(n88) );
  MUX2_X1 U266 ( .A(n351), .B(n243), .S(n247), .Z(n392) );
  FA_X1 U267 ( .A(n246), .B(n245), .CI(n244), .CO(n248), .S(n175) );
  MUX2_X1 U268 ( .A(n353), .B(n248), .S(n247), .Z(n396) );
  MUX2_X1 U269 ( .A(product[0]), .B(n516), .S(n21), .Z(n408) );
  MUX2_X1 U270 ( .A(n516), .B(n517), .S(n188), .Z(n410) );
  AND2_X1 U271 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n249) );
  MUX2_X1 U272 ( .A(n517), .B(n249), .S(n21), .Z(n412) );
  MUX2_X1 U273 ( .A(product[1]), .B(n519), .S(n21), .Z(n414) );
  MUX2_X1 U274 ( .A(n519), .B(n520), .S(n22), .Z(n416) );
  OR2_X1 U275 ( .A1(n251), .A2(n250), .ZN(n252) );
  AND2_X1 U276 ( .A1(n252), .A2(n257), .ZN(n253) );
  MUX2_X1 U277 ( .A(n520), .B(n253), .S(n247), .Z(n418) );
  MUX2_X1 U278 ( .A(product[2]), .B(n522), .S(n23), .Z(n420) );
  MUX2_X1 U279 ( .A(n522), .B(n523), .S(n22), .Z(n422) );
  INV_X1 U280 ( .A(n254), .ZN(n256) );
  NAND2_X1 U281 ( .A1(n256), .A2(n255), .ZN(n258) );
  XOR2_X1 U282 ( .A(n258), .B(n257), .Z(n259) );
  MUX2_X1 U283 ( .A(n523), .B(n259), .S(n23), .Z(n424) );
  MUX2_X1 U284 ( .A(product[3]), .B(n525), .S(en), .Z(n426) );
  MUX2_X1 U285 ( .A(n525), .B(n526), .S(n22), .Z(n428) );
  NAND2_X1 U286 ( .A1(n261), .A2(n260), .ZN(n263) );
  XNOR2_X1 U287 ( .A(n263), .B(n262), .ZN(n264) );
  MUX2_X1 U288 ( .A(n526), .B(n264), .S(en), .Z(n430) );
  MUX2_X1 U289 ( .A(product[4]), .B(n528), .S(n23), .Z(n432) );
  MUX2_X1 U290 ( .A(n528), .B(n529), .S(en), .Z(n434) );
  INV_X1 U291 ( .A(n265), .ZN(n267) );
  NAND2_X1 U292 ( .A1(n267), .A2(n266), .ZN(n269) );
  XOR2_X1 U293 ( .A(n269), .B(n268), .Z(n270) );
  MUX2_X1 U294 ( .A(n529), .B(n270), .S(n23), .Z(n436) );
  MUX2_X1 U295 ( .A(product[5]), .B(n531), .S(en), .Z(n438) );
  NAND2_X1 U296 ( .A1(n332), .A2(n342), .ZN(n271) );
  XNOR2_X1 U297 ( .A(n271), .B(n345), .ZN(n272) );
  MUX2_X1 U298 ( .A(n531), .B(n272), .S(n23), .Z(n440) );
  MUX2_X1 U299 ( .A(product[6]), .B(n533), .S(n23), .Z(n442) );
  NAND2_X1 U300 ( .A1(n399), .A2(n341), .ZN(n273) );
  AOI21_X1 U301 ( .B1(n332), .B2(n345), .A(n402), .ZN(n275) );
  XOR2_X1 U302 ( .A(n273), .B(n275), .Z(n274) );
  MUX2_X1 U303 ( .A(n533), .B(n274), .S(n22), .Z(n444) );
  MUX2_X1 U304 ( .A(product[7]), .B(n535), .S(n22), .Z(n446) );
  OAI21_X1 U305 ( .B1(n340), .B2(n275), .A(n341), .ZN(n278) );
  NAND2_X1 U306 ( .A1(n334), .A2(n339), .ZN(n276) );
  XNOR2_X1 U307 ( .A(n278), .B(n276), .ZN(n277) );
  MUX2_X1 U308 ( .A(n535), .B(n277), .S(n22), .Z(n448) );
  MUX2_X1 U309 ( .A(product[8]), .B(n537), .S(n22), .Z(n450) );
  AOI21_X1 U310 ( .B1(n278), .B2(n334), .A(n401), .ZN(n281) );
  NAND2_X1 U311 ( .A1(n403), .A2(n338), .ZN(n279) );
  XOR2_X1 U312 ( .A(n281), .B(n279), .Z(n280) );
  MUX2_X1 U313 ( .A(n537), .B(n280), .S(n23), .Z(n452) );
  MUX2_X1 U314 ( .A(product[9]), .B(n539), .S(n22), .Z(n454) );
  OAI21_X1 U315 ( .B1(n281), .B2(n337), .A(n338), .ZN(n295) );
  INV_X1 U316 ( .A(n295), .ZN(n285) );
  NOR2_X1 U317 ( .A1(n352), .A2(n353), .ZN(n290) );
  INV_X1 U318 ( .A(n290), .ZN(n282) );
  NAND2_X1 U319 ( .A1(n352), .A2(n353), .ZN(n292) );
  NAND2_X1 U320 ( .A1(n282), .A2(n292), .ZN(n283) );
  XOR2_X1 U321 ( .A(n285), .B(n283), .Z(n284) );
  MUX2_X1 U322 ( .A(n539), .B(n284), .S(n23), .Z(n456) );
  MUX2_X1 U323 ( .A(product[10]), .B(n541), .S(n22), .Z(n458) );
  OAI21_X1 U324 ( .B1(n285), .B2(n290), .A(n292), .ZN(n288) );
  NOR2_X1 U325 ( .A1(n350), .A2(n351), .ZN(n293) );
  INV_X1 U326 ( .A(n293), .ZN(n286) );
  NAND2_X1 U327 ( .A1(n350), .A2(n351), .ZN(n291) );
  NAND2_X1 U328 ( .A1(n286), .A2(n291), .ZN(n287) );
  XNOR2_X1 U329 ( .A(n288), .B(n287), .ZN(n289) );
  MUX2_X1 U330 ( .A(n541), .B(n289), .S(n23), .Z(n460) );
  MUX2_X1 U331 ( .A(product[11]), .B(n543), .S(n22), .Z(n462) );
  NOR2_X1 U332 ( .A1(n293), .A2(n290), .ZN(n296) );
  OAI21_X1 U333 ( .B1(n293), .B2(n292), .A(n291), .ZN(n294) );
  AOI21_X1 U334 ( .B1(n296), .B2(n295), .A(n294), .ZN(n326) );
  NOR2_X1 U335 ( .A1(n348), .A2(n349), .ZN(n312) );
  INV_X1 U336 ( .A(n312), .ZN(n302) );
  NAND2_X1 U337 ( .A1(n348), .A2(n349), .ZN(n315) );
  NAND2_X1 U338 ( .A1(n302), .A2(n315), .ZN(n297) );
  XOR2_X1 U339 ( .A(n326), .B(n297), .Z(n298) );
  MUX2_X1 U340 ( .A(n543), .B(n298), .S(n23), .Z(n464) );
  MUX2_X1 U341 ( .A(product[12]), .B(n545), .S(n22), .Z(n466) );
  OAI21_X1 U342 ( .B1(n326), .B2(n312), .A(n315), .ZN(n300) );
  OR2_X1 U343 ( .A1(n346), .A2(n347), .ZN(n304) );
  NAND2_X1 U344 ( .A1(n346), .A2(n347), .ZN(n303) );
  NAND2_X1 U345 ( .A1(n304), .A2(n303), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  MUX2_X1 U347 ( .A(n545), .B(n301), .S(n23), .Z(n468) );
  MUX2_X1 U348 ( .A(product[13]), .B(n547), .S(n22), .Z(n470) );
  NAND2_X1 U349 ( .A1(n302), .A2(n304), .ZN(n307) );
  INV_X1 U350 ( .A(n315), .ZN(n305) );
  INV_X1 U351 ( .A(n303), .ZN(n313) );
  AOI21_X1 U352 ( .B1(n305), .B2(n304), .A(n313), .ZN(n306) );
  OAI21_X1 U353 ( .B1(n326), .B2(n307), .A(n306), .ZN(n309) );
  NAND2_X1 U354 ( .A1(n344), .A2(n343), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U356 ( .A(n547), .B(n310), .S(n23), .Z(n472) );
  MUX2_X1 U357 ( .A(product[14]), .B(n549), .S(n22), .Z(n474) );
  OR2_X1 U358 ( .A1(n346), .A2(n347), .ZN(n311) );
  NAND2_X1 U359 ( .A1(n311), .A2(n344), .ZN(n316) );
  NOR2_X1 U360 ( .A1(n312), .A2(n316), .ZN(n322) );
  INV_X1 U361 ( .A(n322), .ZN(n318) );
  AOI21_X1 U362 ( .B1(n313), .B2(n344), .A(n400), .ZN(n314) );
  OAI21_X1 U363 ( .B1(n316), .B2(n315), .A(n314), .ZN(n323) );
  INV_X1 U364 ( .A(n323), .ZN(n317) );
  OAI21_X1 U365 ( .B1(n326), .B2(n318), .A(n317), .ZN(n320) );
  NAND2_X1 U366 ( .A1(n333), .A2(n336), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U368 ( .A(n549), .B(n321), .S(n23), .Z(n476) );
  MUX2_X1 U369 ( .A(product[15]), .B(n551), .S(n22), .Z(n478) );
  NAND2_X1 U370 ( .A1(n322), .A2(n333), .ZN(n325) );
  AOI21_X1 U371 ( .B1(n323), .B2(n333), .A(n398), .ZN(n324) );
  OAI21_X1 U372 ( .B1(n326), .B2(n325), .A(n324), .ZN(n327) );
  XNOR2_X1 U373 ( .A(n327), .B(n335), .ZN(n328) );
  MUX2_X1 U374 ( .A(n551), .B(n328), .S(n21), .Z(n480) );
  MUX2_X1 U375 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n21), .Z(n482) );
  MUX2_X1 U376 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n21), .Z(n484) );
  MUX2_X1 U377 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n21), .Z(n486) );
  MUX2_X1 U378 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n21), .Z(n488) );
  MUX2_X1 U379 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n21), .Z(n490) );
  MUX2_X1 U380 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n21), .Z(n492) );
  MUX2_X1 U381 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n188), .Z(n494) );
  MUX2_X1 U382 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n21), .Z(n496) );
  MUX2_X1 U383 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n188), .Z(n498) );
  MUX2_X1 U384 ( .A(n24), .B(A_extended[1]), .S(n21), .Z(n500) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n21), .Z(n502) );
  MUX2_X1 U386 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n22), .Z(n504) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n21), .Z(n506) );
  MUX2_X1 U388 ( .A(n25), .B(A_extended[5]), .S(n21), .Z(n508) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n188), .Z(n510) );
  MUX2_X1 U390 ( .A(\mult_x_1/n310 ), .B(A_extended[7]), .S(n23), .Z(n512) );
  OR2_X1 U391 ( .A1(en), .A2(n552), .ZN(n514) );
endmodule


module conv_128_32_DW_mult_pipe_J1_1 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n346, n348, n350,
         n352, n354, n356, n358, n360, n362, n364, n366, n368, n370, n372,
         n374, n376, n378, n380, n382, n384, n386, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n400, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n420, n422, n424, n426, n428,
         n430, n432, n434, n436, n438, n440, n442, n444, n446, n448, n450,
         n452, n454, n456, n458, n460, n462, n464, n466, n468, n470, n472,
         n474, n476, n478, n480, n482, n484, n486, n488, n490, n492, n494,
         n496, n498, n500, n502, n504, n506, n508, n509, n511, n512, n514,
         n515, n517, n518, n520, n521, n523, n525, n527, n529, n531, n533,
         n535, n537, n539, n541, n543, n544, n545, n546;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n396), .SE(n506), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n396), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n22) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n396), .SE(n498), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n396), .SE(n494), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n5) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n396), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n10) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n396), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n14) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n396), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n15) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n397), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n17) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n398), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n16) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n396), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n18) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n396), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n20) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n396), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n19) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n396), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n12) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n396), .SE(n472), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n396), .SE(n470), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n396), .SE(n468), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n396), .SE(n466), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n396), .SE(n464), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n398), .SE(n462), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n396), .SE(n460), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n397), .SE(n458), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n396), .SE(n456), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n396), .SE(n454), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n396), .SE(n452), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n396), .SE(n450), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n396), .SE(n448), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n396), .SE(n446), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n396), .SE(n444), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n398), .SE(n442), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n398), .SE(n440), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n398), .SE(n438), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n398), .SE(n436), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n398), .SE(n434), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n398), .SE(n432), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n398), .SE(n430), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n398), .SE(n428), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n398), .SE(n426), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n398), .SE(n424), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n398), .SE(n422), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n397), .SE(n420), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n397), .SE(n418), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n397), .SE(n416), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n397), .SE(n414), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n397), .SE(n412), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n397), .SE(n410), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n397), .SE(n408), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n397), .SE(n406), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n397), .SE(n404), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n397), .SE(n402), .CK(clk), .Q(n508)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n397), .SE(n400), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n396), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n546), .SE(n386), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2_IP  ( .D(1'b1), .SI(n546), .SE(n384), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n546), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n546), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n546), .SE(n378), .CK(
        clk), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n546), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n546), .SE(n374), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n546), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n336), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n546), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n335), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n546), .SE(n368), .CK(
        clk), .Q(n390), .QN(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n546), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n333), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n546), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n546), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n331), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n546), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n330), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n546), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n546), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n328), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n546), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n327), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n546), .SE(n352), .CK(
        clk), .QN(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n546), .SE(n350), .CK(
        clk), .QN(n325) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n546), .SI(1'b1), .SE(n348), .CK(clk), 
        .Q(n324) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n546), .SI(1'b1), .SE(n346), .CK(clk), 
        .Q(n323) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n546), .SE(n344), .CK(
        clk), .QN(n322) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n396), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n11) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n396), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n23) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n396), .SE(n500), .CK(clk), .Q(n544), 
        .QN(n21) );
  BUF_X1 U2 ( .A(n396), .Z(n397) );
  INV_X2 U3 ( .A(n546), .ZN(n396) );
  INV_X1 U4 ( .A(n36), .ZN(n186) );
  NAND2_X1 U5 ( .A1(n30), .A2(n31), .ZN(n151) );
  INV_X1 U6 ( .A(n23), .ZN(n8) );
  BUF_X2 U7 ( .A(en), .Z(n267) );
  BUF_X1 U8 ( .A(n396), .Z(n398) );
  INV_X1 U9 ( .A(rst_n), .ZN(n546) );
  NAND2_X1 U10 ( .A1(n34), .A2(n35), .ZN(n184) );
  NAND2_X1 U11 ( .A1(n230), .A2(n229), .ZN(n231) );
  INV_X1 U12 ( .A(n236), .ZN(n230) );
  INV_X1 U13 ( .A(n235), .ZN(n229) );
  INV_X1 U14 ( .A(n211), .ZN(n157) );
  NAND2_X1 U15 ( .A1(n211), .A2(n210), .ZN(n159) );
  AND2_X1 U16 ( .A1(n545), .A2(\mult_x_1/n310 ), .ZN(n29) );
  NAND2_X1 U17 ( .A1(n228), .A2(n227), .ZN(n235) );
  NAND2_X1 U18 ( .A1(n224), .A2(n223), .ZN(n228) );
  NAND2_X1 U19 ( .A1(n160), .A2(n159), .ZN(n200) );
  XNOR2_X1 U20 ( .A(n165), .B(n164), .ZN(n166) );
  XNOR2_X1 U21 ( .A(n224), .B(n42), .ZN(n239) );
  NAND2_X1 U22 ( .A1(n233), .A2(n232), .ZN(n234) );
  NAND2_X1 U23 ( .A1(n236), .A2(n235), .ZN(n232) );
  NAND2_X1 U24 ( .A1(n13), .A2(n231), .ZN(n233) );
  XNOR2_X1 U25 ( .A(n13), .B(n237), .ZN(n238) );
  XNOR2_X1 U26 ( .A(n236), .B(n235), .ZN(n237) );
  XNOR2_X1 U27 ( .A(n5), .B(n25), .ZN(n35) );
  OAI22_X1 U28 ( .A1(n184), .A2(n152), .B1(n79), .B2(n186), .ZN(n6) );
  INV_X1 U29 ( .A(n11), .ZN(n7) );
  NAND2_X1 U30 ( .A1(n226), .A2(n225), .ZN(n227) );
  XNOR2_X1 U31 ( .A(n226), .B(n225), .ZN(n42) );
  OR2_X1 U32 ( .A1(n226), .A2(n225), .ZN(n223) );
  INV_X1 U33 ( .A(n21), .ZN(n9) );
  XNOR2_X1 U34 ( .A(n167), .B(n166), .ZN(n198) );
  OAI22_X1 U35 ( .A1(n184), .A2(n152), .B1(n79), .B2(n186), .ZN(n162) );
  INV_X1 U36 ( .A(en), .ZN(n133) );
  INV_X2 U37 ( .A(n133), .ZN(n242) );
  XOR2_X1 U38 ( .A(n219), .B(n218), .Z(n13) );
  AND2_X1 U39 ( .A1(n219), .A2(n218), .ZN(n24) );
  XNOR2_X1 U40 ( .A(\mult_x_1/a[6] ), .B(n544), .ZN(n27) );
  XNOR2_X1 U41 ( .A(\mult_x_1/n310 ), .B(n22), .ZN(n26) );
  NAND2_X1 U42 ( .A1(n27), .A2(n26), .ZN(n146) );
  XNOR2_X1 U43 ( .A(n7), .B(\mult_x_1/n287 ), .ZN(n38) );
  INV_X1 U44 ( .A(n27), .ZN(n28) );
  INV_X2 U45 ( .A(n28), .ZN(n144) );
  XNOR2_X1 U46 ( .A(n7), .B(\mult_x_1/n286 ), .ZN(n145) );
  OAI22_X1 U47 ( .A1(n146), .A2(n38), .B1(n144), .B2(n145), .ZN(n206) );
  NAND2_X1 U48 ( .A1(\mult_x_1/n313 ), .A2(n10), .ZN(n188) );
  XNOR2_X1 U49 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n33) );
  AND2_X1 U50 ( .A1(n545), .A2(\mult_x_1/n281 ), .ZN(n78) );
  XNOR2_X1 U51 ( .A(n78), .B(\mult_x_1/n313 ), .ZN(n141) );
  OAI22_X1 U52 ( .A1(n188), .A2(n33), .B1(n141), .B2(n10), .ZN(n205) );
  XNOR2_X1 U53 ( .A(n29), .B(\mult_x_1/n310 ), .ZN(n147) );
  NOR2_X1 U54 ( .A1(n147), .A2(n12), .ZN(n204) );
  XOR2_X1 U55 ( .A(\mult_x_1/a[4] ), .B(n544), .Z(n30) );
  XNOR2_X1 U56 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n31) );
  XNOR2_X1 U57 ( .A(n9), .B(\mult_x_1/n286 ), .ZN(n95) );
  INV_X1 U58 ( .A(n31), .ZN(n32) );
  INV_X2 U59 ( .A(n32), .ZN(n149) );
  XNOR2_X1 U60 ( .A(n9), .B(\mult_x_1/n285 ), .ZN(n40) );
  OAI22_X1 U61 ( .A1(n151), .A2(n95), .B1(n149), .B2(n40), .ZN(n50) );
  XNOR2_X1 U62 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n43) );
  OAI22_X1 U63 ( .A1(n188), .A2(n43), .B1(n33), .B2(n10), .ZN(n49) );
  XOR2_X1 U64 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n34) );
  XNOR2_X1 U65 ( .A(n8), .B(\mult_x_1/n284 ), .ZN(n45) );
  INV_X1 U66 ( .A(n35), .ZN(n36) );
  XNOR2_X1 U67 ( .A(n8), .B(\mult_x_1/n283 ), .ZN(n41) );
  OAI22_X1 U68 ( .A1(n184), .A2(n45), .B1(n186), .B2(n41), .ZN(n48) );
  OR2_X1 U69 ( .A1(\mult_x_1/n288 ), .A2(n11), .ZN(n37) );
  OAI22_X1 U70 ( .A1(n146), .A2(n11), .B1(n37), .B2(n144), .ZN(n47) );
  XNOR2_X1 U71 ( .A(n7), .B(\mult_x_1/n288 ), .ZN(n39) );
  OAI22_X1 U72 ( .A1(n146), .A2(n39), .B1(n144), .B2(n38), .ZN(n46) );
  XNOR2_X1 U73 ( .A(n544), .B(\mult_x_1/n284 ), .ZN(n150) );
  OAI22_X1 U74 ( .A1(n151), .A2(n40), .B1(n149), .B2(n150), .ZN(n226) );
  XNOR2_X1 U75 ( .A(n8), .B(\mult_x_1/n282 ), .ZN(n153) );
  OAI22_X1 U76 ( .A1(n184), .A2(n41), .B1(n186), .B2(n153), .ZN(n225) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n55) );
  OAI22_X1 U78 ( .A1(n188), .A2(n55), .B1(n43), .B2(n10), .ZN(n99) );
  INV_X1 U79 ( .A(n144), .ZN(n44) );
  AND2_X1 U80 ( .A1(\mult_x_1/n288 ), .A2(n44), .ZN(n98) );
  XNOR2_X1 U81 ( .A(n8), .B(\mult_x_1/n285 ), .ZN(n54) );
  OAI22_X1 U82 ( .A1(n184), .A2(n54), .B1(n186), .B2(n45), .ZN(n97) );
  HA_X1 U83 ( .A(n47), .B(n46), .CO(n224), .S(n91) );
  FA_X1 U84 ( .A(n50), .B(n49), .CI(n48), .CO(n240), .S(n90) );
  NAND2_X1 U85 ( .A1(n119), .A2(n118), .ZN(n51) );
  NAND2_X1 U86 ( .A1(n51), .A2(n242), .ZN(n53) );
  NAND2_X1 U87 ( .A1(n133), .A2(n329), .ZN(n52) );
  NAND2_X1 U88 ( .A1(n53), .A2(n52), .ZN(n358) );
  XNOR2_X1 U111 ( .A(n8), .B(\mult_x_1/n286 ), .ZN(n60) );
  OAI22_X1 U112 ( .A1(n184), .A2(n60), .B1(n186), .B2(n54), .ZN(n129) );
  XNOR2_X1 U113 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n58) );
  OAI22_X1 U114 ( .A1(n188), .A2(n58), .B1(n55), .B2(n10), .ZN(n128) );
  OR2_X1 U115 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n56) );
  OAI22_X1 U116 ( .A1(n151), .A2(n21), .B1(n56), .B2(n149), .ZN(n94) );
  XNOR2_X1 U117 ( .A(n9), .B(\mult_x_1/n288 ), .ZN(n57) );
  XNOR2_X1 U118 ( .A(n9), .B(\mult_x_1/n287 ), .ZN(n96) );
  OAI22_X1 U119 ( .A1(n151), .A2(n57), .B1(n149), .B2(n96), .ZN(n93) );
  XNOR2_X1 U120 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n180) );
  OAI22_X1 U121 ( .A1(n188), .A2(n180), .B1(n58), .B2(n10), .ZN(n177) );
  INV_X1 U122 ( .A(n149), .ZN(n59) );
  AND2_X1 U123 ( .A1(\mult_x_1/n288 ), .A2(n59), .ZN(n176) );
  XNOR2_X1 U124 ( .A(n8), .B(\mult_x_1/n287 ), .ZN(n178) );
  OAI22_X1 U125 ( .A1(n184), .A2(n178), .B1(n186), .B2(n60), .ZN(n175) );
  NOR2_X1 U126 ( .A1(n136), .A2(n135), .ZN(n62) );
  NAND2_X1 U127 ( .A1(n133), .A2(n322), .ZN(n61) );
  OAI21_X1 U128 ( .B1(n133), .B2(n62), .A(n61), .ZN(n344) );
  NOR2_X1 U129 ( .A1(n15), .A2(n147), .ZN(n103) );
  XNOR2_X1 U130 ( .A(n7), .B(\mult_x_1/n281 ), .ZN(n63) );
  XNOR2_X1 U131 ( .A(n78), .B(n7), .ZN(n104) );
  OAI22_X1 U132 ( .A1(n146), .A2(n63), .B1(n104), .B2(n144), .ZN(n109) );
  INV_X1 U133 ( .A(n109), .ZN(n102) );
  XNOR2_X1 U134 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n66) );
  OAI22_X1 U135 ( .A1(n146), .A2(n66), .B1(n144), .B2(n63), .ZN(n69) );
  XNOR2_X1 U136 ( .A(n78), .B(n544), .ZN(n65) );
  AOI21_X1 U137 ( .B1(n149), .B2(n151), .A(n65), .ZN(n64) );
  INV_X1 U138 ( .A(n64), .ZN(n68) );
  XNOR2_X1 U139 ( .A(n9), .B(\mult_x_1/n281 ), .ZN(n82) );
  OAI22_X1 U140 ( .A1(n151), .A2(n82), .B1(n65), .B2(n149), .ZN(n67) );
  NOR2_X1 U141 ( .A1(n16), .A2(n147), .ZN(n76) );
  XNOR2_X1 U142 ( .A(n7), .B(\mult_x_1/n283 ), .ZN(n77) );
  OAI22_X1 U143 ( .A1(n146), .A2(n77), .B1(n144), .B2(n66), .ZN(n75) );
  INV_X1 U144 ( .A(n67), .ZN(n74) );
  NOR2_X1 U145 ( .A1(n17), .A2(n147), .ZN(n72) );
  FA_X1 U146 ( .A(n69), .B(n67), .CI(n68), .CO(n101), .S(n71) );
  OR2_X1 U147 ( .A1(n116), .A2(n115), .ZN(n70) );
  MUX2_X1 U148 ( .A(n323), .B(n70), .S(n267), .Z(n346) );
  FA_X1 U149 ( .A(n73), .B(n72), .CI(n71), .CO(n115), .S(n170) );
  FA_X1 U150 ( .A(n76), .B(n75), .CI(n74), .CO(n73), .S(n140) );
  XNOR2_X1 U151 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n81) );
  OAI22_X1 U152 ( .A1(n146), .A2(n81), .B1(n144), .B2(n77), .ZN(n163) );
  XNOR2_X1 U153 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n152) );
  XNOR2_X1 U154 ( .A(n78), .B(\mult_x_1/n312 ), .ZN(n79) );
  AOI21_X1 U155 ( .B1(n186), .B2(n184), .A(n79), .ZN(n80) );
  INV_X1 U156 ( .A(n80), .ZN(n161) );
  XNOR2_X1 U157 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n143) );
  OAI22_X1 U158 ( .A1(n146), .A2(n143), .B1(n144), .B2(n81), .ZN(n209) );
  XNOR2_X1 U159 ( .A(n544), .B(\mult_x_1/n283 ), .ZN(n148) );
  XNOR2_X1 U160 ( .A(n9), .B(\mult_x_1/n282 ), .ZN(n83) );
  OAI22_X1 U161 ( .A1(n151), .A2(n148), .B1(n149), .B2(n83), .ZN(n208) );
  INV_X1 U162 ( .A(n162), .ZN(n207) );
  NOR2_X1 U163 ( .A1(n18), .A2(n147), .ZN(n165) );
  INV_X1 U164 ( .A(n165), .ZN(n85) );
  OAI22_X1 U165 ( .A1(n151), .A2(n83), .B1(n149), .B2(n82), .ZN(n164) );
  INV_X1 U166 ( .A(n164), .ZN(n84) );
  NAND2_X1 U167 ( .A1(n85), .A2(n84), .ZN(n86) );
  NAND2_X1 U168 ( .A1(n167), .A2(n86), .ZN(n88) );
  NAND2_X1 U169 ( .A1(n165), .A2(n164), .ZN(n87) );
  NAND2_X1 U170 ( .A1(n88), .A2(n87), .ZN(n138) );
  OR2_X1 U171 ( .A1(n170), .A2(n169), .ZN(n89) );
  MUX2_X1 U172 ( .A(n324), .B(n89), .S(n267), .Z(n348) );
  FA_X1 U173 ( .A(n92), .B(n91), .CI(n90), .CO(n118), .S(n122) );
  HA_X1 U174 ( .A(n94), .B(n93), .CO(n126), .S(n127) );
  OAI22_X1 U175 ( .A1(n151), .A2(n96), .B1(n149), .B2(n95), .ZN(n125) );
  FA_X1 U176 ( .A(n99), .B(n98), .CI(n97), .CO(n92), .S(n124) );
  OR2_X1 U177 ( .A1(n122), .A2(n121), .ZN(n100) );
  MUX2_X1 U178 ( .A(n325), .B(n100), .S(n267), .Z(n350) );
  FA_X1 U179 ( .A(n103), .B(n102), .CI(n101), .CO(n111), .S(n116) );
  AOI21_X1 U180 ( .B1(n144), .B2(n146), .A(n104), .ZN(n105) );
  INV_X1 U181 ( .A(n105), .ZN(n107) );
  NOR2_X1 U182 ( .A1(n14), .A2(n147), .ZN(n106) );
  XOR2_X1 U183 ( .A(n107), .B(n106), .Z(n108) );
  XOR2_X1 U184 ( .A(n109), .B(n108), .Z(n110) );
  OR2_X1 U185 ( .A1(n111), .A2(n110), .ZN(n113) );
  NAND2_X1 U186 ( .A1(n111), .A2(n110), .ZN(n112) );
  NAND2_X1 U187 ( .A1(n113), .A2(n112), .ZN(n114) );
  MUX2_X1 U188 ( .A(n326), .B(n114), .S(n267), .Z(n352) );
  NAND2_X1 U189 ( .A1(n116), .A2(n115), .ZN(n117) );
  MUX2_X1 U190 ( .A(n327), .B(n117), .S(n267), .Z(n354) );
  NOR2_X1 U191 ( .A1(n119), .A2(n118), .ZN(n120) );
  MUX2_X1 U192 ( .A(n328), .B(n120), .S(n242), .Z(n356) );
  NAND2_X1 U193 ( .A1(n122), .A2(n121), .ZN(n123) );
  MUX2_X1 U194 ( .A(n330), .B(n123), .S(n267), .Z(n360) );
  FA_X1 U195 ( .A(n126), .B(n125), .CI(n124), .CO(n121), .S(n132) );
  FA_X1 U196 ( .A(n129), .B(n128), .CI(n127), .CO(n131), .S(n136) );
  NOR2_X1 U197 ( .A1(n132), .A2(n131), .ZN(n130) );
  MUX2_X1 U198 ( .A(n331), .B(n130), .S(n314), .Z(n362) );
  NAND2_X1 U199 ( .A1(n132), .A2(n131), .ZN(n134) );
  MUX2_X1 U200 ( .A(n332), .B(n134), .S(n242), .Z(n364) );
  NAND2_X1 U201 ( .A1(n136), .A2(n135), .ZN(n137) );
  MUX2_X1 U202 ( .A(n333), .B(n137), .S(n242), .Z(n366) );
  FA_X1 U203 ( .A(n140), .B(n139), .CI(n138), .CO(n169), .S(n173) );
  AOI21_X1 U204 ( .B1(n188), .B2(n10), .A(n141), .ZN(n142) );
  INV_X1 U205 ( .A(n142), .ZN(n222) );
  OAI22_X1 U206 ( .A1(n146), .A2(n145), .B1(n144), .B2(n143), .ZN(n221) );
  NOR2_X1 U207 ( .A1(n19), .A2(n147), .ZN(n220) );
  NOR2_X1 U208 ( .A1(n20), .A2(n147), .ZN(n211) );
  OAI22_X1 U209 ( .A1(n151), .A2(n150), .B1(n149), .B2(n148), .ZN(n203) );
  INV_X1 U210 ( .A(n203), .ZN(n155) );
  OAI22_X1 U211 ( .A1(n184), .A2(n153), .B1(n186), .B2(n152), .ZN(n202) );
  INV_X1 U212 ( .A(n202), .ZN(n154) );
  NAND2_X1 U213 ( .A1(n155), .A2(n154), .ZN(n210) );
  INV_X1 U214 ( .A(n210), .ZN(n156) );
  NAND2_X1 U215 ( .A1(n157), .A2(n156), .ZN(n158) );
  NAND2_X1 U216 ( .A1(n213), .A2(n158), .ZN(n160) );
  FA_X1 U217 ( .A(n163), .B(n6), .CI(n161), .CO(n139), .S(n199) );
  NOR2_X1 U218 ( .A1(n173), .A2(n172), .ZN(n168) );
  MUX2_X1 U219 ( .A(n334), .B(n168), .S(n242), .Z(n368) );
  NAND2_X1 U220 ( .A1(n170), .A2(n169), .ZN(n171) );
  MUX2_X1 U221 ( .A(n335), .B(n171), .S(n242), .Z(n370) );
  NAND2_X1 U222 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2_X1 U223 ( .A(n336), .B(n174), .S(n242), .Z(n372) );
  FA_X1 U224 ( .A(n177), .B(n176), .CI(n175), .CO(n135), .S(n196) );
  XNOR2_X1 U225 ( .A(n8), .B(\mult_x_1/n288 ), .ZN(n179) );
  OAI22_X1 U226 ( .A1(n184), .A2(n179), .B1(n186), .B2(n178), .ZN(n182) );
  XNOR2_X1 U227 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n185) );
  OAI22_X1 U228 ( .A1(n188), .A2(n185), .B1(n180), .B2(n10), .ZN(n181) );
  NOR2_X1 U229 ( .A1(n196), .A2(n195), .ZN(n260) );
  HA_X1 U230 ( .A(n182), .B(n181), .CO(n195), .S(n193) );
  OR2_X1 U231 ( .A1(\mult_x_1/n288 ), .A2(n23), .ZN(n183) );
  OAI22_X1 U232 ( .A1(n184), .A2(n23), .B1(n183), .B2(n186), .ZN(n192) );
  OR2_X1 U233 ( .A1(n193), .A2(n192), .ZN(n256) );
  XNOR2_X1 U234 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n187) );
  OAI22_X1 U235 ( .A1(n188), .A2(n187), .B1(n185), .B2(n10), .ZN(n191) );
  AND2_X1 U236 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n190) );
  NOR2_X1 U237 ( .A1(n191), .A2(n190), .ZN(n249) );
  OAI22_X1 U238 ( .A1(n188), .A2(\mult_x_1/n288 ), .B1(n187), .B2(n10), .ZN(
        n246) );
  OR2_X1 U239 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n189) );
  NAND2_X1 U240 ( .A1(n189), .A2(n188), .ZN(n245) );
  NAND2_X1 U241 ( .A1(n246), .A2(n245), .ZN(n252) );
  NAND2_X1 U242 ( .A1(n191), .A2(n190), .ZN(n250) );
  OAI21_X1 U243 ( .B1(n249), .B2(n252), .A(n250), .ZN(n257) );
  NAND2_X1 U244 ( .A1(n193), .A2(n192), .ZN(n255) );
  INV_X1 U245 ( .A(n255), .ZN(n194) );
  AOI21_X1 U246 ( .B1(n256), .B2(n257), .A(n194), .ZN(n263) );
  NAND2_X1 U247 ( .A1(n196), .A2(n195), .ZN(n261) );
  OAI21_X1 U248 ( .B1(n260), .B2(n263), .A(n261), .ZN(n197) );
  MUX2_X1 U249 ( .A(n337), .B(n197), .S(n242), .Z(n374) );
  FA_X1 U250 ( .A(n200), .B(n199), .CI(n198), .CO(n172), .S(n201) );
  MUX2_X1 U251 ( .A(n338), .B(n201), .S(n242), .Z(n376) );
  XNOR2_X1 U252 ( .A(n203), .B(n202), .ZN(n219) );
  FA_X1 U253 ( .A(n206), .B(n205), .CI(n204), .CO(n218), .S(n241) );
  FA_X1 U254 ( .A(n209), .B(n208), .CI(n207), .CO(n167), .S(n216) );
  XNOR2_X1 U255 ( .A(n211), .B(n210), .ZN(n212) );
  XNOR2_X1 U256 ( .A(n213), .B(n212), .ZN(n215) );
  MUX2_X1 U257 ( .A(n339), .B(n214), .S(n242), .Z(n378) );
  FA_X1 U258 ( .A(n24), .B(n216), .CI(n215), .CO(n214), .S(n217) );
  MUX2_X1 U259 ( .A(n340), .B(n217), .S(n242), .Z(n380) );
  FA_X1 U260 ( .A(n222), .B(n221), .CI(n220), .CO(n213), .S(n236) );
  MUX2_X1 U261 ( .A(n341), .B(n234), .S(n242), .Z(n382) );
  MUX2_X1 U262 ( .A(n342), .B(n238), .S(n242), .Z(n384) );
  FA_X1 U263 ( .A(n241), .B(n240), .CI(n239), .CO(n243), .S(n119) );
  MUX2_X1 U264 ( .A(n343), .B(n243), .S(n242), .Z(n386) );
  MUX2_X1 U265 ( .A(product[0]), .B(n508), .S(n267), .Z(n400) );
  MUX2_X1 U266 ( .A(n508), .B(n509), .S(n267), .Z(n402) );
  AND2_X1 U267 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n244) );
  MUX2_X1 U268 ( .A(n509), .B(n244), .S(n267), .Z(n404) );
  MUX2_X1 U269 ( .A(product[1]), .B(n511), .S(n267), .Z(n406) );
  MUX2_X1 U270 ( .A(n511), .B(n512), .S(n267), .Z(n408) );
  OR2_X1 U271 ( .A1(n246), .A2(n245), .ZN(n247) );
  AND2_X1 U272 ( .A1(n247), .A2(n252), .ZN(n248) );
  MUX2_X1 U273 ( .A(n512), .B(n248), .S(n267), .Z(n410) );
  MUX2_X1 U274 ( .A(product[2]), .B(n514), .S(n267), .Z(n412) );
  MUX2_X1 U275 ( .A(n514), .B(n515), .S(n267), .Z(n414) );
  INV_X1 U276 ( .A(n249), .ZN(n251) );
  NAND2_X1 U277 ( .A1(n251), .A2(n250), .ZN(n253) );
  XOR2_X1 U278 ( .A(n253), .B(n252), .Z(n254) );
  MUX2_X1 U279 ( .A(n515), .B(n254), .S(n267), .Z(n416) );
  MUX2_X1 U280 ( .A(product[3]), .B(n517), .S(n267), .Z(n418) );
  MUX2_X1 U281 ( .A(n517), .B(n518), .S(n267), .Z(n420) );
  NAND2_X1 U282 ( .A1(n256), .A2(n255), .ZN(n258) );
  XNOR2_X1 U283 ( .A(n258), .B(n257), .ZN(n259) );
  MUX2_X1 U284 ( .A(n518), .B(n259), .S(n267), .Z(n422) );
  MUX2_X1 U285 ( .A(product[4]), .B(n520), .S(n267), .Z(n424) );
  MUX2_X1 U286 ( .A(n520), .B(n521), .S(n267), .Z(n426) );
  INV_X1 U287 ( .A(n260), .ZN(n262) );
  NAND2_X1 U288 ( .A1(n262), .A2(n261), .ZN(n264) );
  XOR2_X1 U289 ( .A(n264), .B(n263), .Z(n265) );
  MUX2_X1 U290 ( .A(n521), .B(n265), .S(n267), .Z(n428) );
  MUX2_X1 U291 ( .A(product[5]), .B(n523), .S(n267), .Z(n430) );
  NAND2_X1 U292 ( .A1(n322), .A2(n333), .ZN(n266) );
  XNOR2_X1 U293 ( .A(n266), .B(n337), .ZN(n268) );
  MUX2_X1 U294 ( .A(n523), .B(n268), .S(n267), .Z(n432) );
  BUF_X4 U295 ( .A(en), .Z(n314) );
  MUX2_X1 U296 ( .A(product[6]), .B(n525), .S(n314), .Z(n434) );
  NAND2_X1 U297 ( .A1(n389), .A2(n332), .ZN(n269) );
  AOI21_X1 U298 ( .B1(n322), .B2(n337), .A(n393), .ZN(n271) );
  XOR2_X1 U299 ( .A(n269), .B(n271), .Z(n270) );
  MUX2_X1 U300 ( .A(n525), .B(n270), .S(n314), .Z(n436) );
  MUX2_X1 U301 ( .A(product[7]), .B(n527), .S(n314), .Z(n438) );
  OAI21_X1 U302 ( .B1(n331), .B2(n271), .A(n332), .ZN(n274) );
  NAND2_X1 U303 ( .A1(n325), .A2(n330), .ZN(n272) );
  XNOR2_X1 U304 ( .A(n274), .B(n272), .ZN(n273) );
  MUX2_X1 U305 ( .A(n527), .B(n273), .S(n314), .Z(n440) );
  MUX2_X1 U306 ( .A(product[8]), .B(n529), .S(n314), .Z(n442) );
  AOI21_X1 U307 ( .B1(n274), .B2(n325), .A(n392), .ZN(n277) );
  NAND2_X1 U308 ( .A1(n394), .A2(n329), .ZN(n275) );
  XOR2_X1 U309 ( .A(n277), .B(n275), .Z(n276) );
  MUX2_X1 U310 ( .A(n529), .B(n276), .S(n314), .Z(n444) );
  MUX2_X1 U311 ( .A(product[9]), .B(n531), .S(n314), .Z(n446) );
  OAI21_X1 U312 ( .B1(n277), .B2(n328), .A(n329), .ZN(n291) );
  INV_X1 U313 ( .A(n291), .ZN(n281) );
  NOR2_X1 U314 ( .A1(n342), .A2(n343), .ZN(n286) );
  INV_X1 U315 ( .A(n286), .ZN(n278) );
  NAND2_X1 U316 ( .A1(n342), .A2(n343), .ZN(n288) );
  NAND2_X1 U317 ( .A1(n278), .A2(n288), .ZN(n279) );
  XOR2_X1 U318 ( .A(n281), .B(n279), .Z(n280) );
  MUX2_X1 U319 ( .A(n531), .B(n280), .S(n314), .Z(n448) );
  MUX2_X1 U320 ( .A(product[10]), .B(n533), .S(n314), .Z(n450) );
  OAI21_X1 U321 ( .B1(n281), .B2(n286), .A(n288), .ZN(n284) );
  NOR2_X1 U322 ( .A1(n340), .A2(n341), .ZN(n289) );
  INV_X1 U323 ( .A(n289), .ZN(n282) );
  NAND2_X1 U324 ( .A1(n340), .A2(n341), .ZN(n287) );
  NAND2_X1 U325 ( .A1(n282), .A2(n287), .ZN(n283) );
  XNOR2_X1 U326 ( .A(n284), .B(n283), .ZN(n285) );
  MUX2_X1 U327 ( .A(n533), .B(n285), .S(n314), .Z(n452) );
  MUX2_X1 U328 ( .A(product[11]), .B(n535), .S(n314), .Z(n454) );
  NOR2_X1 U329 ( .A1(n289), .A2(n286), .ZN(n292) );
  OAI21_X1 U330 ( .B1(n289), .B2(n288), .A(n287), .ZN(n290) );
  AOI21_X1 U331 ( .B1(n292), .B2(n291), .A(n290), .ZN(n319) );
  NOR2_X1 U332 ( .A1(n338), .A2(n339), .ZN(n305) );
  INV_X1 U333 ( .A(n305), .ZN(n298) );
  NAND2_X1 U334 ( .A1(n338), .A2(n339), .ZN(n307) );
  NAND2_X1 U335 ( .A1(n298), .A2(n307), .ZN(n293) );
  XOR2_X1 U336 ( .A(n319), .B(n293), .Z(n294) );
  MUX2_X1 U337 ( .A(n535), .B(n294), .S(n314), .Z(n456) );
  MUX2_X1 U338 ( .A(product[12]), .B(n537), .S(n314), .Z(n458) );
  OAI21_X1 U339 ( .B1(n319), .B2(n305), .A(n307), .ZN(n296) );
  NAND2_X1 U340 ( .A1(n390), .A2(n336), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U342 ( .A(n537), .B(n297), .S(n314), .Z(n460) );
  MUX2_X1 U343 ( .A(product[13]), .B(n539), .S(n314), .Z(n462) );
  NAND2_X1 U344 ( .A1(n298), .A2(n390), .ZN(n301) );
  INV_X1 U345 ( .A(n307), .ZN(n299) );
  AOI21_X1 U346 ( .B1(n299), .B2(n390), .A(n395), .ZN(n300) );
  OAI21_X1 U347 ( .B1(n319), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U348 ( .A1(n324), .A2(n335), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U350 ( .A(n539), .B(n304), .S(n314), .Z(n464) );
  MUX2_X1 U351 ( .A(product[14]), .B(n541), .S(n314), .Z(n466) );
  NAND2_X1 U352 ( .A1(n390), .A2(n324), .ZN(n308) );
  NOR2_X1 U353 ( .A1(n305), .A2(n308), .ZN(n315) );
  INV_X1 U354 ( .A(n315), .ZN(n310) );
  AOI21_X1 U355 ( .B1(n395), .B2(n324), .A(n391), .ZN(n306) );
  OAI21_X1 U356 ( .B1(n308), .B2(n307), .A(n306), .ZN(n316) );
  INV_X1 U357 ( .A(n316), .ZN(n309) );
  OAI21_X1 U358 ( .B1(n319), .B2(n310), .A(n309), .ZN(n312) );
  NAND2_X1 U359 ( .A1(n323), .A2(n327), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U361 ( .A(n541), .B(n313), .S(n314), .Z(n468) );
  MUX2_X1 U362 ( .A(product[15]), .B(n543), .S(n314), .Z(n470) );
  NAND2_X1 U363 ( .A1(n315), .A2(n323), .ZN(n318) );
  AOI21_X1 U364 ( .B1(n316), .B2(n323), .A(n388), .ZN(n317) );
  OAI21_X1 U365 ( .B1(n319), .B2(n318), .A(n317), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n320), .B(n326), .ZN(n321) );
  MUX2_X1 U367 ( .A(n543), .B(n321), .S(n314), .Z(n472) );
  MUX2_X1 U368 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n314), .Z(n474) );
  MUX2_X1 U369 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n314), .Z(n476) );
  MUX2_X1 U370 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n314), .Z(n478) );
  MUX2_X1 U371 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n314), .Z(n480) );
  MUX2_X1 U372 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n314), .Z(n482) );
  MUX2_X1 U373 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n314), .Z(n484) );
  MUX2_X1 U374 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n314), .Z(n486) );
  MUX2_X1 U375 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n314), .Z(n488) );
  MUX2_X1 U376 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n314), .Z(n490) );
  MUX2_X1 U377 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n314), .Z(n492) );
  MUX2_X1 U378 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n314), .Z(n494) );
  MUX2_X1 U379 ( .A(n8), .B(A_extended[3]), .S(n314), .Z(n496) );
  MUX2_X1 U380 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n314), .Z(n498) );
  MUX2_X1 U381 ( .A(n9), .B(A_extended[5]), .S(n314), .Z(n500) );
  MUX2_X1 U382 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n314), .Z(n502) );
  MUX2_X1 U383 ( .A(n7), .B(A_extended[7]), .S(n314), .Z(n504) );
  OR2_X1 U384 ( .A1(n267), .A2(n545), .ZN(n506) );
endmodule


module conv_128_32_DW_mult_pipe_J1_2 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n355, n357, n359, n361, n363,
         n365, n367, n369, n371, n373, n375, n377, n379, n381, n383, n385,
         n387, n389, n391, n393, n395, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n408, n410, n412, n414, n416, n418, n420,
         n422, n424, n426, n428, n430, n432, n434, n436, n438, n440, n442,
         n444, n446, n448, n450, n452, n454, n456, n458, n460, n462, n464,
         n466, n468, n470, n472, n474, n476, n478, n480, n482, n484, n486,
         n488, n490, n492, n494, n496, n498, n500, n502, n504, n506, n508,
         n510, n512, n514, n516, n517, n519, n520, n522, n523, n525, n526,
         n528, n529, n531, n533, n535, n537, n539, n541, n543, n545, n547,
         n549, n551, n552, n553, n554;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n404), .SE(n514), .CK(clk), .Q(n553), 
        .QN(n5) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n404), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n28) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n404), .SE(n506), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n10) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n404), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n11) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n404), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n15) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n404), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n21) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n404), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n27) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n405), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n406), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n22) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n404), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n23) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n404), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n25) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n404), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n24) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n404), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n13) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n404), .SE(n480), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n404), .SE(n478), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n404), .SE(n476), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n404), .SE(n474), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n404), .SE(n472), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n406), .SE(n470), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n404), .SE(n468), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n405), .SE(n466), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n404), .SE(n464), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n404), .SE(n462), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n404), .SE(n460), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n404), .SE(n458), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n404), .SE(n456), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n404), .SE(n454), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n404), .SE(n452), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n406), .SE(n450), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n406), .SE(n448), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n406), .SE(n446), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n406), .SE(n444), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n406), .SE(n442), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n406), .SE(n440), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n406), .SE(n438), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n406), .SE(n436), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n406), .SE(n434), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n406), .SE(n432), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n406), .SE(n430), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n405), .SE(n428), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n405), .SE(n426), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n405), .SE(n424), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n405), .SE(n422), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n405), .SE(n420), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n405), .SE(n418), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n405), .SE(n416), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n405), .SE(n414), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n405), .SE(n412), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n405), .SE(n410), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n405), .SE(n408), .CK(clk), .Q(
        product[0]) );
  SDFF_X2 clk_r_REG41_S1 ( .D(1'b0), .SI(n404), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n16) );
  SDFF_X2 clk_r_REG51_S1 ( .D(1'b0), .SI(n404), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n17) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n554), .SE(n395), .CK(
        clk), .QN(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2_IP  ( .D(1'b1), .SI(n554), .SE(n393), .CK(
        clk), .QN(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n554), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n554), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n554), .SE(n387), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n554), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n554), .SE(n383), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n554), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n554), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n344), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n554), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n343), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n554), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n342), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n554), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n554), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n340), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n554), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n339), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n554), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n554), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n337), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n554), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n336), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n554), .SE(n361), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n554), .SE(n359), .CK(
        clk), .QN(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n554), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n554), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n554), .SE(n353), .CK(
        clk), .QN(n331) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n404), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n18) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n404), .SE(n512), .CK(clk), .Q(n552), 
        .QN(n19) );
  BUF_X4 U2 ( .A(en), .Z(n276) );
  BUF_X1 U3 ( .A(n404), .Z(n406) );
  INV_X2 U4 ( .A(n554), .ZN(n404) );
  BUF_X1 U5 ( .A(n404), .Z(n405) );
  OAI22_X1 U6 ( .A1(n144), .A2(n91), .B1(n37), .B2(n143), .ZN(n87) );
  INV_X1 U7 ( .A(rst_n), .ZN(n554) );
  INV_X1 U8 ( .A(n31), .ZN(n144) );
  NAND2_X1 U9 ( .A1(n7), .A2(n6), .ZN(n143) );
  AND2_X1 U10 ( .A1(n9), .A2(n8), .ZN(n31) );
  NAND2_X1 U11 ( .A1(n8), .A2(n552), .ZN(n6) );
  NAND2_X1 U12 ( .A1(n19), .A2(n9), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n16), .A2(n28), .ZN(n8) );
  OR2_X1 U14 ( .A1(n16), .A2(n28), .ZN(n9) );
  XNOR2_X1 U15 ( .A(n87), .B(n86), .ZN(n41) );
  NOR2_X1 U16 ( .A1(n209), .A2(n22), .ZN(n86) );
  NAND2_X1 U17 ( .A1(n552), .A2(n5), .ZN(n209) );
  OR2_X1 U18 ( .A1(n246), .A2(n245), .ZN(n241) );
  NAND2_X1 U19 ( .A1(n240), .A2(n239), .ZN(n245) );
  NAND2_X1 U20 ( .A1(n236), .A2(n235), .ZN(n240) );
  NAND2_X1 U21 ( .A1(n234), .A2(n233), .ZN(n235) );
  INV_X1 U22 ( .A(n238), .ZN(n234) );
  NAND2_X1 U23 ( .A1(n99), .A2(n98), .ZN(n177) );
  NAND2_X1 U24 ( .A1(n95), .A2(n94), .ZN(n99) );
  NAND2_X1 U25 ( .A1(n90), .A2(n89), .ZN(n124) );
  NAND2_X1 U26 ( .A1(n116), .A2(n345), .ZN(n62) );
  NAND2_X1 U27 ( .A1(n243), .A2(n242), .ZN(n244) );
  NAND2_X1 U28 ( .A1(n246), .A2(n245), .ZN(n242) );
  NAND2_X1 U29 ( .A1(n20), .A2(n241), .ZN(n243) );
  XNOR2_X1 U30 ( .A(n20), .B(n247), .ZN(n248) );
  XNOR2_X1 U31 ( .A(n246), .B(n245), .ZN(n247) );
  XNOR2_X1 U32 ( .A(n17), .B(n10), .ZN(n39) );
  XNOR2_X1 U33 ( .A(n11), .B(n18), .ZN(n33) );
  XNOR2_X1 U34 ( .A(n223), .B(n222), .ZN(n225) );
  XNOR2_X1 U35 ( .A(n221), .B(n220), .ZN(n222) );
  XNOR2_X1 U36 ( .A(n61), .B(n12), .ZN(n203) );
  XNOR2_X1 U37 ( .A(n60), .B(n59), .ZN(n12) );
  NOR2_X1 U38 ( .A1(n60), .A2(n59), .ZN(n14) );
  XOR2_X1 U39 ( .A(n229), .B(n228), .Z(n20) );
  AND2_X1 U40 ( .A1(n229), .A2(n228), .ZN(n29) );
  INV_X1 U41 ( .A(n323), .ZN(n116) );
  NAND2_X1 U42 ( .A1(n60), .A2(n59), .ZN(n30) );
  XNOR2_X1 U43 ( .A(n552), .B(\mult_x_1/n284 ), .ZN(n42) );
  XNOR2_X1 U44 ( .A(n552), .B(\mult_x_1/n283 ), .ZN(n37) );
  OAI22_X1 U45 ( .A1(n143), .A2(n42), .B1(n144), .B2(n37), .ZN(n58) );
  XOR2_X1 U46 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n32) );
  NAND2_X2 U47 ( .A1(n32), .A2(n33), .ZN(n189) );
  XNOR2_X1 U48 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n50) );
  AND2_X1 U49 ( .A1(n553), .A2(\mult_x_1/n281 ), .ZN(n117) );
  XNOR2_X1 U50 ( .A(n117), .B(\mult_x_1/n312 ), .ZN(n35) );
  INV_X1 U51 ( .A(n33), .ZN(n34) );
  INV_X1 U52 ( .A(n34), .ZN(n191) );
  OAI22_X1 U53 ( .A1(n189), .A2(n50), .B1(n35), .B2(n191), .ZN(n57) );
  AOI21_X1 U54 ( .B1(n191), .B2(n189), .A(n35), .ZN(n36) );
  INV_X1 U55 ( .A(n36), .ZN(n56) );
  XNOR2_X1 U56 ( .A(n552), .B(\mult_x_1/n282 ), .ZN(n91) );
  INV_X1 U57 ( .A(n39), .ZN(n38) );
  INV_X2 U58 ( .A(n38), .ZN(n132) );
  XNOR2_X1 U59 ( .A(n117), .B(\mult_x_1/n311 ), .ZN(n92) );
  XOR2_X1 U60 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n40) );
  NAND2_X2 U61 ( .A1(n40), .A2(n39), .ZN(n134) );
  XNOR2_X1 U62 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n43) );
  OAI22_X1 U63 ( .A1(n132), .A2(n92), .B1(n134), .B2(n43), .ZN(n119) );
  INV_X1 U64 ( .A(n119), .ZN(n88) );
  XNOR2_X1 U65 ( .A(n41), .B(n88), .ZN(n97) );
  XNOR2_X1 U66 ( .A(n96), .B(n97), .ZN(n46) );
  XNOR2_X1 U67 ( .A(n552), .B(\mult_x_1/n285 ), .ZN(n48) );
  OAI22_X1 U68 ( .A1(n143), .A2(n48), .B1(n144), .B2(n42), .ZN(n219) );
  XNOR2_X1 U69 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n49) );
  XNOR2_X1 U70 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n44) );
  OAI22_X1 U71 ( .A1(n134), .A2(n49), .B1(n132), .B2(n44), .ZN(n218) );
  INV_X1 U72 ( .A(n57), .ZN(n217) );
  INV_X1 U73 ( .A(n61), .ZN(n45) );
  NOR2_X1 U74 ( .A1(n23), .A2(n209), .ZN(n60) );
  OAI22_X1 U75 ( .A1(n134), .A2(n44), .B1(n132), .B2(n43), .ZN(n59) );
  OAI21_X1 U76 ( .B1(n45), .B2(n14), .A(n30), .ZN(n95) );
  XNOR2_X1 U77 ( .A(n46), .B(n95), .ZN(n103) );
  NAND2_X1 U78 ( .A1(\mult_x_1/n313 ), .A2(n15), .ZN(n193) );
  XNOR2_X1 U79 ( .A(n117), .B(\mult_x_1/n313 ), .ZN(n65) );
  AOI21_X1 U80 ( .B1(n193), .B2(n15), .A(n65), .ZN(n47) );
  INV_X1 U81 ( .A(n47), .ZN(n232) );
  XNOR2_X1 U82 ( .A(n552), .B(\mult_x_1/n286 ), .ZN(n64) );
  OAI22_X1 U83 ( .A1(n143), .A2(n64), .B1(n144), .B2(n48), .ZN(n231) );
  NOR2_X1 U84 ( .A1(n24), .A2(n209), .ZN(n230) );
  INV_X1 U85 ( .A(n223), .ZN(n55) );
  NOR2_X1 U86 ( .A1(n25), .A2(n209), .ZN(n220) );
  INV_X1 U87 ( .A(n220), .ZN(n52) );
  XNOR2_X1 U88 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n73) );
  OAI22_X1 U89 ( .A1(n134), .A2(n73), .B1(n132), .B2(n49), .ZN(n208) );
  XNOR2_X1 U90 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n71) );
  OAI22_X1 U91 ( .A1(n189), .A2(n71), .B1(n191), .B2(n50), .ZN(n207) );
  OR2_X1 U92 ( .A1(n208), .A2(n207), .ZN(n221) );
  INV_X1 U93 ( .A(n221), .ZN(n51) );
  AND2_X1 U94 ( .A1(n52), .A2(n51), .ZN(n54) );
  NAND2_X1 U95 ( .A1(n221), .A2(n220), .ZN(n53) );
  OAI21_X1 U96 ( .B1(n55), .B2(n54), .A(n53), .ZN(n205) );
  FA_X1 U97 ( .A(n58), .B(n57), .CI(n56), .CO(n96), .S(n204) );
  OAI21_X1 U98 ( .B1(n103), .B2(n102), .A(n276), .ZN(n63) );
  NAND2_X1 U99 ( .A1(n63), .A2(n62), .ZN(n381) );
  XNOR2_X1 U100 ( .A(n552), .B(\mult_x_1/n287 ), .ZN(n69) );
  OAI22_X1 U101 ( .A1(n143), .A2(n69), .B1(n144), .B2(n64), .ZN(n212) );
  NOR2_X1 U102 ( .A1(n209), .A2(n13), .ZN(n214) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n67) );
  OAI22_X1 U104 ( .A1(n193), .A2(n67), .B1(n65), .B2(n15), .ZN(n213) );
  XNOR2_X1 U105 ( .A(n214), .B(n213), .ZN(n66) );
  XNOR2_X1 U106 ( .A(n212), .B(n66), .ZN(n251) );
  XNOR2_X1 U107 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n286 ), .ZN(n131) );
  XNOR2_X1 U108 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n285 ), .ZN(n74) );
  OAI22_X1 U109 ( .A1(n134), .A2(n131), .B1(n132), .B2(n74), .ZN(n82) );
  XNOR2_X1 U110 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n76) );
  OAI22_X1 U111 ( .A1(n193), .A2(n76), .B1(n67), .B2(n15), .ZN(n81) );
  XNOR2_X1 U112 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n77) );
  XNOR2_X1 U113 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n72) );
  OAI22_X1 U114 ( .A1(n189), .A2(n77), .B1(n191), .B2(n72), .ZN(n80) );
  OR2_X1 U115 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n68) );
  OAI22_X1 U116 ( .A1(n143), .A2(n19), .B1(n68), .B2(n144), .ZN(n79) );
  XNOR2_X1 U117 ( .A(n552), .B(\mult_x_1/n288 ), .ZN(n70) );
  OAI22_X1 U118 ( .A1(n143), .A2(n70), .B1(n144), .B2(n69), .ZN(n78) );
  OAI22_X1 U119 ( .A1(n189), .A2(n72), .B1(n191), .B2(n71), .ZN(n238) );
  OAI22_X1 U120 ( .A1(n134), .A2(n74), .B1(n132), .B2(n73), .ZN(n237) );
  XNOR2_X1 U121 ( .A(n238), .B(n237), .ZN(n75) );
  XNOR2_X1 U122 ( .A(n236), .B(n75), .ZN(n249) );
  XNOR2_X1 U123 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n108) );
  OAI22_X1 U124 ( .A1(n193), .A2(n108), .B1(n76), .B2(n15), .ZN(n137) );
  AND2_X1 U125 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n136) );
  XNOR2_X1 U126 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n107) );
  OAI22_X1 U127 ( .A1(n189), .A2(n107), .B1(n191), .B2(n77), .ZN(n135) );
  HA_X1 U128 ( .A(n79), .B(n78), .CO(n236), .S(n127) );
  FA_X1 U129 ( .A(n82), .B(n81), .CI(n80), .CO(n250), .S(n126) );
  NAND2_X1 U130 ( .A1(n159), .A2(n158), .ZN(n83) );
  NAND2_X1 U131 ( .A1(n83), .A2(n276), .ZN(n85) );
  NAND2_X1 U132 ( .A1(n116), .A2(n338), .ZN(n84) );
  NAND2_X1 U133 ( .A1(n85), .A2(n84), .ZN(n367) );
  OAI21_X1 U134 ( .B1(n88), .B2(n87), .A(n86), .ZN(n90) );
  NAND2_X1 U135 ( .A1(n88), .A2(n87), .ZN(n89) );
  NOR2_X1 U136 ( .A1(n26), .A2(n209), .ZN(n123) );
  XNOR2_X1 U137 ( .A(n552), .B(\mult_x_1/n281 ), .ZN(n118) );
  OAI22_X1 U138 ( .A1(n143), .A2(n91), .B1(n144), .B2(n118), .ZN(n121) );
  AOI21_X1 U139 ( .B1(n132), .B2(n134), .A(n92), .ZN(n93) );
  INV_X1 U140 ( .A(n93), .ZN(n120) );
  OR2_X1 U141 ( .A1(n97), .A2(n96), .ZN(n94) );
  NAND2_X1 U142 ( .A1(n97), .A2(n96), .ZN(n98) );
  OAI21_X1 U143 ( .B1(n178), .B2(n177), .A(n276), .ZN(n101) );
  NAND2_X1 U144 ( .A1(n116), .A2(n333), .ZN(n100) );
  NAND2_X1 U145 ( .A1(n101), .A2(n100), .ZN(n357) );
  NAND2_X1 U146 ( .A1(n103), .A2(n102), .ZN(n104) );
  NAND2_X1 U147 ( .A1(n104), .A2(n276), .ZN(n106) );
  NAND2_X1 U148 ( .A1(n116), .A2(n344), .ZN(n105) );
  NAND2_X1 U149 ( .A1(n106), .A2(n105), .ZN(n379) );
  XNOR2_X1 U172 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n113) );
  OAI22_X1 U173 ( .A1(n189), .A2(n113), .B1(n191), .B2(n107), .ZN(n169) );
  XNOR2_X1 U174 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n111) );
  OAI22_X1 U175 ( .A1(n193), .A2(n111), .B1(n108), .B2(n15), .ZN(n168) );
  OR2_X1 U176 ( .A1(\mult_x_1/n288 ), .A2(n16), .ZN(n109) );
  OAI22_X1 U177 ( .A1(n134), .A2(n16), .B1(n109), .B2(n132), .ZN(n130) );
  XNOR2_X1 U178 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n288 ), .ZN(n110) );
  XNOR2_X1 U179 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n133) );
  OAI22_X1 U180 ( .A1(n134), .A2(n110), .B1(n132), .B2(n133), .ZN(n129) );
  XNOR2_X1 U181 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n185) );
  OAI22_X1 U182 ( .A1(n193), .A2(n185), .B1(n111), .B2(n15), .ZN(n182) );
  INV_X1 U183 ( .A(n132), .ZN(n112) );
  AND2_X1 U184 ( .A1(\mult_x_1/n288 ), .A2(n112), .ZN(n181) );
  XNOR2_X1 U185 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n183) );
  OAI22_X1 U186 ( .A1(n189), .A2(n183), .B1(n191), .B2(n113), .ZN(n180) );
  NOR2_X1 U187 ( .A1(n175), .A2(n174), .ZN(n115) );
  NAND2_X1 U188 ( .A1(n116), .A2(n331), .ZN(n114) );
  OAI21_X1 U189 ( .B1(n116), .B2(n115), .A(n114), .ZN(n353) );
  NOR2_X1 U190 ( .A1(n27), .A2(n209), .ZN(n141) );
  XNOR2_X1 U191 ( .A(n117), .B(n552), .ZN(n142) );
  OAI22_X1 U192 ( .A1(n143), .A2(n118), .B1(n142), .B2(n144), .ZN(n149) );
  INV_X1 U193 ( .A(n149), .ZN(n140) );
  FA_X1 U194 ( .A(n121), .B(n120), .CI(n119), .CO(n139), .S(n122) );
  FA_X1 U195 ( .A(n124), .B(n123), .CI(n122), .CO(n155), .S(n178) );
  OR2_X1 U196 ( .A1(n156), .A2(n155), .ZN(n125) );
  MUX2_X1 U197 ( .A(n332), .B(n125), .S(n276), .Z(n355) );
  FA_X1 U198 ( .A(n128), .B(n127), .CI(n126), .CO(n158), .S(n162) );
  HA_X1 U199 ( .A(n130), .B(n129), .CO(n166), .S(n167) );
  OAI22_X1 U200 ( .A1(n134), .A2(n133), .B1(n132), .B2(n131), .ZN(n165) );
  FA_X1 U201 ( .A(n137), .B(n136), .CI(n135), .CO(n128), .S(n164) );
  OR2_X1 U202 ( .A1(n162), .A2(n161), .ZN(n138) );
  MUX2_X1 U203 ( .A(n334), .B(n138), .S(n276), .Z(n359) );
  FA_X1 U204 ( .A(n141), .B(n140), .CI(n139), .CO(n151), .S(n156) );
  AOI21_X1 U205 ( .B1(n144), .B2(n143), .A(n142), .ZN(n145) );
  INV_X1 U206 ( .A(n145), .ZN(n147) );
  NOR2_X1 U207 ( .A1(n21), .A2(n209), .ZN(n146) );
  XOR2_X1 U208 ( .A(n147), .B(n146), .Z(n148) );
  XOR2_X1 U209 ( .A(n149), .B(n148), .Z(n150) );
  OR2_X1 U210 ( .A1(n151), .A2(n150), .ZN(n153) );
  NAND2_X1 U211 ( .A1(n151), .A2(n150), .ZN(n152) );
  NAND2_X1 U212 ( .A1(n153), .A2(n152), .ZN(n154) );
  MUX2_X1 U213 ( .A(n335), .B(n154), .S(n276), .Z(n361) );
  NAND2_X1 U214 ( .A1(n156), .A2(n155), .ZN(n157) );
  MUX2_X1 U215 ( .A(n336), .B(n157), .S(n276), .Z(n363) );
  NOR2_X1 U216 ( .A1(n159), .A2(n158), .ZN(n160) );
  MUX2_X1 U217 ( .A(n337), .B(n160), .S(n276), .Z(n365) );
  NAND2_X1 U218 ( .A1(n162), .A2(n161), .ZN(n163) );
  MUX2_X1 U219 ( .A(n339), .B(n163), .S(n276), .Z(n369) );
  FA_X1 U220 ( .A(n166), .B(n165), .CI(n164), .CO(n161), .S(n172) );
  FA_X1 U221 ( .A(n169), .B(n168), .CI(n167), .CO(n171), .S(n175) );
  NOR2_X1 U222 ( .A1(n172), .A2(n171), .ZN(n170) );
  MUX2_X1 U223 ( .A(n340), .B(n170), .S(n276), .Z(n371) );
  NAND2_X1 U224 ( .A1(n172), .A2(n171), .ZN(n173) );
  MUX2_X1 U225 ( .A(n341), .B(n173), .S(n276), .Z(n373) );
  NAND2_X1 U226 ( .A1(n175), .A2(n174), .ZN(n176) );
  MUX2_X1 U227 ( .A(n342), .B(n176), .S(n276), .Z(n375) );
  NAND2_X1 U228 ( .A1(n178), .A2(n177), .ZN(n179) );
  MUX2_X1 U229 ( .A(n343), .B(n179), .S(n276), .Z(n377) );
  FA_X1 U230 ( .A(n182), .B(n181), .CI(n180), .CO(n174), .S(n201) );
  XNOR2_X1 U231 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n184) );
  OAI22_X1 U232 ( .A1(n189), .A2(n184), .B1(n191), .B2(n183), .ZN(n187) );
  XNOR2_X1 U233 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n190) );
  OAI22_X1 U234 ( .A1(n193), .A2(n190), .B1(n185), .B2(n15), .ZN(n186) );
  NOR2_X1 U235 ( .A1(n201), .A2(n200), .ZN(n269) );
  HA_X1 U236 ( .A(n187), .B(n186), .CO(n200), .S(n198) );
  OR2_X1 U237 ( .A1(\mult_x_1/n288 ), .A2(n17), .ZN(n188) );
  OAI22_X1 U238 ( .A1(n189), .A2(n17), .B1(n188), .B2(n191), .ZN(n197) );
  OR2_X1 U239 ( .A1(n198), .A2(n197), .ZN(n265) );
  XNOR2_X1 U240 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n192) );
  OAI22_X1 U241 ( .A1(n193), .A2(n192), .B1(n190), .B2(n15), .ZN(n196) );
  AND2_X1 U242 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n195) );
  NOR2_X1 U243 ( .A1(n196), .A2(n195), .ZN(n258) );
  OAI22_X1 U244 ( .A1(n193), .A2(\mult_x_1/n288 ), .B1(n192), .B2(n15), .ZN(
        n255) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n18), .ZN(n194) );
  NAND2_X1 U246 ( .A1(n194), .A2(n193), .ZN(n254) );
  NAND2_X1 U247 ( .A1(n255), .A2(n254), .ZN(n261) );
  NAND2_X1 U248 ( .A1(n196), .A2(n195), .ZN(n259) );
  OAI21_X1 U249 ( .B1(n258), .B2(n261), .A(n259), .ZN(n266) );
  NAND2_X1 U250 ( .A1(n198), .A2(n197), .ZN(n264) );
  INV_X1 U251 ( .A(n264), .ZN(n199) );
  AOI21_X1 U252 ( .B1(n265), .B2(n266), .A(n199), .ZN(n272) );
  NAND2_X1 U253 ( .A1(n201), .A2(n200), .ZN(n270) );
  OAI21_X1 U254 ( .B1(n269), .B2(n272), .A(n270), .ZN(n202) );
  MUX2_X1 U255 ( .A(n346), .B(n202), .S(n276), .Z(n383) );
  FA_X1 U256 ( .A(n205), .B(n204), .CI(n203), .CO(n102), .S(n206) );
  MUX2_X1 U257 ( .A(n347), .B(n206), .S(n276), .Z(n385) );
  XNOR2_X1 U258 ( .A(n208), .B(n207), .ZN(n229) );
  INV_X1 U259 ( .A(n209), .ZN(n211) );
  AND2_X1 U260 ( .A1(n213), .A2(\mult_x_1/n288 ), .ZN(n210) );
  NAND2_X1 U261 ( .A1(n211), .A2(n210), .ZN(n216) );
  OAI21_X1 U262 ( .B1(n214), .B2(n213), .A(n212), .ZN(n215) );
  NAND2_X1 U263 ( .A1(n216), .A2(n215), .ZN(n228) );
  FA_X1 U264 ( .A(n219), .B(n218), .CI(n217), .CO(n61), .S(n226) );
  MUX2_X1 U265 ( .A(n348), .B(n224), .S(n276), .Z(n387) );
  FA_X1 U266 ( .A(n29), .B(n226), .CI(n225), .CO(n224), .S(n227) );
  MUX2_X1 U267 ( .A(n349), .B(n227), .S(n276), .Z(n389) );
  FA_X1 U268 ( .A(n232), .B(n231), .CI(n230), .CO(n223), .S(n246) );
  INV_X1 U269 ( .A(n237), .ZN(n233) );
  NAND2_X1 U270 ( .A1(n238), .A2(n237), .ZN(n239) );
  MUX2_X1 U271 ( .A(n350), .B(n244), .S(n276), .Z(n391) );
  MUX2_X1 U272 ( .A(n351), .B(n248), .S(n276), .Z(n393) );
  FA_X1 U273 ( .A(n251), .B(n250), .CI(n249), .CO(n252), .S(n159) );
  MUX2_X1 U274 ( .A(n352), .B(n252), .S(n276), .Z(n395) );
  MUX2_X1 U275 ( .A(product[0]), .B(n516), .S(n276), .Z(n408) );
  MUX2_X1 U276 ( .A(n516), .B(n517), .S(n276), .Z(n410) );
  AND2_X1 U277 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n253) );
  MUX2_X1 U278 ( .A(n517), .B(n253), .S(n276), .Z(n412) );
  MUX2_X1 U279 ( .A(product[1]), .B(n519), .S(n276), .Z(n414) );
  MUX2_X1 U280 ( .A(n519), .B(n520), .S(n276), .Z(n416) );
  OR2_X1 U281 ( .A1(n255), .A2(n254), .ZN(n256) );
  AND2_X1 U282 ( .A1(n256), .A2(n261), .ZN(n257) );
  MUX2_X1 U283 ( .A(n520), .B(n257), .S(n276), .Z(n418) );
  MUX2_X1 U284 ( .A(product[2]), .B(n522), .S(n276), .Z(n420) );
  MUX2_X1 U285 ( .A(n522), .B(n523), .S(n276), .Z(n422) );
  INV_X1 U286 ( .A(n258), .ZN(n260) );
  NAND2_X1 U287 ( .A1(n260), .A2(n259), .ZN(n262) );
  XOR2_X1 U288 ( .A(n262), .B(n261), .Z(n263) );
  MUX2_X1 U289 ( .A(n523), .B(n263), .S(n276), .Z(n424) );
  MUX2_X1 U290 ( .A(product[3]), .B(n525), .S(n276), .Z(n426) );
  MUX2_X1 U291 ( .A(n525), .B(n526), .S(n276), .Z(n428) );
  NAND2_X1 U292 ( .A1(n265), .A2(n264), .ZN(n267) );
  XNOR2_X1 U293 ( .A(n267), .B(n266), .ZN(n268) );
  MUX2_X1 U294 ( .A(n526), .B(n268), .S(n276), .Z(n430) );
  MUX2_X1 U295 ( .A(product[4]), .B(n528), .S(n276), .Z(n432) );
  MUX2_X1 U296 ( .A(n528), .B(n529), .S(n276), .Z(n434) );
  INV_X1 U297 ( .A(n269), .ZN(n271) );
  NAND2_X1 U298 ( .A1(n271), .A2(n270), .ZN(n273) );
  XOR2_X1 U299 ( .A(n273), .B(n272), .Z(n274) );
  MUX2_X1 U300 ( .A(n529), .B(n274), .S(n276), .Z(n436) );
  MUX2_X1 U301 ( .A(product[5]), .B(n531), .S(n276), .Z(n438) );
  NAND2_X1 U302 ( .A1(n331), .A2(n342), .ZN(n275) );
  XNOR2_X1 U303 ( .A(n275), .B(n346), .ZN(n277) );
  MUX2_X1 U304 ( .A(n531), .B(n277), .S(n276), .Z(n440) );
  BUF_X4 U305 ( .A(en), .Z(n323) );
  MUX2_X1 U306 ( .A(product[6]), .B(n533), .S(n323), .Z(n442) );
  NAND2_X1 U307 ( .A1(n399), .A2(n341), .ZN(n278) );
  AOI21_X1 U308 ( .B1(n331), .B2(n346), .A(n401), .ZN(n280) );
  XOR2_X1 U309 ( .A(n278), .B(n280), .Z(n279) );
  MUX2_X1 U310 ( .A(n533), .B(n279), .S(n323), .Z(n444) );
  MUX2_X1 U311 ( .A(product[7]), .B(n535), .S(n323), .Z(n446) );
  OAI21_X1 U312 ( .B1(n340), .B2(n280), .A(n341), .ZN(n283) );
  NAND2_X1 U313 ( .A1(n334), .A2(n339), .ZN(n281) );
  XNOR2_X1 U314 ( .A(n283), .B(n281), .ZN(n282) );
  MUX2_X1 U315 ( .A(n535), .B(n282), .S(n323), .Z(n448) );
  MUX2_X1 U316 ( .A(product[8]), .B(n537), .S(n323), .Z(n450) );
  AOI21_X1 U317 ( .B1(n283), .B2(n334), .A(n400), .ZN(n286) );
  NAND2_X1 U318 ( .A1(n402), .A2(n338), .ZN(n284) );
  XOR2_X1 U319 ( .A(n286), .B(n284), .Z(n285) );
  MUX2_X1 U320 ( .A(n537), .B(n285), .S(n323), .Z(n452) );
  MUX2_X1 U321 ( .A(product[9]), .B(n539), .S(n323), .Z(n454) );
  OAI21_X1 U322 ( .B1(n286), .B2(n337), .A(n338), .ZN(n300) );
  INV_X1 U323 ( .A(n300), .ZN(n290) );
  NOR2_X1 U324 ( .A1(n351), .A2(n352), .ZN(n295) );
  INV_X1 U325 ( .A(n295), .ZN(n287) );
  NAND2_X1 U326 ( .A1(n351), .A2(n352), .ZN(n297) );
  NAND2_X1 U327 ( .A1(n287), .A2(n297), .ZN(n288) );
  XOR2_X1 U328 ( .A(n290), .B(n288), .Z(n289) );
  MUX2_X1 U329 ( .A(n539), .B(n289), .S(n323), .Z(n456) );
  MUX2_X1 U330 ( .A(product[10]), .B(n541), .S(n323), .Z(n458) );
  OAI21_X1 U331 ( .B1(n290), .B2(n295), .A(n297), .ZN(n293) );
  NOR2_X1 U332 ( .A1(n349), .A2(n350), .ZN(n298) );
  INV_X1 U333 ( .A(n298), .ZN(n291) );
  NAND2_X1 U334 ( .A1(n349), .A2(n350), .ZN(n296) );
  NAND2_X1 U335 ( .A1(n291), .A2(n296), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  MUX2_X1 U337 ( .A(n541), .B(n294), .S(n323), .Z(n460) );
  MUX2_X1 U338 ( .A(product[11]), .B(n543), .S(n323), .Z(n462) );
  NOR2_X1 U339 ( .A1(n298), .A2(n295), .ZN(n301) );
  OAI21_X1 U340 ( .B1(n298), .B2(n297), .A(n296), .ZN(n299) );
  AOI21_X1 U341 ( .B1(n301), .B2(n300), .A(n299), .ZN(n328) );
  NOR2_X1 U342 ( .A1(n347), .A2(n348), .ZN(n314) );
  INV_X1 U343 ( .A(n314), .ZN(n307) );
  NAND2_X1 U344 ( .A1(n347), .A2(n348), .ZN(n316) );
  NAND2_X1 U345 ( .A1(n307), .A2(n316), .ZN(n302) );
  XOR2_X1 U346 ( .A(n328), .B(n302), .Z(n303) );
  MUX2_X1 U347 ( .A(n543), .B(n303), .S(n323), .Z(n464) );
  MUX2_X1 U348 ( .A(product[12]), .B(n545), .S(n323), .Z(n466) );
  OAI21_X1 U349 ( .B1(n328), .B2(n314), .A(n316), .ZN(n305) );
  NAND2_X1 U350 ( .A1(n345), .A2(n344), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  MUX2_X1 U352 ( .A(n545), .B(n306), .S(n323), .Z(n468) );
  MUX2_X1 U353 ( .A(product[13]), .B(n547), .S(n323), .Z(n470) );
  NAND2_X1 U354 ( .A1(n307), .A2(n345), .ZN(n310) );
  INV_X1 U355 ( .A(n316), .ZN(n308) );
  AOI21_X1 U356 ( .B1(n308), .B2(n345), .A(n403), .ZN(n309) );
  OAI21_X1 U357 ( .B1(n328), .B2(n310), .A(n309), .ZN(n312) );
  NAND2_X1 U358 ( .A1(n333), .A2(n343), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U360 ( .A(n547), .B(n313), .S(n323), .Z(n472) );
  MUX2_X1 U361 ( .A(product[14]), .B(n549), .S(n323), .Z(n474) );
  NAND2_X1 U362 ( .A1(n345), .A2(n333), .ZN(n317) );
  NOR2_X1 U363 ( .A1(n314), .A2(n317), .ZN(n324) );
  INV_X1 U364 ( .A(n324), .ZN(n319) );
  AOI21_X1 U365 ( .B1(n403), .B2(n333), .A(n397), .ZN(n315) );
  OAI21_X1 U366 ( .B1(n317), .B2(n316), .A(n315), .ZN(n325) );
  INV_X1 U367 ( .A(n325), .ZN(n318) );
  OAI21_X1 U368 ( .B1(n328), .B2(n319), .A(n318), .ZN(n321) );
  NAND2_X1 U369 ( .A1(n332), .A2(n336), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U371 ( .A(n549), .B(n322), .S(n323), .Z(n476) );
  MUX2_X1 U372 ( .A(product[15]), .B(n551), .S(n323), .Z(n478) );
  NAND2_X1 U373 ( .A1(n324), .A2(n332), .ZN(n327) );
  AOI21_X1 U374 ( .B1(n325), .B2(n332), .A(n398), .ZN(n326) );
  OAI21_X1 U375 ( .B1(n328), .B2(n327), .A(n326), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n329), .B(n335), .ZN(n330) );
  MUX2_X1 U377 ( .A(n551), .B(n330), .S(n323), .Z(n480) );
  MUX2_X1 U378 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n323), .Z(n482) );
  MUX2_X1 U379 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n323), .Z(n484) );
  MUX2_X1 U380 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n323), .Z(n486) );
  MUX2_X1 U381 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n323), .Z(n488) );
  MUX2_X1 U382 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n323), .Z(n490) );
  MUX2_X1 U383 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n323), .Z(n492) );
  MUX2_X1 U384 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n323), .Z(n494) );
  MUX2_X1 U385 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n323), .Z(n496) );
  MUX2_X1 U386 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n323), .Z(n498) );
  MUX2_X1 U387 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n323), .Z(n500) );
  MUX2_X1 U388 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n323), .Z(n502) );
  MUX2_X1 U389 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n323), .Z(n504) );
  MUX2_X1 U390 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n323), .Z(n506) );
  MUX2_X1 U391 ( .A(\mult_x_1/n311 ), .B(A_extended[5]), .S(n323), .Z(n508) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n323), .Z(n510) );
  MUX2_X1 U393 ( .A(n552), .B(A_extended[7]), .S(n323), .Z(n512) );
  OR2_X1 U394 ( .A1(n323), .A2(n553), .ZN(n514) );
endmodule


module conv_128_32_DW_mult_pipe_J1_3 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n353, n355, n357, n359, n361, n363, n365,
         n367, n369, n371, n373, n375, n377, n379, n381, n383, n385, n387,
         n389, n391, n393, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n405, n407, n409, n411, n413, n415, n417, n419, n421, n423,
         n425, n427, n429, n431, n433, n435, n437, n439, n441, n443, n445,
         n447, n449, n451, n453, n455, n457, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n514, n516, n517, n519, n520, n522, n523, n525, n526, n528,
         n530, n532, n534, n536, n538, n540, n542, n544, n546, n548, n549,
         n550, n551;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n401), .SE(n511), .CK(clk), .Q(n550), 
        .QN(n50) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n401), .SE(n503), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n401), .SE(n499), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n47) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n401), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n37) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n401), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n40) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n401), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n46) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n402), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n42) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n403), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n41) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n401), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n43) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n401), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n44) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n401), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n45) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n401), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n401), .SE(n477), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n401), .SE(n475), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n401), .SE(n473), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n401), .SE(n471), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n401), .SE(n469), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n403), .SE(n467), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n401), .SE(n465), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n402), .SE(n463), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n401), .SE(n461), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n401), .SE(n459), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n401), .SE(n457), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n401), .SE(n455), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n401), .SE(n453), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n401), .SE(n451), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n401), .SE(n449), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n403), .SE(n447), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n403), .SE(n445), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n403), .SE(n443), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n403), .SE(n441), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n403), .SE(n439), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n403), .SE(n437), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n403), .SE(n435), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n403), .SE(n433), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n403), .SE(n431), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n403), .SE(n429), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n403), .SE(n427), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n402), .SE(n425), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n402), .SE(n423), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n402), .SE(n421), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n402), .SE(n419), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n402), .SE(n417), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n402), .SE(n415), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n402), .SE(n413), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n402), .SE(n411), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n402), .SE(n409), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n402), .SE(n407), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n402), .SE(n405), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2  ( .D(n551), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n551), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n551), .SE(n357), .CK(
        clk), .Q(n5), .QN(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n551), .SE(n359), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n551), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n337), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n551), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n335), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n551), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n338), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n551), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n334), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n551), .SE(n393), .CK(
        clk), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n551), .SE(n391), .CK(
        clk), .Q(n328), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n551), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n551), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n347), .QN(n53) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n551), .SE(n385), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n551), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n551), .SE(n381), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n551), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n551), .SE(n377), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n551), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n341), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n551), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n340), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n551), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n551), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n551), .SE(n351), .CK(
        clk), .QN(n329) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n401), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n327) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n401), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n39) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n401), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n38) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n401), .SE(n507), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n48) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n401), .SE(n497), .CK(clk), .Q(n549), 
        .QN(n51) );
  BUF_X1 U2 ( .A(n401), .Z(n402) );
  INV_X2 U3 ( .A(n551), .ZN(n401) );
  INV_X1 U4 ( .A(n31), .ZN(n7) );
  OR2_X1 U5 ( .A1(n269), .A2(n5), .ZN(n8) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(n245) );
  NAND2_X1 U7 ( .A1(n23), .A2(n22), .ZN(n238) );
  XNOR2_X1 U8 ( .A(n122), .B(n19), .ZN(n195) );
  NAND2_X1 U9 ( .A1(n242), .A2(n12), .ZN(n11) );
  NAND2_X1 U10 ( .A1(n236), .A2(n24), .ZN(n23) );
  XNOR2_X1 U11 ( .A(n30), .B(n29), .ZN(n232) );
  XNOR2_X1 U12 ( .A(n124), .B(n123), .ZN(n19) );
  OR2_X1 U13 ( .A1(n237), .A2(n49), .ZN(n24) );
  NAND2_X1 U14 ( .A1(n237), .A2(n49), .ZN(n22) );
  NAND2_X1 U15 ( .A1(n14), .A2(n13), .ZN(n12) );
  OR2_X1 U16 ( .A1(n124), .A2(n123), .ZN(n18) );
  NAND2_X1 U17 ( .A1(n124), .A2(n123), .ZN(n16) );
  BUF_X1 U18 ( .A(n401), .Z(n403) );
  INV_X1 U19 ( .A(n243), .ZN(n14) );
  INV_X1 U20 ( .A(n244), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n243), .A2(n244), .ZN(n10) );
  XNOR2_X1 U22 ( .A(n229), .B(n230), .ZN(n30) );
  OR2_X1 U23 ( .A1(n88), .A2(n87), .ZN(n225) );
  INV_X1 U24 ( .A(rst_n), .ZN(n551) );
  NAND2_X1 U25 ( .A1(n55), .A2(n56), .ZN(n147) );
  BUF_X2 U26 ( .A(n72), .Z(n6) );
  NAND2_X1 U27 ( .A1(n67), .A2(n34), .ZN(n206) );
  AND2_X1 U28 ( .A1(n550), .A2(\mult_x_1/n281 ), .ZN(n117) );
  NAND2_X1 U29 ( .A1(n9), .A2(n8), .ZN(n357) );
  OAI21_X1 U30 ( .B1(n179), .B2(n178), .A(n269), .ZN(n9) );
  NAND2_X1 U31 ( .A1(n175), .A2(n176), .ZN(n177) );
  XNOR2_X1 U32 ( .A(n242), .B(n15), .ZN(n176) );
  XNOR2_X1 U33 ( .A(n244), .B(n243), .ZN(n15) );
  NAND2_X1 U34 ( .A1(n17), .A2(n16), .ZN(n159) );
  NAND2_X1 U35 ( .A1(n122), .A2(n18), .ZN(n17) );
  NAND2_X1 U36 ( .A1(n21), .A2(n20), .ZN(n119) );
  INV_X1 U37 ( .A(n61), .ZN(n20) );
  NAND2_X1 U38 ( .A1(n6), .A2(n138), .ZN(n21) );
  XNOR2_X1 U39 ( .A(n236), .B(n25), .ZN(n93) );
  XNOR2_X1 U40 ( .A(n237), .B(n49), .ZN(n25) );
  NAND2_X1 U41 ( .A1(n27), .A2(n26), .ZN(n219) );
  NAND2_X1 U42 ( .A1(n229), .A2(n230), .ZN(n26) );
  NAND2_X1 U43 ( .A1(n29), .A2(n28), .ZN(n27) );
  OR2_X1 U44 ( .A1(n229), .A2(n230), .ZN(n28) );
  NAND2_X1 U45 ( .A1(n77), .A2(n76), .ZN(n29) );
  OAI21_X1 U46 ( .B1(n65), .B2(n63), .A(n62), .ZN(n58) );
  XNOR2_X1 U47 ( .A(n86), .B(n85), .ZN(n237) );
  NAND2_X1 U48 ( .A1(n58), .A2(n57), .ZN(n124) );
  NAND2_X1 U49 ( .A1(n65), .A2(n63), .ZN(n57) );
  XNOR2_X1 U50 ( .A(n65), .B(n64), .ZN(n221) );
  XNOR2_X1 U51 ( .A(n63), .B(n62), .ZN(n64) );
  NAND2_X1 U52 ( .A1(n79), .A2(n78), .ZN(n355) );
  NAND2_X1 U53 ( .A1(n116), .A2(n331), .ZN(n78) );
  OAI21_X1 U54 ( .B1(n195), .B2(n194), .A(n269), .ZN(n79) );
  XOR2_X1 U55 ( .A(n327), .B(n48), .Z(n31) );
  INV_X1 U56 ( .A(n38), .ZN(n32) );
  OAI22_X1 U57 ( .A1(n206), .A2(n81), .B1(n70), .B2(n68), .ZN(n33) );
  XNOR2_X1 U58 ( .A(n47), .B(n51), .ZN(n34) );
  OAI22_X1 U59 ( .A1(n206), .A2(n81), .B1(n70), .B2(n68), .ZN(n227) );
  INV_X1 U60 ( .A(n39), .ZN(n35) );
  OAI22_X1 U61 ( .A1(n6), .A2(n80), .B1(n138), .B2(n74), .ZN(n36) );
  XNOR2_X1 U62 ( .A(n327), .B(n48), .ZN(n56) );
  XNOR2_X1 U63 ( .A(n47), .B(n51), .ZN(n68) );
  AND2_X1 U64 ( .A1(n105), .A2(n104), .ZN(n49) );
  XOR2_X1 U65 ( .A(n105), .B(n104), .Z(n52) );
  XOR2_X1 U66 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n54) );
  XNOR2_X1 U67 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n60) );
  NAND2_X1 U68 ( .A1(n54), .A2(n60), .ZN(n72) );
  XNOR2_X1 U69 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n73) );
  XNOR2_X1 U70 ( .A(n117), .B(\mult_x_1/n311 ), .ZN(n61) );
  OAI22_X1 U71 ( .A1(n72), .A2(n73), .B1(n61), .B2(n60), .ZN(n120) );
  INV_X1 U72 ( .A(n120), .ZN(n65) );
  XNOR2_X1 U73 ( .A(n48), .B(\mult_x_1/n310 ), .ZN(n55) );
  XNOR2_X1 U74 ( .A(n32), .B(\mult_x_1/n283 ), .ZN(n66) );
  XNOR2_X1 U75 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n59) );
  OAI22_X1 U76 ( .A1(n147), .A2(n66), .B1(n7), .B2(n59), .ZN(n63) );
  NAND2_X1 U77 ( .A1(n50), .A2(n32), .ZN(n149) );
  NOR2_X1 U78 ( .A1(n41), .A2(n149), .ZN(n62) );
  NOR2_X1 U79 ( .A1(n42), .A2(n149), .ZN(n123) );
  XNOR2_X1 U80 ( .A(n32), .B(\mult_x_1/n281 ), .ZN(n118) );
  OAI22_X1 U81 ( .A1(n147), .A2(n59), .B1(n7), .B2(n118), .ZN(n121) );
  INV_X1 U82 ( .A(n60), .ZN(n112) );
  INV_X1 U83 ( .A(n112), .ZN(n138) );
  XNOR2_X1 U84 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n75) );
  OAI22_X1 U85 ( .A1(n147), .A2(n75), .B1(n7), .B2(n66), .ZN(n228) );
  XNOR2_X1 U86 ( .A(\mult_x_1/n312 ), .B(n47), .ZN(n67) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n81) );
  XNOR2_X1 U88 ( .A(n117), .B(\mult_x_1/n312 ), .ZN(n70) );
  INV_X1 U89 ( .A(n68), .ZN(n69) );
  AOI21_X1 U90 ( .B1(n68), .B2(n206), .A(n70), .ZN(n71) );
  INV_X1 U91 ( .A(n71), .ZN(n226) );
  NOR2_X1 U92 ( .A1(n43), .A2(n149), .ZN(n230) );
  XNOR2_X1 U93 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n74) );
  OAI22_X1 U94 ( .A1(n6), .A2(n74), .B1(n138), .B2(n73), .ZN(n229) );
  XNOR2_X1 U95 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n80) );
  OAI22_X1 U96 ( .A1(n6), .A2(n80), .B1(n138), .B2(n74), .ZN(n84) );
  XNOR2_X1 U97 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n91) );
  OAI22_X1 U98 ( .A1(n147), .A2(n91), .B1(n7), .B2(n75), .ZN(n83) );
  INV_X1 U99 ( .A(n227), .ZN(n85) );
  OAI21_X1 U100 ( .B1(n84), .B2(n83), .A(n85), .ZN(n77) );
  NAND2_X1 U101 ( .A1(n36), .A2(n83), .ZN(n76) );
  INV_X1 U102 ( .A(en), .ZN(n116) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n99) );
  OAI22_X1 U104 ( .A1(n6), .A2(n99), .B1(n138), .B2(n80), .ZN(n88) );
  XNOR2_X1 U105 ( .A(n35), .B(\mult_x_1/n282 ), .ZN(n100) );
  OAI22_X1 U106 ( .A1(n206), .A2(n100), .B1(n68), .B2(n81), .ZN(n87) );
  XNOR2_X1 U107 ( .A(n88), .B(n87), .ZN(n105) );
  XNOR2_X1 U108 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n102) );
  XNOR2_X1 U109 ( .A(n32), .B(\mult_x_1/n286 ), .ZN(n92) );
  OAI22_X1 U110 ( .A1(n147), .A2(n102), .B1(n7), .B2(n92), .ZN(n164) );
  NAND2_X1 U111 ( .A1(n549), .A2(n37), .ZN(n209) );
  XNOR2_X1 U112 ( .A(n549), .B(\mult_x_1/n281 ), .ZN(n131) );
  XNOR2_X1 U113 ( .A(n117), .B(n549), .ZN(n89) );
  OAI22_X1 U114 ( .A1(n209), .A2(n131), .B1(n89), .B2(n37), .ZN(n163) );
  INV_X1 U115 ( .A(n149), .ZN(n82) );
  AND2_X1 U116 ( .A1(\mult_x_1/n288 ), .A2(n82), .ZN(n162) );
  XNOR2_X1 U117 ( .A(n36), .B(n83), .ZN(n86) );
  NOR2_X1 U118 ( .A1(n44), .A2(n149), .ZN(n224) );
  AOI21_X1 U119 ( .B1(n209), .B2(n37), .A(n89), .ZN(n90) );
  INV_X1 U120 ( .A(n90), .ZN(n98) );
  OAI22_X1 U121 ( .A1(n147), .A2(n92), .B1(n7), .B2(n91), .ZN(n97) );
  NOR2_X1 U122 ( .A1(n45), .A2(n149), .ZN(n96) );
  NAND2_X1 U123 ( .A1(n93), .A2(n269), .ZN(n95) );
  OR2_X1 U124 ( .A1(n269), .A2(n53), .ZN(n94) );
  NAND2_X1 U125 ( .A1(n95), .A2(n94), .ZN(n387) );
  FA_X1 U126 ( .A(n98), .B(n97), .CI(n96), .CO(n223), .S(n240) );
  XNOR2_X1 U127 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n285 ), .ZN(n130) );
  OAI22_X1 U128 ( .A1(n6), .A2(n130), .B1(n138), .B2(n99), .ZN(n170) );
  XNOR2_X1 U129 ( .A(n35), .B(\mult_x_1/n283 ), .ZN(n133) );
  OAI22_X1 U130 ( .A1(n206), .A2(n133), .B1(n68), .B2(n100), .ZN(n169) );
  OR2_X1 U131 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n101) );
  OAI22_X1 U132 ( .A1(n147), .A2(n38), .B1(n101), .B2(n7), .ZN(n129) );
  XNOR2_X1 U133 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n103) );
  OAI22_X1 U134 ( .A1(n147), .A2(n103), .B1(n7), .B2(n102), .ZN(n128) );
  NAND2_X1 U135 ( .A1(n106), .A2(n269), .ZN(n108) );
  OR2_X1 U136 ( .A1(n269), .A2(n328), .ZN(n107) );
  NAND2_X1 U137 ( .A1(n108), .A2(n107), .ZN(n391) );
  XNOR2_X1 U160 ( .A(n35), .B(\mult_x_1/n286 ), .ZN(n113) );
  XNOR2_X1 U161 ( .A(n35), .B(\mult_x_1/n285 ), .ZN(n127) );
  OAI22_X1 U162 ( .A1(n206), .A2(n113), .B1(n68), .B2(n127), .ZN(n186) );
  XNOR2_X1 U163 ( .A(n549), .B(\mult_x_1/n284 ), .ZN(n111) );
  XNOR2_X1 U164 ( .A(n549), .B(\mult_x_1/n283 ), .ZN(n126) );
  OAI22_X1 U165 ( .A1(n209), .A2(n111), .B1(n126), .B2(n37), .ZN(n185) );
  OR2_X1 U166 ( .A1(\mult_x_1/n288 ), .A2(n327), .ZN(n109) );
  OAI22_X1 U167 ( .A1(n6), .A2(n327), .B1(n109), .B2(n138), .ZN(n136) );
  XNOR2_X1 U168 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n288 ), .ZN(n110) );
  XNOR2_X1 U169 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n139) );
  OAI22_X1 U170 ( .A1(n6), .A2(n110), .B1(n138), .B2(n139), .ZN(n135) );
  XNOR2_X1 U171 ( .A(n549), .B(\mult_x_1/n285 ), .ZN(n202) );
  OAI22_X1 U172 ( .A1(n209), .A2(n202), .B1(n111), .B2(n37), .ZN(n199) );
  AND2_X1 U173 ( .A1(\mult_x_1/n288 ), .A2(n112), .ZN(n198) );
  XNOR2_X1 U174 ( .A(n35), .B(\mult_x_1/n287 ), .ZN(n200) );
  OAI22_X1 U175 ( .A1(n206), .A2(n200), .B1(n68), .B2(n113), .ZN(n197) );
  NOR2_X1 U176 ( .A1(n192), .A2(n191), .ZN(n115) );
  NAND2_X1 U177 ( .A1(n116), .A2(n329), .ZN(n114) );
  OAI21_X1 U178 ( .B1(n116), .B2(n115), .A(n114), .ZN(n351) );
  NOR2_X1 U179 ( .A1(n46), .A2(n149), .ZN(n145) );
  XNOR2_X1 U180 ( .A(n117), .B(n32), .ZN(n146) );
  OAI22_X1 U181 ( .A1(n147), .A2(n118), .B1(n146), .B2(n7), .ZN(n153) );
  INV_X1 U182 ( .A(n153), .ZN(n144) );
  FA_X1 U183 ( .A(n121), .B(n120), .CI(n119), .CO(n143), .S(n122) );
  OR2_X1 U184 ( .A1(n160), .A2(n159), .ZN(n125) );
  MUX2_X1 U185 ( .A(n330), .B(n125), .S(n269), .Z(n353) );
  XNOR2_X1 U186 ( .A(n549), .B(\mult_x_1/n282 ), .ZN(n132) );
  OAI22_X1 U187 ( .A1(n209), .A2(n126), .B1(n132), .B2(n37), .ZN(n142) );
  AND2_X1 U188 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n141) );
  XNOR2_X1 U189 ( .A(n35), .B(\mult_x_1/n284 ), .ZN(n134) );
  OAI22_X1 U190 ( .A1(n206), .A2(n127), .B1(n68), .B2(n134), .ZN(n140) );
  HA_X1 U191 ( .A(n129), .B(n128), .CO(n168), .S(n172) );
  XNOR2_X1 U192 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n286 ), .ZN(n137) );
  OAI22_X1 U193 ( .A1(n6), .A2(n137), .B1(n138), .B2(n130), .ZN(n167) );
  OAI22_X1 U194 ( .A1(n209), .A2(n132), .B1(n131), .B2(n37), .ZN(n166) );
  OAI22_X1 U195 ( .A1(n206), .A2(n134), .B1(n68), .B2(n133), .ZN(n165) );
  HA_X1 U196 ( .A(n136), .B(n135), .CO(n183), .S(n184) );
  OAI22_X1 U197 ( .A1(n6), .A2(n139), .B1(n138), .B2(n137), .ZN(n182) );
  FA_X1 U198 ( .A(n142), .B(n141), .CI(n140), .CO(n173), .S(n181) );
  FA_X1 U199 ( .A(n145), .B(n144), .CI(n143), .CO(n155), .S(n160) );
  AOI21_X1 U200 ( .B1(n7), .B2(n147), .A(n146), .ZN(n148) );
  INV_X1 U201 ( .A(n148), .ZN(n151) );
  NOR2_X1 U202 ( .A1(n40), .A2(n149), .ZN(n150) );
  XOR2_X1 U203 ( .A(n151), .B(n150), .Z(n152) );
  XOR2_X1 U204 ( .A(n153), .B(n152), .Z(n154) );
  OR2_X1 U205 ( .A1(n155), .A2(n154), .ZN(n157) );
  NAND2_X1 U206 ( .A1(n155), .A2(n154), .ZN(n156) );
  NAND2_X1 U207 ( .A1(n157), .A2(n156), .ZN(n158) );
  MUX2_X1 U208 ( .A(n333), .B(n158), .S(n269), .Z(n359) );
  NAND2_X1 U209 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2_X1 U210 ( .A(n334), .B(n161), .S(n269), .Z(n361) );
  FA_X1 U211 ( .A(n164), .B(n163), .CI(n162), .CO(n104), .S(n244) );
  FA_X1 U212 ( .A(n165), .B(n166), .CI(n167), .CO(n243), .S(n171) );
  FA_X1 U213 ( .A(n170), .B(n169), .CI(n168), .CO(n239), .S(n242) );
  FA_X1 U214 ( .A(n173), .B(n172), .CI(n171), .CO(n175), .S(n179) );
  NOR2_X1 U215 ( .A1(n176), .A2(n175), .ZN(n174) );
  MUX2_X1 U216 ( .A(n335), .B(n174), .S(n269), .Z(n363) );
  MUX2_X1 U217 ( .A(n336), .B(n177), .S(n269), .Z(n365) );
  NAND2_X1 U218 ( .A1(n179), .A2(n178), .ZN(n180) );
  MUX2_X1 U219 ( .A(n337), .B(n180), .S(n269), .Z(n367) );
  FA_X1 U220 ( .A(n183), .B(n182), .CI(n181), .CO(n178), .S(n189) );
  FA_X1 U221 ( .A(n186), .B(n185), .CI(n184), .CO(n188), .S(n192) );
  NOR2_X1 U222 ( .A1(n189), .A2(n188), .ZN(n187) );
  MUX2_X1 U223 ( .A(n338), .B(n187), .S(n269), .Z(n369) );
  NAND2_X1 U224 ( .A1(n189), .A2(n188), .ZN(n190) );
  MUX2_X1 U225 ( .A(n339), .B(n190), .S(n269), .Z(n371) );
  NAND2_X1 U226 ( .A1(n192), .A2(n191), .ZN(n193) );
  MUX2_X1 U227 ( .A(n340), .B(n193), .S(n269), .Z(n373) );
  NAND2_X1 U228 ( .A1(n195), .A2(n194), .ZN(n196) );
  MUX2_X1 U229 ( .A(n341), .B(n196), .S(n269), .Z(n375) );
  FA_X1 U230 ( .A(n199), .B(n198), .CI(n197), .CO(n191), .S(n217) );
  XNOR2_X1 U231 ( .A(n35), .B(\mult_x_1/n288 ), .ZN(n201) );
  OAI22_X1 U232 ( .A1(n206), .A2(n201), .B1(n68), .B2(n200), .ZN(n204) );
  XNOR2_X1 U233 ( .A(n549), .B(\mult_x_1/n286 ), .ZN(n207) );
  OAI22_X1 U234 ( .A1(n209), .A2(n207), .B1(n202), .B2(n37), .ZN(n203) );
  NOR2_X1 U235 ( .A1(n217), .A2(n216), .ZN(n262) );
  HA_X1 U236 ( .A(n204), .B(n203), .CO(n216), .S(n214) );
  OR2_X1 U237 ( .A1(\mult_x_1/n288 ), .A2(n39), .ZN(n205) );
  OAI22_X1 U238 ( .A1(n206), .A2(n39), .B1(n205), .B2(n68), .ZN(n213) );
  OR2_X1 U239 ( .A1(n214), .A2(n213), .ZN(n258) );
  XNOR2_X1 U240 ( .A(n549), .B(\mult_x_1/n287 ), .ZN(n208) );
  OAI22_X1 U241 ( .A1(n209), .A2(n208), .B1(n207), .B2(n37), .ZN(n212) );
  AND2_X1 U242 ( .A1(\mult_x_1/n288 ), .A2(n69), .ZN(n211) );
  NOR2_X1 U243 ( .A1(n212), .A2(n211), .ZN(n251) );
  OAI22_X1 U244 ( .A1(n209), .A2(\mult_x_1/n288 ), .B1(n208), .B2(n37), .ZN(
        n248) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n51), .ZN(n210) );
  NAND2_X1 U246 ( .A1(n210), .A2(n209), .ZN(n247) );
  NAND2_X1 U247 ( .A1(n248), .A2(n247), .ZN(n254) );
  NAND2_X1 U248 ( .A1(n212), .A2(n211), .ZN(n252) );
  OAI21_X1 U249 ( .B1(n251), .B2(n254), .A(n252), .ZN(n259) );
  NAND2_X1 U250 ( .A1(n214), .A2(n213), .ZN(n257) );
  INV_X1 U251 ( .A(n257), .ZN(n215) );
  AOI21_X1 U252 ( .B1(n258), .B2(n259), .A(n215), .ZN(n265) );
  NAND2_X1 U253 ( .A1(n217), .A2(n216), .ZN(n263) );
  OAI21_X1 U254 ( .B1(n262), .B2(n265), .A(n263), .ZN(n218) );
  MUX2_X1 U255 ( .A(n342), .B(n218), .S(n269), .Z(n377) );
  FA_X1 U256 ( .A(n221), .B(n220), .CI(n219), .CO(n194), .S(n222) );
  MUX2_X1 U257 ( .A(n343), .B(n222), .S(n269), .Z(n379) );
  FA_X1 U258 ( .A(n225), .B(n224), .CI(n223), .CO(n234), .S(n236) );
  FA_X1 U259 ( .A(n228), .B(n33), .CI(n226), .CO(n220), .S(n233) );
  MUX2_X1 U260 ( .A(n344), .B(n231), .S(n269), .Z(n381) );
  FA_X1 U261 ( .A(n234), .B(n233), .CI(n232), .CO(n231), .S(n235) );
  MUX2_X1 U262 ( .A(n345), .B(n235), .S(n269), .Z(n383) );
  MUX2_X1 U263 ( .A(n346), .B(n238), .S(n269), .Z(n385) );
  FA_X1 U264 ( .A(n240), .B(n239), .CI(n52), .CO(n241), .S(n106) );
  MUX2_X1 U265 ( .A(n348), .B(n241), .S(n269), .Z(n389) );
  MUX2_X1 U266 ( .A(n350), .B(n245), .S(n269), .Z(n393) );
  BUF_X4 U267 ( .A(en), .Z(n269) );
  MUX2_X1 U268 ( .A(product[0]), .B(n513), .S(n269), .Z(n405) );
  MUX2_X1 U269 ( .A(n513), .B(n514), .S(n269), .Z(n407) );
  AND2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n246) );
  MUX2_X1 U271 ( .A(n514), .B(n246), .S(n269), .Z(n409) );
  MUX2_X1 U272 ( .A(product[1]), .B(n516), .S(n269), .Z(n411) );
  MUX2_X1 U273 ( .A(n516), .B(n517), .S(n269), .Z(n413) );
  OR2_X1 U274 ( .A1(n248), .A2(n247), .ZN(n249) );
  AND2_X1 U275 ( .A1(n249), .A2(n254), .ZN(n250) );
  MUX2_X1 U276 ( .A(n517), .B(n250), .S(n269), .Z(n415) );
  MUX2_X1 U277 ( .A(product[2]), .B(n519), .S(n269), .Z(n417) );
  MUX2_X1 U278 ( .A(n519), .B(n520), .S(n269), .Z(n419) );
  INV_X1 U279 ( .A(n251), .ZN(n253) );
  NAND2_X1 U280 ( .A1(n253), .A2(n252), .ZN(n255) );
  XOR2_X1 U281 ( .A(n255), .B(n254), .Z(n256) );
  MUX2_X1 U282 ( .A(n520), .B(n256), .S(n269), .Z(n421) );
  MUX2_X1 U283 ( .A(product[3]), .B(n522), .S(n269), .Z(n423) );
  MUX2_X1 U284 ( .A(n522), .B(n523), .S(n269), .Z(n425) );
  NAND2_X1 U285 ( .A1(n258), .A2(n257), .ZN(n260) );
  XNOR2_X1 U286 ( .A(n260), .B(n259), .ZN(n261) );
  MUX2_X1 U287 ( .A(n523), .B(n261), .S(n269), .Z(n427) );
  MUX2_X1 U288 ( .A(product[4]), .B(n525), .S(n269), .Z(n429) );
  MUX2_X1 U289 ( .A(n525), .B(n526), .S(n269), .Z(n431) );
  INV_X1 U290 ( .A(n262), .ZN(n264) );
  NAND2_X1 U291 ( .A1(n264), .A2(n263), .ZN(n266) );
  XOR2_X1 U292 ( .A(n266), .B(n265), .Z(n267) );
  MUX2_X1 U293 ( .A(n526), .B(n267), .S(n269), .Z(n433) );
  MUX2_X1 U294 ( .A(product[5]), .B(n528), .S(n269), .Z(n435) );
  NAND2_X1 U295 ( .A1(n329), .A2(n340), .ZN(n268) );
  XNOR2_X1 U296 ( .A(n268), .B(n342), .ZN(n270) );
  MUX2_X1 U297 ( .A(n528), .B(n270), .S(n269), .Z(n437) );
  CLKBUF_X1 U298 ( .A(en), .Z(n319) );
  MUX2_X1 U299 ( .A(product[6]), .B(n530), .S(n319), .Z(n439) );
  NAND2_X1 U300 ( .A1(n398), .A2(n339), .ZN(n271) );
  AOI21_X1 U301 ( .B1(n329), .B2(n342), .A(n397), .ZN(n273) );
  XOR2_X1 U302 ( .A(n271), .B(n273), .Z(n272) );
  MUX2_X1 U303 ( .A(n530), .B(n272), .S(n319), .Z(n441) );
  MUX2_X1 U304 ( .A(product[7]), .B(n532), .S(n319), .Z(n443) );
  OAI21_X1 U305 ( .B1(n338), .B2(n273), .A(n339), .ZN(n276) );
  NAND2_X1 U306 ( .A1(n332), .A2(n337), .ZN(n274) );
  XNOR2_X1 U307 ( .A(n276), .B(n274), .ZN(n275) );
  MUX2_X1 U308 ( .A(n532), .B(n275), .S(n319), .Z(n445) );
  MUX2_X1 U309 ( .A(product[8]), .B(n534), .S(n319), .Z(n447) );
  AOI21_X1 U310 ( .B1(n276), .B2(n332), .A(n400), .ZN(n279) );
  NAND2_X1 U311 ( .A1(n399), .A2(n336), .ZN(n277) );
  XOR2_X1 U312 ( .A(n279), .B(n277), .Z(n278) );
  MUX2_X1 U313 ( .A(n534), .B(n278), .S(n319), .Z(n449) );
  MUX2_X1 U314 ( .A(product[9]), .B(n536), .S(n319), .Z(n451) );
  OAI21_X1 U315 ( .B1(n279), .B2(n335), .A(n336), .ZN(n293) );
  INV_X1 U316 ( .A(n293), .ZN(n283) );
  NOR2_X1 U317 ( .A1(n349), .A2(n350), .ZN(n288) );
  INV_X1 U318 ( .A(n288), .ZN(n280) );
  NAND2_X1 U319 ( .A1(n349), .A2(n350), .ZN(n290) );
  NAND2_X1 U320 ( .A1(n280), .A2(n290), .ZN(n281) );
  XOR2_X1 U321 ( .A(n283), .B(n281), .Z(n282) );
  MUX2_X1 U322 ( .A(n536), .B(n282), .S(n319), .Z(n453) );
  MUX2_X1 U323 ( .A(product[10]), .B(n538), .S(n319), .Z(n455) );
  OAI21_X1 U324 ( .B1(n283), .B2(n288), .A(n290), .ZN(n286) );
  NOR2_X1 U325 ( .A1(n347), .A2(n348), .ZN(n291) );
  INV_X1 U326 ( .A(n291), .ZN(n284) );
  NAND2_X1 U327 ( .A1(n347), .A2(n348), .ZN(n289) );
  NAND2_X1 U328 ( .A1(n284), .A2(n289), .ZN(n285) );
  XNOR2_X1 U329 ( .A(n286), .B(n285), .ZN(n287) );
  MUX2_X1 U330 ( .A(n538), .B(n287), .S(n319), .Z(n457) );
  MUX2_X1 U331 ( .A(product[11]), .B(n540), .S(n319), .Z(n459) );
  NOR2_X1 U332 ( .A1(n291), .A2(n288), .ZN(n294) );
  OAI21_X1 U333 ( .B1(n291), .B2(n290), .A(n289), .ZN(n292) );
  AOI21_X1 U334 ( .B1(n294), .B2(n293), .A(n292), .ZN(n324) );
  NOR2_X1 U335 ( .A1(n345), .A2(n346), .ZN(n309) );
  INV_X1 U336 ( .A(n309), .ZN(n300) );
  NAND2_X1 U337 ( .A1(n345), .A2(n346), .ZN(n312) );
  NAND2_X1 U338 ( .A1(n300), .A2(n312), .ZN(n295) );
  XOR2_X1 U339 ( .A(n324), .B(n295), .Z(n296) );
  MUX2_X1 U340 ( .A(n540), .B(n296), .S(n319), .Z(n461) );
  MUX2_X1 U341 ( .A(product[12]), .B(n542), .S(n319), .Z(n463) );
  OAI21_X1 U342 ( .B1(n324), .B2(n309), .A(n312), .ZN(n298) );
  OR2_X1 U343 ( .A1(n343), .A2(n344), .ZN(n308) );
  NAND2_X1 U344 ( .A1(n343), .A2(n344), .ZN(n301) );
  NAND2_X1 U345 ( .A1(n308), .A2(n301), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  MUX2_X1 U347 ( .A(n542), .B(n299), .S(n319), .Z(n465) );
  MUX2_X1 U348 ( .A(product[13]), .B(n544), .S(n319), .Z(n467) );
  NAND2_X1 U349 ( .A1(n300), .A2(n308), .ZN(n304) );
  INV_X1 U350 ( .A(n312), .ZN(n302) );
  INV_X1 U351 ( .A(n301), .ZN(n310) );
  AOI21_X1 U352 ( .B1(n302), .B2(n308), .A(n310), .ZN(n303) );
  OAI21_X1 U353 ( .B1(n324), .B2(n304), .A(n303), .ZN(n306) );
  NAND2_X1 U354 ( .A1(n331), .A2(n341), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U356 ( .A(n544), .B(n307), .S(n319), .Z(n469) );
  MUX2_X1 U357 ( .A(product[14]), .B(n546), .S(n319), .Z(n471) );
  NAND2_X1 U358 ( .A1(n308), .A2(n331), .ZN(n313) );
  NOR2_X1 U359 ( .A1(n309), .A2(n313), .ZN(n320) );
  INV_X1 U360 ( .A(n320), .ZN(n315) );
  AOI21_X1 U361 ( .B1(n310), .B2(n331), .A(n395), .ZN(n311) );
  OAI21_X1 U362 ( .B1(n313), .B2(n312), .A(n311), .ZN(n321) );
  INV_X1 U363 ( .A(n321), .ZN(n314) );
  OAI21_X1 U364 ( .B1(n324), .B2(n315), .A(n314), .ZN(n317) );
  NAND2_X1 U365 ( .A1(n330), .A2(n334), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U367 ( .A(n546), .B(n318), .S(n319), .Z(n473) );
  MUX2_X1 U368 ( .A(product[15]), .B(n548), .S(n319), .Z(n475) );
  NAND2_X1 U369 ( .A1(n320), .A2(n330), .ZN(n323) );
  AOI21_X1 U370 ( .B1(n321), .B2(n330), .A(n396), .ZN(n322) );
  OAI21_X1 U371 ( .B1(n324), .B2(n323), .A(n322), .ZN(n325) );
  XNOR2_X1 U372 ( .A(n325), .B(n333), .ZN(n326) );
  MUX2_X1 U373 ( .A(n548), .B(n326), .S(n269), .Z(n477) );
  MUX2_X1 U374 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n269), .Z(n479) );
  MUX2_X1 U375 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n269), .Z(n481) );
  MUX2_X1 U376 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n269), .Z(n483) );
  MUX2_X1 U377 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n269), .Z(n485) );
  MUX2_X1 U378 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n269), .Z(n487) );
  MUX2_X1 U379 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n269), .Z(n489) );
  MUX2_X1 U380 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n269), .Z(n491) );
  MUX2_X1 U381 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n269), .Z(n493) );
  MUX2_X1 U382 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n269), .Z(n495) );
  MUX2_X1 U383 ( .A(n549), .B(A_extended[1]), .S(n269), .Z(n497) );
  MUX2_X1 U384 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n269), .Z(n499) );
  MUX2_X1 U385 ( .A(n35), .B(A_extended[3]), .S(n269), .Z(n501) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n269), .Z(n503) );
  MUX2_X1 U387 ( .A(\mult_x_1/n311 ), .B(A_extended[5]), .S(n269), .Z(n505) );
  MUX2_X1 U388 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n269), .Z(n507) );
  MUX2_X1 U389 ( .A(n32), .B(A_extended[7]), .S(n269), .Z(n509) );
  OR2_X1 U390 ( .A1(n269), .A2(n550), .ZN(n511) );
endmodule


module conv_128_32_DW_mult_pipe_J1_4 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n345, n347, n349, n351, n353, n355, n357, n359, n361, n363,
         n365, n367, n369, n371, n373, n375, n377, n379, n381, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n396,
         n398, n400, n402, n404, n406, n408, n410, n412, n414, n416, n418,
         n420, n422, n424, n426, n428, n430, n432, n434, n436, n438, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n458, n460, n462,
         n464, n466, n468, n470, n472, n474, n476, n478, n480, n482, n484,
         n486, n488, n490, n492, n494, n496, n498, n500, n502, n504, n506,
         n507, n509, n510, n512, n513, n515, n516, n518, n519, n521, n522,
         n524, n526, n528, n530, n532, n534, n536, n538, n540, n542, n543,
         n544, n545, n546, n547;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n394), .SE(n504), .CK(clk), .Q(n546), 
        .QN(n29) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n394), .SE(n502), .CK(clk), .Q(n545), 
        .QN(n32) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n394), .SE(n500), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n394), .SE(n496), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n394), .SE(n492), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n28) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n394), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n30) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n394), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n33) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n394), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n36) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n394), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n38) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n392), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n37) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n393), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n39) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n391), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n41) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n391), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n40) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n391), .SE(n472), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n391), .SE(n470), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n391), .SE(n468), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n391), .SE(n466), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n391), .SE(n464), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n391), .SE(n462), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n394), .SE(n460), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n393), .SE(n458), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n392), .SE(n456), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n391), .SE(n454), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n391), .SE(n452), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n391), .SE(n450), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n391), .SE(n448), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n391), .SE(n446), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n391), .SE(n444), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n391), .SE(n442), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n391), .SE(n440), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n393), .SE(n438), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n393), .SE(n436), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n393), .SE(n434), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n393), .SE(n432), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n393), .SE(n430), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n393), .SE(n428), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n393), .SE(n426), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n393), .SE(n424), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n393), .SE(n422), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n393), .SE(n420), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n393), .SE(n418), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n392), .SE(n416), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n392), .SE(n414), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n392), .SE(n412), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n392), .SE(n410), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n392), .SE(n408), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n392), .SE(n406), .CK(clk), .Q(n510)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n392), .SE(n404), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n392), .SE(n402), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n392), .SE(n400), .CK(clk), .Q(n507)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n392), .SE(n398), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n392), .SE(n396), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n547), .SE(n381), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2  ( .D(n547), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n547), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2_IP  ( .D(1'b1), .SI(n547), .SE(n375), .CK(
        clk), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG15_S2_IP  ( .D(1'b1), .SI(n547), .SE(n373), .CK(
        clk), .Q(n389), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2  ( .D(n547), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n337), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n547), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n547), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n335), .QN(n385) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n547), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n334), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n547), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n333), .QN(n44) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n547), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n332), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n547), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n547), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n330), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n547), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n329), .QN(n383) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n547), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n328), .QN(n384) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n547), .SE(n351), .CK(
        clk), .QN(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n547), .SE(n349), .CK(
        clk), .QN(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n547), .SI(1'b1), .SE(n347), .CK(clk), 
        .Q(n325) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n547), .SI(1'b1), .SE(n345), .CK(clk), 
        .Q(n324) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n547), .SI(1'b1), .SE(n343), .CK(clk), 
        .Q(n323) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n394), .SE(n498), .CK(clk), .Q(n544), 
        .QN(n34) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n394), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n35) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n394), .SE(n490), .CK(clk), .Q(n543), 
        .QN(n43) );
  BUF_X1 U2 ( .A(n391), .Z(n394) );
  BUF_X1 U3 ( .A(n391), .Z(n392) );
  BUF_X1 U4 ( .A(n391), .Z(n393) );
  INV_X1 U5 ( .A(n547), .ZN(n391) );
  NAND2_X1 U6 ( .A1(n13), .A2(n12), .ZN(n151) );
  OAI21_X1 U7 ( .B1(n99), .B2(n98), .A(n14), .ZN(n13) );
  NAND3_X1 U8 ( .A1(n95), .A2(n96), .A3(n94), .ZN(n14) );
  MUX2_X1 U9 ( .A(n332), .B(n175), .S(en), .Z(n361) );
  BUF_X2 U10 ( .A(en), .Z(n279) );
  BUF_X4 U11 ( .A(en), .Z(n322) );
  NAND2_X1 U12 ( .A1(n99), .A2(n98), .ZN(n12) );
  OR2_X1 U13 ( .A1(n21), .A2(n154), .ZN(n198) );
  INV_X1 U14 ( .A(rst_n), .ZN(n547) );
  AND2_X1 U15 ( .A1(n63), .A2(n17), .ZN(n159) );
  INV_X1 U16 ( .A(n17), .ZN(n16) );
  OAI22_X1 U17 ( .A1(n135), .A2(n60), .B1(n136), .B2(n59), .ZN(n17) );
  AND2_X1 U18 ( .A1(n546), .A2(\mult_x_1/n281 ), .ZN(n87) );
  NAND2_X1 U19 ( .A1(n9), .A2(n7), .ZN(n371) );
  NAND2_X1 U20 ( .A1(n8), .A2(n337), .ZN(n7) );
  INV_X1 U21 ( .A(n322), .ZN(n8) );
  NAND2_X1 U22 ( .A1(n10), .A2(n322), .ZN(n9) );
  NAND2_X1 U23 ( .A1(n191), .A2(n190), .ZN(n10) );
  XNOR2_X1 U24 ( .A(n11), .B(n85), .ZN(n99) );
  XNOR2_X1 U25 ( .A(n83), .B(n84), .ZN(n11) );
  XNOR2_X1 U26 ( .A(n15), .B(n14), .ZN(n191) );
  XNOR2_X1 U27 ( .A(n99), .B(n98), .ZN(n15) );
  XNOR2_X1 U28 ( .A(n63), .B(n16), .ZN(n120) );
  INV_X1 U29 ( .A(n200), .ZN(n110) );
  NOR2_X1 U30 ( .A1(n198), .A2(n197), .ZN(n109) );
  NAND2_X1 U31 ( .A1(n198), .A2(n197), .ZN(n108) );
  NAND2_X1 U32 ( .A1(n75), .A2(n74), .ZN(n82) );
  XNOR2_X1 U33 ( .A(n31), .B(n165), .ZN(n171) );
  XNOR2_X1 U34 ( .A(n203), .B(n202), .ZN(n165) );
  NAND2_X1 U35 ( .A1(n205), .A2(n204), .ZN(n207) );
  NAND2_X1 U36 ( .A1(n203), .A2(n202), .ZN(n204) );
  NAND2_X1 U37 ( .A1(n31), .A2(n201), .ZN(n205) );
  OR2_X1 U38 ( .A1(n202), .A2(n203), .ZN(n201) );
  OAI21_X1 U39 ( .B1(n110), .B2(n109), .A(n108), .ZN(n244) );
  NAND2_X2 U40 ( .A1(n54), .A2(n53), .ZN(n88) );
  INV_X1 U41 ( .A(n55), .ZN(n18) );
  INV_X1 U42 ( .A(n55), .ZN(n226) );
  INV_X1 U43 ( .A(n32), .ZN(n19) );
  BUF_X2 U44 ( .A(\mult_x_1/n312 ), .Z(n20) );
  OAI22_X1 U45 ( .A1(n126), .A2(n105), .B1(n214), .B2(n104), .ZN(n21) );
  INV_X2 U46 ( .A(n34), .ZN(n22) );
  XOR2_X1 U47 ( .A(n196), .B(n195), .Z(n23) );
  XOR2_X1 U48 ( .A(n194), .B(n23), .Z(n247) );
  NAND2_X1 U49 ( .A1(n194), .A2(n196), .ZN(n24) );
  NAND2_X1 U50 ( .A1(n194), .A2(n195), .ZN(n25) );
  NAND2_X1 U51 ( .A1(n196), .A2(n195), .ZN(n26) );
  NAND3_X1 U52 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n117) );
  OAI22_X1 U53 ( .A1(n18), .A2(n89), .B1(n88), .B2(n106), .ZN(n27) );
  XNOR2_X1 U54 ( .A(n28), .B(n43), .ZN(n54) );
  NAND2_X1 U55 ( .A1(n85), .A2(n83), .ZN(n74) );
  OAI21_X1 U56 ( .B1(n85), .B2(n83), .A(n84), .ZN(n75) );
  XOR2_X1 U57 ( .A(n193), .B(n192), .Z(n31) );
  AND2_X1 U58 ( .A1(n192), .A2(n193), .ZN(n42) );
  XOR2_X1 U59 ( .A(\mult_x_1/a[6] ), .B(n545), .Z(n45) );
  XNOR2_X1 U60 ( .A(\mult_x_1/a[6] ), .B(n544), .ZN(n46) );
  NAND2_X2 U61 ( .A1(n45), .A2(n46), .ZN(n135) );
  XNOR2_X1 U62 ( .A(n545), .B(\mult_x_1/n287 ), .ZN(n59) );
  INV_X1 U63 ( .A(n46), .ZN(n47) );
  INV_X2 U64 ( .A(n47), .ZN(n136) );
  XNOR2_X1 U65 ( .A(n545), .B(\mult_x_1/n286 ), .ZN(n103) );
  OAI22_X1 U66 ( .A1(n135), .A2(n59), .B1(n136), .B2(n103), .ZN(n158) );
  NAND2_X1 U67 ( .A1(n543), .A2(n30), .ZN(n229) );
  XNOR2_X1 U68 ( .A(n543), .B(\mult_x_1/n281 ), .ZN(n52) );
  XNOR2_X1 U69 ( .A(n87), .B(n543), .ZN(n100) );
  OAI22_X1 U70 ( .A1(n229), .A2(n52), .B1(n100), .B2(n30), .ZN(n157) );
  NAND2_X1 U71 ( .A1(n19), .A2(n29), .ZN(n138) );
  INV_X1 U72 ( .A(n138), .ZN(n48) );
  AND2_X1 U73 ( .A1(\mult_x_1/n288 ), .A2(n48), .ZN(n156) );
  XOR2_X1 U74 ( .A(\mult_x_1/a[4] ), .B(n544), .Z(n49) );
  XNOR2_X1 U75 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n50) );
  NAND2_X1 U76 ( .A1(n49), .A2(n50), .ZN(n126) );
  XNOR2_X1 U77 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n124) );
  INV_X1 U78 ( .A(n50), .ZN(n51) );
  INV_X2 U79 ( .A(n51), .ZN(n214) );
  XNOR2_X1 U80 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n56) );
  OAI22_X1 U81 ( .A1(n126), .A2(n124), .B1(n214), .B2(n56), .ZN(n66) );
  XNOR2_X1 U82 ( .A(n543), .B(\mult_x_1/n282 ), .ZN(n61) );
  OAI22_X1 U83 ( .A1(n229), .A2(n61), .B1(n52), .B2(n30), .ZN(n65) );
  XOR2_X1 U84 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n53) );
  XNOR2_X1 U85 ( .A(n20), .B(\mult_x_1/n284 ), .ZN(n62) );
  INV_X1 U86 ( .A(n54), .ZN(n55) );
  XNOR2_X1 U87 ( .A(n20), .B(\mult_x_1/n283 ), .ZN(n57) );
  OAI22_X1 U88 ( .A1(n88), .A2(n62), .B1(n18), .B2(n57), .ZN(n64) );
  XNOR2_X1 U89 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n105) );
  OAI22_X1 U90 ( .A1(n126), .A2(n56), .B1(n214), .B2(n105), .ZN(n161) );
  XNOR2_X1 U91 ( .A(n20), .B(\mult_x_1/n282 ), .ZN(n107) );
  OAI22_X1 U92 ( .A1(n88), .A2(n57), .B1(n18), .B2(n107), .ZN(n160) );
  OR2_X1 U93 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n58) );
  OAI22_X1 U94 ( .A1(n135), .A2(n32), .B1(n58), .B2(n136), .ZN(n63) );
  XNOR2_X1 U95 ( .A(n19), .B(\mult_x_1/n288 ), .ZN(n60) );
  XNOR2_X1 U96 ( .A(n543), .B(\mult_x_1/n283 ), .ZN(n183) );
  OAI22_X1 U97 ( .A1(n229), .A2(n183), .B1(n61), .B2(n30), .ZN(n129) );
  AND2_X1 U98 ( .A1(\mult_x_1/n288 ), .A2(n47), .ZN(n128) );
  XNOR2_X1 U99 ( .A(n20), .B(\mult_x_1/n285 ), .ZN(n182) );
  OAI22_X1 U100 ( .A1(n88), .A2(n182), .B1(n18), .B2(n62), .ZN(n127) );
  FA_X1 U101 ( .A(n66), .B(n65), .CI(n64), .CO(n167), .S(n119) );
  NAND2_X1 U102 ( .A1(n174), .A2(n173), .ZN(n67) );
  NAND2_X1 U103 ( .A1(n67), .A2(en), .ZN(n69) );
  OR2_X1 U104 ( .A1(n279), .A2(n44), .ZN(n68) );
  NAND2_X1 U105 ( .A1(n69), .A2(n68), .ZN(n363) );
  NOR2_X1 U126 ( .A1(n36), .A2(n138), .ZN(n133) );
  XNOR2_X1 U127 ( .A(n19), .B(\mult_x_1/n281 ), .ZN(n70) );
  XNOR2_X1 U128 ( .A(n87), .B(n19), .ZN(n134) );
  OAI22_X1 U129 ( .A1(n135), .A2(n70), .B1(n134), .B2(n136), .ZN(n142) );
  INV_X1 U130 ( .A(n142), .ZN(n132) );
  XNOR2_X1 U131 ( .A(n545), .B(\mult_x_1/n282 ), .ZN(n73) );
  OAI22_X1 U132 ( .A1(n135), .A2(n73), .B1(n136), .B2(n70), .ZN(n78) );
  XNOR2_X1 U133 ( .A(n87), .B(n22), .ZN(n72) );
  AOI21_X1 U134 ( .B1(n214), .B2(n126), .A(n72), .ZN(n71) );
  INV_X1 U135 ( .A(n71), .ZN(n77) );
  XNOR2_X1 U136 ( .A(n22), .B(\mult_x_1/n281 ), .ZN(n92) );
  OAI22_X1 U137 ( .A1(n126), .A2(n92), .B1(n72), .B2(n214), .ZN(n76) );
  INV_X1 U138 ( .A(n76), .ZN(n85) );
  XNOR2_X1 U139 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n86) );
  OAI22_X1 U140 ( .A1(n135), .A2(n86), .B1(n136), .B2(n73), .ZN(n83) );
  NOR2_X1 U141 ( .A1(n37), .A2(n138), .ZN(n84) );
  NOR2_X1 U142 ( .A1(n38), .A2(n138), .ZN(n81) );
  FA_X1 U143 ( .A(n78), .B(n77), .CI(n76), .CO(n131), .S(n80) );
  OR2_X1 U144 ( .A1(n149), .A2(n148), .ZN(n79) );
  MUX2_X1 U145 ( .A(n323), .B(n79), .S(n279), .Z(n343) );
  FA_X1 U146 ( .A(n82), .B(n81), .CI(n80), .CO(n148), .S(n152) );
  XNOR2_X1 U147 ( .A(n545), .B(\mult_x_1/n284 ), .ZN(n91) );
  OAI22_X1 U148 ( .A1(n135), .A2(n91), .B1(n136), .B2(n86), .ZN(n113) );
  XNOR2_X1 U149 ( .A(n87), .B(n20), .ZN(n89) );
  XNOR2_X1 U150 ( .A(n20), .B(\mult_x_1/n281 ), .ZN(n106) );
  OAI22_X1 U151 ( .A1(n226), .A2(n89), .B1(n88), .B2(n106), .ZN(n112) );
  AOI21_X1 U152 ( .B1(n18), .B2(n88), .A(n89), .ZN(n90) );
  INV_X1 U153 ( .A(n90), .ZN(n111) );
  XNOR2_X1 U154 ( .A(n545), .B(\mult_x_1/n285 ), .ZN(n102) );
  OAI22_X1 U155 ( .A1(n135), .A2(n102), .B1(n136), .B2(n91), .ZN(n196) );
  XNOR2_X1 U156 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n104) );
  XNOR2_X1 U157 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n93) );
  OAI22_X1 U158 ( .A1(n126), .A2(n104), .B1(n214), .B2(n93), .ZN(n195) );
  INV_X1 U159 ( .A(n112), .ZN(n194) );
  OAI22_X1 U160 ( .A1(n126), .A2(n93), .B1(n214), .B2(n92), .ZN(n114) );
  NAND2_X1 U161 ( .A1(n117), .A2(n114), .ZN(n96) );
  NOR2_X1 U162 ( .A1(n39), .A2(n138), .ZN(n115) );
  NAND2_X1 U163 ( .A1(n117), .A2(n115), .ZN(n95) );
  NAND2_X1 U164 ( .A1(n115), .A2(n114), .ZN(n94) );
  OR2_X1 U165 ( .A1(n152), .A2(n151), .ZN(n97) );
  MUX2_X1 U166 ( .A(n324), .B(n97), .S(n279), .Z(n345) );
  AOI21_X1 U167 ( .B1(n229), .B2(n30), .A(n100), .ZN(n101) );
  INV_X1 U168 ( .A(n101), .ZN(n164) );
  OAI22_X1 U169 ( .A1(n135), .A2(n103), .B1(n136), .B2(n102), .ZN(n163) );
  NOR2_X1 U170 ( .A1(n40), .A2(n138), .ZN(n162) );
  OAI22_X1 U171 ( .A1(n126), .A2(n105), .B1(n214), .B2(n104), .ZN(n155) );
  OAI22_X1 U172 ( .A1(n88), .A2(n107), .B1(n226), .B2(n106), .ZN(n154) );
  NOR2_X1 U173 ( .A1(n41), .A2(n138), .ZN(n197) );
  FA_X1 U174 ( .A(n113), .B(n27), .CI(n111), .CO(n98), .S(n243) );
  XOR2_X1 U175 ( .A(n115), .B(n114), .Z(n116) );
  XOR2_X1 U176 ( .A(n117), .B(n116), .Z(n242) );
  OR2_X1 U177 ( .A1(n191), .A2(n190), .ZN(n118) );
  MUX2_X1 U178 ( .A(n325), .B(n118), .S(n279), .Z(n347) );
  FA_X1 U179 ( .A(n121), .B(n120), .CI(n119), .CO(n173), .S(n177) );
  OR2_X1 U180 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n122) );
  OAI22_X1 U181 ( .A1(n126), .A2(n34), .B1(n122), .B2(n214), .ZN(n185) );
  XNOR2_X1 U182 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n123) );
  XNOR2_X1 U183 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n125) );
  OAI22_X1 U184 ( .A1(n126), .A2(n123), .B1(n214), .B2(n125), .ZN(n184) );
  OAI22_X1 U185 ( .A1(n126), .A2(n125), .B1(n214), .B2(n124), .ZN(n180) );
  FA_X1 U186 ( .A(n129), .B(n128), .CI(n127), .CO(n121), .S(n179) );
  OR2_X1 U187 ( .A1(n177), .A2(n176), .ZN(n130) );
  MUX2_X1 U188 ( .A(n326), .B(n130), .S(n322), .Z(n349) );
  FA_X1 U189 ( .A(n133), .B(n132), .CI(n131), .CO(n144), .S(n149) );
  AOI21_X1 U190 ( .B1(n136), .B2(n135), .A(n134), .ZN(n137) );
  INV_X1 U191 ( .A(n137), .ZN(n140) );
  NOR2_X1 U192 ( .A1(n33), .A2(n138), .ZN(n139) );
  XOR2_X1 U193 ( .A(n140), .B(n139), .Z(n141) );
  XOR2_X1 U194 ( .A(n142), .B(n141), .Z(n143) );
  OR2_X1 U195 ( .A1(n144), .A2(n143), .ZN(n146) );
  NAND2_X1 U196 ( .A1(n144), .A2(n143), .ZN(n145) );
  NAND2_X1 U197 ( .A1(n146), .A2(n145), .ZN(n147) );
  MUX2_X1 U198 ( .A(n327), .B(n147), .S(n322), .Z(n351) );
  NAND2_X1 U199 ( .A1(n149), .A2(n148), .ZN(n150) );
  MUX2_X1 U200 ( .A(n328), .B(n150), .S(n279), .Z(n353) );
  NAND2_X1 U201 ( .A1(n152), .A2(n151), .ZN(n153) );
  MUX2_X1 U202 ( .A(n329), .B(n153), .S(n322), .Z(n355) );
  XNOR2_X1 U203 ( .A(n155), .B(n154), .ZN(n193) );
  FA_X1 U204 ( .A(n158), .B(n157), .CI(n156), .CO(n192), .S(n168) );
  FA_X1 U205 ( .A(n161), .B(n160), .CI(n159), .CO(n203), .S(n166) );
  FA_X1 U206 ( .A(n164), .B(n163), .CI(n162), .CO(n200), .S(n202) );
  FA_X1 U207 ( .A(n168), .B(n167), .CI(n166), .CO(n170), .S(n174) );
  NOR2_X1 U208 ( .A1(n171), .A2(n170), .ZN(n169) );
  MUX2_X1 U209 ( .A(n330), .B(n169), .S(en), .Z(n357) );
  NAND2_X1 U210 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U211 ( .A(n331), .B(n172), .S(n279), .Z(n359) );
  NOR2_X1 U212 ( .A1(n174), .A2(n173), .ZN(n175) );
  NAND2_X1 U213 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2_X1 U214 ( .A(n334), .B(n178), .S(en), .Z(n365) );
  FA_X1 U215 ( .A(n181), .B(n180), .CI(n179), .CO(n176), .S(n188) );
  XNOR2_X1 U216 ( .A(n20), .B(\mult_x_1/n286 ), .ZN(n215) );
  OAI22_X1 U217 ( .A1(n88), .A2(n215), .B1(n18), .B2(n182), .ZN(n212) );
  XNOR2_X1 U218 ( .A(n543), .B(\mult_x_1/n284 ), .ZN(n213) );
  OAI22_X1 U219 ( .A1(n229), .A2(n213), .B1(n183), .B2(n30), .ZN(n211) );
  HA_X1 U220 ( .A(n185), .B(n184), .CO(n181), .S(n210) );
  NOR2_X1 U221 ( .A1(n188), .A2(n187), .ZN(n186) );
  MUX2_X1 U222 ( .A(n335), .B(n186), .S(n322), .Z(n367) );
  NAND2_X1 U223 ( .A1(n188), .A2(n187), .ZN(n189) );
  MUX2_X1 U224 ( .A(n336), .B(n189), .S(n322), .Z(n369) );
  XNOR2_X1 U225 ( .A(n198), .B(n197), .ZN(n199) );
  XNOR2_X1 U226 ( .A(n200), .B(n199), .ZN(n246) );
  NOR2_X1 U227 ( .A1(n208), .A2(n207), .ZN(n206) );
  MUX2_X1 U228 ( .A(n338), .B(n206), .S(n322), .Z(n373) );
  NAND2_X1 U229 ( .A1(n208), .A2(n207), .ZN(n209) );
  MUX2_X1 U230 ( .A(n339), .B(n209), .S(n322), .Z(n375) );
  FA_X1 U231 ( .A(n212), .B(n211), .CI(n210), .CO(n187), .S(n239) );
  XNOR2_X1 U232 ( .A(n543), .B(\mult_x_1/n285 ), .ZN(n221) );
  OAI22_X1 U233 ( .A1(n229), .A2(n221), .B1(n213), .B2(n30), .ZN(n218) );
  AND2_X1 U234 ( .A1(\mult_x_1/n288 ), .A2(n51), .ZN(n217) );
  XNOR2_X1 U235 ( .A(n20), .B(\mult_x_1/n287 ), .ZN(n219) );
  OAI22_X1 U236 ( .A1(n88), .A2(n219), .B1(n18), .B2(n215), .ZN(n216) );
  OR2_X1 U237 ( .A1(n239), .A2(n238), .ZN(n272) );
  FA_X1 U238 ( .A(n218), .B(n217), .CI(n216), .CO(n238), .S(n237) );
  XNOR2_X1 U239 ( .A(n20), .B(\mult_x_1/n288 ), .ZN(n220) );
  OAI22_X1 U240 ( .A1(n88), .A2(n220), .B1(n226), .B2(n219), .ZN(n223) );
  XNOR2_X1 U241 ( .A(n543), .B(\mult_x_1/n286 ), .ZN(n225) );
  OAI22_X1 U242 ( .A1(n229), .A2(n225), .B1(n221), .B2(n30), .ZN(n222) );
  NOR2_X1 U243 ( .A1(n237), .A2(n236), .ZN(n265) );
  HA_X1 U244 ( .A(n223), .B(n222), .CO(n236), .S(n234) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n224) );
  OAI22_X1 U246 ( .A1(n88), .A2(n35), .B1(n224), .B2(n18), .ZN(n233) );
  OR2_X1 U247 ( .A1(n234), .A2(n233), .ZN(n261) );
  XNOR2_X1 U248 ( .A(n543), .B(\mult_x_1/n287 ), .ZN(n228) );
  OAI22_X1 U249 ( .A1(n229), .A2(n228), .B1(n225), .B2(n30), .ZN(n232) );
  INV_X1 U250 ( .A(n18), .ZN(n227) );
  AND2_X1 U251 ( .A1(\mult_x_1/n288 ), .A2(n227), .ZN(n231) );
  NOR2_X1 U252 ( .A1(n232), .A2(n231), .ZN(n254) );
  OAI22_X1 U253 ( .A1(n229), .A2(\mult_x_1/n288 ), .B1(n228), .B2(n30), .ZN(
        n251) );
  OR2_X1 U254 ( .A1(\mult_x_1/n288 ), .A2(n43), .ZN(n230) );
  NAND2_X1 U255 ( .A1(n230), .A2(n229), .ZN(n250) );
  NAND2_X1 U256 ( .A1(n251), .A2(n250), .ZN(n257) );
  NAND2_X1 U257 ( .A1(n232), .A2(n231), .ZN(n255) );
  OAI21_X1 U258 ( .B1(n254), .B2(n257), .A(n255), .ZN(n262) );
  NAND2_X1 U259 ( .A1(n234), .A2(n233), .ZN(n260) );
  INV_X1 U260 ( .A(n260), .ZN(n235) );
  AOI21_X1 U261 ( .B1(n261), .B2(n262), .A(n235), .ZN(n268) );
  NAND2_X1 U262 ( .A1(n237), .A2(n236), .ZN(n266) );
  OAI21_X1 U263 ( .B1(n265), .B2(n268), .A(n266), .ZN(n273) );
  NAND2_X1 U264 ( .A1(n239), .A2(n238), .ZN(n271) );
  INV_X1 U265 ( .A(n271), .ZN(n240) );
  AOI21_X1 U266 ( .B1(n272), .B2(n273), .A(n240), .ZN(n241) );
  MUX2_X1 U267 ( .A(n340), .B(n241), .S(n322), .Z(n377) );
  FA_X1 U268 ( .A(n244), .B(n243), .CI(n242), .CO(n190), .S(n245) );
  MUX2_X1 U269 ( .A(n341), .B(n245), .S(n322), .Z(n379) );
  FA_X1 U270 ( .A(n42), .B(n247), .CI(n246), .CO(n248), .S(n208) );
  MUX2_X1 U271 ( .A(n342), .B(n248), .S(n322), .Z(n381) );
  MUX2_X1 U272 ( .A(product[0]), .B(n506), .S(n279), .Z(n396) );
  MUX2_X1 U273 ( .A(n506), .B(n507), .S(n279), .Z(n398) );
  AND2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n249) );
  MUX2_X1 U275 ( .A(n507), .B(n249), .S(n279), .Z(n400) );
  MUX2_X1 U276 ( .A(product[1]), .B(n509), .S(n279), .Z(n402) );
  MUX2_X1 U277 ( .A(n509), .B(n510), .S(n279), .Z(n404) );
  OR2_X1 U278 ( .A1(n251), .A2(n250), .ZN(n252) );
  AND2_X1 U279 ( .A1(n252), .A2(n257), .ZN(n253) );
  MUX2_X1 U280 ( .A(n510), .B(n253), .S(n279), .Z(n406) );
  MUX2_X1 U281 ( .A(product[2]), .B(n512), .S(n279), .Z(n408) );
  MUX2_X1 U282 ( .A(n512), .B(n513), .S(n279), .Z(n410) );
  INV_X1 U283 ( .A(n254), .ZN(n256) );
  NAND2_X1 U284 ( .A1(n256), .A2(n255), .ZN(n258) );
  XOR2_X1 U285 ( .A(n258), .B(n257), .Z(n259) );
  MUX2_X1 U286 ( .A(n513), .B(n259), .S(n279), .Z(n412) );
  MUX2_X1 U287 ( .A(product[3]), .B(n515), .S(n279), .Z(n414) );
  MUX2_X1 U288 ( .A(n515), .B(n516), .S(n279), .Z(n416) );
  NAND2_X1 U289 ( .A1(n261), .A2(n260), .ZN(n263) );
  XNOR2_X1 U290 ( .A(n263), .B(n262), .ZN(n264) );
  MUX2_X1 U291 ( .A(n516), .B(n264), .S(n279), .Z(n418) );
  MUX2_X1 U292 ( .A(product[4]), .B(n518), .S(n279), .Z(n420) );
  MUX2_X1 U293 ( .A(n518), .B(n519), .S(n279), .Z(n422) );
  INV_X1 U294 ( .A(n265), .ZN(n267) );
  NAND2_X1 U295 ( .A1(n267), .A2(n266), .ZN(n269) );
  XOR2_X1 U296 ( .A(n269), .B(n268), .Z(n270) );
  MUX2_X1 U297 ( .A(n519), .B(n270), .S(n279), .Z(n424) );
  MUX2_X1 U298 ( .A(product[5]), .B(n521), .S(n279), .Z(n426) );
  MUX2_X1 U299 ( .A(n521), .B(n522), .S(n279), .Z(n428) );
  NAND2_X1 U300 ( .A1(n272), .A2(n271), .ZN(n274) );
  XNOR2_X1 U301 ( .A(n274), .B(n273), .ZN(n275) );
  MUX2_X1 U302 ( .A(n522), .B(n275), .S(n279), .Z(n430) );
  MUX2_X1 U303 ( .A(product[6]), .B(n524), .S(n279), .Z(n432) );
  NAND2_X1 U304 ( .A1(n385), .A2(n336), .ZN(n276) );
  XOR2_X1 U305 ( .A(n276), .B(n340), .Z(n277) );
  MUX2_X1 U306 ( .A(n524), .B(n277), .S(n279), .Z(n434) );
  MUX2_X1 U307 ( .A(product[7]), .B(n526), .S(n279), .Z(n436) );
  OAI21_X1 U308 ( .B1(n335), .B2(n340), .A(n336), .ZN(n281) );
  NAND2_X1 U309 ( .A1(n326), .A2(n334), .ZN(n278) );
  XNOR2_X1 U310 ( .A(n281), .B(n278), .ZN(n280) );
  MUX2_X1 U311 ( .A(n526), .B(n280), .S(n279), .Z(n438) );
  MUX2_X1 U312 ( .A(product[8]), .B(n528), .S(n322), .Z(n440) );
  AOI21_X1 U313 ( .B1(n281), .B2(n326), .A(n386), .ZN(n284) );
  NAND2_X1 U314 ( .A1(n387), .A2(n333), .ZN(n282) );
  XOR2_X1 U315 ( .A(n284), .B(n282), .Z(n283) );
  MUX2_X1 U316 ( .A(n528), .B(n283), .S(n322), .Z(n442) );
  MUX2_X1 U317 ( .A(product[9]), .B(n530), .S(n322), .Z(n444) );
  OAI21_X1 U318 ( .B1(n284), .B2(n332), .A(n333), .ZN(n292) );
  INV_X1 U319 ( .A(n292), .ZN(n287) );
  NAND2_X1 U320 ( .A1(n388), .A2(n331), .ZN(n285) );
  XOR2_X1 U321 ( .A(n287), .B(n285), .Z(n286) );
  MUX2_X1 U322 ( .A(n530), .B(n286), .S(n322), .Z(n446) );
  MUX2_X1 U323 ( .A(product[10]), .B(n532), .S(n322), .Z(n448) );
  OAI21_X1 U324 ( .B1(n287), .B2(n330), .A(n331), .ZN(n289) );
  NAND2_X1 U325 ( .A1(n389), .A2(n339), .ZN(n288) );
  XNOR2_X1 U326 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U327 ( .A(n532), .B(n290), .S(n322), .Z(n450) );
  MUX2_X1 U328 ( .A(product[11]), .B(n534), .S(n322), .Z(n452) );
  NOR2_X1 U329 ( .A1(n338), .A2(n330), .ZN(n293) );
  OAI21_X1 U330 ( .B1(n338), .B2(n331), .A(n339), .ZN(n291) );
  AOI21_X1 U331 ( .B1(n293), .B2(n292), .A(n291), .ZN(n319) );
  NOR2_X1 U332 ( .A1(n341), .A2(n342), .ZN(n306) );
  INV_X1 U333 ( .A(n306), .ZN(n299) );
  NAND2_X1 U334 ( .A1(n341), .A2(n342), .ZN(n308) );
  NAND2_X1 U335 ( .A1(n299), .A2(n308), .ZN(n294) );
  XOR2_X1 U336 ( .A(n319), .B(n294), .Z(n295) );
  MUX2_X1 U337 ( .A(n534), .B(n295), .S(n322), .Z(n454) );
  MUX2_X1 U338 ( .A(product[12]), .B(n536), .S(n322), .Z(n456) );
  OAI21_X1 U339 ( .B1(n319), .B2(n306), .A(n308), .ZN(n297) );
  NAND2_X1 U340 ( .A1(n325), .A2(n337), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  MUX2_X1 U342 ( .A(n536), .B(n298), .S(n322), .Z(n458) );
  MUX2_X1 U343 ( .A(product[13]), .B(n538), .S(n322), .Z(n460) );
  NAND2_X1 U344 ( .A1(n299), .A2(n325), .ZN(n302) );
  INV_X1 U345 ( .A(n308), .ZN(n300) );
  AOI21_X1 U346 ( .B1(n300), .B2(n325), .A(n390), .ZN(n301) );
  OAI21_X1 U347 ( .B1(n319), .B2(n302), .A(n301), .ZN(n304) );
  NAND2_X1 U348 ( .A1(n324), .A2(n329), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  MUX2_X1 U350 ( .A(n538), .B(n305), .S(n322), .Z(n462) );
  MUX2_X1 U351 ( .A(product[14]), .B(n540), .S(n322), .Z(n464) );
  NAND2_X1 U352 ( .A1(n325), .A2(n324), .ZN(n309) );
  NOR2_X1 U353 ( .A1(n306), .A2(n309), .ZN(n315) );
  INV_X1 U354 ( .A(n315), .ZN(n311) );
  AOI21_X1 U355 ( .B1(n390), .B2(n324), .A(n383), .ZN(n307) );
  OAI21_X1 U356 ( .B1(n309), .B2(n308), .A(n307), .ZN(n316) );
  INV_X1 U357 ( .A(n316), .ZN(n310) );
  OAI21_X1 U358 ( .B1(n319), .B2(n311), .A(n310), .ZN(n313) );
  NAND2_X1 U359 ( .A1(n323), .A2(n328), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  MUX2_X1 U361 ( .A(n540), .B(n314), .S(n322), .Z(n466) );
  MUX2_X1 U362 ( .A(product[15]), .B(n542), .S(n322), .Z(n468) );
  NAND2_X1 U363 ( .A1(n315), .A2(n323), .ZN(n318) );
  AOI21_X1 U364 ( .B1(n316), .B2(n323), .A(n384), .ZN(n317) );
  OAI21_X1 U365 ( .B1(n319), .B2(n318), .A(n317), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n320), .B(n327), .ZN(n321) );
  MUX2_X1 U367 ( .A(n542), .B(n321), .S(n322), .Z(n470) );
  MUX2_X1 U368 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n322), .Z(n472) );
  MUX2_X1 U369 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n322), .Z(n474) );
  MUX2_X1 U370 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n322), .Z(n476) );
  MUX2_X1 U371 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n322), .Z(n478) );
  MUX2_X1 U372 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n322), .Z(n480) );
  MUX2_X1 U373 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n322), .Z(n482) );
  MUX2_X1 U374 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n322), .Z(n484) );
  MUX2_X1 U375 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n322), .Z(n486) );
  MUX2_X1 U376 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n322), .Z(n488) );
  MUX2_X1 U377 ( .A(n543), .B(A_extended[1]), .S(n322), .Z(n490) );
  MUX2_X1 U378 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n322), .Z(n492) );
  MUX2_X1 U379 ( .A(n20), .B(A_extended[3]), .S(n322), .Z(n494) );
  MUX2_X1 U380 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n322), .Z(n496) );
  MUX2_X1 U381 ( .A(n22), .B(A_extended[5]), .S(n322), .Z(n498) );
  MUX2_X1 U382 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n322), .Z(n500) );
  MUX2_X1 U383 ( .A(n19), .B(A_extended[7]), .S(n322), .Z(n502) );
  OR2_X1 U384 ( .A1(n322), .A2(n546), .ZN(n504) );
endmodule


module conv_128_32_DW_mult_pipe_J1_5 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n349, n351, n353,
         n355, n357, n359, n361, n363, n365, n367, n369, n371, n373, n375,
         n377, n379, n381, n383, n385, n387, n389, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n404, n406, n408,
         n410, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n442, n444, n446, n448, n450, n452,
         n454, n456, n458, n460, n462, n464, n466, n468, n470, n472, n474,
         n476, n478, n480, n482, n484, n486, n488, n490, n492, n494, n496,
         n498, n500, n502, n504, n506, n508, n510, n512, n513, n515, n516,
         n518, n519, n521, n522, n524, n525, n527, n529, n531, n533, n535,
         n537, n539, n541, n543, n545, n547, n548, n549, n550, n551;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n402), .SE(n510), .CK(clk), .Q(n550), 
        .QN(n36) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n402), .SE(n506), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n402), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n324) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n402), .SE(n498), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n35) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n402), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n23) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n402), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n27) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n402), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n29) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n400), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n31) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n401), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n400), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n32) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n402), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n28) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n400), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n33) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n400), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n25) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n400), .SE(n476), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n400), .SE(n474), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n400), .SE(n472), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n400), .SE(n470), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n400), .SE(n468), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n401), .SE(n466), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n402), .SE(n464), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n400), .SE(n462), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n400), .SE(n460), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n400), .SE(n458), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n400), .SE(n456), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n400), .SE(n454), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n400), .SE(n452), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n400), .SE(n450), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n400), .SE(n448), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n401), .SE(n446), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n401), .SE(n444), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n401), .SE(n442), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n401), .SE(n440), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n401), .SE(n438), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n401), .SE(n436), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n401), .SE(n434), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n401), .SE(n432), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n401), .SE(n430), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n401), .SE(n428), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n401), .SE(n426), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n400), .SE(n424), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n400), .SE(n422), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n400), .SE(n420), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n400), .SE(n418), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n400), .SE(n416), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n400), .SE(n414), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n400), .SE(n412), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n400), .SE(n410), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n400), .SE(n408), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n400), .SE(n406), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n400), .SE(n404), .CK(clk), .Q(
        product[0]) );
  SDFF_X2 clk_r_REG51_S1 ( .D(1'b0), .SI(n402), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n323) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n551), .SE(n389), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2_IP  ( .D(1'b1), .SI(n551), .SE(n387), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n551), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n551), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n551), .SE(n381), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n551), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n551), .SE(n377), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n551), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n339), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n551), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n338), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n551), .SE(n371), .CK(
        clk), .Q(n398), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n551), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n336), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n551), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n551), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n334), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n551), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n333), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n551), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n551), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n331), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n551), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n330), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n551), .SE(n355), .CK(
        clk), .QN(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n551), .SE(n353), .CK(
        clk), .QN(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n551), .SI(1'b1), .SE(n351), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n551), .SI(1'b1), .SE(n349), .CK(clk), 
        .Q(n326), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n551), .SE(n347), .CK(
        clk), .QN(n325) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n402), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n24) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n402), .SE(n496), .CK(clk), .Q(n548), 
        .QN(n37) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n402), .SE(n504), .CK(clk), .Q(n549), 
        .QN(n34) );
  BUF_X1 U2 ( .A(en), .Z(n19) );
  BUF_X1 U3 ( .A(en), .Z(n18) );
  INV_X2 U4 ( .A(n41), .ZN(n133) );
  BUF_X1 U5 ( .A(n400), .Z(n401) );
  INV_X2 U6 ( .A(n551), .ZN(n400) );
  INV_X1 U7 ( .A(n87), .ZN(n17) );
  XNOR2_X1 U8 ( .A(n14), .B(n12), .ZN(n200) );
  XNOR2_X1 U9 ( .A(n90), .B(n89), .ZN(n14) );
  BUF_X1 U10 ( .A(n400), .Z(n402) );
  NAND2_X1 U11 ( .A1(n9), .A2(n8), .ZN(n128) );
  NAND2_X1 U12 ( .A1(n85), .A2(n86), .ZN(n8) );
  OAI21_X1 U13 ( .B1(n85), .B2(n86), .A(n21), .ZN(n9) );
  OR2_X1 U14 ( .A1(n71), .A2(n70), .ZN(n188) );
  INV_X1 U15 ( .A(rst_n), .ZN(n551) );
  NAND2_X1 U16 ( .A1(n7), .A2(n5), .ZN(n353) );
  NAND2_X1 U17 ( .A1(n6), .A2(n328), .ZN(n5) );
  INV_X1 U18 ( .A(n18), .ZN(n6) );
  OAI21_X1 U19 ( .B1(n166), .B2(n165), .A(n18), .ZN(n7) );
  NAND2_X1 U20 ( .A1(n11), .A2(n10), .ZN(n145) );
  NAND2_X1 U21 ( .A1(n90), .A2(n89), .ZN(n10) );
  OAI21_X1 U22 ( .B1(n90), .B2(n89), .A(n12), .ZN(n11) );
  XNOR2_X1 U23 ( .A(n13), .B(n21), .ZN(n12) );
  XNOR2_X1 U24 ( .A(n85), .B(n86), .ZN(n13) );
  NAND2_X2 U25 ( .A1(n46), .A2(n47), .ZN(n214) );
  NAND2_X1 U26 ( .A1(n16), .A2(n15), .ZN(n85) );
  INV_X1 U27 ( .A(n82), .ZN(n15) );
  NAND2_X1 U28 ( .A1(n122), .A2(n124), .ZN(n16) );
  XNOR2_X1 U29 ( .A(n35), .B(n37), .ZN(n47) );
  OR2_X1 U30 ( .A1(n242), .A2(n241), .ZN(n239) );
  XNOR2_X1 U31 ( .A(n323), .B(n324), .ZN(n44) );
  NAND2_X1 U32 ( .A1(n195), .A2(n194), .ZN(n96) );
  NOR2_X1 U33 ( .A1(n195), .A2(n194), .ZN(n97) );
  NAND2_X1 U34 ( .A1(n186), .A2(n185), .ZN(n190) );
  OR2_X1 U35 ( .A1(n188), .A2(n187), .ZN(n185) );
  NAND2_X1 U36 ( .A1(n188), .A2(n187), .ZN(n189) );
  XNOR2_X1 U37 ( .A(\mult_x_1/n312 ), .B(n35), .ZN(n46) );
  XNOR2_X1 U38 ( .A(n42), .B(n67), .ZN(n237) );
  XNOR2_X1 U39 ( .A(n65), .B(n66), .ZN(n42) );
  NAND2_X1 U40 ( .A1(n244), .A2(n243), .ZN(n245) );
  NAND2_X1 U41 ( .A1(n242), .A2(n241), .ZN(n243) );
  NAND2_X1 U42 ( .A1(n240), .A2(n239), .ZN(n244) );
  NAND2_X1 U43 ( .A1(n190), .A2(n189), .ZN(n230) );
  INV_X1 U44 ( .A(n24), .ZN(n20) );
  OAI22_X1 U45 ( .A1(n124), .A2(n94), .B1(n82), .B2(n122), .ZN(n21) );
  INV_X1 U46 ( .A(n34), .ZN(n22) );
  INV_X2 U47 ( .A(n48), .ZN(n216) );
  MUX2_X1 U48 ( .A(n343), .B(n73), .S(n18), .Z(n383) );
  OAI21_X1 U49 ( .B1(n98), .B2(n97), .A(n96), .ZN(n183) );
  INV_X1 U50 ( .A(n197), .ZN(n98) );
  BUF_X4 U51 ( .A(en), .Z(n322) );
  NAND2_X2 U52 ( .A1(n44), .A2(n43), .ZN(n124) );
  AND2_X1 U53 ( .A1(n61), .A2(n60), .ZN(n26) );
  NAND2_X1 U54 ( .A1(n36), .A2(n20), .ZN(n135) );
  NOR2_X1 U55 ( .A1(n135), .A2(n33), .ZN(n65) );
  NAND2_X1 U56 ( .A1(n548), .A2(n23), .ZN(n218) );
  AND2_X1 U57 ( .A1(n550), .A2(\mult_x_1/n281 ), .ZN(n81) );
  XNOR2_X1 U58 ( .A(n81), .B(n548), .ZN(n53) );
  AOI21_X1 U59 ( .B1(n218), .B2(n23), .A(n53), .ZN(n38) );
  INV_X1 U60 ( .A(n38), .ZN(n66) );
  XOR2_X1 U61 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n39) );
  XNOR2_X1 U62 ( .A(\mult_x_1/a[6] ), .B(n549), .ZN(n40) );
  NAND2_X1 U63 ( .A1(n39), .A2(n40), .ZN(n132) );
  XNOR2_X1 U64 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n51) );
  INV_X1 U65 ( .A(n40), .ZN(n41) );
  XNOR2_X1 U66 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n62) );
  OAI22_X1 U67 ( .A1(n132), .A2(n51), .B1(n133), .B2(n62), .ZN(n67) );
  XOR2_X1 U68 ( .A(\mult_x_1/a[4] ), .B(n549), .Z(n43) );
  XNOR2_X1 U69 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n114) );
  INV_X1 U70 ( .A(n44), .ZN(n45) );
  INV_X2 U71 ( .A(n45), .ZN(n122) );
  XNOR2_X1 U72 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n54) );
  OAI22_X1 U73 ( .A1(n124), .A2(n114), .B1(n122), .B2(n54), .ZN(n150) );
  XNOR2_X1 U74 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n117) );
  INV_X1 U75 ( .A(n47), .ZN(n48) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n55) );
  OAI22_X1 U77 ( .A1(n214), .A2(n117), .B1(n216), .B2(n55), .ZN(n149) );
  OR2_X1 U78 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n49) );
  OAI22_X1 U79 ( .A1(n132), .A2(n24), .B1(n49), .B2(n133), .ZN(n113) );
  XNOR2_X1 U80 ( .A(n20), .B(\mult_x_1/n288 ), .ZN(n50) );
  XNOR2_X1 U81 ( .A(n20), .B(\mult_x_1/n287 ), .ZN(n52) );
  OAI22_X1 U82 ( .A1(n132), .A2(n50), .B1(n133), .B2(n52), .ZN(n112) );
  OAI22_X1 U83 ( .A1(n132), .A2(n52), .B1(n133), .B2(n51), .ZN(n153) );
  XNOR2_X1 U84 ( .A(n548), .B(\mult_x_1/n281 ), .ZN(n115) );
  OAI22_X1 U85 ( .A1(n218), .A2(n115), .B1(n53), .B2(n23), .ZN(n152) );
  NOR2_X1 U86 ( .A1(n135), .A2(n25), .ZN(n151) );
  XNOR2_X1 U87 ( .A(n549), .B(\mult_x_1/n283 ), .ZN(n63) );
  OAI22_X1 U88 ( .A1(n124), .A2(n54), .B1(n122), .B2(n63), .ZN(n71) );
  XNOR2_X1 U89 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n64) );
  OAI22_X1 U90 ( .A1(n214), .A2(n55), .B1(n216), .B2(n64), .ZN(n70) );
  XNOR2_X1 U91 ( .A(n71), .B(n70), .ZN(n60) );
  INV_X1 U92 ( .A(n60), .ZN(n56) );
  XNOR2_X1 U93 ( .A(n61), .B(n56), .ZN(n235) );
  INV_X1 U94 ( .A(en), .ZN(n87) );
  NAND2_X1 U95 ( .A1(n57), .A2(en), .ZN(n59) );
  NAND2_X1 U96 ( .A1(n87), .A2(n345), .ZN(n58) );
  NAND2_X1 U97 ( .A1(n59), .A2(n58), .ZN(n387) );
  XNOR2_X1 U98 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n103) );
  OAI22_X1 U99 ( .A1(n132), .A2(n62), .B1(n133), .B2(n103), .ZN(n93) );
  XNOR2_X1 U100 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n95) );
  OAI22_X1 U101 ( .A1(n124), .A2(n63), .B1(n122), .B2(n95), .ZN(n92) );
  XNOR2_X1 U102 ( .A(n81), .B(\mult_x_1/n312 ), .ZN(n104) );
  OAI22_X1 U103 ( .A1(n214), .A2(n64), .B1(n104), .B2(n216), .ZN(n192) );
  INV_X1 U104 ( .A(n192), .ZN(n91) );
  OAI21_X1 U105 ( .B1(n67), .B2(n66), .A(n65), .ZN(n69) );
  NAND2_X1 U106 ( .A1(n67), .A2(n66), .ZN(n68) );
  NAND2_X1 U107 ( .A1(n69), .A2(n68), .ZN(n186) );
  NOR2_X1 U108 ( .A1(n28), .A2(n135), .ZN(n187) );
  XNOR2_X1 U109 ( .A(n188), .B(n187), .ZN(n72) );
  XNOR2_X1 U110 ( .A(n186), .B(n72), .ZN(n232) );
  XNOR2_X1 U133 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n77) );
  XNOR2_X1 U134 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n111) );
  OAI22_X1 U135 ( .A1(n214), .A2(n77), .B1(n216), .B2(n111), .ZN(n173) );
  XNOR2_X1 U136 ( .A(n548), .B(\mult_x_1/n284 ), .ZN(n76) );
  XNOR2_X1 U137 ( .A(n548), .B(\mult_x_1/n283 ), .ZN(n110) );
  OAI22_X1 U138 ( .A1(n218), .A2(n76), .B1(n110), .B2(n23), .ZN(n172) );
  OR2_X1 U139 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n74) );
  OAI22_X1 U140 ( .A1(n124), .A2(n34), .B1(n74), .B2(n122), .ZN(n120) );
  XNOR2_X1 U141 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n75) );
  XNOR2_X1 U142 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n123) );
  OAI22_X1 U143 ( .A1(n124), .A2(n75), .B1(n122), .B2(n123), .ZN(n119) );
  XNOR2_X1 U144 ( .A(n548), .B(\mult_x_1/n285 ), .ZN(n210) );
  OAI22_X1 U145 ( .A1(n218), .A2(n210), .B1(n76), .B2(n23), .ZN(n207) );
  AND2_X1 U146 ( .A1(\mult_x_1/n288 ), .A2(n45), .ZN(n206) );
  XNOR2_X1 U147 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n208) );
  OAI22_X1 U148 ( .A1(n214), .A2(n208), .B1(n216), .B2(n77), .ZN(n205) );
  NOR2_X1 U149 ( .A1(n179), .A2(n178), .ZN(n79) );
  NAND2_X1 U150 ( .A1(n87), .A2(n325), .ZN(n78) );
  OAI21_X1 U151 ( .B1(n87), .B2(n79), .A(n78), .ZN(n347) );
  NOR2_X1 U152 ( .A1(n29), .A2(n135), .ZN(n130) );
  XNOR2_X1 U153 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n80) );
  XNOR2_X1 U154 ( .A(n81), .B(n20), .ZN(n131) );
  OAI22_X1 U155 ( .A1(n132), .A2(n80), .B1(n131), .B2(n133), .ZN(n139) );
  INV_X1 U156 ( .A(n139), .ZN(n129) );
  XNOR2_X1 U157 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n83) );
  OAI22_X1 U158 ( .A1(n132), .A2(n83), .B1(n133), .B2(n80), .ZN(n86) );
  XNOR2_X1 U159 ( .A(n81), .B(n549), .ZN(n82) );
  XNOR2_X1 U160 ( .A(n549), .B(\mult_x_1/n281 ), .ZN(n94) );
  OAI22_X1 U161 ( .A1(n124), .A2(n94), .B1(n82), .B2(n122), .ZN(n84) );
  NOR2_X1 U162 ( .A1(n30), .A2(n135), .ZN(n101) );
  XNOR2_X1 U163 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n102) );
  OAI22_X1 U164 ( .A1(n132), .A2(n102), .B1(n133), .B2(n83), .ZN(n100) );
  INV_X1 U165 ( .A(n84), .ZN(n99) );
  NOR2_X1 U166 ( .A1(n31), .A2(n135), .ZN(n89) );
  OR2_X1 U167 ( .A1(n146), .A2(n145), .ZN(n88) );
  MUX2_X1 U168 ( .A(n326), .B(n88), .S(n18), .Z(n349) );
  FA_X1 U169 ( .A(n93), .B(n92), .CI(n91), .CO(n197), .S(n233) );
  NOR2_X1 U170 ( .A1(n32), .A2(n135), .ZN(n195) );
  OAI22_X1 U171 ( .A1(n124), .A2(n95), .B1(n122), .B2(n94), .ZN(n194) );
  FA_X1 U172 ( .A(n101), .B(n100), .CI(n99), .CO(n90), .S(n182) );
  NAND2_X1 U173 ( .A1(n183), .A2(n182), .ZN(n108) );
  OAI22_X1 U174 ( .A1(n132), .A2(n103), .B1(n133), .B2(n102), .ZN(n193) );
  AOI21_X1 U175 ( .B1(n216), .B2(n214), .A(n104), .ZN(n105) );
  INV_X1 U176 ( .A(n105), .ZN(n191) );
  NAND2_X1 U177 ( .A1(n183), .A2(n181), .ZN(n107) );
  NAND2_X1 U178 ( .A1(n182), .A2(n181), .ZN(n106) );
  NAND3_X1 U179 ( .A1(n108), .A2(n107), .A3(n106), .ZN(n199) );
  OR2_X1 U180 ( .A1(n200), .A2(n199), .ZN(n109) );
  MUX2_X1 U181 ( .A(n327), .B(n109), .S(n18), .Z(n351) );
  XNOR2_X1 U182 ( .A(n548), .B(\mult_x_1/n282 ), .ZN(n116) );
  OAI22_X1 U183 ( .A1(n218), .A2(n110), .B1(n116), .B2(n23), .ZN(n127) );
  AND2_X1 U184 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n126) );
  XNOR2_X1 U185 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n118) );
  OAI22_X1 U186 ( .A1(n214), .A2(n111), .B1(n216), .B2(n118), .ZN(n125) );
  HA_X1 U187 ( .A(n113), .B(n112), .CO(n148), .S(n159) );
  XNOR2_X1 U188 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n121) );
  OAI22_X1 U189 ( .A1(n124), .A2(n121), .B1(n122), .B2(n114), .ZN(n156) );
  OAI22_X1 U190 ( .A1(n218), .A2(n116), .B1(n115), .B2(n23), .ZN(n155) );
  OAI22_X1 U191 ( .A1(n214), .A2(n118), .B1(n216), .B2(n117), .ZN(n154) );
  HA_X1 U192 ( .A(n120), .B(n119), .CO(n170), .S(n171) );
  OAI22_X1 U193 ( .A1(n124), .A2(n123), .B1(n122), .B2(n121), .ZN(n169) );
  FA_X1 U194 ( .A(n127), .B(n126), .CI(n125), .CO(n160), .S(n168) );
  FA_X1 U195 ( .A(n130), .B(n129), .CI(n128), .CO(n141), .S(n146) );
  AOI21_X1 U196 ( .B1(n133), .B2(n132), .A(n131), .ZN(n134) );
  INV_X1 U197 ( .A(n134), .ZN(n137) );
  NOR2_X1 U198 ( .A1(n27), .A2(n135), .ZN(n136) );
  XOR2_X1 U199 ( .A(n137), .B(n136), .Z(n138) );
  XOR2_X1 U200 ( .A(n139), .B(n138), .Z(n140) );
  OR2_X1 U201 ( .A1(n141), .A2(n140), .ZN(n143) );
  NAND2_X1 U202 ( .A1(n141), .A2(n140), .ZN(n142) );
  NAND2_X1 U203 ( .A1(n143), .A2(n142), .ZN(n144) );
  MUX2_X1 U204 ( .A(n329), .B(n144), .S(n18), .Z(n355) );
  NAND2_X1 U205 ( .A1(n146), .A2(n145), .ZN(n147) );
  MUX2_X1 U206 ( .A(n330), .B(n147), .S(n18), .Z(n357) );
  FA_X1 U207 ( .A(n150), .B(n149), .CI(n148), .CO(n236), .S(n240) );
  FA_X1 U208 ( .A(n151), .B(n152), .CI(n153), .CO(n61), .S(n242) );
  FA_X1 U209 ( .A(n156), .B(n155), .CI(n154), .CO(n241), .S(n158) );
  XNOR2_X1 U210 ( .A(n242), .B(n241), .ZN(n157) );
  XNOR2_X1 U211 ( .A(n240), .B(n157), .ZN(n163) );
  FA_X1 U212 ( .A(n160), .B(n159), .CI(n158), .CO(n162), .S(n166) );
  NOR2_X1 U213 ( .A1(n163), .A2(n162), .ZN(n161) );
  MUX2_X1 U214 ( .A(n331), .B(n161), .S(n18), .Z(n359) );
  NAND2_X1 U215 ( .A1(n163), .A2(n162), .ZN(n164) );
  MUX2_X1 U216 ( .A(n332), .B(n164), .S(n18), .Z(n361) );
  NAND2_X1 U217 ( .A1(n166), .A2(n165), .ZN(n167) );
  MUX2_X1 U218 ( .A(n333), .B(n167), .S(n18), .Z(n363) );
  FA_X1 U219 ( .A(n170), .B(n169), .CI(n168), .CO(n165), .S(n176) );
  FA_X1 U220 ( .A(n173), .B(n172), .CI(n171), .CO(n175), .S(n179) );
  NOR2_X1 U221 ( .A1(n176), .A2(n175), .ZN(n174) );
  MUX2_X1 U222 ( .A(n334), .B(n174), .S(n18), .Z(n365) );
  NAND2_X1 U223 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U224 ( .A(n335), .B(n177), .S(n322), .Z(n367) );
  NAND2_X1 U225 ( .A1(n179), .A2(n178), .ZN(n180) );
  MUX2_X1 U226 ( .A(n336), .B(n180), .S(n322), .Z(n369) );
  XNOR2_X1 U227 ( .A(n182), .B(n181), .ZN(n184) );
  XNOR2_X1 U228 ( .A(n183), .B(n184), .ZN(n202) );
  FA_X1 U229 ( .A(n193), .B(n192), .CI(n191), .CO(n181), .S(n229) );
  XNOR2_X1 U230 ( .A(n195), .B(n194), .ZN(n196) );
  XNOR2_X1 U231 ( .A(n197), .B(n196), .ZN(n228) );
  NOR2_X1 U232 ( .A1(n202), .A2(n203), .ZN(n198) );
  MUX2_X1 U233 ( .A(n337), .B(n198), .S(n322), .Z(n371) );
  NAND2_X1 U234 ( .A1(n200), .A2(n199), .ZN(n201) );
  MUX2_X1 U235 ( .A(n338), .B(n201), .S(n322), .Z(n373) );
  NAND2_X1 U236 ( .A1(n202), .A2(n203), .ZN(n204) );
  MUX2_X1 U237 ( .A(n339), .B(n204), .S(n18), .Z(n375) );
  FA_X1 U238 ( .A(n207), .B(n206), .CI(n205), .CO(n178), .S(n226) );
  XNOR2_X1 U239 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n209) );
  OAI22_X1 U240 ( .A1(n214), .A2(n209), .B1(n216), .B2(n208), .ZN(n212) );
  XNOR2_X1 U241 ( .A(n548), .B(\mult_x_1/n286 ), .ZN(n215) );
  OAI22_X1 U242 ( .A1(n218), .A2(n215), .B1(n210), .B2(n23), .ZN(n211) );
  NOR2_X1 U243 ( .A1(n226), .A2(n225), .ZN(n262) );
  HA_X1 U244 ( .A(n212), .B(n211), .CO(n225), .S(n223) );
  OR2_X1 U245 ( .A1(\mult_x_1/n288 ), .A2(n323), .ZN(n213) );
  OAI22_X1 U246 ( .A1(n214), .A2(n323), .B1(n213), .B2(n216), .ZN(n222) );
  OR2_X1 U247 ( .A1(n223), .A2(n222), .ZN(n258) );
  XNOR2_X1 U248 ( .A(n548), .B(\mult_x_1/n287 ), .ZN(n217) );
  OAI22_X1 U249 ( .A1(n218), .A2(n217), .B1(n215), .B2(n23), .ZN(n221) );
  AND2_X1 U250 ( .A1(\mult_x_1/n288 ), .A2(n48), .ZN(n220) );
  NOR2_X1 U251 ( .A1(n221), .A2(n220), .ZN(n251) );
  OAI22_X1 U252 ( .A1(n218), .A2(\mult_x_1/n288 ), .B1(n217), .B2(n23), .ZN(
        n248) );
  OR2_X1 U253 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n219) );
  NAND2_X1 U254 ( .A1(n219), .A2(n218), .ZN(n247) );
  NAND2_X1 U255 ( .A1(n248), .A2(n247), .ZN(n254) );
  NAND2_X1 U256 ( .A1(n221), .A2(n220), .ZN(n252) );
  OAI21_X1 U257 ( .B1(n251), .B2(n254), .A(n252), .ZN(n259) );
  NAND2_X1 U258 ( .A1(n223), .A2(n222), .ZN(n257) );
  INV_X1 U259 ( .A(n257), .ZN(n224) );
  AOI21_X1 U260 ( .B1(n258), .B2(n259), .A(n224), .ZN(n265) );
  NAND2_X1 U261 ( .A1(n226), .A2(n225), .ZN(n263) );
  OAI21_X1 U262 ( .B1(n262), .B2(n265), .A(n263), .ZN(n227) );
  MUX2_X1 U263 ( .A(n340), .B(n227), .S(n322), .Z(n377) );
  FA_X1 U264 ( .A(n230), .B(n229), .CI(n228), .CO(n203), .S(n231) );
  MUX2_X1 U265 ( .A(n341), .B(n231), .S(n322), .Z(n379) );
  FA_X1 U266 ( .A(n26), .B(n233), .CI(n232), .CO(n234), .S(n73) );
  MUX2_X1 U267 ( .A(n342), .B(n234), .S(en), .Z(n381) );
  FA_X1 U268 ( .A(n237), .B(n236), .CI(n235), .CO(n238), .S(n57) );
  MUX2_X1 U269 ( .A(n344), .B(n238), .S(en), .Z(n385) );
  MUX2_X1 U270 ( .A(n346), .B(n245), .S(en), .Z(n389) );
  MUX2_X1 U271 ( .A(product[0]), .B(n512), .S(n18), .Z(n404) );
  MUX2_X1 U272 ( .A(n512), .B(n513), .S(n18), .Z(n406) );
  AND2_X1 U273 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n246) );
  MUX2_X1 U274 ( .A(n513), .B(n246), .S(n18), .Z(n408) );
  MUX2_X1 U275 ( .A(product[1]), .B(n515), .S(n19), .Z(n410) );
  MUX2_X1 U276 ( .A(n515), .B(n516), .S(n19), .Z(n412) );
  OR2_X1 U277 ( .A1(n248), .A2(n247), .ZN(n249) );
  AND2_X1 U278 ( .A1(n249), .A2(n254), .ZN(n250) );
  MUX2_X1 U279 ( .A(n516), .B(n250), .S(n19), .Z(n414) );
  MUX2_X1 U280 ( .A(product[2]), .B(n518), .S(n19), .Z(n416) );
  MUX2_X1 U281 ( .A(n518), .B(n519), .S(n19), .Z(n418) );
  INV_X1 U282 ( .A(n251), .ZN(n253) );
  NAND2_X1 U283 ( .A1(n253), .A2(n252), .ZN(n255) );
  XOR2_X1 U284 ( .A(n255), .B(n254), .Z(n256) );
  MUX2_X1 U285 ( .A(n519), .B(n256), .S(n19), .Z(n420) );
  MUX2_X1 U286 ( .A(product[3]), .B(n521), .S(n19), .Z(n422) );
  MUX2_X1 U287 ( .A(n521), .B(n522), .S(n19), .Z(n424) );
  NAND2_X1 U288 ( .A1(n258), .A2(n257), .ZN(n260) );
  XNOR2_X1 U289 ( .A(n260), .B(n259), .ZN(n261) );
  MUX2_X1 U290 ( .A(n522), .B(n261), .S(n19), .Z(n426) );
  MUX2_X1 U291 ( .A(product[4]), .B(n524), .S(n19), .Z(n428) );
  MUX2_X1 U292 ( .A(n524), .B(n525), .S(n19), .Z(n430) );
  INV_X1 U293 ( .A(n262), .ZN(n264) );
  NAND2_X1 U294 ( .A1(n264), .A2(n263), .ZN(n266) );
  XOR2_X1 U295 ( .A(n266), .B(n265), .Z(n267) );
  MUX2_X1 U296 ( .A(n525), .B(n267), .S(n19), .Z(n432) );
  MUX2_X1 U297 ( .A(product[5]), .B(n527), .S(n19), .Z(n434) );
  NAND2_X1 U298 ( .A1(n325), .A2(n336), .ZN(n268) );
  XNOR2_X1 U299 ( .A(n268), .B(n340), .ZN(n269) );
  MUX2_X1 U300 ( .A(n527), .B(n269), .S(n19), .Z(n436) );
  MUX2_X1 U301 ( .A(product[6]), .B(n529), .S(n322), .Z(n438) );
  NAND2_X1 U302 ( .A1(n393), .A2(n335), .ZN(n270) );
  AOI21_X1 U303 ( .B1(n325), .B2(n340), .A(n396), .ZN(n272) );
  XOR2_X1 U304 ( .A(n270), .B(n272), .Z(n271) );
  MUX2_X1 U305 ( .A(n529), .B(n271), .S(n322), .Z(n440) );
  MUX2_X1 U306 ( .A(product[7]), .B(n531), .S(n322), .Z(n442) );
  OAI21_X1 U307 ( .B1(n334), .B2(n272), .A(n335), .ZN(n275) );
  NAND2_X1 U308 ( .A1(n328), .A2(n333), .ZN(n273) );
  XNOR2_X1 U309 ( .A(n275), .B(n273), .ZN(n274) );
  MUX2_X1 U310 ( .A(n531), .B(n274), .S(n322), .Z(n444) );
  MUX2_X1 U311 ( .A(product[8]), .B(n533), .S(n322), .Z(n446) );
  AOI21_X1 U312 ( .B1(n275), .B2(n328), .A(n395), .ZN(n278) );
  NAND2_X1 U313 ( .A1(n397), .A2(n332), .ZN(n276) );
  XOR2_X1 U314 ( .A(n278), .B(n276), .Z(n277) );
  MUX2_X1 U315 ( .A(n533), .B(n277), .S(n322), .Z(n448) );
  MUX2_X1 U316 ( .A(product[9]), .B(n535), .S(n322), .Z(n450) );
  OAI21_X1 U317 ( .B1(n278), .B2(n331), .A(n332), .ZN(n292) );
  INV_X1 U318 ( .A(n292), .ZN(n282) );
  NOR2_X1 U319 ( .A1(n345), .A2(n346), .ZN(n287) );
  INV_X1 U320 ( .A(n287), .ZN(n279) );
  NAND2_X1 U321 ( .A1(n345), .A2(n346), .ZN(n289) );
  NAND2_X1 U322 ( .A1(n279), .A2(n289), .ZN(n280) );
  XOR2_X1 U323 ( .A(n282), .B(n280), .Z(n281) );
  MUX2_X1 U324 ( .A(n535), .B(n281), .S(n322), .Z(n452) );
  MUX2_X1 U325 ( .A(product[10]), .B(n537), .S(n322), .Z(n454) );
  OAI21_X1 U326 ( .B1(n282), .B2(n287), .A(n289), .ZN(n285) );
  NOR2_X1 U327 ( .A1(n343), .A2(n344), .ZN(n290) );
  INV_X1 U328 ( .A(n290), .ZN(n283) );
  NAND2_X1 U329 ( .A1(n343), .A2(n344), .ZN(n288) );
  NAND2_X1 U330 ( .A1(n283), .A2(n288), .ZN(n284) );
  XNOR2_X1 U331 ( .A(n285), .B(n284), .ZN(n286) );
  MUX2_X1 U332 ( .A(n537), .B(n286), .S(n322), .Z(n456) );
  MUX2_X1 U333 ( .A(product[11]), .B(n539), .S(n322), .Z(n458) );
  NOR2_X1 U334 ( .A1(n290), .A2(n287), .ZN(n293) );
  OAI21_X1 U335 ( .B1(n290), .B2(n289), .A(n288), .ZN(n291) );
  AOI21_X1 U336 ( .B1(n293), .B2(n292), .A(n291), .ZN(n319) );
  NOR2_X1 U337 ( .A1(n341), .A2(n342), .ZN(n305) );
  INV_X1 U338 ( .A(n305), .ZN(n315) );
  NAND2_X1 U339 ( .A1(n341), .A2(n342), .ZN(n307) );
  NAND2_X1 U340 ( .A1(n315), .A2(n307), .ZN(n294) );
  XOR2_X1 U341 ( .A(n319), .B(n294), .Z(n295) );
  MUX2_X1 U342 ( .A(n539), .B(n295), .S(n322), .Z(n460) );
  MUX2_X1 U343 ( .A(product[12]), .B(n541), .S(n322), .Z(n462) );
  OAI21_X1 U344 ( .B1(n319), .B2(n305), .A(n307), .ZN(n297) );
  NAND2_X1 U345 ( .A1(n398), .A2(n339), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n298) );
  MUX2_X1 U347 ( .A(n541), .B(n298), .S(n322), .Z(n464) );
  MUX2_X1 U348 ( .A(product[13]), .B(n543), .S(n322), .Z(n466) );
  NAND2_X1 U349 ( .A1(n315), .A2(n398), .ZN(n301) );
  INV_X1 U350 ( .A(n307), .ZN(n299) );
  AOI21_X1 U351 ( .B1(n299), .B2(n398), .A(n399), .ZN(n300) );
  OAI21_X1 U352 ( .B1(n319), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U353 ( .A1(n327), .A2(n338), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U355 ( .A(n543), .B(n304), .S(n322), .Z(n468) );
  MUX2_X1 U356 ( .A(product[14]), .B(n545), .S(n322), .Z(n470) );
  NAND2_X1 U357 ( .A1(n398), .A2(n327), .ZN(n313) );
  OR2_X1 U358 ( .A1(n305), .A2(n313), .ZN(n309) );
  AOI21_X1 U359 ( .B1(n399), .B2(n327), .A(n394), .ZN(n306) );
  OAI21_X1 U360 ( .B1(n313), .B2(n307), .A(n306), .ZN(n316) );
  INV_X1 U361 ( .A(n316), .ZN(n308) );
  OAI21_X1 U362 ( .B1(n319), .B2(n309), .A(n308), .ZN(n311) );
  NAND2_X1 U363 ( .A1(n326), .A2(n330), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  MUX2_X1 U365 ( .A(n545), .B(n312), .S(n322), .Z(n472) );
  MUX2_X1 U366 ( .A(product[15]), .B(n547), .S(n17), .Z(n474) );
  NOR2_X1 U367 ( .A1(n313), .A2(n392), .ZN(n314) );
  NAND2_X1 U368 ( .A1(n315), .A2(n314), .ZN(n318) );
  AOI21_X1 U369 ( .B1(n316), .B2(n326), .A(n391), .ZN(n317) );
  OAI21_X1 U370 ( .B1(n319), .B2(n318), .A(n317), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n320), .B(n329), .ZN(n321) );
  MUX2_X1 U372 ( .A(n547), .B(n321), .S(n17), .Z(n476) );
  MUX2_X1 U373 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n322), .Z(n478) );
  MUX2_X1 U374 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n322), .Z(n480) );
  MUX2_X1 U375 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n322), .Z(n482) );
  MUX2_X1 U376 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n322), .Z(n484) );
  MUX2_X1 U377 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n322), .Z(n486) );
  MUX2_X1 U378 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n322), .Z(n488) );
  MUX2_X1 U379 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n322), .Z(n490) );
  MUX2_X1 U380 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n322), .Z(n492) );
  MUX2_X1 U381 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n17), .Z(n494) );
  MUX2_X1 U382 ( .A(n548), .B(A_extended[1]), .S(n322), .Z(n496) );
  MUX2_X1 U383 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n17), .Z(n498) );
  MUX2_X1 U384 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n322), .Z(n500) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n17), .Z(n502) );
  MUX2_X1 U386 ( .A(n22), .B(A_extended[5]), .S(n17), .Z(n504) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n17), .Z(n506) );
  MUX2_X1 U388 ( .A(n20), .B(A_extended[7]), .S(n17), .Z(n508) );
  OR2_X1 U389 ( .A1(n17), .A2(n550), .ZN(n510) );
endmodule


module conv_128_32_DW_mult_pipe_J1_6 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n350,
         n352, n354, n356, n358, n360, n362, n364, n366, n368, n370, n372,
         n374, n376, n378, n380, n382, n384, n386, n388, n390, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n420, n422, n424, n426, n428,
         n430, n432, n434, n436, n438, n440, n442, n444, n446, n448, n450,
         n452, n454, n456, n458, n460, n462, n464, n466, n468, n470, n472,
         n474, n476, n478, n480, n482, n484, n486, n488, n490, n492, n494,
         n496, n498, n500, n502, n504, n506, n508, n510, n512, n513, n515,
         n516, n518, n519, n521, n522, n524, n525, n527, n529, n531, n533,
         n535, n537, n539, n541, n543, n545, n547, n548, n549, n550;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n402), .SE(n510), .CK(clk), .Q(n549), 
        .QN(n323) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n402), .SE(n506), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n19) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n402), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n18) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n402), .SE(n500), .CK(clk), .Q(n548), 
        .QN(n322) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n402), .SE(n498), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n20) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n402), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n21) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n402), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n5) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n402), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n402), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n402), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n402), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(rst_n), .SE(n476), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(rst_n), .SE(n474), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n470), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(rst_n), .SE(n468), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n402), .SE(n466), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n402), .SE(n464), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n402), .SE(n462), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(rst_n), .SE(n460), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(rst_n), .SE(n458), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n456), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n454), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(rst_n), .SE(n450), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n448), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n402), .SE(n446), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n402), .SE(n444), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n402), .SE(n442), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n402), .SE(n440), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n402), .SE(n438), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n402), .SE(n436), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n402), .SE(n434), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n402), .SE(n432), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n402), .SE(n430), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n402), .SE(n428), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n402), .SE(n426), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n402), .SE(n424), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n402), .SE(n422), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n402), .SE(n420), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n402), .SE(n418), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n402), .SE(n416), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n402), .SE(n414), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n402), .SE(n412), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n402), .SE(n410), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n402), .SE(n408), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n402), .SE(n406), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n402), .SE(n404), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n550), .SE(n390), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n550), .SE(n388), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2_IP  ( .D(1'b1), .SI(n550), .SE(n386), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n550), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n550), .SE(n382), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2_IP  ( .D(1'b1), .SI(n550), .SE(n380), .CK(
        clk), .Q(n326), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n550), .SE(n378), .CK(
        clk), .Q(n393), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n550), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n340), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2_IP  ( .D(1'b1), .SI(n550), .SE(n374), .CK(
        clk), .Q(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n550), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n339), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n550), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n550), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n337), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n550), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n336), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n550), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n550), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n334), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n550), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n333), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n550), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n332), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n550), .SE(n356), .CK(
        clk), .QN(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n550), .SE(n354), .CK(
        clk), .QN(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n550), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n329), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n550), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n550), .SE(n348), .CK(
        clk), .QN(n327) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n402), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n325) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n402), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n324) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n402), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  OR2_X4 U2 ( .A1(n15), .A2(n22), .ZN(n207) );
  INV_X2 U3 ( .A(n94), .ZN(n129) );
  INV_X1 U4 ( .A(rst_n), .ZN(n550) );
  INV_X2 U5 ( .A(n27), .ZN(n140) );
  NAND2_X1 U6 ( .A1(n9), .A2(n8), .ZN(n242) );
  INV_X1 U7 ( .A(n111), .ZN(n240) );
  INV_X1 U8 ( .A(n111), .ZN(n244) );
  OAI21_X1 U9 ( .B1(n161), .B2(n160), .A(n11), .ZN(n9) );
  BUF_X4 U10 ( .A(en), .Z(n321) );
  NAND2_X1 U11 ( .A1(n161), .A2(n160), .ZN(n8) );
  CLKBUF_X2 U12 ( .A(rst_n), .Z(n402) );
  NAND2_X1 U13 ( .A1(n26), .A2(n25), .ZN(n139) );
  NAND2_X2 U14 ( .A1(n69), .A2(n120), .ZN(n121) );
  INV_X1 U15 ( .A(n22), .ZN(n209) );
  INV_X1 U16 ( .A(n324), .ZN(n14) );
  INV_X1 U17 ( .A(n325), .ZN(n320) );
  XNOR2_X1 U18 ( .A(n10), .B(n161), .ZN(n87) );
  XNOR2_X1 U19 ( .A(n11), .B(n160), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n84), .A2(n83), .ZN(n11) );
  NOR2_X2 U21 ( .A1(n324), .A2(n323), .ZN(n17) );
  NOR2_X1 U22 ( .A1(n196), .A2(n195), .ZN(n197) );
  XNOR2_X1 U23 ( .A(n39), .B(n226), .ZN(n196) );
  INV_X1 U24 ( .A(n68), .ZN(n70) );
  NAND2_X1 U25 ( .A1(n78), .A2(n77), .ZN(n79) );
  INV_X1 U26 ( .A(n82), .ZN(n78) );
  CLKBUF_X1 U27 ( .A(\mult_x_1/n281 ), .Z(n12) );
  NAND2_X2 U28 ( .A1(n113), .A2(n5), .ZN(n212) );
  OAI22_X1 U29 ( .A1(n207), .A2(n38), .B1(n59), .B2(n209), .ZN(n13) );
  XNOR2_X1 U30 ( .A(\mult_x_1/a[2] ), .B(n548), .ZN(n15) );
  XNOR2_X1 U31 ( .A(n80), .B(n66), .ZN(n222) );
  OAI22_X1 U32 ( .A1(n207), .A2(n38), .B1(n59), .B2(n209), .ZN(n75) );
  XNOR2_X1 U33 ( .A(n142), .B(n46), .ZN(n16) );
  NOR2_X1 U34 ( .A1(n323), .A2(n324), .ZN(n142) );
  XNOR2_X2 U35 ( .A(n322), .B(n18), .ZN(n120) );
  XNOR2_X1 U36 ( .A(n20), .B(\mult_x_1/n313 ), .ZN(n22) );
  XNOR2_X1 U37 ( .A(n548), .B(\mult_x_1/n282 ), .ZN(n44) );
  XNOR2_X1 U38 ( .A(n548), .B(n12), .ZN(n38) );
  OAI22_X1 U39 ( .A1(n207), .A2(n44), .B1(n209), .B2(n38), .ZN(n29) );
  XOR2_X1 U40 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n69) );
  XNOR2_X1 U41 ( .A(n320), .B(\mult_x_1/n284 ), .ZN(n43) );
  INV_X1 U42 ( .A(n120), .ZN(n94) );
  XNOR2_X1 U43 ( .A(n320), .B(\mult_x_1/n283 ), .ZN(n37) );
  OAI22_X1 U44 ( .A1(n121), .A2(n43), .B1(n120), .B2(n37), .ZN(n30) );
  OR2_X1 U45 ( .A1(n29), .A2(n30), .ZN(n57) );
  XNOR2_X1 U46 ( .A(n17), .B(\mult_x_1/n286 ), .ZN(n23) );
  INV_X1 U47 ( .A(\mult_x_1/n310 ), .ZN(n46) );
  XNOR2_X1 U48 ( .A(n17), .B(n46), .ZN(n35) );
  INV_X1 U49 ( .A(n16), .ZN(n143) );
  NOR2_X1 U50 ( .A1(n23), .A2(n143), .ZN(n56) );
  BUF_X2 U51 ( .A(\mult_x_1/n313 ), .Z(n113) );
  AND2_X1 U52 ( .A1(n549), .A2(\mult_x_1/n281 ), .ZN(n99) );
  XNOR2_X1 U53 ( .A(n99), .B(n113), .ZN(n34) );
  AOI21_X1 U54 ( .B1(n212), .B2(n5), .A(n34), .ZN(n24) );
  INV_X1 U55 ( .A(n24), .ZN(n42) );
  XNOR2_X1 U56 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n26) );
  XNOR2_X1 U57 ( .A(\mult_x_1/n310 ), .B(n19), .ZN(n25) );
  XNOR2_X1 U58 ( .A(n14), .B(\mult_x_1/n286 ), .ZN(n33) );
  INV_X1 U59 ( .A(n26), .ZN(n27) );
  XNOR2_X1 U60 ( .A(n14), .B(\mult_x_1/n285 ), .ZN(n36) );
  OAI22_X1 U61 ( .A1(n139), .A2(n33), .B1(n140), .B2(n36), .ZN(n41) );
  XNOR2_X1 U62 ( .A(n17), .B(\mult_x_1/n287 ), .ZN(n28) );
  NOR2_X1 U63 ( .A1(n28), .A2(n143), .ZN(n40) );
  XNOR2_X1 U64 ( .A(n30), .B(n29), .ZN(n51) );
  INV_X1 U65 ( .A(n17), .ZN(n31) );
  OR2_X1 U66 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n32) );
  NOR2_X1 U67 ( .A1(n32), .A2(n143), .ZN(n50) );
  XNOR2_X1 U68 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n47) );
  OAI22_X1 U69 ( .A1(n139), .A2(n47), .B1(n140), .B2(n33), .ZN(n165) );
  XNOR2_X1 U70 ( .A(n113), .B(n12), .ZN(n122) );
  OAI22_X1 U71 ( .A1(n212), .A2(n122), .B1(n34), .B2(n5), .ZN(n164) );
  AND2_X1 U72 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n163) );
  XNOR2_X1 U73 ( .A(n14), .B(\mult_x_1/n284 ), .ZN(n58) );
  OAI22_X1 U74 ( .A1(n139), .A2(n36), .B1(n140), .B2(n58), .ZN(n63) );
  XNOR2_X1 U75 ( .A(n320), .B(\mult_x_1/n282 ), .ZN(n65) );
  OAI22_X1 U76 ( .A1(n121), .A2(n37), .B1(n120), .B2(n65), .ZN(n62) );
  XNOR2_X1 U77 ( .A(n99), .B(n548), .ZN(n59) );
  INV_X1 U78 ( .A(n75), .ZN(n61) );
  XNOR2_X1 U79 ( .A(n228), .B(n227), .ZN(n39) );
  FA_X1 U80 ( .A(n42), .B(n41), .CI(n40), .CO(n55), .S(n235) );
  XNOR2_X1 U81 ( .A(n320), .B(\mult_x_1/n285 ), .ZN(n119) );
  OAI22_X1 U82 ( .A1(n121), .A2(n119), .B1(n129), .B2(n43), .ZN(n171) );
  XNOR2_X1 U83 ( .A(n548), .B(\mult_x_1/n283 ), .ZN(n124) );
  OAI22_X1 U84 ( .A1(n207), .A2(n124), .B1(n209), .B2(n44), .ZN(n170) );
  OR2_X1 U85 ( .A1(\mult_x_1/n288 ), .A2(n46), .ZN(n45) );
  OAI22_X1 U86 ( .A1(n139), .A2(n46), .B1(n45), .B2(n140), .ZN(n118) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n48) );
  OAI22_X1 U88 ( .A1(n139), .A2(n48), .B1(n140), .B2(n47), .ZN(n117) );
  FA_X1 U89 ( .A(n51), .B(n50), .CI(n49), .CO(n228), .S(n233) );
  NAND2_X1 U90 ( .A1(n196), .A2(n195), .ZN(n52) );
  INV_X1 U91 ( .A(en), .ZN(n111) );
  NAND2_X1 U92 ( .A1(n52), .A2(n240), .ZN(n54) );
  OR2_X1 U93 ( .A1(n240), .A2(n326), .ZN(n53) );
  NAND2_X1 U94 ( .A1(n54), .A2(n53), .ZN(n380) );
  FA_X1 U95 ( .A(n57), .B(n56), .CI(n55), .CO(n224), .S(n226) );
  XNOR2_X1 U96 ( .A(n14), .B(\mult_x_1/n283 ), .ZN(n72) );
  OAI22_X1 U97 ( .A1(n139), .A2(n58), .B1(n140), .B2(n72), .ZN(n76) );
  AOI21_X1 U98 ( .B1(n209), .B2(n207), .A(n59), .ZN(n60) );
  INV_X1 U99 ( .A(n60), .ZN(n74) );
  FA_X1 U100 ( .A(n63), .B(n62), .CI(n61), .CO(n80), .S(n227) );
  XNOR2_X1 U101 ( .A(n17), .B(\mult_x_1/n285 ), .ZN(n64) );
  NOR2_X1 U102 ( .A1(n64), .A2(n143), .ZN(n82) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n68) );
  OAI22_X1 U104 ( .A1(n121), .A2(n65), .B1(n129), .B2(n68), .ZN(n81) );
  XNOR2_X1 U105 ( .A(n82), .B(n81), .ZN(n66) );
  INV_X1 U106 ( .A(n86), .ZN(n67) );
  NAND2_X1 U107 ( .A1(n67), .A2(n240), .ZN(n85) );
  XNOR2_X1 U108 ( .A(n99), .B(n320), .ZN(n102) );
  NAND3_X1 U109 ( .A1(n70), .A2(n69), .A3(n120), .ZN(n71) );
  OAI21_X1 U110 ( .B1(n129), .B2(n102), .A(n71), .ZN(n109) );
  INV_X1 U111 ( .A(n109), .ZN(n106) );
  XNOR2_X1 U112 ( .A(n14), .B(\mult_x_1/n282 ), .ZN(n101) );
  OAI22_X1 U113 ( .A1(n139), .A2(n72), .B1(n140), .B2(n101), .ZN(n105) );
  XNOR2_X1 U114 ( .A(n17), .B(\mult_x_1/n284 ), .ZN(n73) );
  NOR2_X1 U115 ( .A1(n73), .A2(n143), .ZN(n104) );
  FA_X1 U116 ( .A(n76), .B(n13), .CI(n74), .CO(n160), .S(n223) );
  INV_X1 U117 ( .A(n81), .ZN(n77) );
  NAND2_X1 U118 ( .A1(n80), .A2(n79), .ZN(n84) );
  NAND2_X1 U119 ( .A1(n82), .A2(n81), .ZN(n83) );
  OAI22_X1 U120 ( .A1(n85), .A2(n87), .B1(n240), .B2(n400), .ZN(n374) );
  NAND2_X1 U121 ( .A1(n87), .A2(n86), .ZN(n88) );
  NAND2_X1 U122 ( .A1(n88), .A2(n240), .ZN(n90) );
  OR2_X1 U123 ( .A1(n240), .A2(n401), .ZN(n89) );
  NAND2_X1 U124 ( .A1(n90), .A2(n89), .ZN(n376) );
  XNOR2_X1 U147 ( .A(n548), .B(\mult_x_1/n286 ), .ZN(n95) );
  XNOR2_X1 U148 ( .A(n548), .B(\mult_x_1/n285 ), .ZN(n116) );
  OAI22_X1 U149 ( .A1(n207), .A2(n95), .B1(n209), .B2(n116), .ZN(n187) );
  XNOR2_X1 U150 ( .A(n113), .B(\mult_x_1/n284 ), .ZN(n93) );
  XNOR2_X1 U151 ( .A(n113), .B(\mult_x_1/n283 ), .ZN(n114) );
  OAI22_X1 U152 ( .A1(n212), .A2(n93), .B1(n114), .B2(n5), .ZN(n186) );
  OR2_X1 U153 ( .A1(\mult_x_1/n288 ), .A2(n325), .ZN(n91) );
  OAI22_X1 U154 ( .A1(n121), .A2(n325), .B1(n91), .B2(n129), .ZN(n127) );
  XNOR2_X1 U155 ( .A(n320), .B(\mult_x_1/n288 ), .ZN(n92) );
  XNOR2_X1 U156 ( .A(n320), .B(\mult_x_1/n287 ), .ZN(n130) );
  OAI22_X1 U157 ( .A1(n121), .A2(n92), .B1(n129), .B2(n130), .ZN(n126) );
  XNOR2_X1 U158 ( .A(n113), .B(\mult_x_1/n285 ), .ZN(n203) );
  OAI22_X1 U159 ( .A1(n212), .A2(n203), .B1(n93), .B2(n5), .ZN(n200) );
  AND2_X1 U160 ( .A1(\mult_x_1/n288 ), .A2(n94), .ZN(n199) );
  XNOR2_X1 U161 ( .A(n548), .B(\mult_x_1/n287 ), .ZN(n201) );
  OAI22_X1 U162 ( .A1(n207), .A2(n201), .B1(n209), .B2(n95), .ZN(n198) );
  NOR2_X1 U163 ( .A1(n193), .A2(n192), .ZN(n97) );
  NAND2_X1 U164 ( .A1(n111), .A2(n327), .ZN(n96) );
  OAI21_X1 U165 ( .B1(n111), .B2(n97), .A(n96), .ZN(n348) );
  XNOR2_X1 U166 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n98) );
  NOR2_X1 U167 ( .A1(n98), .A2(n143), .ZN(n137) );
  XNOR2_X1 U168 ( .A(n14), .B(n12), .ZN(n100) );
  XNOR2_X1 U169 ( .A(n99), .B(n14), .ZN(n138) );
  OAI22_X1 U170 ( .A1(n139), .A2(n100), .B1(n138), .B2(n140), .ZN(n148) );
  INV_X1 U171 ( .A(n148), .ZN(n136) );
  OAI22_X1 U172 ( .A1(n139), .A2(n101), .B1(n140), .B2(n100), .ZN(n110) );
  AOI21_X1 U173 ( .B1(n129), .B2(n121), .A(n102), .ZN(n103) );
  INV_X1 U174 ( .A(n103), .ZN(n108) );
  FA_X1 U175 ( .A(n106), .B(n105), .CI(n104), .CO(n159), .S(n161) );
  XNOR2_X1 U176 ( .A(n17), .B(\mult_x_1/n283 ), .ZN(n107) );
  NOR2_X1 U177 ( .A1(n107), .A2(n143), .ZN(n158) );
  FA_X1 U178 ( .A(n110), .B(n109), .CI(n108), .CO(n135), .S(n157) );
  OR2_X1 U179 ( .A1(n155), .A2(n154), .ZN(n112) );
  MUX2_X1 U180 ( .A(n328), .B(n112), .S(n244), .Z(n350) );
  XNOR2_X1 U181 ( .A(n113), .B(\mult_x_1/n282 ), .ZN(n123) );
  OAI22_X1 U182 ( .A1(n212), .A2(n114), .B1(n123), .B2(n5), .ZN(n133) );
  INV_X1 U183 ( .A(n140), .ZN(n115) );
  AND2_X1 U184 ( .A1(\mult_x_1/n288 ), .A2(n115), .ZN(n132) );
  XNOR2_X1 U185 ( .A(n548), .B(\mult_x_1/n284 ), .ZN(n125) );
  OAI22_X1 U186 ( .A1(n207), .A2(n116), .B1(n209), .B2(n125), .ZN(n131) );
  HA_X1 U187 ( .A(n118), .B(n117), .CO(n169), .S(n173) );
  XNOR2_X1 U188 ( .A(n320), .B(\mult_x_1/n286 ), .ZN(n128) );
  OAI22_X1 U189 ( .A1(n121), .A2(n128), .B1(n129), .B2(n119), .ZN(n168) );
  OAI22_X1 U190 ( .A1(n212), .A2(n123), .B1(n122), .B2(n5), .ZN(n167) );
  OAI22_X1 U191 ( .A1(n207), .A2(n125), .B1(n209), .B2(n124), .ZN(n166) );
  HA_X1 U192 ( .A(n127), .B(n126), .CO(n184), .S(n185) );
  OAI22_X1 U193 ( .A1(n121), .A2(n130), .B1(n129), .B2(n128), .ZN(n183) );
  FA_X1 U194 ( .A(n133), .B(n132), .CI(n131), .CO(n174), .S(n182) );
  OR2_X1 U195 ( .A1(n180), .A2(n179), .ZN(n134) );
  MUX2_X1 U196 ( .A(n330), .B(n134), .S(n244), .Z(n354) );
  FA_X1 U197 ( .A(n137), .B(n136), .CI(n135), .CO(n150), .S(n155) );
  AOI21_X1 U198 ( .B1(n140), .B2(n139), .A(n138), .ZN(n141) );
  INV_X1 U199 ( .A(n141), .ZN(n146) );
  XNOR2_X1 U200 ( .A(n17), .B(n12), .ZN(n144) );
  NOR2_X1 U201 ( .A1(n144), .A2(n143), .ZN(n145) );
  XOR2_X1 U202 ( .A(n146), .B(n145), .Z(n147) );
  XOR2_X1 U203 ( .A(n148), .B(n147), .Z(n149) );
  OR2_X1 U204 ( .A1(n150), .A2(n149), .ZN(n152) );
  NAND2_X1 U205 ( .A1(n150), .A2(n149), .ZN(n151) );
  NAND2_X1 U206 ( .A1(n152), .A2(n151), .ZN(n153) );
  MUX2_X1 U207 ( .A(n331), .B(n153), .S(n244), .Z(n356) );
  NAND2_X1 U208 ( .A1(n155), .A2(n154), .ZN(n156) );
  MUX2_X1 U209 ( .A(n332), .B(n156), .S(n244), .Z(n358) );
  FA_X1 U210 ( .A(n159), .B(n158), .CI(n157), .CO(n154), .S(n243) );
  NAND2_X1 U211 ( .A1(n243), .A2(n242), .ZN(n162) );
  MUX2_X1 U212 ( .A(n333), .B(n162), .S(n244), .Z(n360) );
  FA_X1 U213 ( .A(n163), .B(n164), .CI(n165), .CO(n49), .S(n239) );
  FA_X1 U214 ( .A(n168), .B(n167), .CI(n166), .CO(n238), .S(n172) );
  FA_X1 U215 ( .A(n171), .B(n170), .CI(n169), .CO(n234), .S(n237) );
  FA_X1 U216 ( .A(n174), .B(n173), .CI(n172), .CO(n176), .S(n180) );
  NOR2_X1 U217 ( .A1(n177), .A2(n176), .ZN(n175) );
  MUX2_X1 U218 ( .A(n334), .B(n175), .S(n244), .Z(n362) );
  NAND2_X1 U219 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2_X1 U220 ( .A(n335), .B(n178), .S(n244), .Z(n364) );
  NAND2_X1 U221 ( .A1(n180), .A2(n179), .ZN(n181) );
  MUX2_X1 U222 ( .A(n336), .B(n181), .S(n244), .Z(n366) );
  FA_X1 U223 ( .A(n184), .B(n183), .CI(n182), .CO(n179), .S(n190) );
  FA_X1 U224 ( .A(n187), .B(n186), .CI(n185), .CO(n189), .S(n193) );
  NOR2_X1 U225 ( .A1(n190), .A2(n189), .ZN(n188) );
  MUX2_X1 U226 ( .A(n337), .B(n188), .S(n240), .Z(n368) );
  NAND2_X1 U227 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U228 ( .A(n338), .B(n191), .S(n240), .Z(n370) );
  NAND2_X1 U229 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U230 ( .A(n339), .B(n194), .S(n240), .Z(n372) );
  MUX2_X1 U231 ( .A(n341), .B(n197), .S(n240), .Z(n378) );
  FA_X1 U232 ( .A(n200), .B(n199), .CI(n198), .CO(n192), .S(n220) );
  XNOR2_X1 U233 ( .A(n548), .B(\mult_x_1/n288 ), .ZN(n202) );
  OAI22_X1 U234 ( .A1(n207), .A2(n202), .B1(n209), .B2(n201), .ZN(n205) );
  XNOR2_X1 U235 ( .A(n113), .B(\mult_x_1/n286 ), .ZN(n208) );
  OAI22_X1 U236 ( .A1(n212), .A2(n208), .B1(n203), .B2(n5), .ZN(n204) );
  NOR2_X1 U237 ( .A1(n220), .A2(n219), .ZN(n263) );
  HA_X1 U238 ( .A(n205), .B(n204), .CO(n219), .S(n217) );
  OR2_X1 U239 ( .A1(\mult_x_1/n288 ), .A2(n322), .ZN(n206) );
  OAI22_X1 U240 ( .A1(n207), .A2(n322), .B1(n206), .B2(n209), .ZN(n216) );
  OR2_X1 U241 ( .A1(n217), .A2(n216), .ZN(n259) );
  XNOR2_X1 U242 ( .A(n113), .B(\mult_x_1/n287 ), .ZN(n211) );
  OAI22_X1 U243 ( .A1(n212), .A2(n211), .B1(n208), .B2(n5), .ZN(n215) );
  AND2_X1 U244 ( .A1(\mult_x_1/n288 ), .A2(n22), .ZN(n214) );
  NOR2_X1 U245 ( .A1(n215), .A2(n214), .ZN(n252) );
  OAI22_X1 U246 ( .A1(n212), .A2(\mult_x_1/n288 ), .B1(n211), .B2(n5), .ZN(
        n249) );
  OR2_X1 U247 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n213) );
  NAND2_X1 U248 ( .A1(n213), .A2(n212), .ZN(n248) );
  NAND2_X1 U249 ( .A1(n249), .A2(n248), .ZN(n255) );
  NAND2_X1 U250 ( .A1(n215), .A2(n214), .ZN(n253) );
  OAI21_X1 U251 ( .B1(n252), .B2(n255), .A(n253), .ZN(n260) );
  NAND2_X1 U252 ( .A1(n217), .A2(n216), .ZN(n258) );
  INV_X1 U253 ( .A(n258), .ZN(n218) );
  AOI21_X1 U254 ( .B1(n259), .B2(n260), .A(n218), .ZN(n266) );
  NAND2_X1 U255 ( .A1(n220), .A2(n219), .ZN(n264) );
  OAI21_X1 U256 ( .B1(n263), .B2(n266), .A(n264), .ZN(n221) );
  MUX2_X1 U257 ( .A(n343), .B(n221), .S(n240), .Z(n382) );
  FA_X1 U258 ( .A(n224), .B(n223), .CI(n222), .CO(n86), .S(n225) );
  MUX2_X1 U259 ( .A(n344), .B(n225), .S(n240), .Z(n384) );
  NAND2_X1 U260 ( .A1(n226), .A2(n228), .ZN(n231) );
  NAND2_X1 U261 ( .A1(n226), .A2(n227), .ZN(n230) );
  NAND2_X1 U262 ( .A1(n228), .A2(n227), .ZN(n229) );
  NAND3_X1 U263 ( .A1(n231), .A2(n230), .A3(n229), .ZN(n232) );
  MUX2_X1 U264 ( .A(n345), .B(n232), .S(n240), .Z(n386) );
  FA_X1 U265 ( .A(n235), .B(n234), .CI(n233), .CO(n195), .S(n236) );
  MUX2_X1 U266 ( .A(n346), .B(n236), .S(n240), .Z(n388) );
  FA_X1 U267 ( .A(n239), .B(n238), .CI(n237), .CO(n241), .S(n177) );
  MUX2_X1 U268 ( .A(n347), .B(n241), .S(n240), .Z(n390) );
  OAI21_X1 U269 ( .B1(n243), .B2(n242), .A(n244), .ZN(n246) );
  OR2_X1 U270 ( .A1(n244), .A2(n394), .ZN(n245) );
  NAND2_X1 U271 ( .A1(n246), .A2(n245), .ZN(n352) );
  MUX2_X1 U272 ( .A(product[0]), .B(n512), .S(n321), .Z(n404) );
  MUX2_X1 U273 ( .A(n512), .B(n513), .S(n321), .Z(n406) );
  AND2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n247) );
  MUX2_X1 U275 ( .A(n513), .B(n247), .S(en), .Z(n408) );
  MUX2_X1 U276 ( .A(product[1]), .B(n515), .S(en), .Z(n410) );
  MUX2_X1 U277 ( .A(n515), .B(n516), .S(n321), .Z(n412) );
  OR2_X1 U278 ( .A1(n249), .A2(n248), .ZN(n250) );
  AND2_X1 U279 ( .A1(n250), .A2(n255), .ZN(n251) );
  MUX2_X1 U280 ( .A(n516), .B(n251), .S(n321), .Z(n414) );
  MUX2_X1 U281 ( .A(product[2]), .B(n518), .S(n321), .Z(n416) );
  MUX2_X1 U282 ( .A(n518), .B(n519), .S(n321), .Z(n418) );
  INV_X1 U283 ( .A(n252), .ZN(n254) );
  NAND2_X1 U284 ( .A1(n254), .A2(n253), .ZN(n256) );
  XOR2_X1 U285 ( .A(n256), .B(n255), .Z(n257) );
  MUX2_X1 U286 ( .A(n519), .B(n257), .S(n321), .Z(n420) );
  MUX2_X1 U287 ( .A(product[3]), .B(n521), .S(n321), .Z(n422) );
  MUX2_X1 U288 ( .A(n521), .B(n522), .S(n321), .Z(n424) );
  NAND2_X1 U289 ( .A1(n259), .A2(n258), .ZN(n261) );
  XNOR2_X1 U290 ( .A(n261), .B(n260), .ZN(n262) );
  MUX2_X1 U291 ( .A(n522), .B(n262), .S(n321), .Z(n426) );
  MUX2_X1 U292 ( .A(product[4]), .B(n524), .S(n321), .Z(n428) );
  MUX2_X1 U293 ( .A(n524), .B(n525), .S(n321), .Z(n430) );
  INV_X1 U294 ( .A(n263), .ZN(n265) );
  NAND2_X1 U295 ( .A1(n265), .A2(n264), .ZN(n267) );
  XOR2_X1 U296 ( .A(n267), .B(n266), .Z(n268) );
  MUX2_X1 U297 ( .A(n525), .B(n268), .S(n244), .Z(n432) );
  MUX2_X1 U298 ( .A(product[5]), .B(n527), .S(n321), .Z(n434) );
  NAND2_X1 U299 ( .A1(n327), .A2(n339), .ZN(n269) );
  XNOR2_X1 U300 ( .A(n269), .B(n343), .ZN(n270) );
  MUX2_X1 U301 ( .A(n527), .B(n270), .S(n321), .Z(n436) );
  MUX2_X1 U302 ( .A(product[6]), .B(n529), .S(n321), .Z(n438) );
  NAND2_X1 U303 ( .A1(n395), .A2(n338), .ZN(n271) );
  AOI21_X1 U304 ( .B1(n327), .B2(n343), .A(n398), .ZN(n273) );
  XOR2_X1 U305 ( .A(n271), .B(n273), .Z(n272) );
  MUX2_X1 U306 ( .A(n529), .B(n272), .S(n321), .Z(n440) );
  MUX2_X1 U307 ( .A(product[7]), .B(n531), .S(n321), .Z(n442) );
  OAI21_X1 U308 ( .B1(n337), .B2(n273), .A(n338), .ZN(n276) );
  NAND2_X1 U309 ( .A1(n330), .A2(n336), .ZN(n274) );
  XNOR2_X1 U310 ( .A(n276), .B(n274), .ZN(n275) );
  MUX2_X1 U311 ( .A(n531), .B(n275), .S(n321), .Z(n444) );
  MUX2_X1 U312 ( .A(product[8]), .B(n533), .S(n244), .Z(n446) );
  AOI21_X1 U313 ( .B1(n276), .B2(n330), .A(n397), .ZN(n279) );
  NAND2_X1 U314 ( .A1(n399), .A2(n335), .ZN(n277) );
  XOR2_X1 U315 ( .A(n279), .B(n277), .Z(n278) );
  MUX2_X1 U316 ( .A(n533), .B(n278), .S(n321), .Z(n448) );
  MUX2_X1 U317 ( .A(product[9]), .B(n535), .S(n321), .Z(n450) );
  OAI21_X1 U318 ( .B1(n279), .B2(n334), .A(n335), .ZN(n290) );
  INV_X1 U319 ( .A(n290), .ZN(n283) );
  NOR2_X1 U320 ( .A1(n346), .A2(n347), .ZN(n287) );
  INV_X1 U321 ( .A(n287), .ZN(n280) );
  NAND2_X1 U322 ( .A1(n346), .A2(n347), .ZN(n288) );
  NAND2_X1 U323 ( .A1(n280), .A2(n288), .ZN(n281) );
  XOR2_X1 U324 ( .A(n283), .B(n281), .Z(n282) );
  MUX2_X1 U325 ( .A(n535), .B(n282), .S(n321), .Z(n452) );
  MUX2_X1 U326 ( .A(product[10]), .B(n537), .S(n321), .Z(n454) );
  OAI21_X1 U327 ( .B1(n283), .B2(n287), .A(n288), .ZN(n285) );
  NAND2_X1 U328 ( .A1(n393), .A2(n342), .ZN(n284) );
  XNOR2_X1 U329 ( .A(n285), .B(n284), .ZN(n286) );
  MUX2_X1 U330 ( .A(n537), .B(n286), .S(n321), .Z(n456) );
  MUX2_X1 U331 ( .A(product[11]), .B(n539), .S(n244), .Z(n458) );
  NOR2_X1 U332 ( .A1(n341), .A2(n287), .ZN(n291) );
  OAI21_X1 U333 ( .B1(n341), .B2(n288), .A(n342), .ZN(n289) );
  AOI21_X1 U334 ( .B1(n291), .B2(n290), .A(n289), .ZN(n317) );
  NOR2_X1 U335 ( .A1(n344), .A2(n345), .ZN(n304) );
  INV_X1 U336 ( .A(n304), .ZN(n297) );
  NAND2_X1 U337 ( .A1(n344), .A2(n345), .ZN(n306) );
  NAND2_X1 U338 ( .A1(n297), .A2(n306), .ZN(n292) );
  XOR2_X1 U339 ( .A(n317), .B(n292), .Z(n293) );
  MUX2_X1 U340 ( .A(n539), .B(n293), .S(n321), .Z(n460) );
  MUX2_X1 U341 ( .A(product[12]), .B(n541), .S(n321), .Z(n462) );
  OAI21_X1 U342 ( .B1(n317), .B2(n304), .A(n306), .ZN(n295) );
  NAND2_X1 U343 ( .A1(n400), .A2(n340), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n296) );
  MUX2_X1 U345 ( .A(n541), .B(n296), .S(n321), .Z(n464) );
  MUX2_X1 U346 ( .A(product[13]), .B(n543), .S(n321), .Z(n466) );
  NAND2_X1 U347 ( .A1(n297), .A2(n400), .ZN(n300) );
  INV_X1 U348 ( .A(n306), .ZN(n298) );
  AOI21_X1 U349 ( .B1(n298), .B2(n400), .A(n401), .ZN(n299) );
  OAI21_X1 U350 ( .B1(n317), .B2(n300), .A(n299), .ZN(n302) );
  NAND2_X1 U351 ( .A1(n329), .A2(n333), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  MUX2_X1 U353 ( .A(n543), .B(n303), .S(n244), .Z(n468) );
  MUX2_X1 U354 ( .A(product[14]), .B(n545), .S(n321), .Z(n470) );
  NAND2_X1 U355 ( .A1(n400), .A2(n329), .ZN(n307) );
  NOR2_X1 U356 ( .A1(n304), .A2(n307), .ZN(n313) );
  INV_X1 U357 ( .A(n313), .ZN(n309) );
  AOI21_X1 U358 ( .B1(n401), .B2(n329), .A(n396), .ZN(n305) );
  OAI21_X1 U359 ( .B1(n307), .B2(n306), .A(n305), .ZN(n314) );
  INV_X1 U360 ( .A(n314), .ZN(n308) );
  OAI21_X1 U361 ( .B1(n317), .B2(n309), .A(n308), .ZN(n311) );
  NAND2_X1 U362 ( .A1(n328), .A2(n332), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  MUX2_X1 U364 ( .A(n545), .B(n312), .S(n321), .Z(n472) );
  MUX2_X1 U365 ( .A(product[15]), .B(n547), .S(n321), .Z(n474) );
  NAND2_X1 U366 ( .A1(n313), .A2(n328), .ZN(n316) );
  AOI21_X1 U367 ( .B1(n314), .B2(n328), .A(n392), .ZN(n315) );
  OAI21_X1 U368 ( .B1(n317), .B2(n316), .A(n315), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n318), .B(n331), .ZN(n319) );
  MUX2_X1 U370 ( .A(n547), .B(n319), .S(n321), .Z(n476) );
  MUX2_X1 U371 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n321), .Z(n478) );
  MUX2_X1 U372 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n321), .Z(n480) );
  MUX2_X1 U373 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n321), .Z(n482) );
  MUX2_X1 U374 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n321), .Z(n484) );
  MUX2_X1 U375 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n321), .Z(n486) );
  MUX2_X1 U376 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n321), .Z(n488) );
  MUX2_X1 U377 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n321), .Z(n490) );
  MUX2_X1 U378 ( .A(n12), .B(B_extended[7]), .S(n321), .Z(n492) );
  MUX2_X1 U379 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n321), .Z(n494) );
  MUX2_X1 U380 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n321), .Z(n496) );
  MUX2_X1 U381 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n321), .Z(n498) );
  MUX2_X1 U382 ( .A(n548), .B(A_extended[3]), .S(n321), .Z(n500) );
  MUX2_X1 U383 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n321), .Z(n502) );
  MUX2_X1 U384 ( .A(n320), .B(A_extended[5]), .S(n321), .Z(n504) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n321), .Z(n506) );
  MUX2_X1 U386 ( .A(n14), .B(A_extended[7]), .S(n321), .Z(n508) );
  OR2_X1 U387 ( .A1(n321), .A2(n549), .ZN(n510) );
endmodule


module conv_128_32_DW_mult_pipe_J1_7 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n364, n366, n368, n370, n372, n374, n376,
         n378, n380, n382, n384, n386, n388, n390, n392, n394, n396, n398,
         n400, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n442, n444, n446, n448, n450, n452,
         n454, n456, n458, n460, n462, n464, n466, n468, n470, n472, n474,
         n476, n478, n480, n482, n484, n486, n488, n490, n492, n494, n496,
         n498, n500, n502, n504, n506, n508, n510, n512, n514, n516, n518,
         n520, n522, n524, n526, n527, n529, n530, n532, n533, n535, n536,
         n538, n539, n541, n542, n544, n546, n548, n550, n552, n554, n556,
         n558, n560, n562, n563, n564, n565;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n414), .SE(n524), .CK(clk), .Q(n564), 
        .QN(n5) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n414), .SE(n520), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n414), .SE(n516), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n340) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n414), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n30) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n414), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n33) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n414), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n39) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n412), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n40) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n413), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n38) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n411), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n37) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n414), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n35) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n411), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n36) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n411), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n32) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n411), .SE(n490), .CK(clk), .Q(n562)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n411), .SE(n488), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n411), .SE(n486), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n411), .SE(n484), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n411), .SE(n482), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n413), .SE(n480), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n412), .SE(n478), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n414), .SE(n476), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n411), .SE(n474), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n411), .SE(n472), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n411), .SE(n470), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n411), .SE(n468), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n411), .SE(n466), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n411), .SE(n464), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n411), .SE(n462), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n411), .SE(n460), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n413), .SE(n458), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n413), .SE(n456), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n413), .SE(n454), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n413), .SE(n452), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n413), .SE(n450), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n413), .SE(n448), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n413), .SE(n446), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n413), .SE(n444), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n413), .SE(n442), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n413), .SE(n440), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n413), .SE(n438), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n412), .SE(n436), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n412), .SE(n434), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n412), .SE(n432), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n412), .SE(n430), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n412), .SE(n428), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n412), .SE(n426), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n412), .SE(n424), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n412), .SE(n422), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n412), .SE(n420), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n412), .SE(n418), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n412), .SE(n416), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n565), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n565), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n360), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n565), .SE(n396), .CK(
        clk), .Q(n341), .QN(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n565), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n358), .QN(n43) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n565), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n357), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n565), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n356), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n565), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n355), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n565), .SE(n386), .CK(
        clk), .Q(n338), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n565), .SE(n384), .CK(
        clk), .Q(n409), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n565), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n565), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n351), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n565), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n350), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n565), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n565), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n348), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n565), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n565), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n346), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n565), .SE(n368), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n565), .SE(n366), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n565), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n565), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n342) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n414), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n339) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n414), .SE(n522), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n31) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n414), .SE(n518), .CK(clk), .Q(n563), 
        .QN(n34) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n414), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n414), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n41) );
  BUF_X1 U2 ( .A(n411), .Z(n413) );
  BUF_X1 U3 ( .A(n411), .Z(n412) );
  BUF_X1 U4 ( .A(n411), .Z(n414) );
  INV_X1 U5 ( .A(n565), .ZN(n411) );
  NAND2_X1 U6 ( .A1(n10), .A2(n7), .ZN(n364) );
  OAI21_X1 U7 ( .B1(n227), .B2(n228), .A(n298), .ZN(n7) );
  MUX2_X1 U8 ( .A(n542), .B(n294), .S(n298), .Z(n450) );
  NAND2_X1 U9 ( .A1(n23), .A2(n22), .ZN(n141) );
  NAND2_X1 U10 ( .A1(n25), .A2(n24), .ZN(n23) );
  INV_X1 U11 ( .A(n298), .ZN(n6) );
  NOR2_X1 U12 ( .A1(n104), .A2(n103), .ZN(n101) );
  NAND2_X1 U13 ( .A1(n15), .A2(n14), .ZN(n222) );
  NAND2_X1 U14 ( .A1(n236), .A2(n16), .ZN(n15) );
  INV_X1 U15 ( .A(rst_n), .ZN(n565) );
  NAND2_X1 U16 ( .A1(n114), .A2(n113), .ZN(n22) );
  OR2_X1 U17 ( .A1(n114), .A2(n113), .ZN(n24) );
  OR2_X1 U18 ( .A1(n56), .A2(n55), .ZN(n86) );
  OR2_X1 U19 ( .A1(n238), .A2(n237), .ZN(n16) );
  NAND2_X1 U20 ( .A1(n238), .A2(n237), .ZN(n14) );
  INV_X1 U21 ( .A(n240), .ZN(n157) );
  NOR2_X1 U22 ( .A1(n35), .A2(n106), .ZN(n85) );
  INV_X1 U23 ( .A(n26), .ZN(n253) );
  INV_X1 U24 ( .A(n45), .ZN(n169) );
  NAND2_X1 U25 ( .A1(n5), .A2(\mult_x_1/n310 ), .ZN(n106) );
  OAI21_X1 U26 ( .B1(n101), .B2(n8), .A(n105), .ZN(n230) );
  INV_X1 U27 ( .A(n102), .ZN(n8) );
  XNOR2_X1 U28 ( .A(n25), .B(n9), .ZN(n102) );
  XNOR2_X1 U29 ( .A(n114), .B(n113), .ZN(n9) );
  NAND2_X1 U30 ( .A1(n83), .A2(n82), .ZN(n25) );
  NAND2_X1 U31 ( .A1(n6), .A2(n343), .ZN(n10) );
  OAI21_X1 U32 ( .B1(n226), .B2(n12), .A(n11), .ZN(n384) );
  NAND2_X1 U33 ( .A1(n6), .A2(n353), .ZN(n11) );
  NAND2_X1 U34 ( .A1(n13), .A2(n298), .ZN(n12) );
  INV_X1 U35 ( .A(n225), .ZN(n13) );
  NAND2_X1 U36 ( .A1(n18), .A2(n17), .ZN(n291) );
  INV_X1 U37 ( .A(n264), .ZN(n17) );
  INV_X1 U38 ( .A(n265), .ZN(n18) );
  XNOR2_X1 U39 ( .A(n236), .B(n19), .ZN(n265) );
  XNOR2_X1 U40 ( .A(n238), .B(n237), .ZN(n19) );
  NAND2_X1 U41 ( .A1(n21), .A2(n20), .ZN(n79) );
  INV_X1 U42 ( .A(n81), .ZN(n20) );
  OAI22_X1 U43 ( .A1(n157), .A2(n77), .B1(n159), .B2(n50), .ZN(n81) );
  INV_X1 U44 ( .A(n80), .ZN(n21) );
  NAND2_X1 U45 ( .A1(n230), .A2(n231), .ZN(n232) );
  XNOR2_X1 U46 ( .A(n203), .B(n202), .ZN(n209) );
  XNOR2_X1 U47 ( .A(n201), .B(n200), .ZN(n202) );
  NAND2_X1 U48 ( .A1(n184), .A2(n183), .ZN(n72) );
  OR2_X1 U49 ( .A1(n184), .A2(n183), .ZN(n71) );
  NAND2_X1 U50 ( .A1(n132), .A2(n131), .ZN(n139) );
  XNOR2_X1 U51 ( .A(n184), .B(n183), .ZN(n186) );
  NAND2_X1 U52 ( .A1(n198), .A2(n197), .ZN(n233) );
  NAND2_X1 U53 ( .A1(n201), .A2(n200), .ZN(n197) );
  NAND2_X1 U54 ( .A1(n203), .A2(n196), .ZN(n198) );
  OR2_X1 U55 ( .A1(n201), .A2(n200), .ZN(n196) );
  XNOR2_X1 U56 ( .A(n54), .B(n78), .ZN(n97) );
  NAND2_X1 U57 ( .A1(n46), .A2(n47), .ZN(n159) );
  XNOR2_X1 U58 ( .A(n41), .B(\mult_x_1/a[2] ), .ZN(n26) );
  XNOR2_X1 U59 ( .A(\mult_x_1/a[4] ), .B(n34), .ZN(n46) );
  INV_X1 U60 ( .A(n31), .ZN(n27) );
  CLKBUF_X1 U61 ( .A(\mult_x_1/n312 ), .Z(n28) );
  XNOR2_X1 U62 ( .A(n41), .B(\mult_x_1/a[2] ), .ZN(n51) );
  XNOR2_X1 U63 ( .A(n81), .B(n29), .ZN(n54) );
  XNOR2_X1 U64 ( .A(\mult_x_1/a[6] ), .B(n34), .ZN(n45) );
  OAI22_X1 U65 ( .A1(n168), .A2(n59), .B1(n169), .B2(n90), .ZN(n29) );
  XOR2_X1 U66 ( .A(n56), .B(n55), .Z(n42) );
  XNOR2_X1 U67 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n44) );
  OR2_X2 U68 ( .A1(n44), .A2(n45), .ZN(n168) );
  XNOR2_X1 U69 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n69) );
  XNOR2_X1 U70 ( .A(n27), .B(\mult_x_1/n286 ), .ZN(n60) );
  OAI22_X1 U71 ( .A1(n168), .A2(n69), .B1(n169), .B2(n60), .ZN(n192) );
  NAND2_X1 U72 ( .A1(\mult_x_1/n313 ), .A2(n30), .ZN(n255) );
  XNOR2_X1 U73 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n150) );
  AND2_X1 U74 ( .A1(n564), .A2(\mult_x_1/n281 ), .ZN(n123) );
  XNOR2_X1 U75 ( .A(n123), .B(\mult_x_1/n313 ), .ZN(n57) );
  OAI22_X1 U76 ( .A1(n255), .A2(n150), .B1(n57), .B2(n30), .ZN(n191) );
  NOR2_X1 U77 ( .A1(n106), .A2(n32), .ZN(n190) );
  INV_X1 U78 ( .A(n62), .ZN(n49) );
  XNOR2_X1 U79 ( .A(n339), .B(n340), .ZN(n47) );
  XNOR2_X1 U80 ( .A(n563), .B(\mult_x_1/n284 ), .ZN(n66) );
  INV_X1 U81 ( .A(n47), .ZN(n240) );
  XNOR2_X1 U82 ( .A(n563), .B(\mult_x_1/n283 ), .ZN(n50) );
  OAI22_X1 U83 ( .A1(n159), .A2(n66), .B1(n47), .B2(n50), .ZN(n56) );
  XNOR2_X1 U84 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n48) );
  OR2_X2 U85 ( .A1(n51), .A2(n48), .ZN(n251) );
  XNOR2_X1 U86 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n67) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n94) );
  OAI22_X1 U88 ( .A1(n251), .A2(n67), .B1(n253), .B2(n94), .ZN(n55) );
  NOR2_X1 U89 ( .A1(n49), .A2(n42), .ZN(n98) );
  XNOR2_X1 U90 ( .A(n563), .B(\mult_x_1/n282 ), .ZN(n77) );
  XNOR2_X1 U91 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n59) );
  XNOR2_X1 U92 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n90) );
  OAI22_X1 U93 ( .A1(n168), .A2(n59), .B1(n169), .B2(n90), .ZN(n80) );
  XNOR2_X1 U94 ( .A(n123), .B(\mult_x_1/n312 ), .ZN(n91) );
  INV_X1 U95 ( .A(n91), .ZN(n52) );
  NAND2_X1 U96 ( .A1(n52), .A2(n26), .ZN(n93) );
  OAI21_X1 U97 ( .B1(n251), .B2(n94), .A(n93), .ZN(n53) );
  INV_X1 U98 ( .A(n53), .ZN(n78) );
  XNOR2_X1 U99 ( .A(n86), .B(n85), .ZN(n61) );
  AOI21_X1 U100 ( .B1(n255), .B2(n30), .A(n57), .ZN(n58) );
  INV_X1 U101 ( .A(n58), .ZN(n65) );
  OAI22_X1 U102 ( .A1(n168), .A2(n60), .B1(n169), .B2(n59), .ZN(n64) );
  NOR2_X1 U103 ( .A1(n36), .A2(n106), .ZN(n63) );
  XNOR2_X1 U104 ( .A(n61), .B(n84), .ZN(n96) );
  XNOR2_X1 U105 ( .A(n62), .B(n42), .ZN(n185) );
  FA_X1 U106 ( .A(n65), .B(n64), .CI(n63), .CO(n84), .S(n184) );
  XNOR2_X1 U107 ( .A(n563), .B(\mult_x_1/n285 ), .ZN(n149) );
  OAI22_X1 U108 ( .A1(n159), .A2(n149), .B1(n157), .B2(n66), .ZN(n189) );
  XNOR2_X1 U109 ( .A(n28), .B(\mult_x_1/n283 ), .ZN(n152) );
  OAI22_X1 U110 ( .A1(n251), .A2(n152), .B1(n253), .B2(n67), .ZN(n188) );
  OR2_X1 U111 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n68) );
  OAI22_X1 U112 ( .A1(n168), .A2(n31), .B1(n68), .B2(n169), .ZN(n148) );
  XNOR2_X1 U113 ( .A(n27), .B(\mult_x_1/n288 ), .ZN(n70) );
  OAI22_X1 U114 ( .A1(n168), .A2(n70), .B1(n169), .B2(n69), .ZN(n147) );
  NAND2_X1 U115 ( .A1(n185), .A2(n71), .ZN(n73) );
  NAND2_X1 U116 ( .A1(n73), .A2(n72), .ZN(n225) );
  NAND2_X1 U117 ( .A1(n226), .A2(n225), .ZN(n74) );
  BUF_X4 U118 ( .A(en), .Z(n298) );
  NAND2_X1 U119 ( .A1(n74), .A2(n298), .ZN(n76) );
  OR2_X1 U120 ( .A1(n298), .A2(n338), .ZN(n75) );
  NAND2_X1 U121 ( .A1(n76), .A2(n75), .ZN(n386) );
  NOR2_X1 U122 ( .A1(n37), .A2(n106), .ZN(n114) );
  XNOR2_X1 U123 ( .A(n563), .B(\mult_x_1/n281 ), .ZN(n108) );
  OAI22_X1 U124 ( .A1(n159), .A2(n77), .B1(n157), .B2(n108), .ZN(n113) );
  NAND2_X1 U125 ( .A1(n79), .A2(n78), .ZN(n83) );
  NAND2_X1 U126 ( .A1(n81), .A2(n80), .ZN(n82) );
  NAND2_X1 U127 ( .A1(n86), .A2(n85), .ZN(n89) );
  INV_X1 U128 ( .A(n84), .ZN(n88) );
  NOR2_X1 U129 ( .A1(n86), .A2(n85), .ZN(n87) );
  AOI21_X2 U130 ( .B1(n89), .B2(n88), .A(n87), .ZN(n104) );
  XNOR2_X1 U131 ( .A(n27), .B(\mult_x_1/n283 ), .ZN(n107) );
  OAI22_X1 U132 ( .A1(n168), .A2(n90), .B1(n169), .B2(n107), .ZN(n112) );
  AOI21_X1 U133 ( .B1(n253), .B2(n251), .A(n91), .ZN(n92) );
  INV_X1 U134 ( .A(n92), .ZN(n111) );
  OAI21_X1 U135 ( .B1(n251), .B2(n94), .A(n93), .ZN(n110) );
  XNOR2_X1 U136 ( .A(n104), .B(n103), .ZN(n95) );
  XNOR2_X1 U137 ( .A(n102), .B(n95), .ZN(n119) );
  FA_X1 U138 ( .A(n98), .B(n97), .CI(n96), .CO(n118), .S(n226) );
  INV_X1 U139 ( .A(n118), .ZN(n99) );
  NAND2_X1 U140 ( .A1(n298), .A2(n99), .ZN(n100) );
  OAI22_X1 U141 ( .A1(n119), .A2(n100), .B1(n298), .B2(n341), .ZN(n396) );
  NAND2_X1 U142 ( .A1(n104), .A2(n103), .ZN(n105) );
  NOR2_X1 U143 ( .A1(n38), .A2(n106), .ZN(n128) );
  XNOR2_X1 U144 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n125) );
  OAI22_X1 U145 ( .A1(n168), .A2(n107), .B1(n169), .B2(n125), .ZN(n129) );
  XNOR2_X1 U146 ( .A(n128), .B(n129), .ZN(n109) );
  XNOR2_X1 U147 ( .A(n123), .B(n563), .ZN(n126) );
  OAI22_X1 U148 ( .A1(n159), .A2(n108), .B1(n126), .B2(n157), .ZN(n134) );
  INV_X1 U149 ( .A(n134), .ZN(n130) );
  XNOR2_X1 U150 ( .A(n109), .B(n130), .ZN(n143) );
  FA_X1 U151 ( .A(n112), .B(n111), .CI(n110), .CO(n142), .S(n103) );
  XNOR2_X1 U152 ( .A(n143), .B(n142), .ZN(n115) );
  XNOR2_X1 U153 ( .A(n115), .B(n141), .ZN(n231) );
  OAI21_X1 U154 ( .B1(n230), .B2(n231), .A(n298), .ZN(n117) );
  OR2_X1 U155 ( .A1(n298), .A2(n43), .ZN(n116) );
  NAND2_X1 U156 ( .A1(n117), .A2(n116), .ZN(n394) );
  NAND2_X1 U157 ( .A1(n119), .A2(n118), .ZN(n120) );
  NAND2_X1 U158 ( .A1(n120), .A2(n298), .ZN(n122) );
  OR2_X1 U159 ( .A1(n298), .A2(n403), .ZN(n121) );
  NAND2_X1 U160 ( .A1(n122), .A2(n121), .ZN(n398) );
  NOR2_X1 U181 ( .A1(n39), .A2(n106), .ZN(n166) );
  XNOR2_X1 U182 ( .A(n27), .B(\mult_x_1/n281 ), .ZN(n124) );
  XNOR2_X1 U183 ( .A(n123), .B(n27), .ZN(n167) );
  OAI22_X1 U184 ( .A1(n168), .A2(n124), .B1(n167), .B2(n169), .ZN(n174) );
  INV_X1 U185 ( .A(n174), .ZN(n165) );
  OAI22_X1 U186 ( .A1(n168), .A2(n125), .B1(n169), .B2(n124), .ZN(n135) );
  AOI21_X1 U187 ( .B1(n157), .B2(n159), .A(n126), .ZN(n127) );
  INV_X1 U188 ( .A(n127), .ZN(n133) );
  OAI21_X1 U189 ( .B1(n130), .B2(n129), .A(n128), .ZN(n132) );
  NAND2_X1 U190 ( .A1(n130), .A2(n129), .ZN(n131) );
  NOR2_X1 U191 ( .A1(n40), .A2(n106), .ZN(n138) );
  FA_X1 U192 ( .A(n135), .B(n134), .CI(n133), .CO(n164), .S(n137) );
  OR2_X1 U193 ( .A1(n181), .A2(n180), .ZN(n136) );
  MUX2_X1 U194 ( .A(n342), .B(n136), .S(n298), .Z(n362) );
  FA_X1 U195 ( .A(n139), .B(n138), .CI(n137), .CO(n180), .S(n228) );
  OR2_X1 U196 ( .A1(n143), .A2(n142), .ZN(n140) );
  NAND2_X1 U197 ( .A1(n141), .A2(n140), .ZN(n145) );
  NAND2_X1 U198 ( .A1(n143), .A2(n142), .ZN(n144) );
  NAND2_X1 U199 ( .A1(n145), .A2(n144), .ZN(n227) );
  XNOR2_X1 U200 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n218) );
  XNOR2_X1 U201 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n151) );
  OAI22_X1 U202 ( .A1(n255), .A2(n218), .B1(n151), .B2(n30), .ZN(n162) );
  INV_X1 U203 ( .A(n169), .ZN(n146) );
  AND2_X1 U204 ( .A1(\mult_x_1/n288 ), .A2(n146), .ZN(n161) );
  XNOR2_X1 U205 ( .A(n28), .B(\mult_x_1/n285 ), .ZN(n217) );
  XNOR2_X1 U206 ( .A(n28), .B(\mult_x_1/n284 ), .ZN(n153) );
  OAI22_X1 U207 ( .A1(n251), .A2(n217), .B1(n253), .B2(n153), .ZN(n160) );
  HA_X1 U208 ( .A(n147), .B(n148), .CO(n187), .S(n205) );
  XNOR2_X1 U209 ( .A(n563), .B(\mult_x_1/n286 ), .ZN(n156) );
  OAI22_X1 U210 ( .A1(n159), .A2(n156), .B1(n157), .B2(n149), .ZN(n195) );
  OAI22_X1 U211 ( .A1(n255), .A2(n151), .B1(n150), .B2(n30), .ZN(n194) );
  OAI22_X1 U212 ( .A1(n251), .A2(n153), .B1(n253), .B2(n152), .ZN(n193) );
  OR2_X1 U213 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n154) );
  OAI22_X1 U214 ( .A1(n159), .A2(n34), .B1(n154), .B2(n157), .ZN(n220) );
  XNOR2_X1 U215 ( .A(n563), .B(\mult_x_1/n288 ), .ZN(n155) );
  XNOR2_X1 U216 ( .A(n563), .B(\mult_x_1/n287 ), .ZN(n158) );
  OAI22_X1 U217 ( .A1(n159), .A2(n155), .B1(n157), .B2(n158), .ZN(n219) );
  OAI22_X1 U218 ( .A1(n159), .A2(n158), .B1(n157), .B2(n156), .ZN(n215) );
  FA_X1 U219 ( .A(n162), .B(n161), .CI(n160), .CO(n206), .S(n214) );
  OR2_X1 U220 ( .A1(n212), .A2(n211), .ZN(n163) );
  MUX2_X1 U221 ( .A(n344), .B(n163), .S(n298), .Z(n366) );
  FA_X1 U222 ( .A(n166), .B(n165), .CI(n164), .CO(n176), .S(n181) );
  AOI21_X1 U223 ( .B1(n169), .B2(n168), .A(n167), .ZN(n170) );
  INV_X1 U224 ( .A(n170), .ZN(n172) );
  NOR2_X1 U225 ( .A1(n33), .A2(n106), .ZN(n171) );
  XOR2_X1 U226 ( .A(n172), .B(n171), .Z(n173) );
  XOR2_X1 U227 ( .A(n174), .B(n173), .Z(n175) );
  OR2_X1 U228 ( .A1(n176), .A2(n175), .ZN(n178) );
  NAND2_X1 U229 ( .A1(n176), .A2(n175), .ZN(n177) );
  NAND2_X1 U230 ( .A1(n178), .A2(n177), .ZN(n179) );
  MUX2_X1 U231 ( .A(n345), .B(n179), .S(n298), .Z(n368) );
  NAND2_X1 U232 ( .A1(n181), .A2(n180), .ZN(n182) );
  MUX2_X1 U233 ( .A(n346), .B(n182), .S(n298), .Z(n370) );
  XNOR2_X1 U234 ( .A(n186), .B(n185), .ZN(n234) );
  FA_X1 U235 ( .A(n189), .B(n188), .CI(n187), .CO(n183), .S(n203) );
  FA_X1 U236 ( .A(n192), .B(n191), .CI(n190), .CO(n62), .S(n201) );
  FA_X1 U237 ( .A(n195), .B(n194), .CI(n193), .CO(n200), .S(n204) );
  NAND2_X1 U238 ( .A1(n234), .A2(n233), .ZN(n199) );
  MUX2_X1 U239 ( .A(n347), .B(n199), .S(n298), .Z(n372) );
  FA_X1 U240 ( .A(n206), .B(n205), .CI(n204), .CO(n208), .S(n212) );
  NOR2_X1 U241 ( .A1(n209), .A2(n208), .ZN(n207) );
  MUX2_X1 U242 ( .A(n348), .B(n207), .S(n298), .Z(n374) );
  NAND2_X1 U243 ( .A1(n209), .A2(n208), .ZN(n210) );
  MUX2_X1 U244 ( .A(n349), .B(n210), .S(n298), .Z(n376) );
  NAND2_X1 U245 ( .A1(n212), .A2(n211), .ZN(n213) );
  MUX2_X1 U246 ( .A(n350), .B(n213), .S(n298), .Z(n378) );
  FA_X1 U247 ( .A(n216), .B(n215), .CI(n214), .CO(n211), .S(n223) );
  XNOR2_X1 U248 ( .A(n28), .B(\mult_x_1/n286 ), .ZN(n241) );
  OAI22_X1 U249 ( .A1(n251), .A2(n241), .B1(n253), .B2(n217), .ZN(n238) );
  XNOR2_X1 U250 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n239) );
  OAI22_X1 U251 ( .A1(n255), .A2(n239), .B1(n218), .B2(n30), .ZN(n237) );
  HA_X1 U252 ( .A(n220), .B(n219), .CO(n216), .S(n236) );
  NOR2_X1 U253 ( .A1(n223), .A2(n222), .ZN(n221) );
  MUX2_X1 U254 ( .A(n351), .B(n221), .S(n298), .Z(n380) );
  NAND2_X1 U255 ( .A1(n223), .A2(n222), .ZN(n224) );
  MUX2_X1 U256 ( .A(n352), .B(n224), .S(n298), .Z(n382) );
  NAND2_X1 U257 ( .A1(n228), .A2(n227), .ZN(n229) );
  MUX2_X1 U258 ( .A(n355), .B(n229), .S(n298), .Z(n388) );
  MUX2_X1 U259 ( .A(n356), .B(n232), .S(n298), .Z(n390) );
  NOR2_X1 U260 ( .A1(n234), .A2(n233), .ZN(n235) );
  MUX2_X1 U261 ( .A(n357), .B(n235), .S(n298), .Z(n392) );
  XNOR2_X1 U262 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n247) );
  OAI22_X1 U263 ( .A1(n255), .A2(n247), .B1(n239), .B2(n30), .ZN(n244) );
  AND2_X1 U264 ( .A1(n240), .A2(\mult_x_1/n288 ), .ZN(n243) );
  XNOR2_X1 U265 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n245) );
  OAI22_X1 U266 ( .A1(n251), .A2(n245), .B1(n253), .B2(n241), .ZN(n242) );
  FA_X1 U267 ( .A(n244), .B(n243), .CI(n242), .CO(n264), .S(n263) );
  XNOR2_X1 U268 ( .A(n28), .B(\mult_x_1/n288 ), .ZN(n246) );
  OAI22_X1 U269 ( .A1(n251), .A2(n246), .B1(n253), .B2(n245), .ZN(n249) );
  XNOR2_X1 U270 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n252) );
  OAI22_X1 U271 ( .A1(n255), .A2(n252), .B1(n247), .B2(n30), .ZN(n248) );
  NOR2_X1 U272 ( .A1(n263), .A2(n262), .ZN(n284) );
  HA_X1 U273 ( .A(n249), .B(n248), .CO(n262), .S(n260) );
  OR2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(n339), .ZN(n250) );
  OAI22_X1 U275 ( .A1(n251), .A2(n339), .B1(n250), .B2(n253), .ZN(n259) );
  OR2_X1 U276 ( .A1(n260), .A2(n259), .ZN(n280) );
  XNOR2_X1 U277 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n254) );
  OAI22_X1 U278 ( .A1(n255), .A2(n254), .B1(n252), .B2(n30), .ZN(n258) );
  AND2_X1 U279 ( .A1(\mult_x_1/n288 ), .A2(n51), .ZN(n257) );
  NOR2_X1 U280 ( .A1(n258), .A2(n257), .ZN(n273) );
  OAI22_X1 U281 ( .A1(n255), .A2(\mult_x_1/n288 ), .B1(n254), .B2(n30), .ZN(
        n270) );
  OR2_X1 U282 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n256) );
  NAND2_X1 U283 ( .A1(n256), .A2(n255), .ZN(n269) );
  NAND2_X1 U284 ( .A1(n270), .A2(n269), .ZN(n276) );
  NAND2_X1 U285 ( .A1(n258), .A2(n257), .ZN(n274) );
  OAI21_X1 U286 ( .B1(n273), .B2(n276), .A(n274), .ZN(n281) );
  NAND2_X1 U287 ( .A1(n260), .A2(n259), .ZN(n279) );
  INV_X1 U288 ( .A(n279), .ZN(n261) );
  AOI21_X1 U289 ( .B1(n280), .B2(n281), .A(n261), .ZN(n287) );
  NAND2_X1 U290 ( .A1(n263), .A2(n262), .ZN(n285) );
  OAI21_X1 U291 ( .B1(n284), .B2(n287), .A(n285), .ZN(n292) );
  NAND2_X1 U292 ( .A1(n265), .A2(n264), .ZN(n290) );
  INV_X1 U293 ( .A(n290), .ZN(n266) );
  AOI21_X1 U294 ( .B1(n291), .B2(n292), .A(n266), .ZN(n267) );
  MUX2_X1 U295 ( .A(n361), .B(n267), .S(n298), .Z(n400) );
  MUX2_X1 U296 ( .A(product[0]), .B(n526), .S(n298), .Z(n416) );
  MUX2_X1 U297 ( .A(n526), .B(n527), .S(n298), .Z(n418) );
  AND2_X1 U298 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n268) );
  MUX2_X1 U299 ( .A(n527), .B(n268), .S(n298), .Z(n420) );
  MUX2_X1 U300 ( .A(product[1]), .B(n529), .S(n298), .Z(n422) );
  MUX2_X1 U301 ( .A(n529), .B(n530), .S(n298), .Z(n424) );
  OR2_X1 U302 ( .A1(n270), .A2(n269), .ZN(n271) );
  AND2_X1 U303 ( .A1(n271), .A2(n276), .ZN(n272) );
  MUX2_X1 U304 ( .A(n530), .B(n272), .S(n298), .Z(n426) );
  MUX2_X1 U305 ( .A(product[2]), .B(n532), .S(n298), .Z(n428) );
  MUX2_X1 U306 ( .A(n532), .B(n533), .S(n298), .Z(n430) );
  INV_X1 U307 ( .A(n273), .ZN(n275) );
  NAND2_X1 U308 ( .A1(n275), .A2(n274), .ZN(n277) );
  XOR2_X1 U309 ( .A(n277), .B(n276), .Z(n278) );
  MUX2_X1 U310 ( .A(n533), .B(n278), .S(n298), .Z(n432) );
  MUX2_X1 U311 ( .A(product[3]), .B(n535), .S(n298), .Z(n434) );
  MUX2_X1 U312 ( .A(n535), .B(n536), .S(n298), .Z(n436) );
  NAND2_X1 U313 ( .A1(n280), .A2(n279), .ZN(n282) );
  XNOR2_X1 U314 ( .A(n282), .B(n281), .ZN(n283) );
  MUX2_X1 U315 ( .A(n536), .B(n283), .S(n298), .Z(n438) );
  MUX2_X1 U316 ( .A(product[4]), .B(n538), .S(n298), .Z(n440) );
  MUX2_X1 U317 ( .A(n538), .B(n539), .S(n298), .Z(n442) );
  INV_X1 U318 ( .A(n284), .ZN(n286) );
  NAND2_X1 U319 ( .A1(n286), .A2(n285), .ZN(n288) );
  XOR2_X1 U320 ( .A(n288), .B(n287), .Z(n289) );
  MUX2_X1 U321 ( .A(n539), .B(n289), .S(n298), .Z(n444) );
  MUX2_X1 U322 ( .A(product[5]), .B(n541), .S(n298), .Z(n446) );
  MUX2_X1 U323 ( .A(n541), .B(n542), .S(n298), .Z(n448) );
  NAND2_X1 U324 ( .A1(n291), .A2(n290), .ZN(n293) );
  XNOR2_X1 U325 ( .A(n293), .B(n292), .ZN(n294) );
  MUX2_X1 U326 ( .A(product[6]), .B(n544), .S(n298), .Z(n452) );
  NAND2_X1 U327 ( .A1(n404), .A2(n352), .ZN(n295) );
  XOR2_X1 U328 ( .A(n295), .B(n361), .Z(n296) );
  MUX2_X1 U329 ( .A(n544), .B(n296), .S(n298), .Z(n454) );
  MUX2_X1 U330 ( .A(product[7]), .B(n546), .S(n298), .Z(n456) );
  OAI21_X1 U331 ( .B1(n351), .B2(n361), .A(n352), .ZN(n300) );
  NAND2_X1 U332 ( .A1(n344), .A2(n350), .ZN(n297) );
  XNOR2_X1 U333 ( .A(n300), .B(n297), .ZN(n299) );
  MUX2_X1 U334 ( .A(n546), .B(n299), .S(n298), .Z(n458) );
  BUF_X2 U335 ( .A(en), .Z(n337) );
  MUX2_X1 U336 ( .A(product[8]), .B(n548), .S(n337), .Z(n460) );
  AOI21_X1 U337 ( .B1(n300), .B2(n344), .A(n406), .ZN(n303) );
  NAND2_X1 U338 ( .A1(n407), .A2(n349), .ZN(n301) );
  XOR2_X1 U339 ( .A(n303), .B(n301), .Z(n302) );
  MUX2_X1 U340 ( .A(n548), .B(n302), .S(n337), .Z(n462) );
  MUX2_X1 U341 ( .A(product[9]), .B(n550), .S(n337), .Z(n464) );
  OAI21_X1 U342 ( .B1(n303), .B2(n348), .A(n349), .ZN(n311) );
  INV_X1 U343 ( .A(n311), .ZN(n306) );
  NAND2_X1 U344 ( .A1(n408), .A2(n347), .ZN(n304) );
  XOR2_X1 U345 ( .A(n306), .B(n304), .Z(n305) );
  MUX2_X1 U346 ( .A(n550), .B(n305), .S(n337), .Z(n466) );
  MUX2_X1 U347 ( .A(product[10]), .B(n552), .S(n337), .Z(n468) );
  OAI21_X1 U348 ( .B1(n306), .B2(n357), .A(n347), .ZN(n308) );
  NAND2_X1 U349 ( .A1(n409), .A2(n354), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U351 ( .A(n552), .B(n309), .S(n337), .Z(n470) );
  MUX2_X1 U352 ( .A(product[11]), .B(n554), .S(n337), .Z(n472) );
  NOR2_X1 U353 ( .A1(n353), .A2(n357), .ZN(n312) );
  OAI21_X1 U354 ( .B1(n353), .B2(n347), .A(n354), .ZN(n310) );
  AOI21_X1 U355 ( .B1(n312), .B2(n311), .A(n310), .ZN(n334) );
  NAND2_X1 U356 ( .A1(n341), .A2(n360), .ZN(n313) );
  XOR2_X1 U357 ( .A(n334), .B(n313), .Z(n314) );
  MUX2_X1 U358 ( .A(n554), .B(n314), .S(n337), .Z(n474) );
  MUX2_X1 U359 ( .A(product[12]), .B(n556), .S(n337), .Z(n476) );
  OAI21_X1 U360 ( .B1(n334), .B2(n359), .A(n360), .ZN(n316) );
  NAND2_X1 U361 ( .A1(n358), .A2(n356), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  MUX2_X1 U363 ( .A(n556), .B(n317), .S(n337), .Z(n478) );
  MUX2_X1 U364 ( .A(product[13]), .B(n558), .S(n337), .Z(n480) );
  NAND2_X1 U365 ( .A1(n341), .A2(n358), .ZN(n319) );
  AOI21_X1 U366 ( .B1(n403), .B2(n358), .A(n410), .ZN(n318) );
  OAI21_X1 U367 ( .B1(n334), .B2(n319), .A(n318), .ZN(n321) );
  NAND2_X1 U368 ( .A1(n343), .A2(n355), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  MUX2_X1 U370 ( .A(n558), .B(n322), .S(n337), .Z(n482) );
  MUX2_X1 U371 ( .A(product[14]), .B(n560), .S(n337), .Z(n484) );
  NAND2_X1 U372 ( .A1(n358), .A2(n343), .ZN(n324) );
  NOR2_X1 U373 ( .A1(n359), .A2(n324), .ZN(n330) );
  INV_X1 U374 ( .A(n330), .ZN(n326) );
  AOI21_X1 U375 ( .B1(n410), .B2(n343), .A(n405), .ZN(n323) );
  OAI21_X1 U376 ( .B1(n324), .B2(n360), .A(n323), .ZN(n331) );
  INV_X1 U377 ( .A(n331), .ZN(n325) );
  OAI21_X1 U378 ( .B1(n334), .B2(n326), .A(n325), .ZN(n328) );
  NAND2_X1 U379 ( .A1(n342), .A2(n346), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  MUX2_X1 U381 ( .A(n560), .B(n329), .S(n337), .Z(n486) );
  MUX2_X1 U382 ( .A(product[15]), .B(n562), .S(n337), .Z(n488) );
  NAND2_X1 U383 ( .A1(n330), .A2(n342), .ZN(n333) );
  AOI21_X1 U384 ( .B1(n331), .B2(n342), .A(n402), .ZN(n332) );
  OAI21_X1 U385 ( .B1(n334), .B2(n333), .A(n332), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n335), .B(n345), .ZN(n336) );
  MUX2_X1 U387 ( .A(n562), .B(n336), .S(n337), .Z(n490) );
  MUX2_X1 U388 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n337), .Z(n492) );
  MUX2_X1 U389 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n337), .Z(n494) );
  MUX2_X1 U390 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n337), .Z(n496) );
  MUX2_X1 U391 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n337), .Z(n498) );
  MUX2_X1 U392 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n337), .Z(n500) );
  MUX2_X1 U393 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n337), .Z(n502) );
  MUX2_X1 U394 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n337), .Z(n504) );
  MUX2_X1 U395 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n337), .Z(n506) );
  MUX2_X1 U396 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n337), .Z(n508) );
  MUX2_X1 U397 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n337), .Z(n510) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n337), .Z(n512) );
  MUX2_X1 U399 ( .A(n28), .B(A_extended[3]), .S(n337), .Z(n514) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n337), .Z(n516) );
  MUX2_X1 U401 ( .A(n563), .B(A_extended[5]), .S(n337), .Z(n518) );
  MUX2_X1 U402 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n337), .Z(n520) );
  MUX2_X1 U403 ( .A(n27), .B(A_extended[7]), .S(n337), .Z(n522) );
  OR2_X1 U404 ( .A1(n337), .A2(n564), .ZN(n524) );
endmodule


module conv_128_32_DW_mult_pipe_J1_8 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n348,
         n350, n352, n354, n356, n358, n360, n362, n364, n366, n368, n370,
         n372, n374, n376, n378, n380, n382, n384, n386, n388, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n400, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n420, n422, n424, n426, n428,
         n430, n432, n434, n436, n438, n440, n442, n444, n446, n448, n450,
         n452, n454, n456, n458, n460, n462, n464, n466, n468, n470, n472,
         n474, n476, n478, n480, n482, n484, n486, n488, n490, n492, n494,
         n496, n498, n500, n502, n504, n506, n508, n509, n511, n512, n514,
         n515, n517, n518, n520, n521, n523, n525, n527, n529, n531, n533,
         n535, n537, n539, n541, n543, n544, n545, n546;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n398), .SE(n506), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n398), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n37) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n398), .SE(n494), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n35) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n398), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n23) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n398), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n28) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n398), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n32) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n396), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n30) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n397), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n29) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n396), .SE(n480), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n31) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n398), .SE(n478), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n33) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n396), .SE(n476), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n34) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n396), .SE(n474), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n396), .SE(n472), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n396), .SE(n470), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n396), .SE(n468), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n396), .SE(n466), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n396), .SE(n464), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n397), .SE(n462), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n398), .SE(n460), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n396), .SE(n458), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n396), .SE(n456), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n396), .SE(n454), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n396), .SE(n452), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n396), .SE(n450), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n396), .SE(n448), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n396), .SE(n446), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n396), .SE(n444), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n397), .SE(n442), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n397), .SE(n440), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n397), .SE(n438), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n397), .SE(n436), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n397), .SE(n434), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n397), .SE(n432), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n397), .SE(n430), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n397), .SE(n428), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n397), .SE(n426), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n397), .SE(n424), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n397), .SE(n422), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n396), .SE(n420), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n396), .SE(n418), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n396), .SE(n416), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n396), .SE(n414), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n396), .SE(n412), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n396), .SE(n410), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n396), .SE(n408), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n396), .SE(n406), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n396), .SE(n404), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n396), .SE(n402), .CK(clk), .Q(n508)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n396), .SE(n400), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n398), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n36) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n546), .SE(n388), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2_IP  ( .D(1'b1), .SI(n546), .SE(n386), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n546), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n546), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n546), .SE(n380), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n546), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n546), .SE(n376), .CK(
        clk), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n546), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n546), .SE(n372), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n546), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n336), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n546), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n335), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n546), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n546), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n333), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n546), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n332), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n546), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n546), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n330), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n546), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n329), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n546), .SE(n354), .CK(
        clk), .QN(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n546), .SE(n352), .CK(
        clk), .QN(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n546), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n546), .SI(1'b1), .SE(n348), .CK(clk), 
        .Q(n325) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n546), .SE(n346), .CK(
        clk), .QN(n324) );
  SDFF_X2 clk_r_REG51_S1 ( .D(1'b0), .SI(n398), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n26) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n398), .SE(n500), .CK(clk), .Q(n544), 
        .QN(n27) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n398), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n25) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n398), .SE(n498), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n20) );
  BUF_X1 U2 ( .A(en), .Z(n264) );
  BUF_X1 U3 ( .A(en), .Z(n266) );
  XOR2_X2 U4 ( .A(n39), .B(n25), .Z(n62) );
  INV_X1 U5 ( .A(n93), .ZN(n242) );
  BUF_X1 U6 ( .A(n396), .Z(n397) );
  INV_X2 U7 ( .A(n546), .ZN(n396) );
  NAND2_X1 U8 ( .A1(n12), .A2(n11), .ZN(n236) );
  NAND2_X1 U9 ( .A1(n8), .A2(n7), .ZN(n222) );
  NAND2_X1 U10 ( .A1(n13), .A2(n147), .ZN(n12) );
  BUF_X1 U11 ( .A(n396), .Z(n398) );
  OAI21_X1 U12 ( .B1(n230), .B2(n229), .A(n10), .ZN(n8) );
  NOR2_X1 U13 ( .A1(n198), .A2(n197), .ZN(n260) );
  NAND2_X1 U14 ( .A1(n230), .A2(n229), .ZN(n7) );
  NAND2_X1 U15 ( .A1(n15), .A2(n14), .ZN(n13) );
  INV_X1 U16 ( .A(rst_n), .ZN(n546) );
  NAND2_X1 U17 ( .A1(n149), .A2(n148), .ZN(n11) );
  INV_X1 U18 ( .A(n148), .ZN(n14) );
  INV_X1 U19 ( .A(n149), .ZN(n15) );
  INV_X1 U20 ( .A(n50), .ZN(n188) );
  INV_X1 U21 ( .A(n27), .ZN(n22) );
  NAND2_X1 U22 ( .A1(n41), .A2(n42), .ZN(n126) );
  CLKBUF_X1 U23 ( .A(\mult_x_1/n313 ), .Z(n17) );
  XNOR2_X1 U24 ( .A(n5), .B(n262), .ZN(n263) );
  NOR2_X1 U25 ( .A1(n260), .A2(n6), .ZN(n5) );
  INV_X1 U26 ( .A(n261), .ZN(n6) );
  INV_X1 U27 ( .A(n46), .ZN(n47) );
  XNOR2_X1 U28 ( .A(n26), .B(n20), .ZN(n46) );
  XNOR2_X1 U29 ( .A(n9), .B(n230), .ZN(n232) );
  XNOR2_X1 U30 ( .A(n10), .B(n229), .ZN(n9) );
  NAND2_X1 U31 ( .A1(n211), .A2(n210), .ZN(n10) );
  XNOR2_X1 U32 ( .A(n16), .B(n147), .ZN(n239) );
  XNOR2_X1 U33 ( .A(n149), .B(n148), .ZN(n16) );
  AND2_X1 U34 ( .A1(n545), .A2(\mult_x_1/n310 ), .ZN(n39) );
  XNOR2_X1 U35 ( .A(n44), .B(n209), .ZN(n237) );
  XNOR2_X1 U36 ( .A(n207), .B(n208), .ZN(n44) );
  INV_X1 U37 ( .A(n226), .ZN(n18) );
  INV_X1 U38 ( .A(n25), .ZN(n19) );
  XNOR2_X1 U39 ( .A(\mult_x_1/n312 ), .B(n35), .ZN(n48) );
  OAI22_X1 U40 ( .A1(n117), .A2(n76), .B1(n64), .B2(n115), .ZN(n21) );
  AND2_X1 U41 ( .A1(n225), .A2(n224), .ZN(n24) );
  XOR2_X1 U42 ( .A(n206), .B(n205), .Z(n38) );
  INV_X1 U43 ( .A(n43), .ZN(n127) );
  NOR2_X1 U44 ( .A1(n62), .A2(n34), .ZN(n207) );
  BUF_X1 U45 ( .A(\mult_x_1/n313 ), .Z(n181) );
  NAND2_X1 U46 ( .A1(n181), .A2(n23), .ZN(n190) );
  AND2_X1 U47 ( .A1(n545), .A2(\mult_x_1/n281 ), .ZN(n94) );
  XNOR2_X1 U48 ( .A(n94), .B(n181), .ZN(n57) );
  AOI21_X1 U49 ( .B1(n190), .B2(n23), .A(n57), .ZN(n40) );
  INV_X1 U50 ( .A(n40), .ZN(n208) );
  XNOR2_X1 U51 ( .A(\mult_x_1/n310 ), .B(n37), .ZN(n41) );
  XNOR2_X1 U52 ( .A(\mult_x_1/a[6] ), .B(n544), .ZN(n42) );
  XNOR2_X1 U53 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n55) );
  INV_X1 U54 ( .A(n42), .ZN(n43) );
  XNOR2_X1 U55 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n74) );
  OAI22_X1 U56 ( .A1(n126), .A2(n55), .B1(n42), .B2(n74), .ZN(n209) );
  XOR2_X1 U57 ( .A(\mult_x_1/a[4] ), .B(n544), .Z(n45) );
  NAND2_X1 U58 ( .A1(n45), .A2(n46), .ZN(n117) );
  XNOR2_X1 U59 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n107) );
  INV_X2 U60 ( .A(n47), .ZN(n115) );
  XNOR2_X1 U61 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n53) );
  OAI22_X1 U62 ( .A1(n117), .A2(n107), .B1(n115), .B2(n53), .ZN(n149) );
  XNOR2_X1 U63 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n49) );
  NAND2_X2 U64 ( .A1(n49), .A2(n48), .ZN(n186) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n110) );
  INV_X1 U66 ( .A(n49), .ZN(n50) );
  XNOR2_X1 U67 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n54) );
  OAI22_X1 U68 ( .A1(n186), .A2(n110), .B1(n188), .B2(n54), .ZN(n148) );
  OR2_X1 U69 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n51) );
  OAI22_X1 U70 ( .A1(n126), .A2(n25), .B1(n51), .B2(n127), .ZN(n106) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n52) );
  XNOR2_X1 U72 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n56) );
  OAI22_X1 U73 ( .A1(n126), .A2(n52), .B1(n127), .B2(n56), .ZN(n105) );
  XNOR2_X1 U74 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n75) );
  OAI22_X1 U75 ( .A1(n117), .A2(n53), .B1(n115), .B2(n75), .ZN(n206) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n67) );
  OAI22_X1 U77 ( .A1(n186), .A2(n54), .B1(n188), .B2(n67), .ZN(n205) );
  OAI22_X1 U78 ( .A1(n126), .A2(n56), .B1(n127), .B2(n55), .ZN(n143) );
  XNOR2_X1 U79 ( .A(n181), .B(\mult_x_1/n281 ), .ZN(n108) );
  OAI22_X1 U80 ( .A1(n190), .A2(n108), .B1(n57), .B2(n23), .ZN(n142) );
  INV_X1 U81 ( .A(n62), .ZN(n58) );
  AND2_X1 U82 ( .A1(\mult_x_1/n288 ), .A2(n58), .ZN(n141) );
  XNOR2_X1 U83 ( .A(n38), .B(n225), .ZN(n235) );
  INV_X1 U84 ( .A(en), .ZN(n93) );
  NAND2_X1 U85 ( .A1(n59), .A2(n242), .ZN(n61) );
  NAND2_X1 U86 ( .A1(n93), .A2(n344), .ZN(n60) );
  NAND2_X1 U87 ( .A1(n61), .A2(n60), .ZN(n386) );
  NOR2_X1 U88 ( .A1(n29), .A2(n62), .ZN(n72) );
  XNOR2_X1 U89 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n66) );
  XNOR2_X1 U90 ( .A(n19), .B(\mult_x_1/n282 ), .ZN(n63) );
  OAI22_X1 U91 ( .A1(n126), .A2(n66), .B1(n127), .B2(n63), .ZN(n71) );
  XNOR2_X1 U92 ( .A(n22), .B(\mult_x_1/n281 ), .ZN(n76) );
  XNOR2_X1 U93 ( .A(n94), .B(n22), .ZN(n64) );
  OAI22_X1 U94 ( .A1(n117), .A2(n76), .B1(n64), .B2(n115), .ZN(n96) );
  INV_X1 U95 ( .A(n96), .ZN(n70) );
  NOR2_X1 U96 ( .A1(n30), .A2(n62), .ZN(n100) );
  XNOR2_X1 U97 ( .A(n19), .B(\mult_x_1/n281 ), .ZN(n95) );
  OAI22_X1 U98 ( .A1(n126), .A2(n63), .B1(n127), .B2(n95), .ZN(n98) );
  AOI21_X1 U99 ( .B1(n115), .B2(n117), .A(n64), .ZN(n65) );
  INV_X1 U100 ( .A(n65), .ZN(n97) );
  XNOR2_X1 U101 ( .A(n19), .B(\mult_x_1/n284 ), .ZN(n73) );
  OAI22_X1 U102 ( .A1(n126), .A2(n73), .B1(n127), .B2(n66), .ZN(n214) );
  XNOR2_X1 U103 ( .A(n94), .B(\mult_x_1/n312 ), .ZN(n68) );
  OAI22_X1 U104 ( .A1(n186), .A2(n67), .B1(n68), .B2(n188), .ZN(n213) );
  AOI21_X1 U105 ( .B1(n188), .B2(n186), .A(n68), .ZN(n69) );
  INV_X1 U106 ( .A(n69), .ZN(n212) );
  FA_X1 U107 ( .A(n72), .B(n71), .CI(n70), .CO(n101), .S(n200) );
  NAND2_X1 U108 ( .A1(n201), .A2(n200), .ZN(n82) );
  NOR2_X1 U109 ( .A1(n31), .A2(n62), .ZN(n216) );
  OAI22_X1 U110 ( .A1(n126), .A2(n74), .B1(n127), .B2(n73), .ZN(n228) );
  XNOR2_X1 U111 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n77) );
  OAI22_X1 U112 ( .A1(n117), .A2(n75), .B1(n115), .B2(n77), .ZN(n227) );
  INV_X1 U113 ( .A(n213), .ZN(n226) );
  NAND2_X1 U114 ( .A1(n216), .A2(n217), .ZN(n80) );
  OAI22_X1 U115 ( .A1(n117), .A2(n77), .B1(n115), .B2(n76), .ZN(n215) );
  NAND2_X1 U116 ( .A1(n216), .A2(n215), .ZN(n79) );
  NAND2_X1 U117 ( .A1(n215), .A2(n217), .ZN(n78) );
  NAND3_X1 U118 ( .A1(n80), .A2(n79), .A3(n78), .ZN(n202) );
  OAI21_X1 U119 ( .B1(n200), .B2(n201), .A(n202), .ZN(n81) );
  NAND2_X1 U120 ( .A1(n82), .A2(n81), .ZN(n173) );
  OAI21_X1 U121 ( .B1(n174), .B2(n173), .A(n264), .ZN(n85) );
  INV_X1 U122 ( .A(n264), .ZN(n83) );
  NAND2_X1 U123 ( .A1(n83), .A2(n326), .ZN(n84) );
  NAND2_X1 U124 ( .A1(n85), .A2(n84), .ZN(n350) );
  XNOR2_X1 U147 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n90) );
  XNOR2_X1 U148 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n104) );
  OAI22_X1 U149 ( .A1(n186), .A2(n90), .B1(n188), .B2(n104), .ZN(n165) );
  XNOR2_X1 U150 ( .A(n181), .B(\mult_x_1/n284 ), .ZN(n88) );
  XNOR2_X1 U151 ( .A(n17), .B(\mult_x_1/n283 ), .ZN(n103) );
  OAI22_X1 U152 ( .A1(n190), .A2(n88), .B1(n103), .B2(n23), .ZN(n164) );
  OR2_X1 U153 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n86) );
  OAI22_X1 U154 ( .A1(n117), .A2(n27), .B1(n86), .B2(n115), .ZN(n113) );
  XNOR2_X1 U155 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n87) );
  XNOR2_X1 U156 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n116) );
  OAI22_X1 U157 ( .A1(n117), .A2(n87), .B1(n115), .B2(n116), .ZN(n112) );
  XNOR2_X1 U158 ( .A(n181), .B(\mult_x_1/n285 ), .ZN(n182) );
  OAI22_X1 U159 ( .A1(n190), .A2(n182), .B1(n88), .B2(n23), .ZN(n178) );
  INV_X1 U160 ( .A(n115), .ZN(n89) );
  AND2_X1 U161 ( .A1(\mult_x_1/n288 ), .A2(n89), .ZN(n177) );
  XNOR2_X1 U162 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n179) );
  OAI22_X1 U163 ( .A1(n186), .A2(n179), .B1(n188), .B2(n90), .ZN(n176) );
  NOR2_X1 U164 ( .A1(n171), .A2(n170), .ZN(n92) );
  NAND2_X1 U165 ( .A1(n93), .A2(n324), .ZN(n91) );
  OAI21_X1 U166 ( .B1(n93), .B2(n92), .A(n91), .ZN(n346) );
  NOR2_X1 U167 ( .A1(n32), .A2(n62), .ZN(n124) );
  XNOR2_X1 U168 ( .A(n94), .B(n19), .ZN(n125) );
  OAI22_X1 U169 ( .A1(n126), .A2(n95), .B1(n125), .B2(n127), .ZN(n132) );
  INV_X1 U170 ( .A(n132), .ZN(n123) );
  FA_X1 U171 ( .A(n98), .B(n97), .CI(n21), .CO(n122), .S(n99) );
  FA_X1 U172 ( .A(n101), .B(n100), .CI(n99), .CO(n138), .S(n174) );
  OR2_X1 U173 ( .A1(n139), .A2(n138), .ZN(n102) );
  MUX2_X1 U174 ( .A(n325), .B(n102), .S(n266), .Z(n348) );
  XNOR2_X1 U175 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n109) );
  OAI22_X1 U176 ( .A1(n190), .A2(n103), .B1(n109), .B2(n23), .ZN(n120) );
  AND2_X1 U177 ( .A1(\mult_x_1/n288 ), .A2(n43), .ZN(n119) );
  XNOR2_X1 U178 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n111) );
  OAI22_X1 U179 ( .A1(n186), .A2(n104), .B1(n188), .B2(n111), .ZN(n118) );
  HA_X1 U180 ( .A(n106), .B(n105), .CO(n147), .S(n151) );
  XNOR2_X1 U181 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n114) );
  OAI22_X1 U182 ( .A1(n117), .A2(n114), .B1(n115), .B2(n107), .ZN(n146) );
  OAI22_X1 U183 ( .A1(n190), .A2(n109), .B1(n108), .B2(n23), .ZN(n145) );
  OAI22_X1 U184 ( .A1(n186), .A2(n111), .B1(n188), .B2(n110), .ZN(n144) );
  HA_X1 U185 ( .A(n113), .B(n112), .CO(n162), .S(n163) );
  OAI22_X1 U186 ( .A1(n117), .A2(n116), .B1(n115), .B2(n114), .ZN(n161) );
  FA_X1 U187 ( .A(n120), .B(n119), .CI(n118), .CO(n152), .S(n160) );
  OR2_X1 U188 ( .A1(n158), .A2(n157), .ZN(n121) );
  MUX2_X1 U189 ( .A(n327), .B(n121), .S(n264), .Z(n352) );
  FA_X1 U190 ( .A(n124), .B(n123), .CI(n122), .CO(n134), .S(n139) );
  AOI21_X1 U191 ( .B1(n126), .B2(n127), .A(n125), .ZN(n128) );
  INV_X1 U192 ( .A(n128), .ZN(n130) );
  NOR2_X1 U193 ( .A1(n28), .A2(n62), .ZN(n129) );
  XOR2_X1 U194 ( .A(n130), .B(n129), .Z(n131) );
  XOR2_X1 U195 ( .A(n132), .B(n131), .Z(n133) );
  OR2_X1 U196 ( .A1(n134), .A2(n133), .ZN(n136) );
  NAND2_X1 U197 ( .A1(n134), .A2(n133), .ZN(n135) );
  NAND2_X1 U198 ( .A1(n136), .A2(n135), .ZN(n137) );
  MUX2_X1 U199 ( .A(n328), .B(n137), .S(n316), .Z(n354) );
  NAND2_X1 U200 ( .A1(n139), .A2(n138), .ZN(n140) );
  MUX2_X1 U201 ( .A(n329), .B(n140), .S(n266), .Z(n356) );
  FA_X1 U202 ( .A(n143), .B(n142), .CI(n141), .CO(n225), .S(n241) );
  FA_X1 U203 ( .A(n146), .B(n145), .CI(n144), .CO(n240), .S(n150) );
  FA_X1 U204 ( .A(n152), .B(n151), .CI(n150), .CO(n154), .S(n158) );
  NOR2_X1 U205 ( .A1(n155), .A2(n154), .ZN(n153) );
  MUX2_X1 U206 ( .A(n330), .B(n153), .S(n316), .Z(n358) );
  NAND2_X1 U207 ( .A1(n155), .A2(n154), .ZN(n156) );
  MUX2_X1 U208 ( .A(n331), .B(n156), .S(n316), .Z(n360) );
  NAND2_X1 U209 ( .A1(n158), .A2(n157), .ZN(n159) );
  MUX2_X1 U210 ( .A(n332), .B(n159), .S(n316), .Z(n362) );
  FA_X1 U211 ( .A(n162), .B(n161), .CI(n160), .CO(n157), .S(n168) );
  FA_X1 U212 ( .A(n165), .B(n164), .CI(n163), .CO(n167), .S(n171) );
  NOR2_X1 U213 ( .A1(n168), .A2(n167), .ZN(n166) );
  MUX2_X1 U214 ( .A(n333), .B(n166), .S(n242), .Z(n364) );
  NAND2_X1 U215 ( .A1(n168), .A2(n167), .ZN(n169) );
  MUX2_X1 U216 ( .A(n334), .B(n169), .S(n242), .Z(n366) );
  NAND2_X1 U217 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U218 ( .A(n335), .B(n172), .S(n242), .Z(n368) );
  NAND2_X1 U219 ( .A1(n174), .A2(n173), .ZN(n175) );
  MUX2_X1 U220 ( .A(n336), .B(n175), .S(n242), .Z(n370) );
  FA_X1 U221 ( .A(n178), .B(n177), .CI(n176), .CO(n170), .S(n198) );
  XNOR2_X1 U222 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n180) );
  OAI22_X1 U223 ( .A1(n186), .A2(n180), .B1(n188), .B2(n179), .ZN(n184) );
  XNOR2_X1 U224 ( .A(n181), .B(\mult_x_1/n286 ), .ZN(n187) );
  OAI22_X1 U225 ( .A1(n190), .A2(n187), .B1(n182), .B2(n23), .ZN(n183) );
  HA_X1 U226 ( .A(n184), .B(n183), .CO(n197), .S(n195) );
  OR2_X1 U227 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n185) );
  OAI22_X1 U228 ( .A1(n186), .A2(n26), .B1(n185), .B2(n188), .ZN(n194) );
  OR2_X1 U229 ( .A1(n195), .A2(n194), .ZN(n256) );
  XNOR2_X1 U230 ( .A(n17), .B(\mult_x_1/n287 ), .ZN(n189) );
  OAI22_X1 U231 ( .A1(n190), .A2(n189), .B1(n187), .B2(n23), .ZN(n193) );
  AND2_X1 U232 ( .A1(\mult_x_1/n288 ), .A2(n50), .ZN(n192) );
  NOR2_X1 U233 ( .A1(n193), .A2(n192), .ZN(n249) );
  OAI22_X1 U234 ( .A1(n190), .A2(\mult_x_1/n288 ), .B1(n189), .B2(n23), .ZN(
        n246) );
  OR2_X1 U235 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n191) );
  NAND2_X1 U236 ( .A1(n191), .A2(n190), .ZN(n245) );
  NAND2_X1 U237 ( .A1(n246), .A2(n245), .ZN(n252) );
  NAND2_X1 U238 ( .A1(n193), .A2(n192), .ZN(n250) );
  OAI21_X1 U239 ( .B1(n249), .B2(n252), .A(n250), .ZN(n257) );
  NAND2_X1 U240 ( .A1(n195), .A2(n194), .ZN(n255) );
  INV_X1 U241 ( .A(n255), .ZN(n196) );
  AOI21_X1 U242 ( .B1(n256), .B2(n257), .A(n196), .ZN(n262) );
  NAND2_X1 U243 ( .A1(n198), .A2(n197), .ZN(n261) );
  OAI21_X1 U244 ( .B1(n260), .B2(n262), .A(n261), .ZN(n199) );
  MUX2_X1 U245 ( .A(n337), .B(n199), .S(n242), .Z(n372) );
  XOR2_X1 U246 ( .A(n201), .B(n200), .Z(n203) );
  XOR2_X1 U247 ( .A(n203), .B(n202), .Z(n204) );
  MUX2_X1 U248 ( .A(n338), .B(n204), .S(n242), .Z(n374) );
  OR2_X1 U249 ( .A1(n206), .A2(n205), .ZN(n230) );
  NOR2_X1 U250 ( .A1(n33), .A2(n62), .ZN(n229) );
  OAI21_X1 U251 ( .B1(n209), .B2(n208), .A(n207), .ZN(n211) );
  NAND2_X1 U252 ( .A1(n209), .A2(n208), .ZN(n210) );
  FA_X1 U253 ( .A(n214), .B(n18), .CI(n212), .CO(n201), .S(n221) );
  XOR2_X1 U254 ( .A(n216), .B(n215), .Z(n218) );
  XOR2_X1 U255 ( .A(n218), .B(n217), .Z(n220) );
  MUX2_X1 U256 ( .A(n339), .B(n219), .S(n242), .Z(n376) );
  FA_X1 U257 ( .A(n222), .B(n221), .CI(n220), .CO(n219), .S(n223) );
  MUX2_X1 U258 ( .A(n340), .B(n223), .S(n242), .Z(n378) );
  INV_X1 U259 ( .A(n38), .ZN(n224) );
  FA_X1 U260 ( .A(n228), .B(n227), .CI(n226), .CO(n217), .S(n233) );
  MUX2_X1 U261 ( .A(n341), .B(n231), .S(n242), .Z(n380) );
  FA_X1 U262 ( .A(n24), .B(n233), .CI(n232), .CO(n231), .S(n234) );
  MUX2_X1 U263 ( .A(n342), .B(n234), .S(n242), .Z(n382) );
  FA_X1 U264 ( .A(n237), .B(n236), .CI(n235), .CO(n238), .S(n59) );
  MUX2_X1 U265 ( .A(n343), .B(n238), .S(n242), .Z(n384) );
  FA_X1 U266 ( .A(n241), .B(n240), .CI(n239), .CO(n243), .S(n155) );
  MUX2_X1 U267 ( .A(n345), .B(n243), .S(n242), .Z(n388) );
  MUX2_X1 U268 ( .A(product[0]), .B(n508), .S(n266), .Z(n400) );
  MUX2_X1 U269 ( .A(n508), .B(n509), .S(n264), .Z(n402) );
  AND2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n244) );
  MUX2_X1 U271 ( .A(n509), .B(n244), .S(n266), .Z(n404) );
  MUX2_X1 U272 ( .A(product[1]), .B(n511), .S(n264), .Z(n406) );
  MUX2_X1 U273 ( .A(n511), .B(n512), .S(n266), .Z(n408) );
  OR2_X1 U274 ( .A1(n246), .A2(n245), .ZN(n247) );
  AND2_X1 U275 ( .A1(n247), .A2(n252), .ZN(n248) );
  MUX2_X1 U276 ( .A(n512), .B(n248), .S(n264), .Z(n410) );
  MUX2_X1 U277 ( .A(product[2]), .B(n514), .S(n266), .Z(n412) );
  MUX2_X1 U278 ( .A(n514), .B(n515), .S(n264), .Z(n414) );
  INV_X1 U279 ( .A(n249), .ZN(n251) );
  NAND2_X1 U280 ( .A1(n251), .A2(n250), .ZN(n253) );
  XOR2_X1 U281 ( .A(n253), .B(n252), .Z(n254) );
  MUX2_X1 U282 ( .A(n515), .B(n254), .S(n266), .Z(n416) );
  MUX2_X1 U283 ( .A(product[3]), .B(n517), .S(n264), .Z(n418) );
  MUX2_X1 U284 ( .A(n517), .B(n518), .S(n266), .Z(n420) );
  NAND2_X1 U285 ( .A1(n256), .A2(n255), .ZN(n258) );
  XNOR2_X1 U286 ( .A(n258), .B(n257), .ZN(n259) );
  MUX2_X1 U287 ( .A(n518), .B(n259), .S(n264), .Z(n422) );
  MUX2_X1 U288 ( .A(product[4]), .B(n520), .S(n266), .Z(n424) );
  MUX2_X1 U289 ( .A(n520), .B(n521), .S(n264), .Z(n426) );
  MUX2_X1 U290 ( .A(n521), .B(n263), .S(n266), .Z(n428) );
  MUX2_X1 U291 ( .A(product[5]), .B(n523), .S(n264), .Z(n430) );
  NAND2_X1 U292 ( .A1(n324), .A2(n335), .ZN(n265) );
  XNOR2_X1 U293 ( .A(n265), .B(n337), .ZN(n267) );
  MUX2_X1 U294 ( .A(n523), .B(n267), .S(n266), .Z(n432) );
  BUF_X4 U295 ( .A(en), .Z(n316) );
  MUX2_X1 U296 ( .A(product[6]), .B(n525), .S(n316), .Z(n434) );
  NAND2_X1 U297 ( .A1(n392), .A2(n334), .ZN(n268) );
  AOI21_X1 U298 ( .B1(n324), .B2(n337), .A(n394), .ZN(n270) );
  XOR2_X1 U299 ( .A(n268), .B(n270), .Z(n269) );
  MUX2_X1 U300 ( .A(n525), .B(n269), .S(n316), .Z(n436) );
  MUX2_X1 U301 ( .A(product[7]), .B(n527), .S(n316), .Z(n438) );
  OAI21_X1 U302 ( .B1(n333), .B2(n270), .A(n334), .ZN(n273) );
  NAND2_X1 U303 ( .A1(n327), .A2(n332), .ZN(n271) );
  XNOR2_X1 U304 ( .A(n273), .B(n271), .ZN(n272) );
  MUX2_X1 U305 ( .A(n527), .B(n272), .S(n316), .Z(n440) );
  MUX2_X1 U306 ( .A(product[8]), .B(n529), .S(n316), .Z(n442) );
  AOI21_X1 U307 ( .B1(n273), .B2(n327), .A(n393), .ZN(n276) );
  NAND2_X1 U308 ( .A1(n395), .A2(n331), .ZN(n274) );
  XOR2_X1 U309 ( .A(n276), .B(n274), .Z(n275) );
  MUX2_X1 U310 ( .A(n529), .B(n275), .S(n316), .Z(n444) );
  MUX2_X1 U311 ( .A(product[9]), .B(n531), .S(n316), .Z(n446) );
  OAI21_X1 U312 ( .B1(n276), .B2(n330), .A(n331), .ZN(n290) );
  INV_X1 U313 ( .A(n290), .ZN(n280) );
  NOR2_X1 U314 ( .A1(n344), .A2(n345), .ZN(n285) );
  INV_X1 U315 ( .A(n285), .ZN(n277) );
  NAND2_X1 U316 ( .A1(n344), .A2(n345), .ZN(n287) );
  NAND2_X1 U317 ( .A1(n277), .A2(n287), .ZN(n278) );
  XOR2_X1 U318 ( .A(n280), .B(n278), .Z(n279) );
  MUX2_X1 U319 ( .A(n531), .B(n279), .S(n316), .Z(n448) );
  MUX2_X1 U320 ( .A(product[10]), .B(n533), .S(n316), .Z(n450) );
  OAI21_X1 U321 ( .B1(n280), .B2(n285), .A(n287), .ZN(n283) );
  NOR2_X1 U322 ( .A1(n342), .A2(n343), .ZN(n288) );
  INV_X1 U323 ( .A(n288), .ZN(n281) );
  NAND2_X1 U324 ( .A1(n342), .A2(n343), .ZN(n286) );
  NAND2_X1 U325 ( .A1(n281), .A2(n286), .ZN(n282) );
  XNOR2_X1 U326 ( .A(n283), .B(n282), .ZN(n284) );
  MUX2_X1 U327 ( .A(n533), .B(n284), .S(n316), .Z(n452) );
  MUX2_X1 U328 ( .A(product[11]), .B(n535), .S(n316), .Z(n454) );
  NOR2_X1 U329 ( .A1(n288), .A2(n285), .ZN(n291) );
  OAI21_X1 U330 ( .B1(n288), .B2(n287), .A(n286), .ZN(n289) );
  AOI21_X1 U331 ( .B1(n291), .B2(n290), .A(n289), .ZN(n321) );
  NOR2_X1 U332 ( .A1(n340), .A2(n341), .ZN(n306) );
  INV_X1 U333 ( .A(n306), .ZN(n297) );
  NAND2_X1 U334 ( .A1(n340), .A2(n341), .ZN(n309) );
  NAND2_X1 U335 ( .A1(n297), .A2(n309), .ZN(n292) );
  XOR2_X1 U336 ( .A(n321), .B(n292), .Z(n293) );
  MUX2_X1 U337 ( .A(n535), .B(n293), .S(n316), .Z(n456) );
  MUX2_X1 U338 ( .A(product[12]), .B(n537), .S(n316), .Z(n458) );
  OAI21_X1 U339 ( .B1(n321), .B2(n306), .A(n309), .ZN(n295) );
  OR2_X1 U340 ( .A1(n338), .A2(n339), .ZN(n305) );
  NAND2_X1 U341 ( .A1(n338), .A2(n339), .ZN(n298) );
  NAND2_X1 U342 ( .A1(n305), .A2(n298), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  MUX2_X1 U344 ( .A(n537), .B(n296), .S(n316), .Z(n460) );
  MUX2_X1 U345 ( .A(product[13]), .B(n539), .S(n316), .Z(n462) );
  NAND2_X1 U346 ( .A1(n297), .A2(n305), .ZN(n301) );
  INV_X1 U347 ( .A(n309), .ZN(n299) );
  INV_X1 U348 ( .A(n298), .ZN(n307) );
  AOI21_X1 U349 ( .B1(n299), .B2(n305), .A(n307), .ZN(n300) );
  OAI21_X1 U350 ( .B1(n321), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U351 ( .A1(n326), .A2(n336), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U353 ( .A(n539), .B(n304), .S(n316), .Z(n464) );
  MUX2_X1 U354 ( .A(product[14]), .B(n541), .S(n316), .Z(n466) );
  NAND2_X1 U355 ( .A1(n305), .A2(n326), .ZN(n310) );
  NOR2_X1 U356 ( .A1(n306), .A2(n310), .ZN(n317) );
  INV_X1 U357 ( .A(n317), .ZN(n312) );
  AOI21_X1 U358 ( .B1(n307), .B2(n326), .A(n390), .ZN(n308) );
  OAI21_X1 U359 ( .B1(n310), .B2(n309), .A(n308), .ZN(n318) );
  INV_X1 U360 ( .A(n318), .ZN(n311) );
  OAI21_X1 U361 ( .B1(n321), .B2(n312), .A(n311), .ZN(n314) );
  NAND2_X1 U362 ( .A1(n325), .A2(n329), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U364 ( .A(n541), .B(n315), .S(n316), .Z(n468) );
  MUX2_X1 U365 ( .A(product[15]), .B(n543), .S(n316), .Z(n470) );
  NAND2_X1 U366 ( .A1(n317), .A2(n325), .ZN(n320) );
  AOI21_X1 U367 ( .B1(n318), .B2(n325), .A(n391), .ZN(n319) );
  OAI21_X1 U368 ( .B1(n321), .B2(n320), .A(n319), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n322), .B(n328), .ZN(n323) );
  MUX2_X1 U370 ( .A(n543), .B(n323), .S(n316), .Z(n472) );
  MUX2_X1 U371 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n316), .Z(n474) );
  MUX2_X1 U372 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n316), .Z(n476) );
  MUX2_X1 U373 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n316), .Z(n478) );
  MUX2_X1 U374 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n316), .Z(n480) );
  MUX2_X1 U375 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n266), .Z(n482) );
  MUX2_X1 U376 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n264), .Z(n484) );
  MUX2_X1 U377 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n264), .Z(n486) );
  MUX2_X1 U378 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n316), .Z(n488) );
  MUX2_X1 U379 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n316), .Z(n490) );
  MUX2_X1 U380 ( .A(n17), .B(A_extended[1]), .S(n316), .Z(n492) );
  MUX2_X1 U381 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n264), .Z(n494) );
  MUX2_X1 U382 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n316), .Z(n496) );
  MUX2_X1 U383 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n266), .Z(n498) );
  MUX2_X1 U384 ( .A(n22), .B(A_extended[5]), .S(n266), .Z(n500) );
  MUX2_X1 U385 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n316), .Z(n502) );
  MUX2_X1 U386 ( .A(n19), .B(A_extended[7]), .S(n316), .Z(n504) );
  OR2_X1 U387 ( .A1(n264), .A2(n545), .ZN(n506) );
endmodule


module conv_128_32_DW_mult_pipe_J1_9 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n366, n368, n370, n372, n374,
         n376, n378, n380, n382, n384, n386, n388, n390, n392, n394, n396,
         n398, n400, n402, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n419, n421, n423, n425, n427,
         n429, n431, n433, n435, n437, n439, n441, n443, n445, n447, n449,
         n451, n453, n455, n457, n459, n461, n463, n465, n467, n469, n471,
         n473, n475, n477, n479, n481, n483, n485, n487, n489, n491, n493,
         n495, n497, n499, n501, n503, n505, n507, n509, n511, n513, n515,
         n517, n519, n521, n523, n525, n527, n529, n530, n532, n533, n535,
         n536, n538, n539, n541, n542, n544, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n566, n567, n568;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n417), .SE(n527), .CK(clk), .Q(n567), 
        .QN(n342) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n417), .SE(n523), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n21) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n417), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n417), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n23) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n417), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n18) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n417), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n417), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n415), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n416), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n414), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n417), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n414), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n414), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n20) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n414), .SE(n493), .CK(clk), .Q(n565)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n414), .SE(n491), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n414), .SE(n489), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n414), .SE(n487), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n414), .SE(n485), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n416), .SE(n483), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n415), .SE(n481), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n417), .SE(n479), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n414), .SE(n477), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n414), .SE(n475), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n414), .SE(n473), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n414), .SE(n471), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n414), .SE(n469), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n414), .SE(n467), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n414), .SE(n465), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n414), .SE(n463), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n416), .SE(n461), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n416), .SE(n459), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n416), .SE(n457), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n416), .SE(n455), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n416), .SE(n453), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n416), .SE(n451), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n416), .SE(n449), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n416), .SE(n447), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n416), .SE(n445), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n416), .SE(n443), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n416), .SE(n441), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n415), .SE(n439), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n415), .SE(n437), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n415), .SE(n435), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n415), .SE(n433), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n415), .SE(n431), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n415), .SE(n429), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n415), .SE(n427), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n415), .SE(n425), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n415), .SE(n423), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n415), .SE(n421), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n415), .SE(n419), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n568), .SI(1'b1), .SE(n402), .CK(clk), 
        .Q(n363) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n568), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n362), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n568), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n361), .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n568), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n360), .QN(n413) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n568), .SE(n394), .CK(
        clk), .Q(n343), .QN(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n568), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n357), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n568), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n568), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n355), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n568), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n354), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n568), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n568), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n352), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n568), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n349), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n568), .SE(n372), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n568), .SE(n370), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n568), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n346), .QN(n22) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n568), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n568), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n344) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n417), .SE(n525), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n341) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n417), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n340) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n417), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n19) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n417), .SE(n513), .CK(clk), .Q(n566), 
        .QN(n24) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n568), .SE(n392), .CK(
        clk), .Q(n412), .QN(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n568), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n351), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n568), .SE(n376), .CK(
        clk), .Q(n411), .QN(n350) );
  NOR2_X4 U2 ( .A1(n341), .A2(n342), .ZN(n211) );
  BUF_X1 U3 ( .A(en), .Z(n299) );
  BUF_X1 U4 ( .A(n414), .Z(n417) );
  BUF_X1 U5 ( .A(n414), .Z(n415) );
  BUF_X1 U6 ( .A(n414), .Z(n416) );
  INV_X1 U7 ( .A(n568), .ZN(n414) );
  INV_X1 U8 ( .A(n27), .ZN(n186) );
  INV_X1 U9 ( .A(n11), .ZN(n5) );
  BUF_X1 U10 ( .A(n339), .Z(n268) );
  INV_X1 U11 ( .A(rst_n), .ZN(n568) );
  INV_X1 U12 ( .A(n64), .ZN(n209) );
  NAND2_X1 U13 ( .A1(n138), .A2(n139), .ZN(n117) );
  INV_X1 U14 ( .A(n339), .ZN(n10) );
  BUF_X1 U15 ( .A(en), .Z(n339) );
  NAND2_X1 U16 ( .A1(n100), .A2(n99), .ZN(n101) );
  INV_X1 U17 ( .A(n105), .ZN(n100) );
  XNOR2_X1 U18 ( .A(n141), .B(n140), .ZN(n230) );
  XNOR2_X1 U19 ( .A(n139), .B(n138), .ZN(n140) );
  AND2_X1 U20 ( .A1(n147), .A2(n146), .ZN(n26) );
  NAND2_X1 U21 ( .A1(n145), .A2(n144), .ZN(n146) );
  OR2_X1 U22 ( .A1(n145), .A2(n144), .ZN(n142) );
  NAND3_X1 U23 ( .A1(n124), .A2(n123), .A3(n122), .ZN(n128) );
  INV_X1 U24 ( .A(n150), .ZN(n85) );
  OR2_X2 U25 ( .A1(n27), .A2(n6), .ZN(n188) );
  XOR2_X1 U26 ( .A(\mult_x_1/n312 ), .B(n23), .Z(n6) );
  XNOR2_X1 U27 ( .A(n211), .B(\mult_x_1/n310 ), .ZN(n7) );
  XNOR2_X1 U28 ( .A(n211), .B(\mult_x_1/n310 ), .ZN(n212) );
  INV_X1 U29 ( .A(n19), .ZN(n8) );
  MUX2_X1 U30 ( .A(n180), .B(n345), .S(n5), .Z(n366) );
  OR2_X1 U31 ( .A1(n37), .A2(n36), .ZN(n9) );
  INV_X1 U32 ( .A(n10), .ZN(n11) );
  INV_X2 U33 ( .A(n10), .ZN(n12) );
  INV_X2 U34 ( .A(n10), .ZN(n13) );
  NAND2_X1 U35 ( .A1(n37), .A2(n36), .ZN(n260) );
  OR2_X1 U36 ( .A1(n37), .A2(n36), .ZN(n263) );
  NAND2_X1 U37 ( .A1(n143), .A2(n142), .ZN(n147) );
  NAND2_X1 U38 ( .A1(n103), .A2(n102), .ZN(n175) );
  NAND2_X1 U39 ( .A1(n26), .A2(n13), .ZN(n14) );
  OAI22_X1 U40 ( .A1(n199), .A2(n98), .B1(n197), .B2(n97), .ZN(n104) );
  XNOR2_X1 U41 ( .A(n105), .B(n104), .ZN(n106) );
  NAND2_X1 U42 ( .A1(n105), .A2(n104), .ZN(n102) );
  INV_X1 U43 ( .A(n104), .ZN(n99) );
  NAND2_X1 U44 ( .A1(n118), .A2(n117), .ZN(n15) );
  BUF_X2 U45 ( .A(\mult_x_1/n310 ), .Z(n16) );
  XNOR2_X1 U46 ( .A(\mult_x_1/a[2] ), .B(n24), .ZN(n27) );
  OAI22_X1 U47 ( .A1(n188), .A2(n90), .B1(n91), .B2(n186), .ZN(n17) );
  XNOR2_X1 U48 ( .A(n8), .B(\mult_x_1/n286 ), .ZN(n35) );
  XNOR2_X1 U49 ( .A(n8), .B(\mult_x_1/n285 ), .ZN(n187) );
  OAI22_X1 U50 ( .A1(n188), .A2(n35), .B1(n186), .B2(n187), .ZN(n252) );
  NAND2_X1 U51 ( .A1(n566), .A2(n18), .ZN(n183) );
  XNOR2_X1 U52 ( .A(n566), .B(\mult_x_1/n284 ), .ZN(n33) );
  XNOR2_X1 U53 ( .A(n566), .B(\mult_x_1/n283 ), .ZN(n182) );
  OAI22_X1 U54 ( .A1(n183), .A2(n33), .B1(n182), .B2(n18), .ZN(n251) );
  XOR2_X1 U55 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n28) );
  XNOR2_X1 U56 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n29) );
  NAND2_X1 U57 ( .A1(n28), .A2(n29), .ZN(n199) );
  OR2_X1 U58 ( .A1(\mult_x_1/n288 ), .A2(n340), .ZN(n31) );
  INV_X1 U59 ( .A(n29), .ZN(n30) );
  INV_X2 U60 ( .A(n30), .ZN(n197) );
  OAI22_X1 U61 ( .A1(n199), .A2(n340), .B1(n31), .B2(n197), .ZN(n195) );
  INV_X1 U62 ( .A(n340), .ZN(n338) );
  XNOR2_X1 U63 ( .A(n338), .B(\mult_x_1/n288 ), .ZN(n32) );
  XNOR2_X1 U64 ( .A(n338), .B(\mult_x_1/n287 ), .ZN(n198) );
  OAI22_X1 U65 ( .A1(n199), .A2(n32), .B1(n197), .B2(n198), .ZN(n194) );
  XNOR2_X1 U66 ( .A(n566), .B(\mult_x_1/n285 ), .ZN(n40) );
  OAI22_X1 U67 ( .A1(n183), .A2(n40), .B1(n33), .B2(n18), .ZN(n52) );
  INV_X1 U68 ( .A(n197), .ZN(n34) );
  AND2_X1 U69 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n51) );
  XNOR2_X1 U70 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n38) );
  OAI22_X1 U71 ( .A1(n188), .A2(n38), .B1(n186), .B2(n35), .ZN(n50) );
  NAND2_X1 U72 ( .A1(n9), .A2(n260), .ZN(n58) );
  XNOR2_X1 U73 ( .A(n8), .B(\mult_x_1/n288 ), .ZN(n39) );
  OAI22_X1 U74 ( .A1(n188), .A2(n39), .B1(n186), .B2(n38), .ZN(n54) );
  XNOR2_X1 U75 ( .A(n566), .B(\mult_x_1/n286 ), .ZN(n42) );
  OAI22_X1 U76 ( .A1(n183), .A2(n42), .B1(n40), .B2(n18), .ZN(n53) );
  OR2_X1 U77 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n41) );
  OAI22_X1 U78 ( .A1(n188), .A2(n19), .B1(n41), .B2(n186), .ZN(n47) );
  OR2_X1 U79 ( .A1(n48), .A2(n47), .ZN(n286) );
  XNOR2_X1 U80 ( .A(n566), .B(\mult_x_1/n287 ), .ZN(n43) );
  OAI22_X1 U81 ( .A1(n183), .A2(n43), .B1(n42), .B2(n18), .ZN(n46) );
  AND2_X1 U82 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n45) );
  NOR2_X1 U83 ( .A1(n46), .A2(n45), .ZN(n279) );
  OAI22_X1 U84 ( .A1(n183), .A2(\mult_x_1/n288 ), .B1(n43), .B2(n18), .ZN(n276) );
  OR2_X1 U85 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n44) );
  NAND2_X1 U86 ( .A1(n44), .A2(n183), .ZN(n275) );
  NAND2_X1 U87 ( .A1(n276), .A2(n275), .ZN(n282) );
  NAND2_X1 U88 ( .A1(n46), .A2(n45), .ZN(n280) );
  OAI21_X1 U89 ( .B1(n279), .B2(n282), .A(n280), .ZN(n287) );
  NAND2_X1 U90 ( .A1(n48), .A2(n47), .ZN(n285) );
  INV_X1 U91 ( .A(n285), .ZN(n49) );
  AOI21_X1 U92 ( .B1(n286), .B2(n287), .A(n49), .ZN(n293) );
  FA_X1 U93 ( .A(n52), .B(n51), .CI(n50), .CO(n36), .S(n56) );
  HA_X1 U94 ( .A(n54), .B(n53), .CO(n55), .S(n48) );
  NOR2_X1 U95 ( .A1(n56), .A2(n55), .ZN(n290) );
  NAND2_X1 U96 ( .A1(n56), .A2(n55), .ZN(n291) );
  OAI21_X1 U97 ( .B1(n293), .B2(n290), .A(n291), .ZN(n262) );
  INV_X1 U98 ( .A(n262), .ZN(n57) );
  XNOR2_X1 U99 ( .A(n58), .B(n57), .ZN(n60) );
  NAND2_X1 U100 ( .A1(n5), .A2(n545), .ZN(n59) );
  OAI21_X1 U101 ( .B1(n60), .B2(n265), .A(n59), .ZN(n453) );
  XNOR2_X1 U102 ( .A(n338), .B(\mult_x_1/n284 ), .ZN(n69) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n95) );
  OAI22_X1 U104 ( .A1(n199), .A2(n69), .B1(n197), .B2(n95), .ZN(n113) );
  XNOR2_X1 U105 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n70) );
  XNOR2_X1 U106 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n90) );
  OAI22_X1 U107 ( .A1(n188), .A2(n70), .B1(n186), .B2(n90), .ZN(n112) );
  XNOR2_X1 U108 ( .A(n113), .B(n112), .ZN(n134) );
  INV_X1 U109 ( .A(n211), .ZN(n61) );
  OR2_X1 U110 ( .A1(\mult_x_1/n288 ), .A2(n61), .ZN(n62) );
  NOR2_X1 U111 ( .A1(n62), .A2(n7), .ZN(n133) );
  XNOR2_X1 U112 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n63) );
  XNOR2_X1 U113 ( .A(\mult_x_1/n311 ), .B(n21), .ZN(n64) );
  OR2_X2 U114 ( .A1(n63), .A2(n64), .ZN(n208) );
  XNOR2_X1 U115 ( .A(n16), .B(\mult_x_1/n287 ), .ZN(n73) );
  XNOR2_X1 U116 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n67) );
  OAI22_X1 U117 ( .A1(n208), .A2(n73), .B1(n209), .B2(n67), .ZN(n78) );
  XNOR2_X1 U118 ( .A(n566), .B(\mult_x_1/n281 ), .ZN(n80) );
  AND2_X1 U119 ( .A1(n567), .A2(\mult_x_1/n281 ), .ZN(n156) );
  XNOR2_X1 U120 ( .A(n156), .B(n566), .ZN(n65) );
  OAI22_X1 U121 ( .A1(n183), .A2(n80), .B1(n65), .B2(n18), .ZN(n77) );
  NOR2_X1 U122 ( .A1(n212), .A2(n20), .ZN(n76) );
  AOI21_X1 U123 ( .B1(n183), .B2(n18), .A(n65), .ZN(n66) );
  INV_X1 U124 ( .A(n66), .ZN(n110) );
  XNOR2_X1 U125 ( .A(n16), .B(\mult_x_1/n285 ), .ZN(n94) );
  OAI22_X1 U126 ( .A1(n208), .A2(n67), .B1(n209), .B2(n94), .ZN(n109) );
  XNOR2_X1 U127 ( .A(n211), .B(\mult_x_1/n287 ), .ZN(n68) );
  NOR2_X1 U128 ( .A1(n68), .A2(n7), .ZN(n108) );
  XNOR2_X1 U129 ( .A(n338), .B(\mult_x_1/n285 ), .ZN(n79) );
  OAI22_X1 U130 ( .A1(n199), .A2(n79), .B1(n197), .B2(n69), .ZN(n84) );
  XNOR2_X1 U131 ( .A(n8), .B(\mult_x_1/n283 ), .ZN(n81) );
  OAI22_X1 U132 ( .A1(n188), .A2(n81), .B1(n186), .B2(n70), .ZN(n83) );
  INV_X1 U133 ( .A(\mult_x_1/n310 ), .ZN(n72) );
  OR2_X1 U134 ( .A1(\mult_x_1/n288 ), .A2(n72), .ZN(n71) );
  OAI22_X1 U135 ( .A1(n208), .A2(n72), .B1(n71), .B2(n209), .ZN(n190) );
  XNOR2_X1 U136 ( .A(n16), .B(\mult_x_1/n288 ), .ZN(n74) );
  OAI22_X1 U137 ( .A1(n208), .A2(n74), .B1(n209), .B2(n73), .ZN(n189) );
  XNOR2_X1 U138 ( .A(n145), .B(n144), .ZN(n75) );
  XNOR2_X1 U139 ( .A(n143), .B(n75), .ZN(n151) );
  FA_X1 U140 ( .A(n78), .B(n77), .CI(n76), .CO(n132), .S(n236) );
  XNOR2_X1 U141 ( .A(n338), .B(\mult_x_1/n286 ), .ZN(n196) );
  OAI22_X1 U142 ( .A1(n199), .A2(n196), .B1(n197), .B2(n79), .ZN(n193) );
  XNOR2_X1 U143 ( .A(n566), .B(\mult_x_1/n282 ), .ZN(n181) );
  OAI22_X1 U144 ( .A1(n183), .A2(n181), .B1(n80), .B2(n18), .ZN(n192) );
  XNOR2_X1 U145 ( .A(n8), .B(\mult_x_1/n284 ), .ZN(n185) );
  OAI22_X1 U146 ( .A1(n188), .A2(n185), .B1(n186), .B2(n81), .ZN(n191) );
  FA_X1 U147 ( .A(n84), .B(n83), .CI(n82), .CO(n144), .S(n234) );
  NAND2_X1 U148 ( .A1(n85), .A2(n11), .ZN(n86) );
  OAI22_X1 U149 ( .A1(n86), .A2(n151), .B1(n13), .B2(n410), .ZN(n400) );
  XNOR2_X1 U150 ( .A(n338), .B(\mult_x_1/n281 ), .ZN(n97) );
  XNOR2_X1 U151 ( .A(n156), .B(n338), .ZN(n159) );
  OAI22_X1 U152 ( .A1(n199), .A2(n97), .B1(n159), .B2(n197), .ZN(n168) );
  INV_X1 U153 ( .A(n168), .ZN(n161) );
  XNOR2_X1 U154 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n89) );
  XNOR2_X1 U155 ( .A(n16), .B(\mult_x_1/n282 ), .ZN(n158) );
  OAI22_X1 U156 ( .A1(n208), .A2(n89), .B1(n209), .B2(n158), .ZN(n163) );
  XNOR2_X1 U157 ( .A(n211), .B(\mult_x_1/n284 ), .ZN(n87) );
  NOR2_X1 U158 ( .A1(n87), .A2(n212), .ZN(n162) );
  XNOR2_X1 U159 ( .A(n163), .B(n162), .ZN(n88) );
  XNOR2_X1 U160 ( .A(n161), .B(n88), .ZN(n177) );
  XNOR2_X1 U161 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n93) );
  OAI22_X1 U162 ( .A1(n208), .A2(n93), .B1(n209), .B2(n89), .ZN(n121) );
  XNOR2_X1 U163 ( .A(n156), .B(\mult_x_1/n312 ), .ZN(n91) );
  OAI22_X1 U164 ( .A1(n188), .A2(n90), .B1(n91), .B2(n186), .ZN(n120) );
  AOI21_X1 U165 ( .B1(n186), .B2(n188), .A(n91), .ZN(n92) );
  INV_X1 U166 ( .A(n92), .ZN(n119) );
  OAI22_X1 U167 ( .A1(n208), .A2(n94), .B1(n209), .B2(n93), .ZN(n137) );
  XNOR2_X1 U168 ( .A(n338), .B(\mult_x_1/n282 ), .ZN(n98) );
  OAI22_X1 U169 ( .A1(n199), .A2(n95), .B1(n197), .B2(n98), .ZN(n136) );
  INV_X1 U170 ( .A(n120), .ZN(n135) );
  XNOR2_X1 U171 ( .A(n211), .B(\mult_x_1/n285 ), .ZN(n96) );
  NOR2_X1 U172 ( .A1(n96), .A2(n7), .ZN(n105) );
  NAND2_X1 U173 ( .A1(n107), .A2(n101), .ZN(n103) );
  XNOR2_X1 U174 ( .A(n107), .B(n106), .ZN(n228) );
  FA_X1 U175 ( .A(n110), .B(n109), .CI(n108), .CO(n141), .S(n145) );
  XNOR2_X1 U176 ( .A(n211), .B(\mult_x_1/n286 ), .ZN(n111) );
  NOR2_X1 U177 ( .A1(n111), .A2(n7), .ZN(n139) );
  INV_X1 U178 ( .A(n139), .ZN(n115) );
  OR2_X1 U179 ( .A1(n113), .A2(n112), .ZN(n138) );
  INV_X1 U180 ( .A(n138), .ZN(n114) );
  NAND2_X1 U181 ( .A1(n115), .A2(n114), .ZN(n116) );
  NAND2_X1 U182 ( .A1(n141), .A2(n116), .ZN(n118) );
  NAND2_X1 U183 ( .A1(n118), .A2(n117), .ZN(n227) );
  NAND2_X1 U184 ( .A1(n228), .A2(n15), .ZN(n124) );
  FA_X1 U185 ( .A(n121), .B(n17), .CI(n119), .CO(n176), .S(n226) );
  NAND2_X1 U186 ( .A1(n228), .A2(n226), .ZN(n123) );
  NAND2_X1 U187 ( .A1(n15), .A2(n226), .ZN(n122) );
  NAND2_X1 U188 ( .A1(n129), .A2(n128), .ZN(n125) );
  NAND2_X1 U189 ( .A1(n125), .A2(n13), .ZN(n127) );
  OR2_X1 U190 ( .A1(n11), .A2(n413), .ZN(n126) );
  NAND2_X1 U191 ( .A1(n127), .A2(n126), .ZN(n396) );
  OAI21_X1 U192 ( .B1(n129), .B2(n128), .A(n268), .ZN(n131) );
  OR2_X1 U193 ( .A1(n268), .A2(n22), .ZN(n130) );
  NAND2_X1 U194 ( .A1(n131), .A2(n130), .ZN(n368) );
  FA_X1 U195 ( .A(n132), .B(n133), .CI(n134), .CO(n232), .S(n143) );
  FA_X1 U196 ( .A(n137), .B(n136), .CI(n135), .CO(n107), .S(n231) );
  OR2_X1 U197 ( .A1(n11), .A2(n343), .ZN(n149) );
  NAND2_X1 U198 ( .A1(n26), .A2(n12), .ZN(n148) );
  OAI211_X1 U199 ( .C1(n273), .C2(n5), .A(n149), .B(n14), .ZN(n394) );
  NAND2_X1 U200 ( .A1(n151), .A2(n150), .ZN(n152) );
  NAND2_X1 U201 ( .A1(n152), .A2(n12), .ZN(n154) );
  OR2_X1 U202 ( .A1(n11), .A2(n25), .ZN(n153) );
  NAND2_X1 U203 ( .A1(n154), .A2(n153), .ZN(n398) );
  XNOR2_X1 U224 ( .A(n211), .B(\mult_x_1/n282 ), .ZN(n155) );
  NOR2_X1 U225 ( .A1(n155), .A2(n7), .ZN(n206) );
  XNOR2_X1 U226 ( .A(n16), .B(\mult_x_1/n281 ), .ZN(n157) );
  XNOR2_X1 U227 ( .A(n156), .B(n16), .ZN(n207) );
  OAI22_X1 U228 ( .A1(n208), .A2(n157), .B1(n207), .B2(n209), .ZN(n217) );
  INV_X1 U229 ( .A(n217), .ZN(n205) );
  OAI22_X1 U230 ( .A1(n208), .A2(n158), .B1(n209), .B2(n157), .ZN(n170) );
  AOI21_X1 U231 ( .B1(n197), .B2(n199), .A(n159), .ZN(n160) );
  INV_X1 U232 ( .A(n160), .ZN(n169) );
  NAND2_X1 U233 ( .A1(n161), .A2(n163), .ZN(n166) );
  NAND2_X1 U234 ( .A1(n161), .A2(n162), .ZN(n165) );
  NAND2_X1 U235 ( .A1(n163), .A2(n162), .ZN(n164) );
  NAND3_X1 U236 ( .A1(n166), .A2(n165), .A3(n164), .ZN(n174) );
  XNOR2_X1 U237 ( .A(n211), .B(\mult_x_1/n283 ), .ZN(n167) );
  NOR2_X1 U238 ( .A1(n167), .A2(n7), .ZN(n173) );
  FA_X1 U239 ( .A(n170), .B(n168), .CI(n169), .CO(n204), .S(n172) );
  OR2_X1 U240 ( .A1(n224), .A2(n223), .ZN(n171) );
  MUX2_X1 U241 ( .A(n344), .B(n171), .S(n268), .Z(n364) );
  FA_X1 U242 ( .A(n174), .B(n173), .CI(n172), .CO(n223), .S(n258) );
  INV_X1 U243 ( .A(n258), .ZN(n179) );
  FA_X1 U244 ( .A(n177), .B(n176), .CI(n175), .CO(n257), .S(n129) );
  INV_X1 U245 ( .A(n257), .ZN(n178) );
  NAND2_X1 U246 ( .A1(n179), .A2(n178), .ZN(n180) );
  OAI22_X1 U247 ( .A1(n183), .A2(n182), .B1(n181), .B2(n18), .ZN(n202) );
  INV_X1 U248 ( .A(n209), .ZN(n184) );
  AND2_X1 U249 ( .A1(\mult_x_1/n288 ), .A2(n184), .ZN(n201) );
  OAI22_X1 U250 ( .A1(n188), .A2(n187), .B1(n186), .B2(n185), .ZN(n200) );
  HA_X1 U251 ( .A(n190), .B(n189), .CO(n82), .S(n238) );
  FA_X1 U252 ( .A(n193), .B(n192), .CI(n191), .CO(n235), .S(n237) );
  HA_X1 U253 ( .A(n195), .B(n194), .CO(n249), .S(n250) );
  OAI22_X1 U254 ( .A1(n199), .A2(n198), .B1(n197), .B2(n196), .ZN(n248) );
  FA_X1 U255 ( .A(n202), .B(n201), .CI(n200), .CO(n239), .S(n247) );
  OR2_X1 U256 ( .A1(n245), .A2(n244), .ZN(n203) );
  MUX2_X1 U257 ( .A(n347), .B(n203), .S(n268), .Z(n370) );
  FA_X1 U258 ( .A(n206), .B(n205), .CI(n204), .CO(n219), .S(n224) );
  AOI21_X1 U259 ( .B1(n209), .B2(n208), .A(n207), .ZN(n210) );
  INV_X1 U260 ( .A(n210), .ZN(n215) );
  XNOR2_X1 U261 ( .A(n211), .B(\mult_x_1/n281 ), .ZN(n213) );
  NOR2_X1 U262 ( .A1(n213), .A2(n7), .ZN(n214) );
  XOR2_X1 U263 ( .A(n215), .B(n214), .Z(n216) );
  XOR2_X1 U264 ( .A(n217), .B(n216), .Z(n218) );
  OR2_X1 U265 ( .A1(n219), .A2(n218), .ZN(n221) );
  NAND2_X1 U266 ( .A1(n219), .A2(n218), .ZN(n220) );
  NAND2_X1 U267 ( .A1(n221), .A2(n220), .ZN(n222) );
  MUX2_X1 U268 ( .A(n348), .B(n222), .S(n268), .Z(n372) );
  NAND2_X1 U269 ( .A1(n224), .A2(n223), .ZN(n225) );
  MUX2_X1 U270 ( .A(n349), .B(n225), .S(n268), .Z(n374) );
  XNOR2_X1 U271 ( .A(n227), .B(n226), .ZN(n229) );
  XNOR2_X1 U272 ( .A(n229), .B(n228), .ZN(n266) );
  FA_X1 U273 ( .A(n232), .B(n231), .CI(n230), .CO(n267), .S(n273) );
  NOR2_X1 U274 ( .A1(n266), .A2(n267), .ZN(n233) );
  MUX2_X1 U275 ( .A(n350), .B(n233), .S(n268), .Z(n376) );
  FA_X1 U276 ( .A(n236), .B(n235), .CI(n234), .CO(n150), .S(n242) );
  FA_X1 U277 ( .A(n239), .B(n238), .CI(n237), .CO(n241), .S(n245) );
  NOR2_X1 U278 ( .A1(n242), .A2(n241), .ZN(n240) );
  MUX2_X1 U279 ( .A(n352), .B(n240), .S(n268), .Z(n380) );
  NAND2_X1 U280 ( .A1(n242), .A2(n241), .ZN(n243) );
  MUX2_X1 U281 ( .A(n353), .B(n243), .S(n268), .Z(n382) );
  NAND2_X1 U282 ( .A1(n245), .A2(n244), .ZN(n246) );
  MUX2_X1 U283 ( .A(n354), .B(n246), .S(n268), .Z(n384) );
  FA_X1 U284 ( .A(n249), .B(n248), .CI(n247), .CO(n244), .S(n255) );
  FA_X1 U285 ( .A(n252), .B(n251), .CI(n250), .CO(n254), .S(n37) );
  NOR2_X1 U286 ( .A1(n255), .A2(n254), .ZN(n253) );
  MUX2_X1 U287 ( .A(n355), .B(n253), .S(n268), .Z(n386) );
  NAND2_X1 U288 ( .A1(n255), .A2(n254), .ZN(n256) );
  MUX2_X1 U289 ( .A(n356), .B(n256), .S(n12), .Z(n388) );
  NAND2_X1 U290 ( .A1(n258), .A2(n257), .ZN(n259) );
  MUX2_X1 U291 ( .A(n357), .B(n259), .S(n13), .Z(n390) );
  INV_X1 U292 ( .A(n260), .ZN(n261) );
  AOI21_X1 U293 ( .B1(n263), .B2(n262), .A(n261), .ZN(n264) );
  MUX2_X1 U294 ( .A(n363), .B(n264), .S(n12), .Z(n402) );
  INV_X1 U295 ( .A(n268), .ZN(n265) );
  NAND2_X1 U296 ( .A1(n351), .A2(n265), .ZN(n271) );
  NAND2_X1 U297 ( .A1(n266), .A2(n267), .ZN(n269) );
  NAND2_X1 U298 ( .A1(n269), .A2(n268), .ZN(n270) );
  NAND2_X1 U299 ( .A1(n270), .A2(n271), .ZN(n378) );
  NAND2_X1 U300 ( .A1(n5), .A2(n358), .ZN(n272) );
  OAI21_X1 U301 ( .B1(n148), .B2(n273), .A(n272), .ZN(n392) );
  MUX2_X1 U302 ( .A(product[0]), .B(n529), .S(n299), .Z(n419) );
  MUX2_X1 U303 ( .A(n529), .B(n530), .S(n299), .Z(n421) );
  AND2_X1 U304 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n274) );
  MUX2_X1 U305 ( .A(n530), .B(n274), .S(n299), .Z(n423) );
  MUX2_X1 U306 ( .A(product[1]), .B(n532), .S(n299), .Z(n425) );
  MUX2_X1 U307 ( .A(n532), .B(n533), .S(n299), .Z(n427) );
  OR2_X1 U308 ( .A1(n276), .A2(n275), .ZN(n277) );
  AND2_X1 U309 ( .A1(n277), .A2(n282), .ZN(n278) );
  MUX2_X1 U310 ( .A(n533), .B(n278), .S(n299), .Z(n429) );
  MUX2_X1 U311 ( .A(product[2]), .B(n535), .S(n299), .Z(n431) );
  MUX2_X1 U312 ( .A(n535), .B(n536), .S(n299), .Z(n433) );
  INV_X1 U313 ( .A(n279), .ZN(n281) );
  NAND2_X1 U314 ( .A1(n281), .A2(n280), .ZN(n283) );
  XOR2_X1 U315 ( .A(n283), .B(n282), .Z(n284) );
  MUX2_X1 U316 ( .A(n536), .B(n284), .S(n299), .Z(n435) );
  MUX2_X1 U317 ( .A(product[3]), .B(n538), .S(n299), .Z(n437) );
  MUX2_X1 U318 ( .A(n538), .B(n539), .S(n299), .Z(n439) );
  NAND2_X1 U319 ( .A1(n286), .A2(n285), .ZN(n288) );
  XNOR2_X1 U320 ( .A(n288), .B(n287), .ZN(n289) );
  MUX2_X1 U321 ( .A(n539), .B(n289), .S(n299), .Z(n441) );
  MUX2_X1 U322 ( .A(product[4]), .B(n541), .S(n299), .Z(n443) );
  MUX2_X1 U323 ( .A(n541), .B(n542), .S(n299), .Z(n445) );
  INV_X1 U324 ( .A(n290), .ZN(n292) );
  NAND2_X1 U325 ( .A1(n292), .A2(n291), .ZN(n294) );
  XOR2_X1 U326 ( .A(n294), .B(n293), .Z(n295) );
  MUX2_X1 U327 ( .A(n542), .B(n295), .S(n299), .Z(n447) );
  MUX2_X1 U328 ( .A(product[5]), .B(n544), .S(n299), .Z(n449) );
  MUX2_X1 U329 ( .A(n544), .B(n545), .S(n299), .Z(n451) );
  MUX2_X1 U330 ( .A(product[6]), .B(n547), .S(n299), .Z(n455) );
  NAND2_X1 U331 ( .A1(n407), .A2(n356), .ZN(n296) );
  XOR2_X1 U332 ( .A(n296), .B(n363), .Z(n297) );
  MUX2_X1 U333 ( .A(n547), .B(n297), .S(n299), .Z(n457) );
  MUX2_X1 U334 ( .A(product[7]), .B(n549), .S(n299), .Z(n459) );
  OAI21_X1 U335 ( .B1(n355), .B2(n363), .A(n356), .ZN(n301) );
  NAND2_X1 U336 ( .A1(n347), .A2(n354), .ZN(n298) );
  XNOR2_X1 U337 ( .A(n301), .B(n298), .ZN(n300) );
  MUX2_X1 U338 ( .A(n549), .B(n300), .S(n299), .Z(n461) );
  MUX2_X1 U339 ( .A(product[8]), .B(n551), .S(n13), .Z(n463) );
  AOI21_X1 U340 ( .B1(n301), .B2(n347), .A(n408), .ZN(n304) );
  NAND2_X1 U341 ( .A1(n409), .A2(n353), .ZN(n302) );
  XOR2_X1 U342 ( .A(n304), .B(n302), .Z(n303) );
  MUX2_X1 U343 ( .A(n551), .B(n303), .S(n12), .Z(n465) );
  MUX2_X1 U344 ( .A(product[9]), .B(n553), .S(n13), .Z(n467) );
  OAI21_X1 U345 ( .B1(n304), .B2(n352), .A(n353), .ZN(n312) );
  INV_X1 U346 ( .A(n312), .ZN(n307) );
  NAND2_X1 U347 ( .A1(n410), .A2(n361), .ZN(n305) );
  XOR2_X1 U348 ( .A(n307), .B(n305), .Z(n306) );
  MUX2_X1 U349 ( .A(n553), .B(n306), .S(n12), .Z(n469) );
  MUX2_X1 U350 ( .A(product[10]), .B(n555), .S(n13), .Z(n471) );
  OAI21_X1 U351 ( .B1(n307), .B2(n362), .A(n361), .ZN(n309) );
  NAND2_X1 U352 ( .A1(n412), .A2(n359), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U354 ( .A(n555), .B(n310), .S(n12), .Z(n473) );
  MUX2_X1 U355 ( .A(product[11]), .B(n557), .S(n13), .Z(n475) );
  NOR2_X1 U356 ( .A1(n358), .A2(n362), .ZN(n313) );
  OAI21_X1 U357 ( .B1(n358), .B2(n361), .A(n359), .ZN(n311) );
  AOI21_X1 U358 ( .B1(n313), .B2(n312), .A(n311), .ZN(n335) );
  NAND2_X1 U359 ( .A1(n411), .A2(n351), .ZN(n314) );
  XOR2_X1 U360 ( .A(n335), .B(n314), .Z(n315) );
  MUX2_X1 U361 ( .A(n557), .B(n315), .S(n12), .Z(n477) );
  MUX2_X1 U362 ( .A(product[12]), .B(n559), .S(n13), .Z(n479) );
  OAI21_X1 U363 ( .B1(n335), .B2(n350), .A(n351), .ZN(n317) );
  NAND2_X1 U364 ( .A1(n346), .A2(n360), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U366 ( .A(n559), .B(n318), .S(n12), .Z(n481) );
  MUX2_X1 U367 ( .A(product[13]), .B(n561), .S(n13), .Z(n483) );
  NAND2_X1 U368 ( .A1(n411), .A2(n346), .ZN(n320) );
  AOI21_X1 U369 ( .B1(n406), .B2(n346), .A(n413), .ZN(n319) );
  OAI21_X1 U370 ( .B1(n335), .B2(n320), .A(n319), .ZN(n322) );
  NAND2_X1 U371 ( .A1(n345), .A2(n357), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U373 ( .A(n561), .B(n323), .S(n12), .Z(n485) );
  MUX2_X1 U374 ( .A(product[14]), .B(n563), .S(n13), .Z(n487) );
  NAND2_X1 U375 ( .A1(n346), .A2(n345), .ZN(n325) );
  NOR2_X1 U376 ( .A1(n350), .A2(n325), .ZN(n331) );
  INV_X1 U377 ( .A(n331), .ZN(n327) );
  AOI21_X1 U378 ( .B1(n413), .B2(n345), .A(n405), .ZN(n324) );
  OAI21_X1 U379 ( .B1(n325), .B2(n351), .A(n324), .ZN(n332) );
  INV_X1 U380 ( .A(n332), .ZN(n326) );
  OAI21_X1 U381 ( .B1(n335), .B2(n327), .A(n326), .ZN(n329) );
  NAND2_X1 U382 ( .A1(n344), .A2(n349), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  MUX2_X1 U384 ( .A(n563), .B(n330), .S(n12), .Z(n489) );
  MUX2_X1 U385 ( .A(product[15]), .B(n565), .S(n12), .Z(n491) );
  NAND2_X1 U386 ( .A1(n331), .A2(n344), .ZN(n334) );
  AOI21_X1 U387 ( .B1(n332), .B2(n344), .A(n404), .ZN(n333) );
  OAI21_X1 U388 ( .B1(n335), .B2(n334), .A(n333), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n336), .B(n348), .ZN(n337) );
  MUX2_X1 U390 ( .A(n565), .B(n337), .S(n12), .Z(n493) );
  MUX2_X1 U391 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n12), .Z(n495) );
  MUX2_X1 U392 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n13), .Z(n497) );
  MUX2_X1 U393 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n13), .Z(n499) );
  MUX2_X1 U394 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n13), .Z(n501) );
  MUX2_X1 U395 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n13), .Z(n503) );
  MUX2_X1 U396 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n12), .Z(n505) );
  MUX2_X1 U397 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n13), .Z(n507) );
  MUX2_X1 U398 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n12), .Z(n509) );
  MUX2_X1 U399 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n13), .Z(n511) );
  MUX2_X1 U400 ( .A(n566), .B(A_extended[1]), .S(n13), .Z(n513) );
  MUX2_X1 U401 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n12), .Z(n515) );
  MUX2_X1 U402 ( .A(n8), .B(A_extended[3]), .S(n12), .Z(n517) );
  MUX2_X1 U403 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n13), .Z(n519) );
  MUX2_X1 U404 ( .A(n338), .B(A_extended[5]), .S(n12), .Z(n521) );
  MUX2_X1 U405 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n13), .Z(n523) );
  MUX2_X1 U406 ( .A(n16), .B(A_extended[7]), .S(n12), .Z(n525) );
  OR2_X1 U407 ( .A1(n13), .A2(n567), .ZN(n527) );
endmodule


module conv_128_32_DW_mult_pipe_J1_10 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n353, n355, n357, n359, n361, n363,
         n365, n367, n369, n371, n373, n375, n377, n379, n381, n383, n385,
         n387, n389, n391, n393, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n408, n410, n412, n414, n416, n418,
         n420, n422, n424, n426, n428, n430, n432, n434, n436, n438, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n458, n460, n462,
         n464, n466, n468, n470, n472, n474, n476, n478, n480, n482, n484,
         n486, n488, n490, n492, n494, n496, n498, n500, n502, n504, n506,
         n508, n510, n512, n514, n516, n517, n519, n520, n522, n523, n525,
         n526, n528, n529, n531, n533, n535, n537, n539, n541, n543, n545,
         n547, n549, n551, n552, n553;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n406), .SE(n514), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n406), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n23) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n406), .SE(n506), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n327) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n406), .SE(n502), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n20) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n406), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n25) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n406), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n406), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n35) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n405), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n31) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n404), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n404), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n32) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n406), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n34) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n404), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n33) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n404), .SE(n482), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n27) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n404), .SE(n480), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n404), .SE(n478), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n404), .SE(n476), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n404), .SE(n474), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n404), .SE(n472), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n404), .SE(n470), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n406), .SE(n468), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n405), .SE(n466), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n404), .SE(n464), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n404), .SE(n462), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n404), .SE(n460), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n404), .SE(n458), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n404), .SE(n456), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n404), .SE(n454), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n404), .SE(n452), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n404), .SE(n450), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n404), .SE(n448), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n404), .SE(n446), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n404), .SE(n444), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n404), .SE(n442), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n404), .SE(n440), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n404), .SE(n438), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n404), .SE(n436), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n404), .SE(n434), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n404), .SE(n432), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n404), .SE(n430), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n405), .SE(n428), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n405), .SE(n426), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n405), .SE(n424), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n405), .SE(n422), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n405), .SE(n420), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n405), .SE(n418), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n405), .SE(n416), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n405), .SE(n414), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n405), .SE(n412), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n405), .SE(n410), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n405), .SE(n408), .CK(clk), .Q(
        product[0]) );
  SDFF_X2 clk_r_REG51_S1 ( .D(1'b0), .SI(n406), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n326) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n553), .SE(n393), .CK(
        clk), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2_IP  ( .D(1'b1), .SI(n553), .SE(n391), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n553), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n553), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n553), .SE(n385), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n553), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n553), .SE(n381), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n553), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n343), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n553), .SE(n377), .CK(
        clk), .Q(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n553), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n341), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n553), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n553), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n339), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n553), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n338), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n553), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n553), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n336), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n553), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n335), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n553), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n334), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n553), .SE(n359), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n553), .SE(n357), .CK(
        clk), .QN(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n553), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n331), .QN(n5) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n553), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n553), .SE(n351), .CK(
        clk), .Q(n397), .QN(n329) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n406), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n328) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n406), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n26) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n406), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n36) );
  BUF_X4 U2 ( .A(en), .Z(n317) );
  INV_X2 U3 ( .A(n41), .ZN(n177) );
  BUF_X1 U4 ( .A(n404), .Z(n405) );
  INV_X2 U5 ( .A(n553), .ZN(n404) );
  OR2_X1 U6 ( .A1(n206), .A2(n205), .ZN(n214) );
  BUF_X1 U7 ( .A(n49), .Z(n24) );
  OR2_X1 U8 ( .A1(n270), .A2(n5), .ZN(n63) );
  INV_X1 U9 ( .A(n270), .ZN(n7) );
  BUF_X1 U10 ( .A(n404), .Z(n406) );
  NOR2_X1 U11 ( .A1(n214), .A2(n213), .ZN(n19) );
  OAI21_X1 U12 ( .B1(n13), .B2(n97), .A(n12), .ZN(n102) );
  INV_X1 U13 ( .A(rst_n), .ZN(n553) );
  NOR2_X1 U14 ( .A1(n45), .A2(n46), .ZN(n13) );
  NAND2_X1 U15 ( .A1(n46), .A2(n45), .ZN(n12) );
  NAND2_X1 U16 ( .A1(n39), .A2(n40), .ZN(n147) );
  NAND2_X1 U17 ( .A1(n10), .A2(n9), .ZN(n379) );
  NAND2_X1 U18 ( .A1(n7), .A2(n343), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n11), .A2(n270), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n181), .A2(n180), .ZN(n11) );
  XNOR2_X1 U21 ( .A(n15), .B(n14), .ZN(n85) );
  INV_X1 U22 ( .A(n97), .ZN(n14) );
  XNOR2_X1 U23 ( .A(n46), .B(n45), .ZN(n15) );
  NAND2_X1 U24 ( .A1(n17), .A2(n16), .ZN(n357) );
  NAND2_X1 U25 ( .A1(n7), .A2(n332), .ZN(n16) );
  OAI21_X1 U26 ( .B1(n160), .B2(n159), .A(n270), .ZN(n17) );
  XNOR2_X2 U27 ( .A(n328), .B(n23), .ZN(n136) );
  OAI21_X1 U28 ( .B1(n19), .B2(n18), .A(n69), .ZN(n82) );
  INV_X1 U29 ( .A(n216), .ZN(n18) );
  NAND2_X1 U30 ( .A1(n74), .A2(n73), .ZN(n59) );
  NAND2_X1 U31 ( .A1(n57), .A2(n56), .ZN(n58) );
  XNOR2_X1 U32 ( .A(n76), .B(n75), .ZN(n80) );
  XNOR2_X1 U33 ( .A(n74), .B(n73), .ZN(n75) );
  NAND2_X1 U34 ( .A1(n230), .A2(n229), .ZN(n231) );
  INV_X1 U35 ( .A(n236), .ZN(n230) );
  INV_X1 U36 ( .A(n235), .ZN(n229) );
  INV_X1 U37 ( .A(n73), .ZN(n56) );
  INV_X1 U38 ( .A(n74), .ZN(n57) );
  NAND2_X1 U39 ( .A1(n214), .A2(n213), .ZN(n69) );
  CLKBUF_X1 U40 ( .A(n53), .Z(n71) );
  AND2_X1 U41 ( .A1(n552), .A2(\mult_x_1/n310 ), .ZN(n38) );
  NAND2_X1 U42 ( .A1(n62), .A2(n61), .ZN(n180) );
  NAND2_X1 U43 ( .A1(n85), .A2(n84), .ZN(n61) );
  OAI21_X1 U44 ( .B1(n85), .B2(n84), .A(n86), .ZN(n62) );
  NAND2_X1 U45 ( .A1(n233), .A2(n232), .ZN(n234) );
  NAND2_X1 U46 ( .A1(n236), .A2(n235), .ZN(n232) );
  NAND2_X1 U47 ( .A1(n28), .A2(n231), .ZN(n233) );
  XNOR2_X1 U48 ( .A(n28), .B(n237), .ZN(n238) );
  XNOR2_X1 U49 ( .A(n236), .B(n235), .ZN(n237) );
  XNOR2_X1 U50 ( .A(n20), .B(n36), .ZN(n49) );
  XNOR2_X1 U51 ( .A(n328), .B(n23), .ZN(n21) );
  INV_X1 U52 ( .A(n26), .ZN(n22) );
  XOR2_X1 U53 ( .A(n222), .B(n221), .Z(n28) );
  INV_X1 U54 ( .A(n328), .ZN(n325) );
  BUF_X4 U55 ( .A(en), .Z(n270) );
  AND2_X1 U56 ( .A1(n222), .A2(n221), .ZN(n37) );
  XNOR2_X1 U57 ( .A(n38), .B(\mult_x_1/n310 ), .ZN(n141) );
  NOR2_X1 U58 ( .A1(n30), .A2(n141), .ZN(n46) );
  XOR2_X1 U59 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n105) );
  NAND2_X1 U60 ( .A1(n105), .A2(n21), .ZN(n96) );
  XNOR2_X1 U61 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n47) );
  XNOR2_X1 U62 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n42) );
  OAI22_X1 U63 ( .A1(n96), .A2(n47), .B1(n136), .B2(n42), .ZN(n45) );
  XOR2_X1 U64 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n39) );
  XNOR2_X1 U65 ( .A(n326), .B(n327), .ZN(n40) );
  XNOR2_X1 U66 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n54) );
  AND2_X1 U67 ( .A1(n552), .A2(\mult_x_1/n281 ), .ZN(n94) );
  XNOR2_X1 U68 ( .A(n94), .B(\mult_x_1/n311 ), .ZN(n43) );
  INV_X1 U69 ( .A(n40), .ZN(n41) );
  OAI22_X1 U70 ( .A1(n147), .A2(n54), .B1(n43), .B2(n177), .ZN(n97) );
  NOR2_X1 U71 ( .A1(n31), .A2(n141), .ZN(n101) );
  NAND2_X1 U72 ( .A1(n105), .A2(n21), .ZN(n138) );
  XNOR2_X1 U73 ( .A(n22), .B(\mult_x_1/n281 ), .ZN(n95) );
  OAI22_X1 U74 ( .A1(n138), .A2(n42), .B1(n136), .B2(n95), .ZN(n99) );
  AOI21_X1 U75 ( .B1(n177), .B2(n147), .A(n43), .ZN(n44) );
  INV_X1 U76 ( .A(n44), .ZN(n98) );
  XNOR2_X1 U77 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n52) );
  OAI22_X1 U78 ( .A1(n96), .A2(n52), .B1(n136), .B2(n47), .ZN(n72) );
  XOR2_X1 U79 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n48) );
  NAND2_X2 U80 ( .A1(n48), .A2(n49), .ZN(n191) );
  XNOR2_X1 U81 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n68) );
  XNOR2_X1 U82 ( .A(n94), .B(\mult_x_1/n312 ), .ZN(n50) );
  OAI22_X1 U83 ( .A1(n191), .A2(n68), .B1(n50), .B2(n24), .ZN(n53) );
  AOI21_X1 U84 ( .B1(n24), .B2(n191), .A(n50), .ZN(n51) );
  INV_X1 U85 ( .A(n51), .ZN(n70) );
  XNOR2_X1 U86 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n66) );
  OAI22_X1 U87 ( .A1(n96), .A2(n66), .B1(n136), .B2(n52), .ZN(n212) );
  XNOR2_X1 U88 ( .A(n325), .B(\mult_x_1/n283 ), .ZN(n67) );
  XNOR2_X1 U89 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n55) );
  OAI22_X1 U90 ( .A1(n147), .A2(n67), .B1(n177), .B2(n55), .ZN(n211) );
  INV_X1 U91 ( .A(n53), .ZN(n210) );
  NOR2_X1 U92 ( .A1(n32), .A2(n141), .ZN(n74) );
  OAI22_X1 U93 ( .A1(n147), .A2(n55), .B1(n177), .B2(n54), .ZN(n73) );
  NAND2_X1 U94 ( .A1(n76), .A2(n58), .ZN(n60) );
  NAND2_X1 U95 ( .A1(n60), .A2(n59), .ZN(n86) );
  OAI21_X1 U96 ( .B1(n181), .B2(n180), .A(n270), .ZN(n64) );
  NAND2_X1 U97 ( .A1(n64), .A2(n63), .ZN(n355) );
  NAND2_X1 U98 ( .A1(\mult_x_1/n313 ), .A2(n25), .ZN(n195) );
  XNOR2_X1 U99 ( .A(n94), .B(\mult_x_1/n313 ), .ZN(n139) );
  AOI21_X1 U100 ( .B1(n195), .B2(n25), .A(n139), .ZN(n65) );
  INV_X1 U101 ( .A(n65), .ZN(n225) );
  XNOR2_X1 U102 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n135) );
  OAI22_X1 U103 ( .A1(n138), .A2(n135), .B1(n136), .B2(n66), .ZN(n224) );
  NOR2_X1 U104 ( .A1(n33), .A2(n141), .ZN(n223) );
  XNOR2_X1 U105 ( .A(n325), .B(\mult_x_1/n284 ), .ZN(n145) );
  OAI22_X1 U106 ( .A1(n147), .A2(n145), .B1(n177), .B2(n67), .ZN(n206) );
  XNOR2_X1 U107 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n148) );
  OAI22_X1 U108 ( .A1(n191), .A2(n148), .B1(n24), .B2(n68), .ZN(n205) );
  NOR2_X1 U109 ( .A1(n34), .A2(n141), .ZN(n213) );
  FA_X1 U110 ( .A(n72), .B(n71), .CI(n70), .CO(n84), .S(n81) );
  NAND2_X1 U111 ( .A1(n77), .A2(n270), .ZN(n79) );
  NAND2_X1 U112 ( .A1(n7), .A2(n345), .ZN(n78) );
  NAND2_X1 U113 ( .A1(n79), .A2(n78), .ZN(n383) );
  FA_X1 U114 ( .A(n82), .B(n81), .CI(n80), .CO(n89), .S(n77) );
  INV_X1 U115 ( .A(n89), .ZN(n83) );
  NAND2_X1 U116 ( .A1(n83), .A2(n270), .ZN(n88) );
  XNOR2_X1 U117 ( .A(n85), .B(n84), .ZN(n87) );
  XNOR2_X1 U118 ( .A(n87), .B(n86), .ZN(n90) );
  OAI22_X1 U119 ( .A1(n88), .A2(n90), .B1(n270), .B2(n402), .ZN(n377) );
  NAND2_X1 U120 ( .A1(n90), .A2(n89), .ZN(n91) );
  NAND2_X1 U121 ( .A1(n91), .A2(n270), .ZN(n93) );
  NAND2_X1 U122 ( .A1(n7), .A2(n335), .ZN(n92) );
  NAND2_X1 U123 ( .A1(n93), .A2(n92), .ZN(n363) );
  NOR2_X1 U146 ( .A1(n35), .A2(n141), .ZN(n120) );
  XNOR2_X1 U147 ( .A(n94), .B(n22), .ZN(n121) );
  OAI22_X1 U148 ( .A1(n96), .A2(n95), .B1(n121), .B2(n136), .ZN(n126) );
  INV_X1 U149 ( .A(n126), .ZN(n119) );
  FA_X1 U150 ( .A(n99), .B(n98), .CI(n97), .CO(n118), .S(n100) );
  FA_X1 U151 ( .A(n102), .B(n101), .CI(n100), .CO(n132), .S(n181) );
  OR2_X1 U152 ( .A1(n133), .A2(n132), .ZN(n103) );
  MUX2_X1 U153 ( .A(n330), .B(n103), .S(n270), .Z(n353) );
  XNOR2_X1 U154 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n166) );
  XNOR2_X1 U155 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n109) );
  OAI22_X1 U156 ( .A1(n195), .A2(n166), .B1(n109), .B2(n25), .ZN(n117) );
  INV_X1 U157 ( .A(n136), .ZN(n104) );
  AND2_X1 U158 ( .A1(\mult_x_1/n288 ), .A2(n104), .ZN(n116) );
  XNOR2_X1 U159 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n165) );
  XNOR2_X1 U160 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n110) );
  OAI22_X1 U161 ( .A1(n191), .A2(n165), .B1(n24), .B2(n110), .ZN(n115) );
  NAND2_X1 U162 ( .A1(n105), .A2(n21), .ZN(n108) );
  OR2_X1 U163 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n106) );
  OAI22_X1 U164 ( .A1(n108), .A2(n26), .B1(n106), .B2(n136), .ZN(n151) );
  XNOR2_X1 U165 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n107) );
  XNOR2_X1 U166 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n137) );
  OAI22_X1 U167 ( .A1(n108), .A2(n107), .B1(n136), .B2(n137), .ZN(n150) );
  XNOR2_X1 U168 ( .A(n325), .B(\mult_x_1/n286 ), .ZN(n113) );
  XNOR2_X1 U169 ( .A(n325), .B(\mult_x_1/n285 ), .ZN(n146) );
  OAI22_X1 U170 ( .A1(n147), .A2(n113), .B1(n177), .B2(n146), .ZN(n144) );
  XNOR2_X1 U171 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n140) );
  OAI22_X1 U172 ( .A1(n195), .A2(n109), .B1(n140), .B2(n25), .ZN(n143) );
  XNOR2_X1 U173 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n149) );
  OAI22_X1 U174 ( .A1(n191), .A2(n110), .B1(n24), .B2(n149), .ZN(n142) );
  OR2_X1 U175 ( .A1(\mult_x_1/n288 ), .A2(n328), .ZN(n111) );
  OAI22_X1 U176 ( .A1(n147), .A2(n328), .B1(n111), .B2(n177), .ZN(n168) );
  XNOR2_X1 U177 ( .A(n325), .B(\mult_x_1/n288 ), .ZN(n112) );
  XNOR2_X1 U178 ( .A(n325), .B(\mult_x_1/n287 ), .ZN(n114) );
  OAI22_X1 U179 ( .A1(n147), .A2(n112), .B1(n177), .B2(n114), .ZN(n167) );
  OAI22_X1 U180 ( .A1(n147), .A2(n114), .B1(n177), .B2(n113), .ZN(n163) );
  FA_X1 U181 ( .A(n117), .B(n116), .CI(n115), .CO(n154), .S(n162) );
  FA_X1 U182 ( .A(n120), .B(n119), .CI(n118), .CO(n128), .S(n133) );
  AOI21_X1 U183 ( .B1(n136), .B2(n138), .A(n121), .ZN(n122) );
  INV_X1 U184 ( .A(n122), .ZN(n124) );
  NOR2_X1 U185 ( .A1(n29), .A2(n141), .ZN(n123) );
  XOR2_X1 U186 ( .A(n124), .B(n123), .Z(n125) );
  XOR2_X1 U187 ( .A(n126), .B(n125), .Z(n127) );
  OR2_X1 U188 ( .A1(n128), .A2(n127), .ZN(n130) );
  NAND2_X1 U189 ( .A1(n128), .A2(n127), .ZN(n129) );
  NAND2_X1 U190 ( .A1(n130), .A2(n129), .ZN(n131) );
  MUX2_X1 U191 ( .A(n333), .B(n131), .S(n270), .Z(n359) );
  NAND2_X1 U192 ( .A1(n133), .A2(n132), .ZN(n134) );
  MUX2_X1 U193 ( .A(n334), .B(n134), .S(n270), .Z(n361) );
  OAI22_X1 U194 ( .A1(n138), .A2(n137), .B1(n136), .B2(n135), .ZN(n209) );
  OAI22_X1 U195 ( .A1(n195), .A2(n140), .B1(n139), .B2(n25), .ZN(n208) );
  NOR2_X1 U196 ( .A1(n141), .A2(n27), .ZN(n207) );
  FA_X1 U197 ( .A(n144), .B(n143), .CI(n142), .CO(n240), .S(n152) );
  OAI22_X1 U198 ( .A1(n147), .A2(n146), .B1(n177), .B2(n145), .ZN(n228) );
  OAI22_X1 U199 ( .A1(n191), .A2(n149), .B1(n24), .B2(n148), .ZN(n227) );
  HA_X1 U200 ( .A(n151), .B(n150), .CO(n226), .S(n153) );
  FA_X1 U201 ( .A(n154), .B(n153), .CI(n152), .CO(n156), .S(n160) );
  NOR2_X1 U202 ( .A1(n157), .A2(n156), .ZN(n155) );
  MUX2_X1 U203 ( .A(n336), .B(n155), .S(n270), .Z(n365) );
  NAND2_X1 U204 ( .A1(n157), .A2(n156), .ZN(n158) );
  MUX2_X1 U205 ( .A(n337), .B(n158), .S(n270), .Z(n367) );
  NAND2_X1 U206 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2_X1 U207 ( .A(n338), .B(n161), .S(n270), .Z(n369) );
  FA_X1 U208 ( .A(n164), .B(n163), .CI(n162), .CO(n159), .S(n171) );
  XNOR2_X1 U209 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n178) );
  OAI22_X1 U210 ( .A1(n191), .A2(n178), .B1(n24), .B2(n165), .ZN(n175) );
  XNOR2_X1 U211 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n176) );
  OAI22_X1 U212 ( .A1(n195), .A2(n176), .B1(n166), .B2(n25), .ZN(n174) );
  HA_X1 U213 ( .A(n168), .B(n167), .CO(n164), .S(n173) );
  NOR2_X1 U214 ( .A1(n171), .A2(n170), .ZN(n169) );
  MUX2_X1 U215 ( .A(n339), .B(n169), .S(n270), .Z(n371) );
  NAND2_X1 U216 ( .A1(n171), .A2(n170), .ZN(n172) );
  MUX2_X1 U217 ( .A(n340), .B(n172), .S(n270), .Z(n373) );
  FA_X1 U218 ( .A(n175), .B(n174), .CI(n173), .CO(n170), .S(n244) );
  XNOR2_X1 U219 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n187) );
  OAI22_X1 U220 ( .A1(n195), .A2(n187), .B1(n176), .B2(n25), .ZN(n184) );
  AND2_X1 U221 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n183) );
  XNOR2_X1 U222 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n185) );
  OAI22_X1 U223 ( .A1(n191), .A2(n185), .B1(n24), .B2(n178), .ZN(n182) );
  NAND2_X1 U224 ( .A1(n244), .A2(n243), .ZN(n179) );
  MUX2_X1 U225 ( .A(n341), .B(n179), .S(n270), .Z(n375) );
  FA_X1 U226 ( .A(n184), .B(n183), .CI(n182), .CO(n243), .S(n203) );
  XNOR2_X1 U227 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n186) );
  OAI22_X1 U228 ( .A1(n191), .A2(n186), .B1(n24), .B2(n185), .ZN(n189) );
  XNOR2_X1 U229 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n192) );
  OAI22_X1 U230 ( .A1(n195), .A2(n192), .B1(n187), .B2(n25), .ZN(n188) );
  NOR2_X1 U231 ( .A1(n203), .A2(n202), .ZN(n263) );
  HA_X1 U232 ( .A(n189), .B(n188), .CO(n202), .S(n200) );
  OR2_X1 U233 ( .A1(\mult_x_1/n288 ), .A2(n326), .ZN(n190) );
  OAI22_X1 U234 ( .A1(n191), .A2(n326), .B1(n190), .B2(n24), .ZN(n199) );
  OR2_X1 U235 ( .A1(n200), .A2(n199), .ZN(n259) );
  XNOR2_X1 U236 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n194) );
  OAI22_X1 U237 ( .A1(n195), .A2(n194), .B1(n192), .B2(n25), .ZN(n198) );
  INV_X1 U238 ( .A(n24), .ZN(n193) );
  AND2_X1 U239 ( .A1(\mult_x_1/n288 ), .A2(n193), .ZN(n197) );
  NOR2_X1 U240 ( .A1(n198), .A2(n197), .ZN(n252) );
  OAI22_X1 U241 ( .A1(n195), .A2(\mult_x_1/n288 ), .B1(n194), .B2(n25), .ZN(
        n249) );
  OR2_X1 U242 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n196) );
  NAND2_X1 U243 ( .A1(n196), .A2(n195), .ZN(n248) );
  NAND2_X1 U244 ( .A1(n249), .A2(n248), .ZN(n255) );
  NAND2_X1 U245 ( .A1(n198), .A2(n197), .ZN(n253) );
  OAI21_X1 U246 ( .B1(n252), .B2(n255), .A(n253), .ZN(n260) );
  NAND2_X1 U247 ( .A1(n200), .A2(n199), .ZN(n258) );
  INV_X1 U248 ( .A(n258), .ZN(n201) );
  AOI21_X1 U249 ( .B1(n259), .B2(n260), .A(n201), .ZN(n266) );
  NAND2_X1 U250 ( .A1(n203), .A2(n202), .ZN(n264) );
  OAI21_X1 U251 ( .B1(n263), .B2(n266), .A(n264), .ZN(n204) );
  MUX2_X1 U252 ( .A(n344), .B(n204), .S(n270), .Z(n381) );
  XNOR2_X1 U253 ( .A(n206), .B(n205), .ZN(n222) );
  FA_X1 U254 ( .A(n209), .B(n208), .CI(n207), .CO(n221), .S(n241) );
  FA_X1 U255 ( .A(n212), .B(n211), .CI(n210), .CO(n76), .S(n219) );
  XNOR2_X1 U256 ( .A(n214), .B(n213), .ZN(n215) );
  XNOR2_X1 U257 ( .A(n215), .B(n216), .ZN(n218) );
  MUX2_X1 U258 ( .A(n346), .B(n217), .S(n270), .Z(n385) );
  FA_X1 U259 ( .A(n37), .B(n219), .CI(n218), .CO(n217), .S(n220) );
  MUX2_X1 U260 ( .A(n347), .B(n220), .S(n270), .Z(n387) );
  FA_X1 U261 ( .A(n225), .B(n224), .CI(n223), .CO(n216), .S(n236) );
  FA_X1 U262 ( .A(n228), .B(n227), .CI(n226), .CO(n235), .S(n239) );
  MUX2_X1 U263 ( .A(n348), .B(n234), .S(n270), .Z(n389) );
  MUX2_X1 U264 ( .A(n349), .B(n238), .S(n270), .Z(n391) );
  FA_X1 U265 ( .A(n241), .B(n240), .CI(n239), .CO(n242), .S(n157) );
  MUX2_X1 U266 ( .A(n350), .B(n242), .S(n270), .Z(n393) );
  NOR2_X1 U267 ( .A1(n244), .A2(n243), .ZN(n246) );
  OR2_X1 U268 ( .A1(n270), .A2(n397), .ZN(n245) );
  OAI21_X1 U269 ( .B1(n246), .B2(n7), .A(n245), .ZN(n351) );
  MUX2_X1 U270 ( .A(product[0]), .B(n516), .S(n270), .Z(n408) );
  MUX2_X1 U271 ( .A(n516), .B(n517), .S(n270), .Z(n410) );
  AND2_X1 U272 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n247) );
  MUX2_X1 U273 ( .A(n517), .B(n247), .S(n270), .Z(n412) );
  MUX2_X1 U274 ( .A(product[1]), .B(n519), .S(n270), .Z(n414) );
  MUX2_X1 U275 ( .A(n519), .B(n520), .S(n270), .Z(n416) );
  OR2_X1 U276 ( .A1(n249), .A2(n248), .ZN(n250) );
  AND2_X1 U277 ( .A1(n250), .A2(n255), .ZN(n251) );
  MUX2_X1 U278 ( .A(n520), .B(n251), .S(n270), .Z(n418) );
  MUX2_X1 U279 ( .A(product[2]), .B(n522), .S(n270), .Z(n420) );
  MUX2_X1 U280 ( .A(n522), .B(n523), .S(n270), .Z(n422) );
  INV_X1 U281 ( .A(n252), .ZN(n254) );
  NAND2_X1 U282 ( .A1(n254), .A2(n253), .ZN(n256) );
  XOR2_X1 U283 ( .A(n256), .B(n255), .Z(n257) );
  MUX2_X1 U284 ( .A(n523), .B(n257), .S(n270), .Z(n424) );
  MUX2_X1 U285 ( .A(product[3]), .B(n525), .S(n270), .Z(n426) );
  MUX2_X1 U286 ( .A(n525), .B(n526), .S(n270), .Z(n428) );
  NAND2_X1 U287 ( .A1(n259), .A2(n258), .ZN(n261) );
  XNOR2_X1 U288 ( .A(n261), .B(n260), .ZN(n262) );
  MUX2_X1 U289 ( .A(n526), .B(n262), .S(n270), .Z(n430) );
  MUX2_X1 U290 ( .A(product[4]), .B(n528), .S(n270), .Z(n432) );
  MUX2_X1 U291 ( .A(n528), .B(n529), .S(n270), .Z(n434) );
  INV_X1 U292 ( .A(n263), .ZN(n265) );
  NAND2_X1 U293 ( .A1(n265), .A2(n264), .ZN(n267) );
  XOR2_X1 U294 ( .A(n267), .B(n266), .Z(n268) );
  MUX2_X1 U295 ( .A(n529), .B(n268), .S(n270), .Z(n436) );
  MUX2_X1 U296 ( .A(product[5]), .B(n531), .S(n270), .Z(n438) );
  NAND2_X1 U297 ( .A1(n329), .A2(n341), .ZN(n269) );
  XNOR2_X1 U298 ( .A(n269), .B(n344), .ZN(n271) );
  MUX2_X1 U299 ( .A(n531), .B(n271), .S(n270), .Z(n440) );
  MUX2_X1 U300 ( .A(product[6]), .B(n533), .S(n317), .Z(n442) );
  NAND2_X1 U301 ( .A1(n398), .A2(n340), .ZN(n272) );
  AOI21_X1 U302 ( .B1(n329), .B2(n344), .A(n400), .ZN(n274) );
  XOR2_X1 U303 ( .A(n272), .B(n274), .Z(n273) );
  MUX2_X1 U304 ( .A(n533), .B(n273), .S(n317), .Z(n444) );
  MUX2_X1 U305 ( .A(product[7]), .B(n535), .S(n317), .Z(n446) );
  OAI21_X1 U306 ( .B1(n339), .B2(n274), .A(n340), .ZN(n277) );
  NAND2_X1 U307 ( .A1(n332), .A2(n338), .ZN(n275) );
  XNOR2_X1 U308 ( .A(n277), .B(n275), .ZN(n276) );
  MUX2_X1 U309 ( .A(n535), .B(n276), .S(n317), .Z(n448) );
  MUX2_X1 U310 ( .A(product[8]), .B(n537), .S(n317), .Z(n450) );
  AOI21_X1 U311 ( .B1(n277), .B2(n332), .A(n399), .ZN(n280) );
  NAND2_X1 U312 ( .A1(n401), .A2(n337), .ZN(n278) );
  XOR2_X1 U313 ( .A(n280), .B(n278), .Z(n279) );
  MUX2_X1 U314 ( .A(n537), .B(n279), .S(n317), .Z(n452) );
  MUX2_X1 U315 ( .A(product[9]), .B(n539), .S(n317), .Z(n454) );
  OAI21_X1 U316 ( .B1(n280), .B2(n336), .A(n337), .ZN(n294) );
  INV_X1 U317 ( .A(n294), .ZN(n284) );
  NOR2_X1 U318 ( .A1(n349), .A2(n350), .ZN(n289) );
  INV_X1 U319 ( .A(n289), .ZN(n281) );
  NAND2_X1 U320 ( .A1(n349), .A2(n350), .ZN(n291) );
  NAND2_X1 U321 ( .A1(n281), .A2(n291), .ZN(n282) );
  XOR2_X1 U322 ( .A(n284), .B(n282), .Z(n283) );
  MUX2_X1 U323 ( .A(n539), .B(n283), .S(n317), .Z(n456) );
  MUX2_X1 U324 ( .A(product[10]), .B(n541), .S(n317), .Z(n458) );
  OAI21_X1 U325 ( .B1(n284), .B2(n289), .A(n291), .ZN(n287) );
  NOR2_X1 U326 ( .A1(n347), .A2(n348), .ZN(n292) );
  INV_X1 U327 ( .A(n292), .ZN(n285) );
  NAND2_X1 U328 ( .A1(n347), .A2(n348), .ZN(n290) );
  NAND2_X1 U329 ( .A1(n285), .A2(n290), .ZN(n286) );
  XNOR2_X1 U330 ( .A(n287), .B(n286), .ZN(n288) );
  MUX2_X1 U331 ( .A(n541), .B(n288), .S(n317), .Z(n460) );
  MUX2_X1 U332 ( .A(product[11]), .B(n543), .S(n317), .Z(n462) );
  NOR2_X1 U333 ( .A1(n292), .A2(n289), .ZN(n295) );
  OAI21_X1 U334 ( .B1(n292), .B2(n291), .A(n290), .ZN(n293) );
  AOI21_X1 U335 ( .B1(n295), .B2(n294), .A(n293), .ZN(n322) );
  NOR2_X1 U336 ( .A1(n345), .A2(n346), .ZN(n308) );
  INV_X1 U337 ( .A(n308), .ZN(n301) );
  NAND2_X1 U338 ( .A1(n345), .A2(n346), .ZN(n310) );
  NAND2_X1 U339 ( .A1(n301), .A2(n310), .ZN(n296) );
  XOR2_X1 U340 ( .A(n322), .B(n296), .Z(n297) );
  MUX2_X1 U341 ( .A(n543), .B(n297), .S(n317), .Z(n464) );
  MUX2_X1 U342 ( .A(product[12]), .B(n545), .S(n317), .Z(n466) );
  OAI21_X1 U343 ( .B1(n322), .B2(n308), .A(n310), .ZN(n299) );
  NAND2_X1 U344 ( .A1(n402), .A2(n335), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U346 ( .A(n545), .B(n300), .S(n317), .Z(n468) );
  MUX2_X1 U347 ( .A(product[13]), .B(n547), .S(n317), .Z(n470) );
  NAND2_X1 U348 ( .A1(n301), .A2(n402), .ZN(n304) );
  INV_X1 U349 ( .A(n310), .ZN(n302) );
  AOI21_X1 U350 ( .B1(n302), .B2(n402), .A(n403), .ZN(n303) );
  OAI21_X1 U351 ( .B1(n322), .B2(n304), .A(n303), .ZN(n306) );
  NAND2_X1 U352 ( .A1(n331), .A2(n343), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U354 ( .A(n547), .B(n307), .S(n317), .Z(n472) );
  MUX2_X1 U355 ( .A(product[14]), .B(n549), .S(n317), .Z(n474) );
  NAND2_X1 U356 ( .A1(n402), .A2(n331), .ZN(n311) );
  NOR2_X1 U357 ( .A1(n308), .A2(n311), .ZN(n318) );
  INV_X1 U358 ( .A(n318), .ZN(n313) );
  AOI21_X1 U359 ( .B1(n403), .B2(n331), .A(n396), .ZN(n309) );
  OAI21_X1 U360 ( .B1(n311), .B2(n310), .A(n309), .ZN(n319) );
  INV_X1 U361 ( .A(n319), .ZN(n312) );
  OAI21_X1 U362 ( .B1(n322), .B2(n313), .A(n312), .ZN(n315) );
  NAND2_X1 U363 ( .A1(n330), .A2(n334), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U365 ( .A(n549), .B(n316), .S(n317), .Z(n476) );
  MUX2_X1 U366 ( .A(product[15]), .B(n551), .S(n317), .Z(n478) );
  NAND2_X1 U367 ( .A1(n318), .A2(n330), .ZN(n321) );
  AOI21_X1 U368 ( .B1(n319), .B2(n330), .A(n395), .ZN(n320) );
  OAI21_X1 U369 ( .B1(n322), .B2(n321), .A(n320), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n323), .B(n333), .ZN(n324) );
  MUX2_X1 U371 ( .A(n551), .B(n324), .S(n317), .Z(n480) );
  MUX2_X1 U372 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n317), .Z(n482) );
  MUX2_X1 U373 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n317), .Z(n484) );
  MUX2_X1 U374 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n317), .Z(n486) );
  MUX2_X1 U375 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n317), .Z(n488) );
  MUX2_X1 U376 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n317), .Z(n490) );
  MUX2_X1 U377 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n317), .Z(n492) );
  MUX2_X1 U378 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n317), .Z(n494) );
  MUX2_X1 U379 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n317), .Z(n496) );
  MUX2_X1 U380 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n317), .Z(n498) );
  MUX2_X1 U381 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n317), .Z(n500) );
  MUX2_X1 U382 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n317), .Z(n502) );
  MUX2_X1 U383 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n317), .Z(n504) );
  MUX2_X1 U384 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n317), .Z(n506) );
  MUX2_X1 U385 ( .A(n325), .B(A_extended[5]), .S(n317), .Z(n508) );
  MUX2_X1 U386 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n317), .Z(n510) );
  MUX2_X1 U387 ( .A(n22), .B(A_extended[7]), .S(n317), .Z(n512) );
  OR2_X1 U388 ( .A1(n317), .A2(n552), .ZN(n514) );
endmodule


module conv_128_32_DW_mult_pipe_J1_11 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n344, n346, n348, n350, n352,
         n354, n356, n358, n360, n362, n364, n366, n368, n370, n372, n374,
         n376, n378, n380, n382, n384, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n397, n399, n401, n403, n405, n407, n409,
         n411, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n487, n489, n491, n493, n495, n497,
         n499, n501, n503, n505, n506, n508, n509, n511, n512, n514, n515,
         n517, n518, n520, n522, n524, n526, n528, n530, n532, n534, n536,
         n538, n540, n541, n542, n543;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n395), .SE(n503), .CK(clk), .Q(n542), 
        .QN(n38) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n395), .SE(n499), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n17) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n395), .SE(n497), .CK(clk), .Q(n541), 
        .QN(n28) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n395), .SE(n491), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n395), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n24) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n395), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n29) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n395), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n33) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n393), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n31) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n394), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n30) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n393), .SE(n477), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n32) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n395), .SE(n475), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n34) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n393), .SE(n473), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n35) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n393), .SE(n471), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n26) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n393), .SE(n469), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n393), .SE(n467), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n393), .SE(n465), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n393), .SE(n463), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n393), .SE(n461), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n394), .SE(n459), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG11_S3 ( .D(1'b0), .SI(n395), .SE(n457), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG12_S4 ( .D(1'b0), .SI(n393), .SE(n455), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n393), .SE(n453), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n393), .SE(n451), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n393), .SE(n449), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n393), .SE(n447), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG7_S3 ( .D(1'b0), .SI(n393), .SE(n445), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG8_S4 ( .D(1'b0), .SI(n393), .SE(n443), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG3_S3 ( .D(1'b0), .SI(n393), .SE(n441), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG4_S4 ( .D(1'b0), .SI(n394), .SE(n439), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n394), .SE(n437), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n394), .SE(n435), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n394), .SE(n433), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n394), .SE(n431), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n394), .SE(n429), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n394), .SE(n427), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n394), .SE(n425), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n394), .SE(n423), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n394), .SE(n421), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n394), .SE(n419), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n393), .SE(n417), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n393), .SE(n415), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n393), .SE(n413), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n393), .SE(n411), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n393), .SE(n409), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n393), .SE(n407), .CK(clk), .Q(n509)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n393), .SE(n405), .CK(clk), .Q(n508)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n393), .SE(n403), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n393), .SE(n401), .CK(clk), .Q(n506)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n393), .SE(n399), .CK(clk), .Q(n505)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n393), .SE(n397), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n395), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n37) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n543), .SE(n384), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n543), .SE(n382), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n543), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n543), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n543), .SE(n376), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n543), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2_IP  ( .D(1'b1), .SI(n543), .SE(n372), .CK(
        clk), .QN(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n543), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n334), .QN(n5) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n543), .SE(n368), .CK(
        clk), .QN(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n543), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n332), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n543), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n331), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n543), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n543), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n329), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n543), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n328), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG2_S2  ( .D(n543), .SI(1'b1), .SE(n356), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n543), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n326), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n543), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n325), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n543), .SE(n350), .CK(
        clk), .QN(n324) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n543), .SI(1'b1), .SE(n348), .CK(clk), 
        .Q(n323) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n543), .SE(n346), .CK(
        clk), .QN(n322) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n543), .SI(1'b1), .SE(n344), .CK(clk), 
        .Q(n321), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n543), .SE(n342), .CK(
        clk), .QN(n320) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n395), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n36) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n395), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n25) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n395), .SE(n495), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n18) );
  INV_X2 U2 ( .A(n42), .ZN(n188) );
  BUF_X2 U3 ( .A(en), .Z(n262) );
  BUF_X1 U4 ( .A(n393), .Z(n394) );
  INV_X2 U5 ( .A(n543), .ZN(n393) );
  CLKBUF_X1 U6 ( .A(n541), .Z(n23) );
  INV_X1 U7 ( .A(n262), .ZN(n6) );
  OAI21_X1 U8 ( .B1(n10), .B2(n9), .A(n8), .ZN(n144) );
  BUF_X1 U9 ( .A(n393), .Z(n395) );
  NAND2_X1 U10 ( .A1(n170), .A2(n169), .ZN(n8) );
  INV_X1 U11 ( .A(n168), .ZN(n10) );
  NOR2_X1 U12 ( .A1(n170), .A2(n169), .ZN(n9) );
  INV_X1 U13 ( .A(rst_n), .ZN(n543) );
  OAI22_X1 U14 ( .A1(n181), .A2(n178), .B1(n71), .B2(n179), .ZN(n194) );
  INV_X1 U15 ( .A(n83), .ZN(n175) );
  NAND2_X1 U16 ( .A1(n40), .A2(n41), .ZN(n190) );
  NAND2_X1 U17 ( .A1(n44), .A2(n45), .ZN(n177) );
  BUF_X1 U18 ( .A(\mult_x_1/n313 ), .Z(n156) );
  AND2_X1 U19 ( .A1(n542), .A2(\mult_x_1/n281 ), .ZN(n87) );
  XNOR2_X1 U20 ( .A(n234), .B(n7), .ZN(n125) );
  XNOR2_X1 U21 ( .A(n236), .B(n235), .ZN(n7) );
  OAI21_X1 U22 ( .B1(n237), .B2(n5), .A(n11), .ZN(n370) );
  NAND2_X1 U23 ( .A1(n12), .A2(n237), .ZN(n11) );
  XNOR2_X1 U24 ( .A(n168), .B(n13), .ZN(n12) );
  XNOR2_X1 U25 ( .A(n170), .B(n169), .ZN(n13) );
  NAND2_X1 U26 ( .A1(n38), .A2(\mult_x_1/n310 ), .ZN(n185) );
  CLKBUF_X1 U27 ( .A(\mult_x_1/n313 ), .Z(n43) );
  INV_X1 U28 ( .A(n45), .ZN(n83) );
  INV_X1 U29 ( .A(n15), .ZN(n16) );
  INV_X1 U30 ( .A(n48), .ZN(n179) );
  XNOR2_X1 U31 ( .A(n222), .B(n221), .ZN(n232) );
  XNOR2_X1 U32 ( .A(n220), .B(n219), .ZN(n222) );
  INV_X1 U33 ( .A(n25), .ZN(n14) );
  INV_X1 U34 ( .A(n177), .ZN(n15) );
  XNOR2_X1 U35 ( .A(n17), .B(n28), .ZN(n41) );
  XNOR2_X1 U36 ( .A(n36), .B(n18), .ZN(n45) );
  NAND2_X1 U37 ( .A1(n234), .A2(n235), .ZN(n19) );
  NAND2_X1 U38 ( .A1(n234), .A2(n236), .ZN(n20) );
  NAND2_X1 U39 ( .A1(n235), .A2(n236), .ZN(n21) );
  NAND3_X1 U40 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n238) );
  OAI22_X1 U41 ( .A1(n175), .A2(n65), .B1(n177), .B2(n73), .ZN(n22) );
  INV_X1 U42 ( .A(en), .ZN(n139) );
  INV_X2 U43 ( .A(n139), .ZN(n237) );
  AND2_X1 U44 ( .A1(n227), .A2(n226), .ZN(n27) );
  OR2_X1 U45 ( .A1(n200), .A2(n199), .ZN(n39) );
  XOR2_X1 U46 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n40) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n52) );
  INV_X1 U48 ( .A(n41), .ZN(n42) );
  XNOR2_X1 U49 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n189) );
  OAI22_X1 U50 ( .A1(n190), .A2(n52), .B1(n41), .B2(n189), .ZN(n206) );
  NAND2_X1 U51 ( .A1(n43), .A2(n24), .ZN(n183) );
  XNOR2_X1 U52 ( .A(n43), .B(\mult_x_1/n281 ), .ZN(n46) );
  XNOR2_X1 U53 ( .A(n87), .B(n156), .ZN(n182) );
  OAI22_X1 U54 ( .A1(n183), .A2(n46), .B1(n182), .B2(n24), .ZN(n205) );
  NOR2_X1 U55 ( .A1(n185), .A2(n26), .ZN(n204) );
  XOR2_X1 U56 ( .A(\mult_x_1/a[4] ), .B(n541), .Z(n44) );
  XNOR2_X1 U57 ( .A(n541), .B(\mult_x_1/n286 ), .ZN(n101) );
  XNOR2_X1 U58 ( .A(n541), .B(\mult_x_1/n285 ), .ZN(n49) );
  OAI22_X1 U59 ( .A1(n177), .A2(n101), .B1(n175), .B2(n49), .ZN(n60) );
  XNOR2_X1 U60 ( .A(n156), .B(\mult_x_1/n282 ), .ZN(n54) );
  OAI22_X1 U61 ( .A1(n183), .A2(n54), .B1(n46), .B2(n24), .ZN(n59) );
  XNOR2_X1 U62 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n47) );
  XOR2_X1 U63 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .Z(n48) );
  OR2_X2 U64 ( .A1(n47), .A2(n48), .ZN(n181) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n55) );
  XNOR2_X1 U66 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n50) );
  OAI22_X1 U67 ( .A1(n181), .A2(n55), .B1(n179), .B2(n50), .ZN(n58) );
  XNOR2_X1 U68 ( .A(n541), .B(\mult_x_1/n284 ), .ZN(n176) );
  OAI22_X1 U69 ( .A1(n16), .A2(n49), .B1(n175), .B2(n176), .ZN(n225) );
  XNOR2_X1 U70 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n180) );
  OAI22_X1 U71 ( .A1(n181), .A2(n50), .B1(n179), .B2(n180), .ZN(n224) );
  OR2_X1 U72 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n51) );
  OAI22_X1 U73 ( .A1(n190), .A2(n25), .B1(n51), .B2(n188), .ZN(n57) );
  XNOR2_X1 U74 ( .A(n14), .B(\mult_x_1/n288 ), .ZN(n53) );
  OAI22_X1 U75 ( .A1(n190), .A2(n53), .B1(n188), .B2(n52), .ZN(n56) );
  XNOR2_X1 U76 ( .A(n156), .B(\mult_x_1/n283 ), .ZN(n79) );
  OAI22_X1 U77 ( .A1(n183), .A2(n79), .B1(n54), .B2(n24), .ZN(n105) );
  AND2_X1 U78 ( .A1(\mult_x_1/n288 ), .A2(n42), .ZN(n104) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n78) );
  OAI22_X1 U80 ( .A1(n181), .A2(n78), .B1(n179), .B2(n55), .ZN(n103) );
  HA_X1 U81 ( .A(n57), .B(n56), .CO(n223), .S(n97) );
  FA_X1 U82 ( .A(n60), .B(n59), .CI(n58), .CO(n235), .S(n96) );
  NAND2_X1 U83 ( .A1(n125), .A2(n124), .ZN(n61) );
  NAND2_X1 U84 ( .A1(n61), .A2(n262), .ZN(n63) );
  NAND2_X1 U85 ( .A1(n6), .A2(n327), .ZN(n62) );
  NAND2_X1 U86 ( .A1(n63), .A2(n62), .ZN(n356) );
  XNOR2_X1 U87 ( .A(n87), .B(n541), .ZN(n65) );
  XNOR2_X1 U88 ( .A(n541), .B(\mult_x_1/n281 ), .ZN(n73) );
  OAI22_X1 U89 ( .A1(n175), .A2(n65), .B1(n177), .B2(n73), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n69) );
  XNOR2_X1 U91 ( .A(n14), .B(\mult_x_1/n283 ), .ZN(n70) );
  XNOR2_X1 U92 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n64) );
  OAI22_X1 U93 ( .A1(n190), .A2(n70), .B1(n188), .B2(n64), .ZN(n68) );
  NOR2_X1 U94 ( .A1(n30), .A2(n185), .ZN(n67) );
  NOR2_X1 U95 ( .A1(n31), .A2(n185), .ZN(n93) );
  XNOR2_X1 U96 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n88) );
  OAI22_X1 U97 ( .A1(n190), .A2(n64), .B1(n188), .B2(n88), .ZN(n91) );
  AOI21_X1 U98 ( .B1(n175), .B2(n177), .A(n65), .ZN(n66) );
  INV_X1 U99 ( .A(n66), .ZN(n89) );
  FA_X1 U100 ( .A(n69), .B(n68), .CI(n67), .CO(n94), .S(n170) );
  XNOR2_X1 U101 ( .A(n14), .B(\mult_x_1/n284 ), .ZN(n74) );
  OAI22_X1 U102 ( .A1(n190), .A2(n74), .B1(n188), .B2(n70), .ZN(n195) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n178) );
  XNOR2_X1 U104 ( .A(n87), .B(\mult_x_1/n312 ), .ZN(n71) );
  AOI21_X1 U105 ( .B1(n179), .B2(n181), .A(n71), .ZN(n72) );
  INV_X1 U106 ( .A(n72), .ZN(n193) );
  NOR2_X1 U107 ( .A1(n32), .A2(n185), .ZN(n173) );
  XNOR2_X1 U108 ( .A(n541), .B(\mult_x_1/n282 ), .ZN(n75) );
  OAI22_X1 U109 ( .A1(n16), .A2(n75), .B1(n175), .B2(n73), .ZN(n172) );
  XNOR2_X1 U110 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n187) );
  OAI22_X1 U111 ( .A1(n190), .A2(n187), .B1(n188), .B2(n74), .ZN(n211) );
  XNOR2_X1 U112 ( .A(n541), .B(\mult_x_1/n283 ), .ZN(n174) );
  OAI22_X1 U113 ( .A1(n177), .A2(n174), .B1(n175), .B2(n75), .ZN(n210) );
  INV_X1 U114 ( .A(n194), .ZN(n209) );
  OAI21_X1 U115 ( .B1(n145), .B2(n144), .A(n237), .ZN(n77) );
  NAND2_X1 U116 ( .A1(n6), .A2(n323), .ZN(n76) );
  NAND2_X1 U117 ( .A1(n77), .A2(n76), .ZN(n348) );
  XNOR2_X1 U140 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n84) );
  OAI22_X1 U141 ( .A1(n181), .A2(n84), .B1(n179), .B2(n78), .ZN(n135) );
  XNOR2_X1 U142 ( .A(n156), .B(\mult_x_1/n284 ), .ZN(n82) );
  OAI22_X1 U143 ( .A1(n183), .A2(n82), .B1(n79), .B2(n24), .ZN(n134) );
  OR2_X1 U144 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n80) );
  OAI22_X1 U145 ( .A1(n16), .A2(n28), .B1(n80), .B2(n175), .ZN(n100) );
  XNOR2_X1 U146 ( .A(n23), .B(\mult_x_1/n288 ), .ZN(n81) );
  XNOR2_X1 U147 ( .A(n23), .B(\mult_x_1/n287 ), .ZN(n102) );
  OAI22_X1 U148 ( .A1(n16), .A2(n81), .B1(n175), .B2(n102), .ZN(n99) );
  XNOR2_X1 U149 ( .A(n156), .B(\mult_x_1/n285 ), .ZN(n152) );
  OAI22_X1 U150 ( .A1(n183), .A2(n152), .B1(n82), .B2(n24), .ZN(n149) );
  AND2_X1 U151 ( .A1(n83), .A2(\mult_x_1/n288 ), .ZN(n148) );
  XNOR2_X1 U152 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n150) );
  OAI22_X1 U153 ( .A1(n181), .A2(n150), .B1(n179), .B2(n84), .ZN(n147) );
  NOR2_X1 U154 ( .A1(n142), .A2(n141), .ZN(n86) );
  NAND2_X1 U155 ( .A1(n139), .A2(n320), .ZN(n85) );
  OAI21_X1 U156 ( .B1(n139), .B2(n86), .A(n85), .ZN(n342) );
  NOR2_X1 U157 ( .A1(n33), .A2(n185), .ZN(n109) );
  XNOR2_X1 U158 ( .A(n87), .B(n14), .ZN(n110) );
  OAI22_X1 U159 ( .A1(n190), .A2(n88), .B1(n110), .B2(n188), .ZN(n115) );
  INV_X1 U160 ( .A(n115), .ZN(n108) );
  FA_X1 U161 ( .A(n91), .B(n22), .CI(n89), .CO(n107), .S(n92) );
  FA_X1 U162 ( .A(n94), .B(n93), .CI(n92), .CO(n121), .S(n145) );
  OR2_X1 U163 ( .A1(n122), .A2(n121), .ZN(n95) );
  MUX2_X1 U164 ( .A(n321), .B(n95), .S(n262), .Z(n344) );
  FA_X1 U165 ( .A(n98), .B(n97), .CI(n96), .CO(n124), .S(n128) );
  HA_X1 U166 ( .A(n100), .B(n99), .CO(n132), .S(n133) );
  OAI22_X1 U167 ( .A1(n16), .A2(n102), .B1(n175), .B2(n101), .ZN(n131) );
  FA_X1 U168 ( .A(n105), .B(n104), .CI(n103), .CO(n98), .S(n130) );
  OR2_X1 U169 ( .A1(n128), .A2(n127), .ZN(n106) );
  MUX2_X1 U170 ( .A(n322), .B(n106), .S(n262), .Z(n346) );
  FA_X1 U171 ( .A(n109), .B(n108), .CI(n107), .CO(n117), .S(n122) );
  AOI21_X1 U172 ( .B1(n188), .B2(n190), .A(n110), .ZN(n111) );
  INV_X1 U173 ( .A(n111), .ZN(n113) );
  NOR2_X1 U174 ( .A1(n29), .A2(n185), .ZN(n112) );
  XOR2_X1 U175 ( .A(n113), .B(n112), .Z(n114) );
  XOR2_X1 U176 ( .A(n115), .B(n114), .Z(n116) );
  OR2_X1 U177 ( .A1(n117), .A2(n116), .ZN(n119) );
  NAND2_X1 U178 ( .A1(n117), .A2(n116), .ZN(n118) );
  NAND2_X1 U179 ( .A1(n119), .A2(n118), .ZN(n120) );
  MUX2_X1 U180 ( .A(n324), .B(n120), .S(n262), .Z(n350) );
  NAND2_X1 U181 ( .A1(n122), .A2(n121), .ZN(n123) );
  MUX2_X1 U182 ( .A(n325), .B(n123), .S(n262), .Z(n352) );
  NOR2_X1 U183 ( .A1(n125), .A2(n124), .ZN(n126) );
  MUX2_X1 U184 ( .A(n326), .B(n126), .S(n237), .Z(n354) );
  NAND2_X1 U185 ( .A1(n128), .A2(n127), .ZN(n129) );
  MUX2_X1 U186 ( .A(n328), .B(n129), .S(n262), .Z(n358) );
  FA_X1 U187 ( .A(n132), .B(n131), .CI(n130), .CO(n127), .S(n138) );
  FA_X1 U188 ( .A(n135), .B(n134), .CI(n133), .CO(n137), .S(n142) );
  NOR2_X1 U189 ( .A1(n138), .A2(n137), .ZN(n136) );
  MUX2_X1 U190 ( .A(n329), .B(n136), .S(n310), .Z(n360) );
  NAND2_X1 U191 ( .A1(n138), .A2(n137), .ZN(n140) );
  MUX2_X1 U192 ( .A(n330), .B(n140), .S(n237), .Z(n362) );
  NAND2_X1 U193 ( .A1(n142), .A2(n141), .ZN(n143) );
  MUX2_X1 U194 ( .A(n331), .B(n143), .S(n237), .Z(n364) );
  NAND2_X1 U195 ( .A1(n145), .A2(n144), .ZN(n146) );
  MUX2_X1 U196 ( .A(n332), .B(n146), .S(n237), .Z(n366) );
  FA_X1 U197 ( .A(n149), .B(n148), .CI(n147), .CO(n141), .S(n166) );
  XNOR2_X1 U198 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n151) );
  OAI22_X1 U199 ( .A1(n181), .A2(n151), .B1(n179), .B2(n150), .ZN(n154) );
  XNOR2_X1 U200 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n157) );
  OAI22_X1 U201 ( .A1(n183), .A2(n157), .B1(n152), .B2(n24), .ZN(n153) );
  NOR2_X1 U202 ( .A1(n166), .A2(n165), .ZN(n255) );
  HA_X1 U203 ( .A(n154), .B(n153), .CO(n165), .S(n163) );
  OR2_X1 U204 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n155) );
  OAI22_X1 U205 ( .A1(n181), .A2(n36), .B1(n155), .B2(n179), .ZN(n162) );
  OR2_X1 U206 ( .A1(n163), .A2(n162), .ZN(n251) );
  XNOR2_X1 U207 ( .A(n156), .B(\mult_x_1/n287 ), .ZN(n158) );
  OAI22_X1 U208 ( .A1(n183), .A2(n158), .B1(n157), .B2(n24), .ZN(n161) );
  AND2_X1 U209 ( .A1(\mult_x_1/n288 ), .A2(n48), .ZN(n160) );
  NOR2_X1 U210 ( .A1(n161), .A2(n160), .ZN(n244) );
  OAI22_X1 U211 ( .A1(n183), .A2(\mult_x_1/n288 ), .B1(n158), .B2(n24), .ZN(
        n241) );
  OR2_X1 U212 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n159) );
  NAND2_X1 U213 ( .A1(n159), .A2(n183), .ZN(n240) );
  NAND2_X1 U214 ( .A1(n241), .A2(n240), .ZN(n247) );
  NAND2_X1 U215 ( .A1(n161), .A2(n160), .ZN(n245) );
  OAI21_X1 U216 ( .B1(n244), .B2(n247), .A(n245), .ZN(n252) );
  NAND2_X1 U217 ( .A1(n163), .A2(n162), .ZN(n250) );
  INV_X1 U218 ( .A(n250), .ZN(n164) );
  AOI21_X1 U219 ( .B1(n251), .B2(n252), .A(n164), .ZN(n258) );
  NAND2_X1 U220 ( .A1(n166), .A2(n165), .ZN(n256) );
  OAI21_X1 U221 ( .B1(n255), .B2(n258), .A(n256), .ZN(n167) );
  MUX2_X1 U222 ( .A(n333), .B(n167), .S(n237), .Z(n368) );
  FA_X1 U223 ( .A(n173), .B(n172), .CI(n171), .CO(n168), .S(n202) );
  OAI22_X1 U224 ( .A1(n177), .A2(n176), .B1(n175), .B2(n174), .ZN(n208) );
  OAI22_X1 U225 ( .A1(n181), .A2(n180), .B1(n179), .B2(n178), .ZN(n207) );
  OR2_X1 U226 ( .A1(n208), .A2(n207), .ZN(n214) );
  NOR2_X1 U227 ( .A1(n34), .A2(n185), .ZN(n213) );
  OAI22_X1 U228 ( .A1(n190), .A2(n189), .B1(n188), .B2(n187), .ZN(n186) );
  AOI21_X1 U229 ( .B1(n183), .B2(n24), .A(n182), .ZN(n184) );
  INV_X1 U230 ( .A(n184), .ZN(n219) );
  NOR2_X1 U231 ( .A1(n35), .A2(n185), .ZN(n220) );
  OAI21_X1 U232 ( .B1(n186), .B2(n219), .A(n220), .ZN(n192) );
  OAI22_X1 U233 ( .A1(n190), .A2(n189), .B1(n188), .B2(n187), .ZN(n221) );
  NAND2_X1 U234 ( .A1(n221), .A2(n219), .ZN(n191) );
  NAND2_X1 U235 ( .A1(n192), .A2(n191), .ZN(n212) );
  FA_X1 U236 ( .A(n195), .B(n194), .CI(n193), .CO(n169), .S(n199) );
  NAND2_X1 U237 ( .A1(n202), .A2(n39), .ZN(n197) );
  NAND2_X1 U238 ( .A1(n200), .A2(n199), .ZN(n196) );
  NAND2_X1 U239 ( .A1(n197), .A2(n196), .ZN(n198) );
  MUX2_X1 U240 ( .A(n335), .B(n198), .S(n237), .Z(n372) );
  XNOR2_X1 U241 ( .A(n200), .B(n199), .ZN(n201) );
  XNOR2_X1 U242 ( .A(n202), .B(n201), .ZN(n203) );
  MUX2_X1 U243 ( .A(n336), .B(n203), .S(n237), .Z(n374) );
  FA_X1 U244 ( .A(n206), .B(n205), .CI(n204), .CO(n227), .S(n236) );
  XNOR2_X1 U245 ( .A(n208), .B(n207), .ZN(n226) );
  FA_X1 U246 ( .A(n211), .B(n210), .CI(n209), .CO(n171), .S(n217) );
  FA_X1 U247 ( .A(n214), .B(n213), .CI(n212), .CO(n200), .S(n216) );
  MUX2_X1 U248 ( .A(n337), .B(n215), .S(n237), .Z(n376) );
  FA_X1 U249 ( .A(n27), .B(n217), .CI(n216), .CO(n215), .S(n218) );
  MUX2_X1 U250 ( .A(n338), .B(n218), .S(n237), .Z(n378) );
  FA_X1 U251 ( .A(n225), .B(n224), .CI(n223), .CO(n231), .S(n234) );
  INV_X1 U252 ( .A(n226), .ZN(n228) );
  XNOR2_X1 U253 ( .A(n228), .B(n227), .ZN(n230) );
  MUX2_X1 U254 ( .A(n339), .B(n229), .S(n237), .Z(n380) );
  FA_X1 U255 ( .A(n232), .B(n231), .CI(n230), .CO(n229), .S(n233) );
  MUX2_X1 U256 ( .A(n340), .B(n233), .S(n237), .Z(n382) );
  MUX2_X1 U257 ( .A(n341), .B(n238), .S(n237), .Z(n384) );
  MUX2_X1 U258 ( .A(product[0]), .B(n505), .S(n262), .Z(n397) );
  MUX2_X1 U259 ( .A(n505), .B(n506), .S(n262), .Z(n399) );
  AND2_X1 U260 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n239) );
  MUX2_X1 U261 ( .A(n506), .B(n239), .S(n262), .Z(n401) );
  MUX2_X1 U262 ( .A(product[1]), .B(n508), .S(n262), .Z(n403) );
  MUX2_X1 U263 ( .A(n508), .B(n509), .S(n262), .Z(n405) );
  OR2_X1 U264 ( .A1(n241), .A2(n240), .ZN(n242) );
  AND2_X1 U265 ( .A1(n242), .A2(n247), .ZN(n243) );
  MUX2_X1 U266 ( .A(n509), .B(n243), .S(n262), .Z(n407) );
  MUX2_X1 U267 ( .A(product[2]), .B(n511), .S(n262), .Z(n409) );
  MUX2_X1 U268 ( .A(n511), .B(n512), .S(n262), .Z(n411) );
  INV_X1 U269 ( .A(n244), .ZN(n246) );
  NAND2_X1 U270 ( .A1(n246), .A2(n245), .ZN(n248) );
  XOR2_X1 U271 ( .A(n248), .B(n247), .Z(n249) );
  MUX2_X1 U272 ( .A(n512), .B(n249), .S(n262), .Z(n413) );
  MUX2_X1 U273 ( .A(product[3]), .B(n514), .S(n262), .Z(n415) );
  MUX2_X1 U274 ( .A(n514), .B(n515), .S(n262), .Z(n417) );
  NAND2_X1 U275 ( .A1(n251), .A2(n250), .ZN(n253) );
  XNOR2_X1 U276 ( .A(n253), .B(n252), .ZN(n254) );
  MUX2_X1 U277 ( .A(n515), .B(n254), .S(n262), .Z(n419) );
  MUX2_X1 U278 ( .A(product[4]), .B(n517), .S(n262), .Z(n421) );
  MUX2_X1 U279 ( .A(n517), .B(n518), .S(n262), .Z(n423) );
  INV_X1 U280 ( .A(n255), .ZN(n257) );
  NAND2_X1 U281 ( .A1(n257), .A2(n256), .ZN(n259) );
  XOR2_X1 U282 ( .A(n259), .B(n258), .Z(n260) );
  MUX2_X1 U283 ( .A(n518), .B(n260), .S(n262), .Z(n425) );
  MUX2_X1 U284 ( .A(product[5]), .B(n520), .S(n262), .Z(n427) );
  NAND2_X1 U285 ( .A1(n320), .A2(n331), .ZN(n261) );
  XNOR2_X1 U286 ( .A(n261), .B(n333), .ZN(n263) );
  MUX2_X1 U287 ( .A(n520), .B(n263), .S(n262), .Z(n429) );
  BUF_X4 U288 ( .A(en), .Z(n310) );
  MUX2_X1 U289 ( .A(product[6]), .B(n522), .S(n310), .Z(n431) );
  NAND2_X1 U290 ( .A1(n389), .A2(n330), .ZN(n264) );
  AOI21_X1 U291 ( .B1(n320), .B2(n333), .A(n391), .ZN(n266) );
  XOR2_X1 U292 ( .A(n264), .B(n266), .Z(n265) );
  MUX2_X1 U293 ( .A(n522), .B(n265), .S(n310), .Z(n433) );
  MUX2_X1 U294 ( .A(product[7]), .B(n524), .S(n310), .Z(n435) );
  OAI21_X1 U295 ( .B1(n329), .B2(n266), .A(n330), .ZN(n269) );
  NAND2_X1 U296 ( .A1(n322), .A2(n328), .ZN(n267) );
  XNOR2_X1 U297 ( .A(n269), .B(n267), .ZN(n268) );
  MUX2_X1 U298 ( .A(n524), .B(n268), .S(n310), .Z(n437) );
  MUX2_X1 U299 ( .A(product[8]), .B(n526), .S(n310), .Z(n439) );
  AOI21_X1 U300 ( .B1(n269), .B2(n322), .A(n390), .ZN(n272) );
  NAND2_X1 U301 ( .A1(n392), .A2(n327), .ZN(n270) );
  XOR2_X1 U302 ( .A(n272), .B(n270), .Z(n271) );
  MUX2_X1 U303 ( .A(n526), .B(n271), .S(n310), .Z(n441) );
  MUX2_X1 U304 ( .A(product[9]), .B(n528), .S(n310), .Z(n443) );
  OAI21_X1 U305 ( .B1(n272), .B2(n326), .A(n327), .ZN(n286) );
  INV_X1 U306 ( .A(n286), .ZN(n276) );
  NOR2_X1 U307 ( .A1(n340), .A2(n341), .ZN(n281) );
  INV_X1 U308 ( .A(n281), .ZN(n273) );
  NAND2_X1 U309 ( .A1(n340), .A2(n341), .ZN(n283) );
  NAND2_X1 U310 ( .A1(n273), .A2(n283), .ZN(n274) );
  XOR2_X1 U311 ( .A(n276), .B(n274), .Z(n275) );
  MUX2_X1 U312 ( .A(n528), .B(n275), .S(n310), .Z(n445) );
  MUX2_X1 U313 ( .A(product[10]), .B(n530), .S(n310), .Z(n447) );
  OAI21_X1 U314 ( .B1(n276), .B2(n281), .A(n283), .ZN(n279) );
  NOR2_X1 U315 ( .A1(n338), .A2(n339), .ZN(n284) );
  INV_X1 U316 ( .A(n284), .ZN(n277) );
  NAND2_X1 U317 ( .A1(n338), .A2(n339), .ZN(n282) );
  NAND2_X1 U318 ( .A1(n277), .A2(n282), .ZN(n278) );
  XNOR2_X1 U319 ( .A(n279), .B(n278), .ZN(n280) );
  MUX2_X1 U320 ( .A(n530), .B(n280), .S(n310), .Z(n449) );
  MUX2_X1 U321 ( .A(product[11]), .B(n532), .S(n310), .Z(n451) );
  NOR2_X1 U322 ( .A1(n284), .A2(n281), .ZN(n287) );
  OAI21_X1 U323 ( .B1(n284), .B2(n283), .A(n282), .ZN(n285) );
  AOI21_X1 U324 ( .B1(n287), .B2(n286), .A(n285), .ZN(n317) );
  NOR2_X1 U325 ( .A1(n336), .A2(n337), .ZN(n301) );
  INV_X1 U326 ( .A(n301), .ZN(n313) );
  NAND2_X1 U327 ( .A1(n336), .A2(n337), .ZN(n304) );
  NAND2_X1 U328 ( .A1(n313), .A2(n304), .ZN(n288) );
  XOR2_X1 U329 ( .A(n317), .B(n288), .Z(n289) );
  MUX2_X1 U330 ( .A(n532), .B(n289), .S(n310), .Z(n453) );
  MUX2_X1 U331 ( .A(product[12]), .B(n534), .S(n310), .Z(n455) );
  OAI21_X1 U332 ( .B1(n317), .B2(n301), .A(n304), .ZN(n291) );
  OR2_X1 U333 ( .A1(n334), .A2(n335), .ZN(n300) );
  NAND2_X1 U334 ( .A1(n334), .A2(n335), .ZN(n293) );
  NAND2_X1 U335 ( .A1(n300), .A2(n293), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n292) );
  MUX2_X1 U337 ( .A(n534), .B(n292), .S(n310), .Z(n457) );
  MUX2_X1 U338 ( .A(product[13]), .B(n536), .S(n310), .Z(n459) );
  NAND2_X1 U339 ( .A1(n313), .A2(n300), .ZN(n296) );
  INV_X1 U340 ( .A(n304), .ZN(n294) );
  INV_X1 U341 ( .A(n293), .ZN(n302) );
  AOI21_X1 U342 ( .B1(n294), .B2(n300), .A(n302), .ZN(n295) );
  OAI21_X1 U343 ( .B1(n317), .B2(n296), .A(n295), .ZN(n298) );
  NAND2_X1 U344 ( .A1(n323), .A2(n332), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  MUX2_X1 U346 ( .A(n536), .B(n299), .S(n310), .Z(n461) );
  MUX2_X1 U347 ( .A(product[14]), .B(n538), .S(n310), .Z(n463) );
  NAND2_X1 U348 ( .A1(n300), .A2(n323), .ZN(n311) );
  OR2_X1 U349 ( .A1(n301), .A2(n311), .ZN(n306) );
  AOI21_X1 U350 ( .B1(n302), .B2(n323), .A(n387), .ZN(n303) );
  OAI21_X1 U351 ( .B1(n311), .B2(n304), .A(n303), .ZN(n314) );
  INV_X1 U352 ( .A(n314), .ZN(n305) );
  OAI21_X1 U353 ( .B1(n317), .B2(n306), .A(n305), .ZN(n308) );
  NAND2_X1 U354 ( .A1(n321), .A2(n325), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U356 ( .A(n538), .B(n309), .S(n310), .Z(n465) );
  MUX2_X1 U357 ( .A(product[15]), .B(n540), .S(n310), .Z(n467) );
  NOR2_X1 U358 ( .A1(n311), .A2(n388), .ZN(n312) );
  NAND2_X1 U359 ( .A1(n313), .A2(n312), .ZN(n316) );
  AOI21_X1 U360 ( .B1(n314), .B2(n321), .A(n386), .ZN(n315) );
  OAI21_X1 U361 ( .B1(n317), .B2(n316), .A(n315), .ZN(n318) );
  XNOR2_X1 U362 ( .A(n318), .B(n324), .ZN(n319) );
  MUX2_X1 U363 ( .A(n540), .B(n319), .S(n310), .Z(n469) );
  MUX2_X1 U364 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n310), .Z(n471) );
  MUX2_X1 U365 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n310), .Z(n473) );
  MUX2_X1 U366 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n310), .Z(n475) );
  MUX2_X1 U367 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n310), .Z(n477) );
  MUX2_X1 U368 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n310), .Z(n479) );
  MUX2_X1 U369 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n310), .Z(n481) );
  MUX2_X1 U370 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n310), .Z(n483) );
  MUX2_X1 U371 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n310), .Z(n485) );
  MUX2_X1 U372 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n310), .Z(n487) );
  MUX2_X1 U373 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n310), .Z(n489) );
  MUX2_X1 U374 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n310), .Z(n491) );
  MUX2_X1 U375 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n310), .Z(n493) );
  MUX2_X1 U376 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n310), .Z(n495) );
  MUX2_X1 U377 ( .A(n23), .B(A_extended[5]), .S(n310), .Z(n497) );
  MUX2_X1 U378 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n310), .Z(n499) );
  MUX2_X1 U379 ( .A(n14), .B(A_extended[7]), .S(n310), .Z(n501) );
  OR2_X1 U380 ( .A1(n262), .A2(n542), .ZN(n503) );
endmodule


module conv_128_32_DW_mult_pipe_J1_12 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n357, n359, n361, n363, n365, n367, n369, n370,
         n372, n374, n376, n378, n380, n382, n384, n386, n388, n390, n392,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n409, n411, n413, n415, n417, n419, n421, n423,
         n425, n427, n429, n431, n433, n435, n437, n439, n441, n443, n445,
         n447, n449, n451, n453, n455, n457, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n515, n517, n519, n520, n522, n523, n525, n526, n528, n529,
         n531, n532, n534, n535, n537, n539, n541, n543, n545, n547, n549,
         n551, n553, n555, n556, n557, n558, n559;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n407), .SE(n513), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n18) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n407), .SE(n511), .CK(clk), .Q(n557), 
        .QN(n27) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n407), .SE(n509), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n332) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n407), .SE(n505), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n19) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n407), .SE(n503), .CK(clk), .Q(n556), 
        .QN(n28) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n407), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n26) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n407), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n407), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n405), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n406), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n404), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n407), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n404), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n404), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n404), .SE(n483), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n404), .SE(n481), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n404), .SE(n479), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n404), .SE(n477), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n404), .SE(n475), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n406), .SE(n473), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n405), .SE(n471), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n407), .SE(n469), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n404), .SE(n467), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n404), .SE(n465), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n404), .SE(n463), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n404), .SE(n461), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n404), .SE(n459), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n404), .SE(n457), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n404), .SE(n455), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n404), .SE(n453), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n406), .SE(n451), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n406), .SE(n449), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n406), .SE(n447), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n406), .SE(n445), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n406), .SE(n443), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n406), .SE(n441), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n406), .SE(n439), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n406), .SE(n437), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n406), .SE(n435), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n406), .SE(n433), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n406), .SE(n431), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n405), .SE(n429), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n405), .SE(n427), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n405), .SE(n425), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n405), .SE(n423), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n405), .SE(n421), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n405), .SE(n419), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n405), .SE(n417), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n405), .SE(n415), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n405), .SE(n413), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n405), .SE(n411), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n405), .SE(n409), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n559), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2_IP  ( .D(1'b1), .SI(n559), .SE(n390), .CK(
        clk), .Q(n402), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n559), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n352), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2  ( .D(n559), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n559), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2_IP  ( .D(1'b1), .SI(n559), .SE(n382), .CK(
        clk), .Q(n401), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n559), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n348), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n559), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n559), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n346), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n559), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n345), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n559), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n559), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n343), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n559), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n341), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n559), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n340), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n559), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n339), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n559), .SE(n361), .CK(
        clk), .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n559), .SE(n359), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n559), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n559), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n335) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n407), .SE(n517), .CK(clk), .Q(n558), 
        .QN(n333) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n407), .SE(n515), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n334) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n407), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n559), .SE(n369), .CK(
        clk), .QN(n342) );
  BUF_X1 U2 ( .A(n404), .Z(n406) );
  BUF_X1 U3 ( .A(n404), .Z(n405) );
  BUF_X1 U4 ( .A(n404), .Z(n407) );
  INV_X1 U5 ( .A(n559), .ZN(n404) );
  INV_X1 U6 ( .A(n46), .ZN(n245) );
  NOR2_X1 U7 ( .A1(n334), .A2(n333), .ZN(n22) );
  BUF_X1 U8 ( .A(en), .Z(n219) );
  BUF_X2 U9 ( .A(en), .Z(n24) );
  OAI21_X1 U10 ( .B1(n16), .B2(n15), .A(n14), .ZN(n138) );
  AND3_X1 U11 ( .A1(n121), .A2(n120), .A3(n119), .ZN(n124) );
  INV_X1 U12 ( .A(n96), .ZN(n16) );
  NAND2_X1 U13 ( .A1(n7), .A2(n6), .ZN(n221) );
  NAND2_X1 U14 ( .A1(n98), .A2(n97), .ZN(n14) );
  NAND2_X1 U15 ( .A1(n227), .A2(n8), .ZN(n7) );
  NOR2_X1 U16 ( .A1(n97), .A2(n98), .ZN(n15) );
  NAND2_X1 U17 ( .A1(n229), .A2(n228), .ZN(n6) );
  OR2_X1 U18 ( .A1(n229), .A2(n228), .ZN(n8) );
  INV_X1 U19 ( .A(rst_n), .ZN(n559) );
  INV_X1 U20 ( .A(n31), .ZN(n231) );
  NAND2_X1 U21 ( .A1(n29), .A2(n30), .ZN(n172) );
  NAND2_X1 U22 ( .A1(n32), .A2(n33), .ZN(n181) );
  AND2_X1 U23 ( .A1(n558), .A2(\mult_x_1/n281 ), .ZN(n152) );
  XNOR2_X1 U24 ( .A(n227), .B(n9), .ZN(n258) );
  XNOR2_X1 U25 ( .A(n229), .B(n228), .ZN(n9) );
  OAI21_X1 U26 ( .B1(n12), .B2(n11), .A(n10), .ZN(n443) );
  NAND2_X1 U27 ( .A1(n11), .A2(n535), .ZN(n10) );
  INV_X1 U28 ( .A(n329), .ZN(n11) );
  XNOR2_X1 U29 ( .A(n286), .B(n13), .ZN(n12) );
  INV_X1 U30 ( .A(n285), .ZN(n13) );
  XNOR2_X1 U31 ( .A(\mult_x_1/a[4] ), .B(n331), .ZN(n31) );
  XNOR2_X1 U32 ( .A(n96), .B(n17), .ZN(n92) );
  XNOR2_X1 U33 ( .A(n98), .B(n97), .ZN(n17) );
  NOR2_X1 U34 ( .A1(n334), .A2(n333), .ZN(n35) );
  CLKBUF_X1 U35 ( .A(n331), .Z(n20) );
  XNOR2_X1 U36 ( .A(n105), .B(n104), .ZN(n136) );
  XNOR2_X1 U37 ( .A(n103), .B(n102), .ZN(n104) );
  NAND2_X1 U38 ( .A1(n146), .A2(n145), .ZN(n384) );
  NAND2_X1 U39 ( .A1(n128), .A2(n350), .ZN(n145) );
  OAI21_X1 U40 ( .B1(n144), .B2(n143), .A(n24), .ZN(n146) );
  NAND2_X1 U41 ( .A1(n124), .A2(n24), .ZN(n122) );
  NAND2_X1 U42 ( .A1(n140), .A2(n352), .ZN(n125) );
  NAND2_X1 U43 ( .A1(n124), .A2(n24), .ZN(n126) );
  XNOR2_X1 U44 ( .A(n18), .B(n27), .ZN(n33) );
  XNOR2_X1 U45 ( .A(\mult_x_1/a[2] ), .B(n331), .ZN(n48) );
  XNOR2_X1 U46 ( .A(n19), .B(n28), .ZN(n47) );
  BUF_X1 U47 ( .A(\mult_x_1/n310 ), .Z(n21) );
  CLKBUF_X1 U48 ( .A(n184), .Z(n23) );
  XNOR2_X1 U49 ( .A(n35), .B(\mult_x_1/n310 ), .ZN(n184) );
  INV_X1 U50 ( .A(n81), .ZN(n25) );
  CLKBUF_X1 U51 ( .A(n238), .Z(n243) );
  OAI22_X1 U52 ( .A1(n245), .A2(n49), .B1(n238), .B2(n69), .ZN(n100) );
  BUF_X4 U53 ( .A(en), .Z(n329) );
  XOR2_X1 U55 ( .A(\mult_x_1/a[4] ), .B(n557), .Z(n29) );
  XNOR2_X1 U56 ( .A(n331), .B(n332), .ZN(n30) );
  BUF_X1 U57 ( .A(n557), .Z(n328) );
  XNOR2_X1 U58 ( .A(n328), .B(\mult_x_1/n281 ), .ZN(n53) );
  XNOR2_X1 U59 ( .A(n152), .B(n328), .ZN(n39) );
  OAI22_X1 U60 ( .A1(n172), .A2(n53), .B1(n39), .B2(n231), .ZN(n41) );
  INV_X1 U61 ( .A(n41), .ZN(n44) );
  XOR2_X1 U62 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n32) );
  XNOR2_X1 U63 ( .A(n21), .B(\mult_x_1/n283 ), .ZN(n45) );
  INV_X1 U64 ( .A(n33), .ZN(n34) );
  INV_X2 U65 ( .A(n34), .ZN(n182) );
  XNOR2_X1 U66 ( .A(n21), .B(\mult_x_1/n282 ), .ZN(n38) );
  OAI22_X1 U67 ( .A1(n181), .A2(n45), .B1(n182), .B2(n38), .ZN(n43) );
  XNOR2_X1 U68 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n36) );
  NOR2_X1 U69 ( .A1(n36), .A2(n23), .ZN(n42) );
  XNOR2_X1 U70 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n37) );
  NOR2_X1 U71 ( .A1(n37), .A2(n23), .ZN(n157) );
  XNOR2_X1 U72 ( .A(n21), .B(\mult_x_1/n281 ), .ZN(n153) );
  OAI22_X1 U73 ( .A1(n181), .A2(n38), .B1(n182), .B2(n153), .ZN(n155) );
  AOI21_X1 U74 ( .B1(n231), .B2(n172), .A(n39), .ZN(n40) );
  INV_X1 U75 ( .A(n40), .ZN(n154) );
  FA_X1 U76 ( .A(n44), .B(n43), .CI(n42), .CO(n158), .S(n135) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n51) );
  OAI22_X1 U78 ( .A1(n181), .A2(n51), .B1(n182), .B2(n45), .ZN(n101) );
  INV_X1 U79 ( .A(n47), .ZN(n46) );
  XNOR2_X1 U80 ( .A(n152), .B(\mult_x_1/n312 ), .ZN(n49) );
  NAND2_X1 U81 ( .A1(n48), .A2(n47), .ZN(n238) );
  XNOR2_X1 U82 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n69) );
  AOI21_X1 U83 ( .B1(n245), .B2(n243), .A(n49), .ZN(n50) );
  INV_X1 U84 ( .A(n50), .ZN(n99) );
  XNOR2_X1 U85 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n64) );
  OAI22_X1 U86 ( .A1(n181), .A2(n64), .B1(n182), .B2(n51), .ZN(n83) );
  XNOR2_X1 U87 ( .A(n557), .B(\mult_x_1/n283 ), .ZN(n67) );
  XNOR2_X1 U88 ( .A(n557), .B(\mult_x_1/n282 ), .ZN(n54) );
  OAI22_X1 U89 ( .A1(n172), .A2(n67), .B1(n231), .B2(n54), .ZN(n82) );
  INV_X1 U90 ( .A(n100), .ZN(n81) );
  XNOR2_X1 U91 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n52) );
  NOR2_X1 U92 ( .A1(n52), .A2(n23), .ZN(n103) );
  INV_X1 U93 ( .A(n103), .ZN(n56) );
  OAI22_X1 U94 ( .A1(n172), .A2(n54), .B1(n231), .B2(n53), .ZN(n102) );
  INV_X1 U95 ( .A(n102), .ZN(n55) );
  NAND2_X1 U96 ( .A1(n56), .A2(n55), .ZN(n57) );
  AOI22_X1 U97 ( .A1(n105), .A2(n57), .B1(n102), .B2(n103), .ZN(n58) );
  INV_X1 U98 ( .A(n58), .ZN(n133) );
  OR2_X1 U99 ( .A1(n225), .A2(n224), .ZN(n59) );
  NAND2_X1 U100 ( .A1(n59), .A2(n24), .ZN(n61) );
  NAND2_X1 U101 ( .A1(n128), .A2(n336), .ZN(n60) );
  NAND2_X1 U102 ( .A1(n61), .A2(n60), .ZN(n357) );
  NAND2_X1 U103 ( .A1(n556), .A2(n26), .ZN(n248) );
  XNOR2_X1 U104 ( .A(n152), .B(n556), .ZN(n74) );
  AOI21_X1 U105 ( .B1(n248), .B2(n26), .A(n74), .ZN(n62) );
  INV_X1 U106 ( .A(n62), .ZN(n89) );
  XNOR2_X1 U107 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n63) );
  NOR2_X1 U108 ( .A1(n63), .A2(n184), .ZN(n88) );
  XNOR2_X1 U109 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n75) );
  OAI22_X1 U110 ( .A1(n181), .A2(n75), .B1(n182), .B2(n64), .ZN(n87) );
  XNOR2_X1 U111 ( .A(n328), .B(\mult_x_1/n285 ), .ZN(n116) );
  XNOR2_X1 U112 ( .A(n328), .B(\mult_x_1/n284 ), .ZN(n68) );
  OAI22_X1 U113 ( .A1(n172), .A2(n116), .B1(n231), .B2(n68), .ZN(n112) );
  XNOR2_X1 U114 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n118) );
  XNOR2_X1 U115 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n70) );
  OAI22_X1 U116 ( .A1(n238), .A2(n118), .B1(n245), .B2(n70), .ZN(n111) );
  XNOR2_X1 U117 ( .A(n21), .B(\mult_x_1/n288 ), .ZN(n65) );
  XNOR2_X1 U118 ( .A(n21), .B(\mult_x_1/n287 ), .ZN(n76) );
  OAI22_X1 U119 ( .A1(n181), .A2(n65), .B1(n182), .B2(n76), .ZN(n164) );
  OR2_X1 U120 ( .A1(\mult_x_1/n288 ), .A2(n334), .ZN(n66) );
  OAI22_X1 U121 ( .A1(n181), .A2(n334), .B1(n66), .B2(n182), .ZN(n163) );
  OAI22_X1 U122 ( .A1(n172), .A2(n68), .B1(n231), .B2(n67), .ZN(n85) );
  OAI22_X1 U123 ( .A1(n238), .A2(n70), .B1(n245), .B2(n69), .ZN(n84) );
  XNOR2_X1 U124 ( .A(n85), .B(n84), .ZN(n80) );
  INV_X1 U125 ( .A(n22), .ZN(n71) );
  OR2_X1 U126 ( .A1(\mult_x_1/n288 ), .A2(n71), .ZN(n72) );
  NOR2_X1 U127 ( .A1(n72), .A2(n23), .ZN(n79) );
  INV_X1 U128 ( .A(n184), .ZN(n73) );
  AND2_X1 U129 ( .A1(\mult_x_1/n288 ), .A2(n73), .ZN(n115) );
  XNOR2_X1 U130 ( .A(n556), .B(\mult_x_1/n281 ), .ZN(n117) );
  OAI22_X1 U131 ( .A1(n248), .A2(n117), .B1(n74), .B2(n26), .ZN(n114) );
  OAI22_X1 U132 ( .A1(n181), .A2(n76), .B1(n182), .B2(n75), .ZN(n113) );
  INV_X1 U133 ( .A(n77), .ZN(n129) );
  NAND2_X1 U134 ( .A1(n129), .A2(n24), .ZN(n91) );
  FA_X1 U135 ( .A(n80), .B(n79), .CI(n78), .CO(n94), .S(n107) );
  FA_X1 U136 ( .A(n83), .B(n82), .CI(n81), .CO(n105), .S(n93) );
  OR2_X1 U137 ( .A1(n85), .A2(n84), .ZN(n98) );
  XNOR2_X1 U138 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n86) );
  NOR2_X1 U139 ( .A1(n86), .A2(n23), .ZN(n97) );
  FA_X1 U140 ( .A(n89), .B(n88), .CI(n87), .CO(n96), .S(n109) );
  NAND2_X1 U141 ( .A1(n140), .A2(n349), .ZN(n90) );
  OAI21_X1 U142 ( .B1(n91), .B2(n132), .A(n90), .ZN(n382) );
  FA_X1 U143 ( .A(n94), .B(n93), .CI(n92), .CO(n95), .S(n132) );
  INV_X1 U144 ( .A(n95), .ZN(n147) );
  NAND2_X1 U145 ( .A1(n147), .A2(n329), .ZN(n106) );
  FA_X1 U146 ( .A(n101), .B(n25), .CI(n99), .CO(n134), .S(n137) );
  OAI22_X1 U147 ( .A1(n106), .A2(n150), .B1(n329), .B2(n402), .ZN(n390) );
  FA_X1 U148 ( .A(n109), .B(n108), .CI(n107), .CO(n77), .S(n127) );
  NAND2_X1 U149 ( .A1(n140), .A2(n351), .ZN(n123) );
  FA_X1 U150 ( .A(n112), .B(n111), .CI(n110), .CO(n108), .S(n201) );
  FA_X1 U151 ( .A(n115), .B(n114), .CI(n113), .CO(n78), .S(n199) );
  NAND2_X1 U152 ( .A1(n201), .A2(n199), .ZN(n121) );
  XNOR2_X1 U153 ( .A(n328), .B(\mult_x_1/n286 ), .ZN(n170) );
  OAI22_X1 U154 ( .A1(n172), .A2(n170), .B1(n231), .B2(n116), .ZN(n167) );
  XNOR2_X1 U155 ( .A(n556), .B(\mult_x_1/n282 ), .ZN(n160) );
  OAI22_X1 U156 ( .A1(n248), .A2(n160), .B1(n117), .B2(n26), .ZN(n166) );
  XNOR2_X1 U157 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n162) );
  OAI22_X1 U158 ( .A1(n238), .A2(n162), .B1(n245), .B2(n118), .ZN(n165) );
  NAND2_X1 U159 ( .A1(n201), .A2(n198), .ZN(n120) );
  NAND2_X1 U160 ( .A1(n199), .A2(n198), .ZN(n119) );
  OAI211_X1 U161 ( .C1(n127), .C2(n140), .A(n123), .B(n122), .ZN(n386) );
  OAI21_X1 U162 ( .B1(n127), .B2(n126), .A(n125), .ZN(n388) );
  INV_X1 U163 ( .A(n219), .ZN(n128) );
  NAND2_X1 U164 ( .A1(n128), .A2(n342), .ZN(n131) );
  NAND2_X1 U165 ( .A1(n129), .A2(n24), .ZN(n130) );
  OAI211_X1 U166 ( .C1(n132), .C2(n128), .A(n131), .B(n130), .ZN(n369) );
  FA_X1 U167 ( .A(n135), .B(n134), .CI(n133), .CO(n224), .S(n144) );
  FA_X1 U168 ( .A(n138), .B(n137), .CI(n136), .CO(n143), .S(n150) );
  NAND2_X1 U169 ( .A1(n144), .A2(n143), .ZN(n139) );
  NAND2_X1 U170 ( .A1(n139), .A2(n329), .ZN(n142) );
  INV_X1 U171 ( .A(n219), .ZN(n140) );
  NAND2_X1 U172 ( .A1(n140), .A2(n340), .ZN(n141) );
  NAND2_X1 U173 ( .A1(n142), .A2(n141), .ZN(n365) );
  NAND2_X1 U174 ( .A1(n128), .A2(n341), .ZN(n149) );
  NAND2_X1 U175 ( .A1(n147), .A2(n329), .ZN(n148) );
  OAI211_X1 U176 ( .C1(n150), .C2(n140), .A(n149), .B(n148), .ZN(n367) );
  XNOR2_X1 U196 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n151) );
  NOR2_X1 U197 ( .A1(n151), .A2(n23), .ZN(n179) );
  XNOR2_X1 U198 ( .A(n152), .B(n21), .ZN(n180) );
  OAI22_X1 U199 ( .A1(n181), .A2(n153), .B1(n180), .B2(n182), .ZN(n189) );
  INV_X1 U200 ( .A(n189), .ZN(n178) );
  FA_X1 U201 ( .A(n155), .B(n154), .CI(n41), .CO(n177), .S(n156) );
  FA_X1 U202 ( .A(n158), .B(n157), .CI(n156), .CO(n195), .S(n225) );
  OR2_X1 U203 ( .A1(n196), .A2(n195), .ZN(n159) );
  MUX2_X1 U204 ( .A(n335), .B(n159), .S(n329), .Z(n355) );
  XNOR2_X1 U205 ( .A(n556), .B(\mult_x_1/n283 ), .ZN(n216) );
  OAI22_X1 U206 ( .A1(n248), .A2(n216), .B1(n160), .B2(n26), .ZN(n175) );
  INV_X1 U207 ( .A(n182), .ZN(n161) );
  AND2_X1 U208 ( .A1(\mult_x_1/n288 ), .A2(n161), .ZN(n174) );
  XNOR2_X1 U209 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n215) );
  OAI22_X1 U210 ( .A1(n243), .A2(n215), .B1(n245), .B2(n162), .ZN(n173) );
  HA_X1 U211 ( .A(n164), .B(n163), .CO(n110), .S(n203) );
  FA_X1 U212 ( .A(n167), .B(n166), .CI(n165), .CO(n198), .S(n202) );
  OR2_X1 U213 ( .A1(\mult_x_1/n288 ), .A2(n27), .ZN(n168) );
  OAI22_X1 U214 ( .A1(n172), .A2(n27), .B1(n168), .B2(n231), .ZN(n218) );
  XNOR2_X1 U215 ( .A(n328), .B(\mult_x_1/n288 ), .ZN(n169) );
  XNOR2_X1 U216 ( .A(n557), .B(\mult_x_1/n287 ), .ZN(n171) );
  OAI22_X1 U217 ( .A1(n172), .A2(n169), .B1(n231), .B2(n171), .ZN(n217) );
  OAI22_X1 U218 ( .A1(n172), .A2(n171), .B1(n231), .B2(n170), .ZN(n213) );
  FA_X1 U219 ( .A(n175), .B(n174), .CI(n173), .CO(n204), .S(n212) );
  OR2_X1 U220 ( .A1(n210), .A2(n209), .ZN(n176) );
  MUX2_X1 U221 ( .A(n337), .B(n176), .S(n219), .Z(n359) );
  FA_X1 U222 ( .A(n179), .B(n178), .CI(n177), .CO(n191), .S(n196) );
  AOI21_X1 U223 ( .B1(n182), .B2(n181), .A(n180), .ZN(n183) );
  INV_X1 U224 ( .A(n183), .ZN(n187) );
  XNOR2_X1 U225 ( .A(n22), .B(\mult_x_1/n281 ), .ZN(n185) );
  NOR2_X1 U226 ( .A1(n185), .A2(n23), .ZN(n186) );
  XOR2_X1 U227 ( .A(n187), .B(n186), .Z(n188) );
  XOR2_X1 U228 ( .A(n189), .B(n188), .Z(n190) );
  OR2_X1 U229 ( .A1(n191), .A2(n190), .ZN(n193) );
  NAND2_X1 U230 ( .A1(n191), .A2(n190), .ZN(n192) );
  NAND2_X1 U231 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U232 ( .A(n338), .B(n194), .S(n219), .Z(n361) );
  NAND2_X1 U233 ( .A1(n196), .A2(n195), .ZN(n197) );
  MUX2_X1 U234 ( .A(n339), .B(n197), .S(n329), .Z(n363) );
  XOR2_X1 U235 ( .A(n199), .B(n198), .Z(n200) );
  XOR2_X1 U236 ( .A(n201), .B(n200), .Z(n207) );
  FA_X1 U237 ( .A(n204), .B(n203), .CI(n202), .CO(n206), .S(n210) );
  NOR2_X1 U238 ( .A1(n207), .A2(n206), .ZN(n205) );
  MUX2_X1 U239 ( .A(n343), .B(n205), .S(n24), .Z(n370) );
  NAND2_X1 U240 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U241 ( .A(n344), .B(n208), .S(n329), .Z(n372) );
  NAND2_X1 U242 ( .A1(n210), .A2(n209), .ZN(n211) );
  MUX2_X1 U243 ( .A(n345), .B(n211), .S(n24), .Z(n374) );
  FA_X1 U244 ( .A(n214), .B(n213), .CI(n212), .CO(n209), .S(n222) );
  XNOR2_X1 U245 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n232) );
  OAI22_X1 U246 ( .A1(n243), .A2(n232), .B1(n245), .B2(n215), .ZN(n229) );
  XNOR2_X1 U247 ( .A(n556), .B(\mult_x_1/n284 ), .ZN(n230) );
  OAI22_X1 U248 ( .A1(n248), .A2(n230), .B1(n216), .B2(n26), .ZN(n228) );
  HA_X1 U249 ( .A(n218), .B(n217), .CO(n214), .S(n227) );
  NOR2_X1 U250 ( .A1(n222), .A2(n221), .ZN(n220) );
  MUX2_X1 U251 ( .A(n346), .B(n220), .S(n329), .Z(n376) );
  NAND2_X1 U252 ( .A1(n222), .A2(n221), .ZN(n223) );
  MUX2_X1 U253 ( .A(n347), .B(n223), .S(n329), .Z(n378) );
  NAND2_X1 U254 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U255 ( .A(n348), .B(n226), .S(n329), .Z(n380) );
  XNOR2_X1 U256 ( .A(n556), .B(\mult_x_1/n285 ), .ZN(n239) );
  OAI22_X1 U257 ( .A1(n248), .A2(n239), .B1(n230), .B2(n26), .ZN(n235) );
  AND2_X1 U258 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n234) );
  XNOR2_X1 U259 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n236) );
  OAI22_X1 U260 ( .A1(n243), .A2(n236), .B1(n245), .B2(n232), .ZN(n233) );
  OR2_X1 U261 ( .A1(n258), .A2(n257), .ZN(n284) );
  FA_X1 U262 ( .A(n235), .B(n234), .CI(n233), .CO(n257), .S(n256) );
  XNOR2_X1 U263 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n237) );
  OAI22_X1 U264 ( .A1(n238), .A2(n237), .B1(n245), .B2(n236), .ZN(n241) );
  XNOR2_X1 U265 ( .A(n556), .B(\mult_x_1/n286 ), .ZN(n244) );
  OAI22_X1 U266 ( .A1(n248), .A2(n244), .B1(n239), .B2(n26), .ZN(n240) );
  NOR2_X1 U267 ( .A1(n256), .A2(n255), .ZN(n277) );
  HA_X1 U268 ( .A(n241), .B(n240), .CO(n255), .S(n253) );
  OR2_X1 U269 ( .A1(\mult_x_1/n288 ), .A2(n20), .ZN(n242) );
  OAI22_X1 U270 ( .A1(n243), .A2(n20), .B1(n242), .B2(n245), .ZN(n252) );
  OR2_X1 U271 ( .A1(n253), .A2(n252), .ZN(n273) );
  XNOR2_X1 U272 ( .A(n556), .B(\mult_x_1/n287 ), .ZN(n247) );
  OAI22_X1 U273 ( .A1(n248), .A2(n247), .B1(n244), .B2(n26), .ZN(n251) );
  INV_X1 U274 ( .A(n245), .ZN(n246) );
  AND2_X1 U275 ( .A1(\mult_x_1/n288 ), .A2(n246), .ZN(n250) );
  NOR2_X1 U276 ( .A1(n251), .A2(n250), .ZN(n266) );
  OAI22_X1 U277 ( .A1(n248), .A2(\mult_x_1/n288 ), .B1(n247), .B2(n26), .ZN(
        n263) );
  OR2_X1 U278 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n249) );
  NAND2_X1 U279 ( .A1(n249), .A2(n248), .ZN(n262) );
  NAND2_X1 U280 ( .A1(n263), .A2(n262), .ZN(n269) );
  NAND2_X1 U281 ( .A1(n251), .A2(n250), .ZN(n267) );
  OAI21_X1 U282 ( .B1(n266), .B2(n269), .A(n267), .ZN(n274) );
  NAND2_X1 U283 ( .A1(n253), .A2(n252), .ZN(n272) );
  INV_X1 U284 ( .A(n272), .ZN(n254) );
  AOI21_X1 U285 ( .B1(n273), .B2(n274), .A(n254), .ZN(n280) );
  NAND2_X1 U286 ( .A1(n256), .A2(n255), .ZN(n278) );
  OAI21_X1 U287 ( .B1(n277), .B2(n280), .A(n278), .ZN(n285) );
  NAND2_X1 U288 ( .A1(n258), .A2(n257), .ZN(n283) );
  INV_X1 U289 ( .A(n283), .ZN(n259) );
  AOI21_X1 U290 ( .B1(n284), .B2(n285), .A(n259), .ZN(n260) );
  MUX2_X1 U291 ( .A(n354), .B(n260), .S(n329), .Z(n392) );
  MUX2_X1 U292 ( .A(product[0]), .B(n519), .S(en), .Z(n409) );
  MUX2_X1 U293 ( .A(n519), .B(n520), .S(en), .Z(n411) );
  AND2_X1 U294 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n261) );
  MUX2_X1 U295 ( .A(n520), .B(n261), .S(en), .Z(n413) );
  MUX2_X1 U296 ( .A(product[1]), .B(n522), .S(en), .Z(n415) );
  MUX2_X1 U297 ( .A(n522), .B(n523), .S(n329), .Z(n417) );
  OR2_X1 U298 ( .A1(n263), .A2(n262), .ZN(n264) );
  AND2_X1 U299 ( .A1(n264), .A2(n269), .ZN(n265) );
  MUX2_X1 U300 ( .A(n523), .B(n265), .S(n329), .Z(n419) );
  MUX2_X1 U301 ( .A(product[2]), .B(n525), .S(n329), .Z(n421) );
  MUX2_X1 U302 ( .A(n525), .B(n526), .S(n329), .Z(n423) );
  INV_X1 U303 ( .A(n266), .ZN(n268) );
  NAND2_X1 U304 ( .A1(n268), .A2(n267), .ZN(n270) );
  XOR2_X1 U305 ( .A(n270), .B(n269), .Z(n271) );
  MUX2_X1 U306 ( .A(n526), .B(n271), .S(n329), .Z(n425) );
  MUX2_X1 U307 ( .A(product[3]), .B(n528), .S(n329), .Z(n427) );
  MUX2_X1 U308 ( .A(n528), .B(n529), .S(n24), .Z(n429) );
  NAND2_X1 U309 ( .A1(n273), .A2(n272), .ZN(n275) );
  XNOR2_X1 U310 ( .A(n275), .B(n274), .ZN(n276) );
  MUX2_X1 U311 ( .A(n529), .B(n276), .S(n329), .Z(n431) );
  MUX2_X1 U312 ( .A(product[4]), .B(n531), .S(n24), .Z(n433) );
  MUX2_X1 U313 ( .A(n531), .B(n532), .S(n329), .Z(n435) );
  INV_X1 U314 ( .A(n277), .ZN(n279) );
  NAND2_X1 U315 ( .A1(n279), .A2(n278), .ZN(n281) );
  XOR2_X1 U316 ( .A(n281), .B(n280), .Z(n282) );
  MUX2_X1 U317 ( .A(n532), .B(n282), .S(n24), .Z(n437) );
  MUX2_X1 U318 ( .A(product[5]), .B(n534), .S(n329), .Z(n439) );
  MUX2_X1 U319 ( .A(n534), .B(n535), .S(n24), .Z(n441) );
  NAND2_X1 U320 ( .A1(n284), .A2(n283), .ZN(n286) );
  MUX2_X1 U321 ( .A(product[6]), .B(n537), .S(n329), .Z(n445) );
  NAND2_X1 U322 ( .A1(n397), .A2(n347), .ZN(n287) );
  XOR2_X1 U323 ( .A(n287), .B(n354), .Z(n288) );
  MUX2_X1 U324 ( .A(n537), .B(n288), .S(n24), .Z(n447) );
  MUX2_X1 U325 ( .A(product[7]), .B(n539), .S(n24), .Z(n449) );
  OAI21_X1 U326 ( .B1(n346), .B2(n354), .A(n347), .ZN(n291) );
  NAND2_X1 U327 ( .A1(n337), .A2(n345), .ZN(n289) );
  XNOR2_X1 U328 ( .A(n291), .B(n289), .ZN(n290) );
  MUX2_X1 U329 ( .A(n539), .B(n290), .S(n24), .Z(n451) );
  MUX2_X1 U330 ( .A(product[8]), .B(n541), .S(n24), .Z(n453) );
  AOI21_X1 U331 ( .B1(n291), .B2(n337), .A(n398), .ZN(n294) );
  NAND2_X1 U332 ( .A1(n399), .A2(n344), .ZN(n292) );
  XOR2_X1 U333 ( .A(n294), .B(n292), .Z(n293) );
  MUX2_X1 U334 ( .A(n541), .B(n293), .S(n329), .Z(n455) );
  MUX2_X1 U335 ( .A(product[9]), .B(n543), .S(n24), .Z(n457) );
  OAI21_X1 U336 ( .B1(n294), .B2(n343), .A(n344), .ZN(n302) );
  INV_X1 U337 ( .A(n302), .ZN(n297) );
  NAND2_X1 U338 ( .A1(n400), .A2(n351), .ZN(n295) );
  XOR2_X1 U339 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U340 ( .A(n543), .B(n296), .S(n329), .Z(n459) );
  MUX2_X1 U341 ( .A(product[10]), .B(n545), .S(n329), .Z(n461) );
  OAI21_X1 U342 ( .B1(n297), .B2(n352), .A(n351), .ZN(n299) );
  NAND2_X1 U343 ( .A1(n401), .A2(n342), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U345 ( .A(n545), .B(n300), .S(n24), .Z(n463) );
  MUX2_X1 U346 ( .A(product[11]), .B(n547), .S(n329), .Z(n465) );
  NOR2_X1 U347 ( .A1(n349), .A2(n352), .ZN(n303) );
  OAI21_X1 U348 ( .B1(n349), .B2(n351), .A(n342), .ZN(n301) );
  AOI21_X1 U349 ( .B1(n303), .B2(n302), .A(n301), .ZN(n325) );
  NAND2_X1 U350 ( .A1(n402), .A2(n341), .ZN(n304) );
  XOR2_X1 U351 ( .A(n325), .B(n304), .Z(n305) );
  MUX2_X1 U352 ( .A(n547), .B(n305), .S(n24), .Z(n467) );
  MUX2_X1 U353 ( .A(product[12]), .B(n549), .S(n329), .Z(n469) );
  OAI21_X1 U354 ( .B1(n325), .B2(n353), .A(n341), .ZN(n307) );
  NAND2_X1 U355 ( .A1(n350), .A2(n340), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  MUX2_X1 U357 ( .A(n549), .B(n308), .S(n329), .Z(n471) );
  MUX2_X1 U358 ( .A(product[13]), .B(n551), .S(n24), .Z(n473) );
  NAND2_X1 U359 ( .A1(n402), .A2(n350), .ZN(n310) );
  AOI21_X1 U360 ( .B1(n396), .B2(n350), .A(n403), .ZN(n309) );
  OAI21_X1 U361 ( .B1(n325), .B2(n310), .A(n309), .ZN(n312) );
  NAND2_X1 U362 ( .A1(n336), .A2(n348), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U364 ( .A(n551), .B(n313), .S(n329), .Z(n475) );
  MUX2_X1 U365 ( .A(product[14]), .B(n553), .S(n24), .Z(n477) );
  NAND2_X1 U366 ( .A1(n350), .A2(n336), .ZN(n315) );
  NOR2_X1 U367 ( .A1(n353), .A2(n315), .ZN(n321) );
  INV_X1 U368 ( .A(n321), .ZN(n317) );
  AOI21_X1 U369 ( .B1(n403), .B2(n336), .A(n394), .ZN(n314) );
  OAI21_X1 U370 ( .B1(n315), .B2(n341), .A(n314), .ZN(n322) );
  INV_X1 U371 ( .A(n322), .ZN(n316) );
  OAI21_X1 U372 ( .B1(n325), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U373 ( .A1(n335), .A2(n339), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U375 ( .A(n553), .B(n320), .S(n329), .Z(n479) );
  MUX2_X1 U376 ( .A(product[15]), .B(n555), .S(n219), .Z(n481) );
  NAND2_X1 U377 ( .A1(n321), .A2(n335), .ZN(n324) );
  AOI21_X1 U378 ( .B1(n322), .B2(n335), .A(n395), .ZN(n323) );
  OAI21_X1 U379 ( .B1(n325), .B2(n324), .A(n323), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n326), .B(n338), .ZN(n327) );
  MUX2_X1 U381 ( .A(n555), .B(n327), .S(n329), .Z(n483) );
  MUX2_X1 U382 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n219), .Z(n485) );
  MUX2_X1 U383 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n24), .Z(n487) );
  MUX2_X1 U384 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n329), .Z(n489) );
  MUX2_X1 U385 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n219), .Z(n491) );
  MUX2_X1 U386 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n24), .Z(n493) );
  MUX2_X1 U387 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n329), .Z(n495) );
  MUX2_X1 U388 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n219), .Z(n497) );
  MUX2_X1 U389 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n329), .Z(n499) );
  MUX2_X1 U390 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n24), .Z(n501) );
  MUX2_X1 U391 ( .A(n556), .B(A_extended[1]), .S(n329), .Z(n503) );
  MUX2_X1 U392 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n219), .Z(n505) );
  MUX2_X1 U393 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n219), .Z(n507) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n24), .Z(n509) );
  MUX2_X1 U395 ( .A(n328), .B(A_extended[5]), .S(n329), .Z(n511) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n329), .Z(n513) );
  MUX2_X1 U397 ( .A(n21), .B(A_extended[7]), .S(n219), .Z(n515) );
  OR2_X1 U398 ( .A1(n219), .A2(n558), .ZN(n517) );
endmodule


module conv_128_32_DW_mult_pipe_J1_13 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n363, n365,
         n367, n369, n371, n373, n375, n377, n379, n381, n383, n385, n387,
         n389, n391, n393, n395, n397, n399, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n414, n416, n418, n420,
         n422, n424, n426, n428, n430, n432, n434, n436, n438, n440, n442,
         n444, n446, n448, n450, n452, n454, n456, n458, n460, n462, n464,
         n466, n468, n470, n472, n474, n476, n478, n480, n482, n484, n486,
         n488, n490, n492, n494, n496, n498, n500, n502, n504, n506, n508,
         n510, n512, n514, n516, n518, n520, n522, n524, n525, n527, n528,
         n530, n531, n533, n534, n536, n537, n539, n540, n542, n544, n546,
         n548, n550, n552, n554, n556, n558, n560, n561, n562, n563, n564,
         n565;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n412), .SE(n522), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n412), .SE(n518), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n6) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n412), .SE(n516), .CK(clk), .Q(n562), 
        .QN(n46) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n412), .SE(n514), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n412), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n43) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n412), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n45) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n412), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n38) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n412), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n410), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n411), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n409), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n412), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n409), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n409), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n5) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n409), .SE(n488), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n409), .SE(n486), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n409), .SE(n484), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n409), .SE(n482), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n409), .SE(n480), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n411), .SE(n478), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n410), .SE(n476), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n412), .SE(n474), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n409), .SE(n472), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n409), .SE(n470), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n409), .SE(n468), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n409), .SE(n466), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n409), .SE(n464), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n409), .SE(n462), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n409), .SE(n460), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n409), .SE(n458), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n411), .SE(n456), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n411), .SE(n454), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n411), .SE(n452), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n411), .SE(n450), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n411), .SE(n448), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n411), .SE(n446), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n411), .SE(n444), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n411), .SE(n442), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n411), .SE(n440), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n411), .SE(n438), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n411), .SE(n436), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n410), .SE(n434), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n410), .SE(n432), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n410), .SE(n430), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n410), .SE(n428), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n410), .SE(n426), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n410), .SE(n424), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n410), .SE(n422), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n410), .SE(n420), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n410), .SE(n418), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n410), .SE(n416), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n410), .SE(n414), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n412), .SE(n520), .CK(clk), .Q(n563), 
        .QN(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n565), .SE(n399), .CK(
        clk), .QN(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n565), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n565), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n565), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n357), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n565), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n356), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n565), .SE(n389), .CK(
        clk), .Q(n340), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n565), .SE(n387), .CK(
        clk), .Q(n407), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n565), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n565), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n352), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n565), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n351), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n565), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n565), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n349), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n565), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n348), .QN(n48) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n565), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n347), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n565), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n346), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n565), .SE(n369), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n565), .SE(n367), .CK(
        clk), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n565), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n343), .QN(n47) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n565), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n565), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n341) );
  SDFF_X2 clk_r_REG58_S1 ( .D(1'b0), .SI(n412), .SE(n508), .CK(clk), .Q(n561), 
        .QN(n44) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n412), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n339) );
  BUF_X1 U2 ( .A(n563), .Z(n336) );
  BUF_X1 U3 ( .A(n409), .Z(n412) );
  BUF_X1 U4 ( .A(n409), .Z(n411) );
  BUF_X1 U5 ( .A(n409), .Z(n410) );
  INV_X1 U6 ( .A(n565), .ZN(n409) );
  NAND2_X1 U7 ( .A1(n18), .A2(n17), .ZN(n177) );
  NAND2_X1 U8 ( .A1(n561), .A2(n45), .ZN(n243) );
  AND2_X1 U9 ( .A1(n564), .A2(\mult_x_1/n281 ), .ZN(n136) );
  XNOR2_X1 U10 ( .A(n26), .B(n155), .ZN(n132) );
  XNOR2_X1 U11 ( .A(n153), .B(n154), .ZN(n26) );
  INV_X1 U12 ( .A(n214), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n155), .A2(n154), .ZN(n24) );
  XNOR2_X1 U14 ( .A(n23), .B(n21), .ZN(n125) );
  XNOR2_X1 U15 ( .A(n115), .B(n116), .ZN(n23) );
  OAI21_X1 U16 ( .B1(n28), .B2(n29), .A(n27), .ZN(n216) );
  XNOR2_X1 U17 ( .A(n30), .B(n29), .ZN(n253) );
  XNOR2_X1 U18 ( .A(n213), .B(n212), .ZN(n29) );
  INV_X1 U19 ( .A(rst_n), .ZN(n565) );
  NOR2_X1 U20 ( .A1(n225), .A2(n224), .ZN(n28) );
  NAND2_X1 U21 ( .A1(n225), .A2(n224), .ZN(n27) );
  XNOR2_X1 U22 ( .A(n225), .B(n31), .ZN(n30) );
  NOR2_X1 U23 ( .A1(n181), .A2(n8), .ZN(n116) );
  INV_X1 U24 ( .A(n58), .ZN(n36) );
  INV_X1 U25 ( .A(n224), .ZN(n31) );
  NAND2_X1 U26 ( .A1(n180), .A2(n5), .ZN(n8) );
  INV_X1 U27 ( .A(n52), .ZN(n227) );
  INV_X1 U28 ( .A(n178), .ZN(n37) );
  NAND2_X1 U29 ( .A1(n9), .A2(n12), .ZN(n387) );
  NAND2_X1 U30 ( .A1(n11), .A2(n10), .ZN(n9) );
  NOR2_X1 U31 ( .A1(n219), .A2(n13), .ZN(n10) );
  INV_X1 U32 ( .A(n220), .ZN(n11) );
  NAND2_X1 U33 ( .A1(n13), .A2(n354), .ZN(n12) );
  INV_X1 U34 ( .A(n214), .ZN(n13) );
  NAND2_X1 U35 ( .A1(n15), .A2(n14), .ZN(n379) );
  NAND2_X1 U36 ( .A1(n7), .A2(n350), .ZN(n14) );
  NAND2_X1 U37 ( .A1(n16), .A2(n214), .ZN(n15) );
  NAND2_X1 U38 ( .A1(n203), .A2(n202), .ZN(n16) );
  OAI21_X1 U39 ( .B1(n46), .B2(n563), .A(\mult_x_1/a[6] ), .ZN(n17) );
  OAI21_X1 U40 ( .B1(n338), .B2(n562), .A(n6), .ZN(n18) );
  NAND2_X1 U41 ( .A1(n20), .A2(n19), .ZN(n262) );
  NAND2_X1 U42 ( .A1(n115), .A2(n116), .ZN(n19) );
  OAI21_X1 U43 ( .B1(n115), .B2(n116), .A(n21), .ZN(n20) );
  XNOR2_X1 U44 ( .A(n96), .B(n22), .ZN(n21) );
  OAI22_X1 U45 ( .A1(n240), .A2(n72), .B1(n93), .B2(n238), .ZN(n22) );
  NAND2_X1 U46 ( .A1(n57), .A2(n56), .ZN(n238) );
  XNOR2_X2 U47 ( .A(n562), .B(\mult_x_1/a[6] ), .ZN(n178) );
  NAND2_X1 U48 ( .A1(n25), .A2(n24), .ZN(n221) );
  OAI21_X1 U49 ( .B1(n155), .B2(n154), .A(n153), .ZN(n25) );
  OAI21_X1 U50 ( .B1(n33), .B2(n13), .A(n32), .ZN(n448) );
  NAND2_X1 U51 ( .A1(n13), .A2(n540), .ZN(n32) );
  XNOR2_X1 U52 ( .A(n289), .B(n34), .ZN(n33) );
  INV_X1 U53 ( .A(n288), .ZN(n34) );
  INV_X1 U54 ( .A(n100), .ZN(n181) );
  OR2_X1 U55 ( .A1(n42), .A2(n96), .ZN(n122) );
  NAND2_X1 U56 ( .A1(n81), .A2(n80), .ZN(n85) );
  INV_X1 U57 ( .A(n123), .ZN(n76) );
  NOR2_X1 U58 ( .A1(n122), .A2(n121), .ZN(n75) );
  AOI21_X1 U59 ( .B1(n81), .B2(n49), .A(n67), .ZN(n153) );
  NOR2_X1 U60 ( .A1(n83), .A2(n82), .ZN(n67) );
  OAI21_X1 U61 ( .B1(n76), .B2(n75), .A(n74), .ZN(n258) );
  NAND2_X1 U62 ( .A1(n122), .A2(n121), .ZN(n74) );
  XNOR2_X1 U63 ( .A(n120), .B(n119), .ZN(n261) );
  NAND2_X1 U64 ( .A1(n134), .A2(n133), .ZN(n365) );
  OR2_X1 U65 ( .A1(n214), .A2(n47), .ZN(n133) );
  OAI21_X1 U66 ( .B1(n132), .B2(n131), .A(n214), .ZN(n134) );
  INV_X1 U67 ( .A(n111), .ZN(n112) );
  OAI21_X1 U68 ( .B1(n113), .B2(n7), .A(n110), .ZN(n111) );
  OAI22_X1 U69 ( .A1(n114), .A2(n50), .B1(n337), .B2(n406), .ZN(n393) );
  XNOR2_X1 U70 ( .A(n136), .B(n561), .ZN(n35) );
  INV_X1 U71 ( .A(n58), .ZN(n240) );
  INV_X1 U72 ( .A(n38), .ZN(n39) );
  OR2_X2 U73 ( .A1(n52), .A2(n51), .ZN(n40) );
  OR2_X1 U74 ( .A1(n52), .A2(n51), .ZN(n168) );
  INV_X1 U75 ( .A(n339), .ZN(n41) );
  OAI22_X1 U76 ( .A1(n238), .A2(n93), .B1(n240), .B2(n72), .ZN(n42) );
  XNOR2_X1 U77 ( .A(n43), .B(n44), .ZN(n57) );
  BUF_X4 U78 ( .A(en), .Z(n337) );
  BUF_X2 U79 ( .A(n562), .Z(n335) );
  AND2_X1 U80 ( .A1(n66), .A2(n80), .ZN(n49) );
  OR2_X1 U81 ( .A1(n113), .A2(n7), .ZN(n50) );
  XNOR2_X1 U82 ( .A(n339), .B(\mult_x_1/a[4] ), .ZN(n52) );
  XNOR2_X1 U83 ( .A(\mult_x_1/a[4] ), .B(n562), .ZN(n51) );
  XNOR2_X1 U84 ( .A(n335), .B(\mult_x_1/n281 ), .ZN(n63) );
  XNOR2_X1 U85 ( .A(n136), .B(n335), .ZN(n139) );
  OAI22_X1 U86 ( .A1(n40), .A2(n63), .B1(n139), .B2(n227), .ZN(n141) );
  INV_X1 U87 ( .A(n141), .ZN(n144) );
  XNOR2_X1 U88 ( .A(n336), .B(\mult_x_1/n283 ), .ZN(n55) );
  XNOR2_X1 U89 ( .A(n336), .B(\mult_x_1/n282 ), .ZN(n138) );
  OAI22_X1 U90 ( .A1(n177), .A2(n55), .B1(n178), .B2(n138), .ZN(n143) );
  AND2_X1 U91 ( .A1(n564), .A2(n563), .ZN(n53) );
  BUF_X1 U92 ( .A(n53), .Z(n180) );
  XNOR2_X1 U93 ( .A(n180), .B(\mult_x_1/n284 ), .ZN(n54) );
  XNOR2_X1 U94 ( .A(n53), .B(n338), .ZN(n100) );
  NOR2_X1 U95 ( .A1(n54), .A2(n181), .ZN(n142) );
  XNOR2_X1 U96 ( .A(n336), .B(\mult_x_1/n284 ), .ZN(n61) );
  OAI22_X1 U97 ( .A1(n177), .A2(n61), .B1(n178), .B2(n55), .ZN(n79) );
  XOR2_X1 U98 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n56) );
  XNOR2_X1 U99 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n72) );
  XNOR2_X1 U100 ( .A(n136), .B(n41), .ZN(n59) );
  INV_X1 U101 ( .A(n57), .ZN(n58) );
  OAI22_X1 U102 ( .A1(n238), .A2(n72), .B1(n59), .B2(n240), .ZN(n78) );
  AOI21_X1 U103 ( .B1(n36), .B2(n238), .A(n59), .ZN(n60) );
  INV_X1 U104 ( .A(n60), .ZN(n77) );
  XNOR2_X1 U105 ( .A(n335), .B(\mult_x_1/n283 ), .ZN(n71) );
  XNOR2_X1 U106 ( .A(n335), .B(\mult_x_1/n282 ), .ZN(n64) );
  OAI22_X1 U107 ( .A1(n40), .A2(n71), .B1(n227), .B2(n64), .ZN(n118) );
  XNOR2_X1 U108 ( .A(n336), .B(\mult_x_1/n285 ), .ZN(n69) );
  OAI22_X1 U109 ( .A1(n177), .A2(n69), .B1(n178), .B2(n61), .ZN(n117) );
  OR2_X1 U110 ( .A1(n118), .A2(n117), .ZN(n62) );
  INV_X1 U111 ( .A(n78), .ZN(n119) );
  NAND2_X1 U112 ( .A1(n62), .A2(n119), .ZN(n81) );
  OAI22_X1 U113 ( .A1(n40), .A2(n64), .B1(n227), .B2(n63), .ZN(n83) );
  XNOR2_X1 U114 ( .A(n180), .B(\mult_x_1/n285 ), .ZN(n65) );
  NOR2_X1 U115 ( .A1(n65), .A2(n181), .ZN(n82) );
  NAND2_X1 U116 ( .A1(n83), .A2(n82), .ZN(n66) );
  NAND2_X1 U117 ( .A1(n118), .A2(n117), .ZN(n80) );
  XNOR2_X1 U118 ( .A(n136), .B(n561), .ZN(n99) );
  AOI21_X1 U119 ( .B1(n243), .B2(n45), .A(n99), .ZN(n68) );
  INV_X1 U120 ( .A(n68), .ZN(n91) );
  XNOR2_X1 U121 ( .A(n336), .B(\mult_x_1/n286 ), .ZN(n97) );
  OAI22_X1 U122 ( .A1(n177), .A2(n97), .B1(n178), .B2(n69), .ZN(n90) );
  XNOR2_X1 U123 ( .A(n180), .B(\mult_x_1/n287 ), .ZN(n70) );
  NOR2_X1 U124 ( .A1(n70), .A2(n181), .ZN(n89) );
  XNOR2_X1 U125 ( .A(n335), .B(\mult_x_1/n284 ), .ZN(n92) );
  OAI22_X1 U126 ( .A1(n168), .A2(n92), .B1(n227), .B2(n71), .ZN(n96) );
  XNOR2_X1 U127 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n93) );
  XNOR2_X1 U128 ( .A(n180), .B(\mult_x_1/n286 ), .ZN(n73) );
  NOR2_X1 U129 ( .A1(n73), .A2(n181), .ZN(n121) );
  FA_X1 U130 ( .A(n79), .B(n78), .CI(n77), .CO(n154), .S(n257) );
  XOR2_X1 U131 ( .A(n83), .B(n82), .Z(n84) );
  XOR2_X1 U132 ( .A(n85), .B(n84), .Z(n256) );
  NAND2_X1 U133 ( .A1(n132), .A2(n131), .ZN(n86) );
  BUF_X2 U134 ( .A(en), .Z(n214) );
  NAND2_X1 U135 ( .A1(n86), .A2(n214), .ZN(n88) );
  OR2_X1 U136 ( .A1(n214), .A2(n408), .ZN(n87) );
  NAND2_X1 U137 ( .A1(n88), .A2(n87), .ZN(n373) );
  FA_X1 U138 ( .A(n91), .B(n90), .CI(n89), .CO(n123), .S(n127) );
  XNOR2_X1 U139 ( .A(n335), .B(\mult_x_1/n285 ), .ZN(n104) );
  OAI22_X1 U140 ( .A1(n40), .A2(n104), .B1(n227), .B2(n92), .ZN(n109) );
  XNOR2_X1 U141 ( .A(n41), .B(\mult_x_1/n283 ), .ZN(n106) );
  OAI22_X1 U142 ( .A1(n238), .A2(n106), .B1(n36), .B2(n93), .ZN(n108) );
  OR2_X1 U143 ( .A1(\mult_x_1/n288 ), .A2(n338), .ZN(n94) );
  OAI22_X1 U144 ( .A1(n177), .A2(n338), .B1(n94), .B2(n178), .ZN(n160) );
  XNOR2_X1 U145 ( .A(n336), .B(\mult_x_1/n288 ), .ZN(n95) );
  XNOR2_X1 U146 ( .A(n336), .B(\mult_x_1/n287 ), .ZN(n98) );
  OAI22_X1 U147 ( .A1(n177), .A2(n95), .B1(n178), .B2(n98), .ZN(n159) );
  OAI22_X1 U148 ( .A1(n177), .A2(n98), .B1(n178), .B2(n97), .ZN(n103) );
  XNOR2_X1 U149 ( .A(n561), .B(\mult_x_1/n281 ), .ZN(n105) );
  OAI22_X1 U150 ( .A1(n243), .A2(n105), .B1(n35), .B2(n45), .ZN(n102) );
  AND2_X1 U151 ( .A1(\mult_x_1/n288 ), .A2(n100), .ZN(n101) );
  FA_X1 U152 ( .A(n102), .B(n101), .CI(n103), .CO(n115), .S(n197) );
  XNOR2_X1 U153 ( .A(n335), .B(\mult_x_1/n286 ), .ZN(n166) );
  OAI22_X1 U154 ( .A1(n40), .A2(n166), .B1(n227), .B2(n104), .ZN(n163) );
  XNOR2_X1 U155 ( .A(n561), .B(\mult_x_1/n282 ), .ZN(n157) );
  OAI22_X1 U156 ( .A1(n243), .A2(n157), .B1(n105), .B2(n45), .ZN(n162) );
  XNOR2_X1 U157 ( .A(n41), .B(\mult_x_1/n284 ), .ZN(n158) );
  OAI22_X1 U158 ( .A1(n238), .A2(n158), .B1(n36), .B2(n106), .ZN(n161) );
  FA_X1 U159 ( .A(n109), .B(n108), .CI(n107), .CO(n126), .S(n195) );
  OR2_X1 U160 ( .A1(n214), .A2(n48), .ZN(n110) );
  OAI21_X1 U161 ( .B1(n114), .B2(n7), .A(n112), .ZN(n375) );
  XNOR2_X1 U162 ( .A(n118), .B(n117), .ZN(n120) );
  XNOR2_X1 U163 ( .A(n122), .B(n121), .ZN(n124) );
  XNOR2_X1 U164 ( .A(n124), .B(n123), .ZN(n260) );
  FA_X1 U165 ( .A(n127), .B(n126), .CI(n125), .CO(n219), .S(n114) );
  NAND2_X1 U166 ( .A1(n220), .A2(n219), .ZN(n128) );
  NAND2_X1 U167 ( .A1(n128), .A2(n337), .ZN(n130) );
  OR2_X1 U168 ( .A1(n214), .A2(n340), .ZN(n129) );
  NAND2_X1 U169 ( .A1(n130), .A2(n129), .ZN(n389) );
  XNOR2_X1 U190 ( .A(n180), .B(\mult_x_1/n282 ), .ZN(n135) );
  NOR2_X1 U191 ( .A1(n135), .A2(n181), .ZN(n175) );
  XNOR2_X1 U192 ( .A(n336), .B(n39), .ZN(n137) );
  XNOR2_X1 U193 ( .A(n136), .B(n336), .ZN(n176) );
  OAI22_X1 U194 ( .A1(n177), .A2(n137), .B1(n176), .B2(n178), .ZN(n186) );
  INV_X1 U195 ( .A(n186), .ZN(n174) );
  OAI22_X1 U196 ( .A1(n177), .A2(n138), .B1(n178), .B2(n137), .ZN(n148) );
  AOI21_X1 U197 ( .B1(n227), .B2(n168), .A(n139), .ZN(n140) );
  INV_X1 U198 ( .A(n140), .ZN(n147) );
  BUF_X1 U199 ( .A(n141), .Z(n146) );
  FA_X1 U200 ( .A(n144), .B(n143), .CI(n142), .CO(n152), .S(n155) );
  XNOR2_X1 U201 ( .A(n180), .B(\mult_x_1/n283 ), .ZN(n145) );
  NOR2_X1 U202 ( .A1(n145), .A2(n181), .ZN(n151) );
  FA_X1 U203 ( .A(n148), .B(n147), .CI(n146), .CO(n173), .S(n150) );
  OR2_X1 U204 ( .A1(n193), .A2(n192), .ZN(n149) );
  MUX2_X1 U205 ( .A(n341), .B(n149), .S(n214), .Z(n361) );
  FA_X1 U206 ( .A(n152), .B(n151), .CI(n150), .CO(n192), .S(n222) );
  OR2_X1 U207 ( .A1(n222), .A2(n221), .ZN(n156) );
  MUX2_X1 U208 ( .A(n342), .B(n156), .S(n214), .Z(n363) );
  XNOR2_X1 U209 ( .A(n561), .B(\mult_x_1/n283 ), .ZN(n211) );
  OAI22_X1 U210 ( .A1(n243), .A2(n211), .B1(n157), .B2(n45), .ZN(n171) );
  AND2_X1 U211 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n170) );
  XNOR2_X1 U212 ( .A(n41), .B(\mult_x_1/n285 ), .ZN(n210) );
  OAI22_X1 U213 ( .A1(n238), .A2(n210), .B1(n36), .B2(n158), .ZN(n169) );
  HA_X1 U214 ( .A(n160), .B(n159), .CO(n107), .S(n199) );
  FA_X1 U215 ( .A(n163), .B(n162), .CI(n161), .CO(n196), .S(n198) );
  OR2_X1 U216 ( .A1(\mult_x_1/n288 ), .A2(n46), .ZN(n164) );
  OAI22_X1 U217 ( .A1(n40), .A2(n46), .B1(n164), .B2(n227), .ZN(n213) );
  XNOR2_X1 U218 ( .A(n335), .B(\mult_x_1/n288 ), .ZN(n165) );
  XNOR2_X1 U219 ( .A(n335), .B(\mult_x_1/n287 ), .ZN(n167) );
  OAI22_X1 U220 ( .A1(n168), .A2(n165), .B1(n227), .B2(n167), .ZN(n212) );
  AND2_X1 U221 ( .A1(n213), .A2(n212), .ZN(n209) );
  OAI22_X1 U222 ( .A1(n40), .A2(n167), .B1(n227), .B2(n166), .ZN(n208) );
  FA_X1 U223 ( .A(n171), .B(n170), .CI(n169), .CO(n200), .S(n207) );
  OR2_X1 U224 ( .A1(n205), .A2(n204), .ZN(n172) );
  MUX2_X1 U225 ( .A(n344), .B(n172), .S(n214), .Z(n367) );
  FA_X1 U226 ( .A(n175), .B(n174), .CI(n173), .CO(n188), .S(n193) );
  AOI21_X1 U227 ( .B1(n178), .B2(n177), .A(n176), .ZN(n179) );
  INV_X1 U228 ( .A(n179), .ZN(n184) );
  XNOR2_X1 U229 ( .A(n180), .B(n39), .ZN(n182) );
  NOR2_X1 U230 ( .A1(n182), .A2(n181), .ZN(n183) );
  XOR2_X1 U231 ( .A(n184), .B(n183), .Z(n185) );
  XOR2_X1 U232 ( .A(n186), .B(n185), .Z(n187) );
  OR2_X1 U233 ( .A1(n188), .A2(n187), .ZN(n190) );
  NAND2_X1 U234 ( .A1(n188), .A2(n187), .ZN(n189) );
  NAND2_X1 U235 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U236 ( .A(n345), .B(n191), .S(n214), .Z(n369) );
  NAND2_X1 U237 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U238 ( .A(n346), .B(n194), .S(n214), .Z(n371) );
  FA_X1 U239 ( .A(n197), .B(n196), .CI(n195), .CO(n113), .S(n203) );
  FA_X1 U240 ( .A(n200), .B(n199), .CI(n198), .CO(n202), .S(n205) );
  NOR2_X1 U241 ( .A1(n203), .A2(n202), .ZN(n201) );
  MUX2_X1 U242 ( .A(n349), .B(n201), .S(n214), .Z(n377) );
  NAND2_X1 U243 ( .A1(n205), .A2(n204), .ZN(n206) );
  MUX2_X1 U244 ( .A(n351), .B(n206), .S(n214), .Z(n381) );
  FA_X1 U245 ( .A(n209), .B(n208), .CI(n207), .CO(n204), .S(n217) );
  XNOR2_X1 U246 ( .A(n41), .B(\mult_x_1/n286 ), .ZN(n228) );
  OAI22_X1 U247 ( .A1(n238), .A2(n228), .B1(n36), .B2(n210), .ZN(n225) );
  XNOR2_X1 U248 ( .A(n561), .B(\mult_x_1/n284 ), .ZN(n226) );
  OAI22_X1 U249 ( .A1(n243), .A2(n226), .B1(n211), .B2(n45), .ZN(n224) );
  NOR2_X1 U250 ( .A1(n217), .A2(n216), .ZN(n215) );
  MUX2_X1 U251 ( .A(n352), .B(n215), .S(n214), .Z(n383) );
  NAND2_X1 U252 ( .A1(n217), .A2(n216), .ZN(n218) );
  MUX2_X1 U253 ( .A(n353), .B(n218), .S(n214), .Z(n385) );
  NAND2_X1 U254 ( .A1(n222), .A2(n221), .ZN(n223) );
  MUX2_X1 U255 ( .A(n356), .B(n223), .S(n214), .Z(n391) );
  XNOR2_X1 U256 ( .A(n561), .B(\mult_x_1/n285 ), .ZN(n234) );
  OAI22_X1 U257 ( .A1(n243), .A2(n234), .B1(n226), .B2(n45), .ZN(n231) );
  AND2_X1 U258 ( .A1(n52), .A2(\mult_x_1/n288 ), .ZN(n230) );
  XNOR2_X1 U259 ( .A(n41), .B(\mult_x_1/n287 ), .ZN(n232) );
  OAI22_X1 U260 ( .A1(n238), .A2(n232), .B1(n36), .B2(n228), .ZN(n229) );
  OR2_X1 U261 ( .A1(n253), .A2(n252), .ZN(n287) );
  FA_X1 U262 ( .A(n231), .B(n230), .CI(n229), .CO(n252), .S(n251) );
  XNOR2_X1 U263 ( .A(n41), .B(\mult_x_1/n288 ), .ZN(n233) );
  OAI22_X1 U264 ( .A1(n238), .A2(n233), .B1(n36), .B2(n232), .ZN(n236) );
  XNOR2_X1 U265 ( .A(n561), .B(\mult_x_1/n286 ), .ZN(n239) );
  OAI22_X1 U266 ( .A1(n243), .A2(n239), .B1(n234), .B2(n45), .ZN(n235) );
  NOR2_X1 U267 ( .A1(n251), .A2(n250), .ZN(n280) );
  HA_X1 U268 ( .A(n236), .B(n235), .CO(n250), .S(n248) );
  OR2_X1 U269 ( .A1(\mult_x_1/n288 ), .A2(n339), .ZN(n237) );
  OAI22_X1 U270 ( .A1(n238), .A2(n339), .B1(n237), .B2(n36), .ZN(n247) );
  OR2_X1 U271 ( .A1(n248), .A2(n247), .ZN(n276) );
  XNOR2_X1 U272 ( .A(n561), .B(\mult_x_1/n287 ), .ZN(n241) );
  OAI22_X1 U273 ( .A1(n243), .A2(n241), .B1(n239), .B2(n45), .ZN(n246) );
  AND2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(n58), .ZN(n245) );
  NOR2_X1 U275 ( .A1(n246), .A2(n245), .ZN(n269) );
  OAI22_X1 U276 ( .A1(n243), .A2(\mult_x_1/n288 ), .B1(n241), .B2(n45), .ZN(
        n266) );
  INV_X1 U277 ( .A(n561), .ZN(n242) );
  OR2_X1 U278 ( .A1(\mult_x_1/n288 ), .A2(n242), .ZN(n244) );
  NAND2_X1 U279 ( .A1(n244), .A2(n243), .ZN(n265) );
  NAND2_X1 U280 ( .A1(n266), .A2(n265), .ZN(n272) );
  NAND2_X1 U281 ( .A1(n246), .A2(n245), .ZN(n270) );
  OAI21_X1 U282 ( .B1(n269), .B2(n272), .A(n270), .ZN(n277) );
  NAND2_X1 U283 ( .A1(n248), .A2(n247), .ZN(n275) );
  INV_X1 U284 ( .A(n275), .ZN(n249) );
  AOI21_X1 U285 ( .B1(n276), .B2(n277), .A(n249), .ZN(n283) );
  NAND2_X1 U286 ( .A1(n251), .A2(n250), .ZN(n281) );
  OAI21_X1 U287 ( .B1(n280), .B2(n283), .A(n281), .ZN(n288) );
  NAND2_X1 U288 ( .A1(n253), .A2(n252), .ZN(n286) );
  INV_X1 U289 ( .A(n286), .ZN(n254) );
  AOI21_X1 U290 ( .B1(n287), .B2(n288), .A(n254), .ZN(n255) );
  MUX2_X1 U291 ( .A(n358), .B(n255), .S(n337), .Z(n395) );
  FA_X1 U292 ( .A(n258), .B(n257), .CI(n256), .CO(n131), .S(n259) );
  MUX2_X1 U293 ( .A(n359), .B(n259), .S(n214), .Z(n397) );
  FA_X1 U294 ( .A(n262), .B(n261), .CI(n260), .CO(n263), .S(n220) );
  MUX2_X1 U295 ( .A(n360), .B(n263), .S(n337), .Z(n399) );
  MUX2_X1 U296 ( .A(product[0]), .B(n524), .S(n337), .Z(n414) );
  MUX2_X1 U297 ( .A(n524), .B(n525), .S(n337), .Z(n416) );
  AND2_X1 U298 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n264) );
  MUX2_X1 U299 ( .A(n525), .B(n264), .S(n337), .Z(n418) );
  MUX2_X1 U300 ( .A(product[1]), .B(n527), .S(n337), .Z(n420) );
  MUX2_X1 U301 ( .A(n527), .B(n528), .S(n337), .Z(n422) );
  OR2_X1 U302 ( .A1(n266), .A2(n265), .ZN(n267) );
  AND2_X1 U303 ( .A1(n267), .A2(n272), .ZN(n268) );
  MUX2_X1 U304 ( .A(n528), .B(n268), .S(n337), .Z(n424) );
  MUX2_X1 U305 ( .A(product[2]), .B(n530), .S(n337), .Z(n426) );
  MUX2_X1 U306 ( .A(n530), .B(n531), .S(n337), .Z(n428) );
  INV_X1 U307 ( .A(n269), .ZN(n271) );
  NAND2_X1 U308 ( .A1(n271), .A2(n270), .ZN(n273) );
  XOR2_X1 U309 ( .A(n273), .B(n272), .Z(n274) );
  MUX2_X1 U310 ( .A(n531), .B(n274), .S(n337), .Z(n430) );
  MUX2_X1 U311 ( .A(product[3]), .B(n533), .S(n337), .Z(n432) );
  MUX2_X1 U312 ( .A(n533), .B(n534), .S(n337), .Z(n434) );
  NAND2_X1 U313 ( .A1(n276), .A2(n275), .ZN(n278) );
  XNOR2_X1 U314 ( .A(n278), .B(n277), .ZN(n279) );
  MUX2_X1 U315 ( .A(n534), .B(n279), .S(n337), .Z(n436) );
  MUX2_X1 U316 ( .A(product[4]), .B(n536), .S(n337), .Z(n438) );
  MUX2_X1 U317 ( .A(n536), .B(n537), .S(n337), .Z(n440) );
  INV_X1 U318 ( .A(n280), .ZN(n282) );
  NAND2_X1 U319 ( .A1(n282), .A2(n281), .ZN(n284) );
  XOR2_X1 U320 ( .A(n284), .B(n283), .Z(n285) );
  MUX2_X1 U321 ( .A(n537), .B(n285), .S(n337), .Z(n442) );
  MUX2_X1 U322 ( .A(product[5]), .B(n539), .S(n337), .Z(n444) );
  MUX2_X1 U323 ( .A(n539), .B(n540), .S(n337), .Z(n446) );
  NAND2_X1 U324 ( .A1(n287), .A2(n286), .ZN(n289) );
  MUX2_X1 U325 ( .A(product[6]), .B(n542), .S(n337), .Z(n450) );
  NAND2_X1 U326 ( .A1(n403), .A2(n353), .ZN(n290) );
  XOR2_X1 U327 ( .A(n290), .B(n358), .Z(n291) );
  MUX2_X1 U328 ( .A(n542), .B(n291), .S(n337), .Z(n452) );
  MUX2_X1 U329 ( .A(product[7]), .B(n544), .S(n337), .Z(n454) );
  OAI21_X1 U330 ( .B1(n352), .B2(n358), .A(n353), .ZN(n294) );
  NAND2_X1 U331 ( .A1(n344), .A2(n351), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n294), .B(n292), .ZN(n293) );
  MUX2_X1 U333 ( .A(n544), .B(n293), .S(n337), .Z(n456) );
  MUX2_X1 U334 ( .A(product[8]), .B(n546), .S(n337), .Z(n458) );
  AOI21_X1 U335 ( .B1(n294), .B2(n344), .A(n404), .ZN(n297) );
  NAND2_X1 U336 ( .A1(n405), .A2(n350), .ZN(n295) );
  XOR2_X1 U337 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U338 ( .A(n546), .B(n296), .S(n337), .Z(n460) );
  MUX2_X1 U339 ( .A(product[9]), .B(n548), .S(n337), .Z(n462) );
  OAI21_X1 U340 ( .B1(n297), .B2(n349), .A(n350), .ZN(n305) );
  INV_X1 U341 ( .A(n305), .ZN(n300) );
  NAND2_X1 U342 ( .A1(n406), .A2(n348), .ZN(n298) );
  XOR2_X1 U343 ( .A(n300), .B(n298), .Z(n299) );
  MUX2_X1 U344 ( .A(n548), .B(n299), .S(n337), .Z(n464) );
  MUX2_X1 U345 ( .A(product[10]), .B(n550), .S(n337), .Z(n466) );
  OAI21_X1 U346 ( .B1(n300), .B2(n357), .A(n348), .ZN(n302) );
  NAND2_X1 U347 ( .A1(n407), .A2(n355), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  MUX2_X1 U349 ( .A(n550), .B(n303), .S(n337), .Z(n468) );
  MUX2_X1 U350 ( .A(product[11]), .B(n552), .S(n337), .Z(n470) );
  NOR2_X1 U351 ( .A1(n354), .A2(n357), .ZN(n306) );
  OAI21_X1 U352 ( .B1(n354), .B2(n348), .A(n355), .ZN(n304) );
  AOI21_X1 U353 ( .B1(n306), .B2(n305), .A(n304), .ZN(n332) );
  NOR2_X1 U354 ( .A1(n359), .A2(n360), .ZN(n319) );
  INV_X1 U355 ( .A(n319), .ZN(n312) );
  NAND2_X1 U356 ( .A1(n359), .A2(n360), .ZN(n321) );
  NAND2_X1 U357 ( .A1(n312), .A2(n321), .ZN(n307) );
  XOR2_X1 U358 ( .A(n332), .B(n307), .Z(n308) );
  MUX2_X1 U359 ( .A(n552), .B(n308), .S(n337), .Z(n472) );
  MUX2_X1 U360 ( .A(product[12]), .B(n554), .S(n337), .Z(n474) );
  OAI21_X1 U361 ( .B1(n332), .B2(n319), .A(n321), .ZN(n310) );
  NAND2_X1 U362 ( .A1(n343), .A2(n347), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  MUX2_X1 U364 ( .A(n554), .B(n311), .S(n337), .Z(n476) );
  MUX2_X1 U365 ( .A(product[13]), .B(n556), .S(n337), .Z(n478) );
  NAND2_X1 U366 ( .A1(n312), .A2(n343), .ZN(n315) );
  INV_X1 U367 ( .A(n321), .ZN(n313) );
  AOI21_X1 U368 ( .B1(n313), .B2(n343), .A(n408), .ZN(n314) );
  OAI21_X1 U369 ( .B1(n332), .B2(n315), .A(n314), .ZN(n317) );
  NAND2_X1 U370 ( .A1(n342), .A2(n356), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  MUX2_X1 U372 ( .A(n556), .B(n318), .S(n337), .Z(n480) );
  MUX2_X1 U373 ( .A(product[14]), .B(n558), .S(n337), .Z(n482) );
  NAND2_X1 U374 ( .A1(n343), .A2(n342), .ZN(n322) );
  NOR2_X1 U375 ( .A1(n319), .A2(n322), .ZN(n328) );
  INV_X1 U376 ( .A(n328), .ZN(n324) );
  AOI21_X1 U377 ( .B1(n408), .B2(n342), .A(n402), .ZN(n320) );
  OAI21_X1 U378 ( .B1(n322), .B2(n321), .A(n320), .ZN(n329) );
  INV_X1 U379 ( .A(n329), .ZN(n323) );
  OAI21_X1 U380 ( .B1(n332), .B2(n324), .A(n323), .ZN(n326) );
  NAND2_X1 U381 ( .A1(n341), .A2(n346), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  MUX2_X1 U383 ( .A(n558), .B(n327), .S(n337), .Z(n484) );
  MUX2_X1 U384 ( .A(product[15]), .B(n560), .S(n337), .Z(n486) );
  NAND2_X1 U385 ( .A1(n328), .A2(n341), .ZN(n331) );
  AOI21_X1 U386 ( .B1(n329), .B2(n341), .A(n401), .ZN(n330) );
  OAI21_X1 U387 ( .B1(n332), .B2(n331), .A(n330), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n333), .B(n345), .ZN(n334) );
  MUX2_X1 U389 ( .A(n560), .B(n334), .S(n337), .Z(n488) );
  MUX2_X1 U390 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n337), .Z(n490) );
  MUX2_X1 U391 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n337), .Z(n492) );
  MUX2_X1 U392 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n337), .Z(n494) );
  MUX2_X1 U393 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n337), .Z(n496) );
  MUX2_X1 U394 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n337), .Z(n498) );
  MUX2_X1 U395 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n337), .Z(n500) );
  MUX2_X1 U396 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n337), .Z(n502) );
  MUX2_X1 U397 ( .A(n39), .B(B_extended[7]), .S(n337), .Z(n504) );
  MUX2_X1 U398 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n337), .Z(n506) );
  MUX2_X1 U399 ( .A(n561), .B(A_extended[1]), .S(n337), .Z(n508) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n337), .Z(n510) );
  MUX2_X1 U401 ( .A(n41), .B(A_extended[3]), .S(n337), .Z(n512) );
  MUX2_X1 U402 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n337), .Z(n514) );
  MUX2_X1 U403 ( .A(n335), .B(A_extended[5]), .S(n337), .Z(n516) );
  MUX2_X1 U404 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n337), .Z(n518) );
  MUX2_X1 U405 ( .A(n336), .B(A_extended[7]), .S(n337), .Z(n520) );
  OR2_X1 U406 ( .A1(n337), .A2(n564), .ZN(n522) );
endmodule


module conv_128_32_DW_mult_pipe_J1_14 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n363,
         n365, n367, n369, n371, n373, n375, n377, n379, n381, n383, n385,
         n387, n389, n391, n393, n395, n397, n399, n401, n403, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n417, n419,
         n421, n423, n425, n427, n429, n431, n433, n435, n437, n439, n441,
         n443, n445, n447, n449, n451, n453, n455, n457, n459, n461, n463,
         n465, n467, n469, n471, n473, n475, n477, n479, n481, n483, n485,
         n487, n489, n491, n493, n495, n497, n499, n501, n503, n505, n507,
         n509, n511, n513, n515, n517, n519, n521, n523, n525, n526, n528,
         n529, n531, n532, n534, n535, n537, n538, n540, n542, n544, n546,
         n548, n550, n552, n554, n556, n558, n560, n561, n562, n563, n564;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n415), .SE(n523), .CK(clk), .Q(n563), 
        .QN(n16) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n415), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n15) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n415), .SE(n517), .CK(clk), .Q(n562), 
        .QN(n18) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n415), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n20) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n415), .SE(n511), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n14) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n415), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n17) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n415), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n19) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n415), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n25) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n414), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n26) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n413), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n23) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n413), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n415), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n22) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n413), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n21) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n413), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n413), .SE(n489), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n413), .SE(n487), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n413), .SE(n485), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n413), .SE(n483), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n413), .SE(n481), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n413), .SE(n479), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n415), .SE(n477), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n414), .SE(n475), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n413), .SE(n473), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n413), .SE(n471), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n413), .SE(n469), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n413), .SE(n467), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n413), .SE(n465), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n413), .SE(n463), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n413), .SE(n461), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n413), .SE(n459), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n413), .SE(n457), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n413), .SE(n455), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n413), .SE(n453), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n413), .SE(n451), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n413), .SE(n449), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n413), .SE(n447), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n413), .SE(n445), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n413), .SE(n443), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n413), .SE(n441), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n413), .SE(n439), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n414), .SE(n437), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n414), .SE(n435), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n414), .SE(n433), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n414), .SE(n431), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n414), .SE(n429), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n414), .SE(n427), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n414), .SE(n425), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n414), .SE(n423), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n414), .SE(n421), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n414), .SE(n419), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n414), .SE(n417), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2_IP  ( .D(1'b1), .SI(n564), .SE(n403), .CK(
        clk), .QN(n360) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n564), .SI(1'b1), .SE(n401), .CK(clk), 
        .Q(n359), .QN(n30) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n564), .SE(n399), .CK(
        clk), .QN(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n564), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2  ( .D(n564), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n356), .QN(n29) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n564), .SE(n393), .CK(
        clk), .Q(n338), .QN(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2_IP  ( .D(1'b1), .SI(n564), .SE(n391), .CK(
        clk), .Q(n337), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n564), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n353), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n564), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n352), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n564), .SE(n385), .CK(
        clk), .Q(n411), .QN(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n564), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n564), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n564), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n348), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n564), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n347), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n564), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n564), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n345), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n564), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n344), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n564), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n343), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n564), .SE(n367), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n564), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n564), .SE(n363), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n564), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n339) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n415), .SE(n521), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n335) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n415), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n336) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n415), .SE(n509), .CK(clk), .Q(n561), 
        .QN(n28) );
  AND2_X1 U2 ( .A1(n55), .A2(n56), .ZN(n262) );
  INV_X2 U3 ( .A(n33), .ZN(n177) );
  BUF_X1 U4 ( .A(en), .Z(n223) );
  BUF_X1 U5 ( .A(n413), .Z(n414) );
  INV_X2 U6 ( .A(n564), .ZN(n413) );
  BUF_X2 U7 ( .A(en), .Z(n12) );
  BUF_X2 U8 ( .A(en), .Z(n11) );
  BUF_X2 U9 ( .A(en), .Z(n334) );
  NAND2_X1 U10 ( .A1(n6), .A2(n5), .ZN(n121) );
  BUF_X1 U11 ( .A(n413), .Z(n415) );
  NAND2_X1 U12 ( .A1(n191), .A2(n7), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n193), .A2(n192), .ZN(n5) );
  OR2_X1 U14 ( .A1(n193), .A2(n192), .ZN(n7) );
  INV_X1 U15 ( .A(rst_n), .ZN(n564) );
  OAI22_X1 U16 ( .A1(n177), .A2(n46), .B1(n176), .B2(n335), .ZN(n149) );
  INV_X1 U17 ( .A(n335), .ZN(n333) );
  NAND2_X1 U18 ( .A1(n199), .A2(n198), .ZN(n200) );
  XNOR2_X1 U19 ( .A(n191), .B(n8), .ZN(n199) );
  XNOR2_X1 U20 ( .A(n193), .B(n192), .ZN(n8) );
  XNOR2_X1 U21 ( .A(n336), .B(\mult_x_1/a[4] ), .ZN(n9) );
  INV_X1 U22 ( .A(n98), .ZN(n50) );
  XNOR2_X1 U23 ( .A(n84), .B(n83), .ZN(n85) );
  NAND2_X1 U24 ( .A1(n90), .A2(n27), .ZN(n94) );
  INV_X1 U25 ( .A(n121), .ZN(n111) );
  XOR2_X1 U26 ( .A(n336), .B(\mult_x_1/a[4] ), .Z(n43) );
  XNOR2_X1 U27 ( .A(n139), .B(n69), .ZN(n167) );
  NAND2_X1 U28 ( .A1(n84), .A2(n83), .ZN(n79) );
  NOR2_X1 U29 ( .A1(n84), .A2(n83), .ZN(n80) );
  NAND2_X1 U30 ( .A1(n53), .A2(n52), .ZN(n126) );
  NAND2_X1 U31 ( .A1(n100), .A2(n51), .ZN(n53) );
  NAND2_X1 U32 ( .A1(n50), .A2(n49), .ZN(n51) );
  NAND2_X1 U33 ( .A1(n94), .A2(n93), .ZN(n115) );
  NAND2_X1 U34 ( .A1(n92), .A2(n91), .ZN(n93) );
  NAND2_X1 U35 ( .A1(n112), .A2(n344), .ZN(n113) );
  NAND2_X1 U36 ( .A1(n111), .A2(n223), .ZN(n114) );
  INV_X1 U37 ( .A(n223), .ZN(n112) );
  NAND2_X1 U38 ( .A1(n122), .A2(n121), .ZN(n123) );
  XNOR2_X1 U39 ( .A(n86), .B(n85), .ZN(n117) );
  BUF_X1 U40 ( .A(n176), .Z(n10) );
  NAND2_X1 U41 ( .A1(n31), .A2(n32), .ZN(n176) );
  INV_X1 U42 ( .A(n38), .ZN(n243) );
  NAND2_X1 U43 ( .A1(n141), .A2(n140), .ZN(n164) );
  OR2_X1 U44 ( .A1(n63), .A2(n62), .ZN(n92) );
  OAI21_X1 U45 ( .B1(n81), .B2(n80), .A(n79), .ZN(n165) );
  INV_X1 U46 ( .A(n86), .ZN(n81) );
  NAND2_X1 U47 ( .A1(n43), .A2(n35), .ZN(n13) );
  NAND2_X1 U48 ( .A1(n43), .A2(n35), .ZN(n157) );
  XOR2_X1 U49 ( .A(n14), .B(n336), .Z(n36) );
  XNOR2_X1 U50 ( .A(n15), .B(n18), .ZN(n32) );
  XNOR2_X1 U51 ( .A(n28), .B(\mult_x_1/a[2] ), .ZN(n38) );
  NAND2_X1 U52 ( .A1(n98), .A2(n99), .ZN(n52) );
  XNOR2_X1 U53 ( .A(n99), .B(n98), .ZN(n101) );
  INV_X1 U54 ( .A(n99), .ZN(n49) );
  OR2_X1 U55 ( .A1(n92), .A2(n91), .ZN(n27) );
  INV_X1 U56 ( .A(n55), .ZN(n58) );
  XOR2_X1 U57 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n31) );
  XNOR2_X1 U58 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n47) );
  INV_X1 U59 ( .A(n32), .ZN(n33) );
  XNOR2_X1 U60 ( .A(n333), .B(\mult_x_1/n286 ), .ZN(n42) );
  OAI22_X1 U61 ( .A1(n176), .A2(n47), .B1(n177), .B2(n42), .ZN(n104) );
  NAND2_X1 U62 ( .A1(n561), .A2(n17), .ZN(n246) );
  XNOR2_X1 U63 ( .A(n561), .B(\mult_x_1/n281 ), .ZN(n106) );
  AND2_X1 U64 ( .A1(n563), .A2(\mult_x_1/n281 ), .ZN(n131) );
  XNOR2_X1 U65 ( .A(n131), .B(n561), .ZN(n39) );
  OAI22_X1 U66 ( .A1(n246), .A2(n106), .B1(n39), .B2(n17), .ZN(n103) );
  NAND2_X1 U67 ( .A1(n16), .A2(\mult_x_1/n310 ), .ZN(n41) );
  INV_X1 U68 ( .A(n41), .ZN(n34) );
  AND2_X1 U69 ( .A1(\mult_x_1/n288 ), .A2(n34), .ZN(n102) );
  XNOR2_X1 U70 ( .A(n562), .B(n20), .ZN(n35) );
  XNOR2_X1 U71 ( .A(n562), .B(\mult_x_1/n284 ), .ZN(n44) );
  XNOR2_X1 U72 ( .A(n562), .B(\mult_x_1/n283 ), .ZN(n60) );
  OAI22_X1 U73 ( .A1(n157), .A2(n44), .B1(n43), .B2(n60), .ZN(n63) );
  INV_X1 U74 ( .A(n38), .ZN(n37) );
  NAND2_X2 U75 ( .A1(n37), .A2(n36), .ZN(n241) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n45) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n61) );
  OAI22_X1 U78 ( .A1(n241), .A2(n45), .B1(n243), .B2(n61), .ZN(n62) );
  XNOR2_X1 U79 ( .A(n63), .B(n62), .ZN(n56) );
  XNOR2_X1 U80 ( .A(n58), .B(n56), .ZN(n100) );
  AOI21_X1 U81 ( .B1(n246), .B2(n17), .A(n39), .ZN(n40) );
  INV_X1 U82 ( .A(n40), .ZN(n66) );
  NOR2_X1 U83 ( .A1(n21), .A2(n41), .ZN(n65) );
  XNOR2_X1 U84 ( .A(n333), .B(\mult_x_1/n285 ), .ZN(n59) );
  OAI22_X1 U85 ( .A1(n176), .A2(n42), .B1(n177), .B2(n59), .ZN(n64) );
  XNOR2_X1 U86 ( .A(n562), .B(\mult_x_1/n285 ), .ZN(n105) );
  INV_X1 U87 ( .A(n9), .ZN(n219) );
  OAI22_X1 U88 ( .A1(n13), .A2(n105), .B1(n219), .B2(n44), .ZN(n110) );
  XNOR2_X1 U89 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n107) );
  OAI22_X1 U90 ( .A1(n241), .A2(n107), .B1(n243), .B2(n45), .ZN(n109) );
  OR2_X1 U91 ( .A1(\mult_x_1/n288 ), .A2(n335), .ZN(n46) );
  XNOR2_X1 U92 ( .A(n333), .B(\mult_x_1/n288 ), .ZN(n48) );
  OAI22_X1 U93 ( .A1(n176), .A2(n48), .B1(n177), .B2(n47), .ZN(n148) );
  INV_X1 U94 ( .A(n126), .ZN(n54) );
  NAND2_X1 U95 ( .A1(n54), .A2(n12), .ZN(n68) );
  XNOR2_X1 U96 ( .A(n333), .B(\mult_x_1/n284 ), .ZN(n71) );
  OAI22_X1 U97 ( .A1(n10), .A2(n59), .B1(n177), .B2(n71), .ZN(n76) );
  XNOR2_X1 U98 ( .A(n562), .B(\mult_x_1/n282 ), .ZN(n78) );
  OAI22_X1 U99 ( .A1(n13), .A2(n60), .B1(n219), .B2(n78), .ZN(n75) );
  XNOR2_X1 U100 ( .A(n131), .B(\mult_x_1/n312 ), .ZN(n72) );
  OAI22_X1 U101 ( .A1(n241), .A2(n61), .B1(n72), .B2(n243), .ZN(n88) );
  INV_X1 U102 ( .A(n88), .ZN(n74) );
  NOR2_X1 U103 ( .A1(n22), .A2(n41), .ZN(n91) );
  XNOR2_X1 U104 ( .A(n92), .B(n91), .ZN(n67) );
  FA_X1 U105 ( .A(n66), .B(n65), .CI(n64), .CO(n90), .S(n98) );
  XNOR2_X1 U106 ( .A(n67), .B(n90), .ZN(n260) );
  OAI22_X1 U107 ( .A1(n68), .A2(n127), .B1(n12), .B2(n337), .ZN(n391) );
  XNOR2_X1 U108 ( .A(n562), .B(\mult_x_1/n281 ), .ZN(n77) );
  XNOR2_X1 U109 ( .A(n131), .B(n562), .ZN(n134) );
  OAI22_X1 U110 ( .A1(n157), .A2(n77), .B1(n134), .B2(n219), .ZN(n142) );
  INV_X1 U111 ( .A(n142), .ZN(n139) );
  XNOR2_X1 U112 ( .A(n333), .B(\mult_x_1/n283 ), .ZN(n70) );
  XNOR2_X1 U113 ( .A(n333), .B(\mult_x_1/n282 ), .ZN(n133) );
  OAI22_X1 U114 ( .A1(n176), .A2(n70), .B1(n177), .B2(n133), .ZN(n138) );
  NOR2_X1 U115 ( .A1(n23), .A2(n41), .ZN(n137) );
  XNOR2_X1 U116 ( .A(n138), .B(n137), .ZN(n69) );
  OAI22_X1 U117 ( .A1(n10), .A2(n71), .B1(n177), .B2(n70), .ZN(n89) );
  AOI21_X1 U118 ( .B1(n243), .B2(n241), .A(n72), .ZN(n73) );
  INV_X1 U119 ( .A(n73), .ZN(n87) );
  XNOR2_X1 U120 ( .A(n167), .B(n166), .ZN(n82) );
  FA_X1 U121 ( .A(n76), .B(n75), .CI(n74), .CO(n86), .S(n261) );
  OAI22_X1 U122 ( .A1(n13), .A2(n78), .B1(n219), .B2(n77), .ZN(n84) );
  NOR2_X1 U123 ( .A1(n24), .A2(n41), .ZN(n83) );
  XNOR2_X1 U124 ( .A(n82), .B(n165), .ZN(n226) );
  FA_X1 U125 ( .A(n89), .B(n88), .CI(n87), .CO(n166), .S(n116) );
  NAND2_X1 U126 ( .A1(n226), .A2(n225), .ZN(n95) );
  NAND2_X1 U127 ( .A1(n95), .A2(n11), .ZN(n97) );
  OR2_X1 U128 ( .A1(n223), .A2(n412), .ZN(n96) );
  NAND2_X1 U129 ( .A1(n97), .A2(n96), .ZN(n389) );
  XNOR2_X1 U130 ( .A(n101), .B(n100), .ZN(n122) );
  FA_X1 U131 ( .A(n104), .B(n103), .CI(n102), .CO(n55), .S(n193) );
  XNOR2_X1 U132 ( .A(n562), .B(\mult_x_1/n286 ), .ZN(n155) );
  OAI22_X1 U133 ( .A1(n13), .A2(n155), .B1(n219), .B2(n105), .ZN(n152) );
  XNOR2_X1 U134 ( .A(n561), .B(\mult_x_1/n282 ), .ZN(n146) );
  OAI22_X1 U135 ( .A1(n246), .A2(n146), .B1(n106), .B2(n17), .ZN(n151) );
  XNOR2_X1 U136 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n147) );
  OAI22_X1 U137 ( .A1(n241), .A2(n147), .B1(n243), .B2(n107), .ZN(n150) );
  FA_X1 U138 ( .A(n110), .B(n109), .CI(n108), .CO(n99), .S(n191) );
  OAI21_X1 U139 ( .B1(n122), .B2(n114), .A(n113), .ZN(n371) );
  FA_X1 U140 ( .A(n117), .B(n116), .CI(n115), .CO(n225), .S(n118) );
  NAND2_X1 U141 ( .A1(n118), .A2(n334), .ZN(n120) );
  OR2_X1 U142 ( .A1(n223), .A2(n30), .ZN(n119) );
  NAND2_X1 U143 ( .A1(n120), .A2(n119), .ZN(n401) );
  NAND2_X1 U144 ( .A1(n123), .A2(n12), .ZN(n125) );
  OR2_X1 U145 ( .A1(n334), .A2(n29), .ZN(n124) );
  NAND2_X1 U146 ( .A1(n125), .A2(n124), .ZN(n395) );
  NAND2_X1 U147 ( .A1(n127), .A2(n126), .ZN(n128) );
  NAND2_X1 U148 ( .A1(n128), .A2(n11), .ZN(n130) );
  OR2_X1 U149 ( .A1(n11), .A2(n338), .ZN(n129) );
  NAND2_X1 U150 ( .A1(n130), .A2(n129), .ZN(n393) );
  NOR2_X1 U173 ( .A1(n25), .A2(n41), .ZN(n174) );
  XNOR2_X1 U174 ( .A(n333), .B(\mult_x_1/n281 ), .ZN(n132) );
  XNOR2_X1 U175 ( .A(n131), .B(n333), .ZN(n175) );
  OAI22_X1 U176 ( .A1(n10), .A2(n132), .B1(n175), .B2(n177), .ZN(n182) );
  INV_X1 U177 ( .A(n182), .ZN(n173) );
  OAI22_X1 U178 ( .A1(n10), .A2(n133), .B1(n177), .B2(n132), .ZN(n144) );
  NAND2_X1 U179 ( .A1(n219), .A2(n157), .ZN(n136) );
  INV_X1 U180 ( .A(n134), .ZN(n135) );
  NAND2_X1 U181 ( .A1(n136), .A2(n135), .ZN(n143) );
  OAI21_X1 U182 ( .B1(n139), .B2(n138), .A(n137), .ZN(n141) );
  NAND2_X1 U183 ( .A1(n139), .A2(n138), .ZN(n140) );
  NOR2_X1 U184 ( .A1(n26), .A2(n41), .ZN(n163) );
  FA_X1 U185 ( .A(n144), .B(n143), .CI(n142), .CO(n172), .S(n162) );
  OR2_X1 U186 ( .A1(n189), .A2(n188), .ZN(n145) );
  MUX2_X1 U187 ( .A(n339), .B(n145), .S(n11), .Z(n361) );
  XNOR2_X1 U188 ( .A(n561), .B(\mult_x_1/n283 ), .ZN(n208) );
  OAI22_X1 U189 ( .A1(n246), .A2(n208), .B1(n146), .B2(n17), .ZN(n160) );
  AND2_X1 U190 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n159) );
  XNOR2_X1 U191 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n207) );
  OAI22_X1 U192 ( .A1(n241), .A2(n207), .B1(n243), .B2(n147), .ZN(n158) );
  HA_X1 U193 ( .A(n149), .B(n148), .CO(n108), .S(n195) );
  FA_X1 U194 ( .A(n152), .B(n151), .CI(n150), .CO(n192), .S(n194) );
  OR2_X1 U195 ( .A1(\mult_x_1/n288 ), .A2(n18), .ZN(n153) );
  OAI22_X1 U196 ( .A1(n13), .A2(n18), .B1(n153), .B2(n219), .ZN(n210) );
  XNOR2_X1 U197 ( .A(n562), .B(\mult_x_1/n288 ), .ZN(n154) );
  XNOR2_X1 U198 ( .A(n562), .B(\mult_x_1/n287 ), .ZN(n156) );
  OAI22_X1 U199 ( .A1(n13), .A2(n154), .B1(n219), .B2(n156), .ZN(n209) );
  OAI22_X1 U200 ( .A1(n13), .A2(n156), .B1(n219), .B2(n155), .ZN(n205) );
  FA_X1 U201 ( .A(n160), .B(n159), .CI(n158), .CO(n196), .S(n204) );
  OR2_X1 U202 ( .A1(n202), .A2(n201), .ZN(n161) );
  MUX2_X1 U203 ( .A(n340), .B(n161), .S(n223), .Z(n363) );
  FA_X1 U204 ( .A(n164), .B(n163), .CI(n162), .CO(n188), .S(n229) );
  NAND2_X1 U205 ( .A1(n165), .A2(n167), .ZN(n170) );
  NAND2_X1 U206 ( .A1(n165), .A2(n166), .ZN(n169) );
  NAND2_X1 U207 ( .A1(n167), .A2(n166), .ZN(n168) );
  NAND3_X1 U208 ( .A1(n170), .A2(n169), .A3(n168), .ZN(n228) );
  OR2_X1 U209 ( .A1(n229), .A2(n228), .ZN(n171) );
  MUX2_X1 U210 ( .A(n341), .B(n171), .S(n223), .Z(n365) );
  FA_X1 U211 ( .A(n174), .B(n173), .CI(n172), .CO(n184), .S(n189) );
  AOI21_X1 U212 ( .B1(n177), .B2(n10), .A(n175), .ZN(n178) );
  INV_X1 U213 ( .A(n178), .ZN(n180) );
  NOR2_X1 U214 ( .A1(n19), .A2(n41), .ZN(n179) );
  XOR2_X1 U215 ( .A(n180), .B(n179), .Z(n181) );
  XOR2_X1 U216 ( .A(n182), .B(n181), .Z(n183) );
  OR2_X1 U217 ( .A1(n184), .A2(n183), .ZN(n186) );
  NAND2_X1 U218 ( .A1(n184), .A2(n183), .ZN(n185) );
  NAND2_X1 U219 ( .A1(n186), .A2(n185), .ZN(n187) );
  MUX2_X1 U220 ( .A(n342), .B(n187), .S(n11), .Z(n367) );
  NAND2_X1 U221 ( .A1(n189), .A2(n188), .ZN(n190) );
  MUX2_X1 U222 ( .A(n343), .B(n190), .S(n334), .Z(n369) );
  FA_X1 U223 ( .A(n196), .B(n195), .CI(n194), .CO(n198), .S(n202) );
  NOR2_X1 U224 ( .A1(n199), .A2(n198), .ZN(n197) );
  MUX2_X1 U225 ( .A(n345), .B(n197), .S(n12), .Z(n373) );
  MUX2_X1 U226 ( .A(n346), .B(n200), .S(n11), .Z(n375) );
  NAND2_X1 U227 ( .A1(n202), .A2(n201), .ZN(n203) );
  MUX2_X1 U228 ( .A(n347), .B(n203), .S(n334), .Z(n377) );
  FA_X1 U229 ( .A(n206), .B(n205), .CI(n204), .CO(n201), .S(n213) );
  XNOR2_X1 U230 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n220) );
  OAI22_X1 U231 ( .A1(n241), .A2(n220), .B1(n243), .B2(n207), .ZN(n217) );
  XNOR2_X1 U232 ( .A(n561), .B(\mult_x_1/n284 ), .ZN(n218) );
  OAI22_X1 U233 ( .A1(n246), .A2(n218), .B1(n208), .B2(n17), .ZN(n216) );
  HA_X1 U234 ( .A(n210), .B(n209), .CO(n206), .S(n215) );
  NOR2_X1 U235 ( .A1(n213), .A2(n212), .ZN(n211) );
  MUX2_X1 U236 ( .A(n348), .B(n211), .S(n12), .Z(n379) );
  NAND2_X1 U237 ( .A1(n213), .A2(n212), .ZN(n214) );
  MUX2_X1 U238 ( .A(n349), .B(n214), .S(n11), .Z(n381) );
  FA_X1 U239 ( .A(n217), .B(n216), .CI(n215), .CO(n212), .S(n222) );
  XNOR2_X1 U240 ( .A(n561), .B(\mult_x_1/n285 ), .ZN(n236) );
  OAI22_X1 U241 ( .A1(n246), .A2(n236), .B1(n218), .B2(n17), .ZN(n233) );
  AND2_X1 U242 ( .A1(\mult_x_1/n288 ), .A2(n9), .ZN(n232) );
  XNOR2_X1 U243 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n234) );
  OAI22_X1 U244 ( .A1(n241), .A2(n234), .B1(n243), .B2(n220), .ZN(n231) );
  OR2_X1 U245 ( .A1(n222), .A2(n221), .ZN(n257) );
  NAND2_X1 U246 ( .A1(n222), .A2(n221), .ZN(n255) );
  NAND2_X1 U247 ( .A1(n257), .A2(n255), .ZN(n224) );
  MUX2_X1 U248 ( .A(n350), .B(n224), .S(n334), .Z(n383) );
  NOR2_X1 U249 ( .A1(n226), .A2(n225), .ZN(n227) );
  MUX2_X1 U250 ( .A(n351), .B(n227), .S(n334), .Z(n385) );
  NAND2_X1 U251 ( .A1(n229), .A2(n228), .ZN(n230) );
  MUX2_X1 U252 ( .A(n352), .B(n230), .S(n12), .Z(n387) );
  FA_X1 U253 ( .A(n233), .B(n232), .CI(n231), .CO(n221), .S(n254) );
  XNOR2_X1 U254 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n235) );
  OAI22_X1 U255 ( .A1(n241), .A2(n235), .B1(n243), .B2(n234), .ZN(n238) );
  XNOR2_X1 U256 ( .A(n561), .B(\mult_x_1/n286 ), .ZN(n242) );
  OAI22_X1 U257 ( .A1(n246), .A2(n242), .B1(n236), .B2(n17), .ZN(n237) );
  NOR2_X1 U258 ( .A1(n254), .A2(n253), .ZN(n280) );
  HA_X1 U259 ( .A(n238), .B(n237), .CO(n253), .S(n251) );
  INV_X1 U260 ( .A(\mult_x_1/n312 ), .ZN(n240) );
  OR2_X1 U261 ( .A1(\mult_x_1/n288 ), .A2(n240), .ZN(n239) );
  OAI22_X1 U262 ( .A1(n241), .A2(n240), .B1(n239), .B2(n243), .ZN(n250) );
  OR2_X1 U263 ( .A1(n251), .A2(n250), .ZN(n276) );
  XNOR2_X1 U264 ( .A(n561), .B(\mult_x_1/n287 ), .ZN(n245) );
  OAI22_X1 U265 ( .A1(n246), .A2(n245), .B1(n242), .B2(n17), .ZN(n249) );
  INV_X1 U266 ( .A(n243), .ZN(n244) );
  AND2_X1 U267 ( .A1(\mult_x_1/n288 ), .A2(n244), .ZN(n248) );
  NOR2_X1 U268 ( .A1(n249), .A2(n248), .ZN(n269) );
  OAI22_X1 U269 ( .A1(n246), .A2(\mult_x_1/n288 ), .B1(n245), .B2(n17), .ZN(
        n266) );
  OR2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n247) );
  NAND2_X1 U271 ( .A1(n247), .A2(n246), .ZN(n265) );
  NAND2_X1 U272 ( .A1(n266), .A2(n265), .ZN(n272) );
  NAND2_X1 U273 ( .A1(n249), .A2(n248), .ZN(n270) );
  OAI21_X1 U274 ( .B1(n269), .B2(n272), .A(n270), .ZN(n277) );
  NAND2_X1 U275 ( .A1(n251), .A2(n250), .ZN(n275) );
  INV_X1 U276 ( .A(n275), .ZN(n252) );
  AOI21_X1 U277 ( .B1(n276), .B2(n277), .A(n252), .ZN(n283) );
  NAND2_X1 U278 ( .A1(n254), .A2(n253), .ZN(n281) );
  OAI21_X1 U279 ( .B1(n280), .B2(n283), .A(n281), .ZN(n259) );
  INV_X1 U280 ( .A(n255), .ZN(n256) );
  AOI21_X1 U281 ( .B1(n257), .B2(n259), .A(n256), .ZN(n258) );
  MUX2_X1 U282 ( .A(n357), .B(n258), .S(n11), .Z(n397) );
  MUX2_X1 U283 ( .A(n358), .B(n259), .S(n334), .Z(n399) );
  FA_X1 U284 ( .A(n262), .B(n261), .CI(n260), .CO(n263), .S(n127) );
  MUX2_X1 U285 ( .A(n360), .B(n263), .S(n12), .Z(n403) );
  MUX2_X1 U286 ( .A(product[0]), .B(n525), .S(n12), .Z(n417) );
  MUX2_X1 U287 ( .A(n525), .B(n526), .S(n334), .Z(n419) );
  AND2_X1 U288 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n264) );
  MUX2_X1 U289 ( .A(n526), .B(n264), .S(n11), .Z(n421) );
  MUX2_X1 U290 ( .A(product[1]), .B(n528), .S(n223), .Z(n423) );
  MUX2_X1 U291 ( .A(n528), .B(n529), .S(n334), .Z(n425) );
  OR2_X1 U292 ( .A1(n266), .A2(n265), .ZN(n267) );
  AND2_X1 U293 ( .A1(n267), .A2(n272), .ZN(n268) );
  MUX2_X1 U294 ( .A(n529), .B(n268), .S(n11), .Z(n427) );
  MUX2_X1 U295 ( .A(product[2]), .B(n531), .S(n12), .Z(n429) );
  MUX2_X1 U296 ( .A(n531), .B(n532), .S(n334), .Z(n431) );
  INV_X1 U297 ( .A(n269), .ZN(n271) );
  NAND2_X1 U298 ( .A1(n271), .A2(n270), .ZN(n273) );
  XOR2_X1 U299 ( .A(n273), .B(n272), .Z(n274) );
  MUX2_X1 U300 ( .A(n532), .B(n274), .S(n11), .Z(n433) );
  MUX2_X1 U301 ( .A(product[3]), .B(n534), .S(n223), .Z(n435) );
  MUX2_X1 U302 ( .A(n534), .B(n535), .S(n12), .Z(n437) );
  NAND2_X1 U303 ( .A1(n276), .A2(n275), .ZN(n278) );
  XNOR2_X1 U304 ( .A(n278), .B(n277), .ZN(n279) );
  MUX2_X1 U305 ( .A(n535), .B(n279), .S(n334), .Z(n439) );
  MUX2_X1 U306 ( .A(product[4]), .B(n537), .S(n11), .Z(n441) );
  MUX2_X1 U307 ( .A(n537), .B(n538), .S(n12), .Z(n443) );
  INV_X1 U308 ( .A(n280), .ZN(n282) );
  NAND2_X1 U309 ( .A1(n282), .A2(n281), .ZN(n284) );
  XOR2_X1 U310 ( .A(n284), .B(n283), .Z(n285) );
  MUX2_X1 U311 ( .A(n538), .B(n285), .S(n12), .Z(n445) );
  MUX2_X1 U312 ( .A(product[5]), .B(n540), .S(n12), .Z(n447) );
  XNOR2_X1 U313 ( .A(n350), .B(n358), .ZN(n286) );
  MUX2_X1 U314 ( .A(n540), .B(n286), .S(n334), .Z(n449) );
  MUX2_X1 U315 ( .A(product[6]), .B(n542), .S(n334), .Z(n451) );
  NAND2_X1 U316 ( .A1(n406), .A2(n349), .ZN(n287) );
  XOR2_X1 U317 ( .A(n287), .B(n357), .Z(n288) );
  MUX2_X1 U318 ( .A(n542), .B(n288), .S(n334), .Z(n453) );
  MUX2_X1 U319 ( .A(product[7]), .B(n544), .S(n11), .Z(n455) );
  OAI21_X1 U320 ( .B1(n348), .B2(n357), .A(n349), .ZN(n291) );
  NAND2_X1 U321 ( .A1(n340), .A2(n347), .ZN(n289) );
  XNOR2_X1 U322 ( .A(n291), .B(n289), .ZN(n290) );
  MUX2_X1 U323 ( .A(n544), .B(n290), .S(n11), .Z(n457) );
  MUX2_X1 U324 ( .A(product[8]), .B(n546), .S(n11), .Z(n459) );
  AOI21_X1 U325 ( .B1(n291), .B2(n340), .A(n408), .ZN(n294) );
  NAND2_X1 U326 ( .A1(n409), .A2(n346), .ZN(n292) );
  XOR2_X1 U327 ( .A(n294), .B(n292), .Z(n293) );
  MUX2_X1 U328 ( .A(n546), .B(n293), .S(n334), .Z(n461) );
  MUX2_X1 U329 ( .A(product[9]), .B(n548), .S(n11), .Z(n463) );
  OAI21_X1 U330 ( .B1(n294), .B2(n345), .A(n346), .ZN(n302) );
  INV_X1 U331 ( .A(n302), .ZN(n297) );
  NAND2_X1 U332 ( .A1(n410), .A2(n356), .ZN(n295) );
  XOR2_X1 U333 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U334 ( .A(n548), .B(n296), .S(n12), .Z(n465) );
  MUX2_X1 U335 ( .A(product[10]), .B(n550), .S(n11), .Z(n467) );
  OAI21_X1 U336 ( .B1(n297), .B2(n344), .A(n356), .ZN(n299) );
  NAND2_X1 U337 ( .A1(n337), .A2(n355), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U339 ( .A(n550), .B(n300), .S(n334), .Z(n469) );
  MUX2_X1 U340 ( .A(product[11]), .B(n552), .S(n12), .Z(n471) );
  NOR2_X1 U341 ( .A1(n354), .A2(n344), .ZN(n303) );
  OAI21_X1 U342 ( .B1(n354), .B2(n356), .A(n355), .ZN(n301) );
  AOI21_X1 U343 ( .B1(n303), .B2(n302), .A(n301), .ZN(n330) );
  OR2_X1 U344 ( .A1(n359), .A2(n360), .ZN(n324) );
  NAND2_X1 U345 ( .A1(n359), .A2(n360), .ZN(n317) );
  NAND2_X1 U346 ( .A1(n324), .A2(n317), .ZN(n304) );
  XOR2_X1 U347 ( .A(n330), .B(n304), .Z(n305) );
  MUX2_X1 U348 ( .A(n552), .B(n305), .S(n223), .Z(n473) );
  MUX2_X1 U349 ( .A(product[12]), .B(n554), .S(n223), .Z(n475) );
  INV_X1 U350 ( .A(n324), .ZN(n306) );
  OAI21_X1 U351 ( .B1(n330), .B2(n306), .A(n317), .ZN(n308) );
  NAND2_X1 U352 ( .A1(n411), .A2(n353), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U354 ( .A(n554), .B(n309), .S(n223), .Z(n477) );
  MUX2_X1 U355 ( .A(product[13]), .B(n556), .S(n223), .Z(n479) );
  NAND2_X1 U356 ( .A1(n324), .A2(n411), .ZN(n312) );
  INV_X1 U357 ( .A(n317), .ZN(n310) );
  AOI21_X1 U358 ( .B1(n310), .B2(n411), .A(n412), .ZN(n311) );
  OAI21_X1 U359 ( .B1(n330), .B2(n312), .A(n311), .ZN(n314) );
  NAND2_X1 U360 ( .A1(n341), .A2(n352), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U362 ( .A(n556), .B(n315), .S(n11), .Z(n481) );
  MUX2_X1 U363 ( .A(product[14]), .B(n558), .S(n334), .Z(n483) );
  AND2_X1 U364 ( .A1(n411), .A2(n341), .ZN(n325) );
  NAND2_X1 U365 ( .A1(n324), .A2(n325), .ZN(n320) );
  NAND2_X1 U366 ( .A1(n411), .A2(n341), .ZN(n318) );
  AOI21_X1 U367 ( .B1(n412), .B2(n341), .A(n407), .ZN(n316) );
  OAI21_X1 U368 ( .B1(n318), .B2(n317), .A(n316), .ZN(n327) );
  INV_X1 U369 ( .A(n327), .ZN(n319) );
  OAI21_X1 U370 ( .B1(n330), .B2(n320), .A(n319), .ZN(n322) );
  NAND2_X1 U371 ( .A1(n339), .A2(n343), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U373 ( .A(n558), .B(n323), .S(n12), .Z(n485) );
  MUX2_X1 U374 ( .A(product[15]), .B(n560), .S(n223), .Z(n487) );
  AND2_X1 U375 ( .A1(n324), .A2(n339), .ZN(n326) );
  NAND2_X1 U376 ( .A1(n326), .A2(n325), .ZN(n329) );
  AOI21_X1 U377 ( .B1(n327), .B2(n339), .A(n405), .ZN(n328) );
  OAI21_X1 U378 ( .B1(n330), .B2(n329), .A(n328), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n331), .B(n342), .ZN(n332) );
  MUX2_X1 U380 ( .A(n560), .B(n332), .S(n11), .Z(n489) );
  MUX2_X1 U381 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n334), .Z(n491) );
  MUX2_X1 U382 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n12), .Z(n493) );
  MUX2_X1 U383 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n334), .Z(n495) );
  MUX2_X1 U384 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n11), .Z(n497) );
  MUX2_X1 U385 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n12), .Z(n499) );
  MUX2_X1 U386 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n223), .Z(n501) );
  MUX2_X1 U387 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n334), .Z(n503) );
  MUX2_X1 U388 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n11), .Z(n505) );
  MUX2_X1 U389 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n334), .Z(n507) );
  MUX2_X1 U390 ( .A(n561), .B(A_extended[1]), .S(n12), .Z(n509) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n12), .Z(n511) );
  MUX2_X1 U392 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n12), .Z(n513) );
  MUX2_X1 U393 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n11), .Z(n515) );
  MUX2_X1 U394 ( .A(n562), .B(A_extended[5]), .S(n11), .Z(n517) );
  MUX2_X1 U395 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n334), .Z(n519) );
  MUX2_X1 U396 ( .A(n333), .B(A_extended[7]), .S(n12), .Z(n521) );
  OR2_X1 U397 ( .A1(n223), .A2(n563), .ZN(n523) );
endmodule


module conv_128_32_DW_mult_pipe_J1_15 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n311 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n360, n362, n364, n366, n368,
         n370, n372, n374, n376, n378, n380, n382, n384, n386, n388, n390,
         n392, n394, n396, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n412, n414, n416, n418, n420, n422,
         n424, n426, n428, n430, n432, n434, n436, n438, n440, n442, n444,
         n446, n448, n450, n452, n454, n456, n458, n460, n462, n464, n466,
         n468, n470, n472, n474, n476, n478, n480, n482, n484, n486, n488,
         n490, n492, n494, n496, n498, n500, n502, n504, n506, n508, n510,
         n512, n514, n516, n518, n520, n522, n523, n525, n526, n528, n529,
         n531, n532, n534, n535, n537, n538, n540, n542, n544, n546, n548,
         n550, n552, n554, n556, n558, n559, n560, n561, n562, n563;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n410), .SE(n520), .CK(clk), .Q(n562), 
        .QN(n41) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n410), .SE(n518), .CK(clk), .Q(n561), 
        .QN(n40) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n410), .SE(n516), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n410), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n42) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n410), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n31) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n410), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n33) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n410), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n37) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n408), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n39) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n409), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n38) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n407), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n36) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n410), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n35) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n407), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n34) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n407), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n407), .SE(n486), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n407), .SE(n484), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n407), .SE(n482), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n407), .SE(n480), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n407), .SE(n478), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n409), .SE(n476), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n408), .SE(n474), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n410), .SE(n472), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n407), .SE(n470), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n407), .SE(n468), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n407), .SE(n466), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n407), .SE(n464), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n407), .SE(n462), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n407), .SE(n460), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n407), .SE(n458), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n407), .SE(n456), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n409), .SE(n454), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n409), .SE(n452), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n409), .SE(n450), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n409), .SE(n448), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n409), .SE(n446), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n409), .SE(n444), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n409), .SE(n442), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n409), .SE(n440), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n409), .SE(n438), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n409), .SE(n436), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n409), .SE(n434), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n408), .SE(n432), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n408), .SE(n430), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n408), .SE(n428), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n408), .SE(n426), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n408), .SE(n424), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n408), .SE(n422), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n408), .SE(n420), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n408), .SE(n418), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n408), .SE(n416), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n408), .SE(n414), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n408), .SE(n412), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n563), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n563), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n356), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n563), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n355), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n563), .SE(n390), .CK(
        clk), .Q(n337), .QN(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n563), .SE(n388), .CK(
        clk), .Q(n336), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n563), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n563), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n351), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n563), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n350), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n563), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n563), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n348), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n563), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n347), .QN(n44) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n563), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n346), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n563), .SE(n372), .CK(
        clk), .Q(n404), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n563), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n344), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n563), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n343), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2_IP  ( .D(1'b1), .SI(n563), .SE(n366), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n563), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n563), .SE(n362), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n563), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n563), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n338) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n410), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n335) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n410), .SE(n510), .CK(clk), .Q(n560), 
        .QN(n32) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n410), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n24) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n410), .SE(n506), .CK(clk), .Q(n559), 
        .QN(n45) );
  AND2_X1 U2 ( .A1(n562), .A2(\mult_x_1/n281 ), .ZN(n120) );
  BUF_X2 U3 ( .A(\mult_x_1/n311 ), .Z(n29) );
  CLKBUF_X1 U4 ( .A(n183), .Z(n5) );
  BUF_X1 U5 ( .A(n183), .Z(n6) );
  BUF_X2 U6 ( .A(n183), .Z(n7) );
  BUF_X1 U7 ( .A(n407), .Z(n408) );
  BUF_X1 U8 ( .A(n407), .Z(n409) );
  BUF_X1 U9 ( .A(n407), .Z(n410) );
  INV_X1 U10 ( .A(n563), .ZN(n407) );
  INV_X1 U11 ( .A(n48), .ZN(n184) );
  NAND2_X1 U12 ( .A1(n46), .A2(n47), .ZN(n183) );
  OR2_X1 U13 ( .A1(n97), .A2(n202), .ZN(n20) );
  NAND2_X1 U14 ( .A1(n14), .A2(n13), .ZN(n231) );
  NAND2_X1 U15 ( .A1(n204), .A2(n15), .ZN(n14) );
  XNOR2_X1 U16 ( .A(n204), .B(n18), .ZN(n212) );
  NAND2_X1 U17 ( .A1(n17), .A2(n16), .ZN(n15) );
  XNOR2_X1 U18 ( .A(n206), .B(n205), .ZN(n18) );
  INV_X1 U19 ( .A(n205), .ZN(n16) );
  NAND2_X1 U20 ( .A1(n206), .A2(n205), .ZN(n13) );
  INV_X1 U21 ( .A(n206), .ZN(n17) );
  INV_X1 U22 ( .A(rst_n), .ZN(n563) );
  NAND2_X1 U23 ( .A1(n561), .A2(n41), .ZN(n186) );
  NAND2_X1 U24 ( .A1(n9), .A2(n8), .ZN(n128) );
  NAND2_X1 U25 ( .A1(n238), .A2(n164), .ZN(n8) );
  INV_X1 U26 ( .A(n121), .ZN(n9) );
  OAI21_X1 U27 ( .B1(n11), .B2(n97), .A(n10), .ZN(n446) );
  NAND2_X1 U28 ( .A1(n97), .A2(n538), .ZN(n10) );
  XNOR2_X1 U29 ( .A(n292), .B(n12), .ZN(n11) );
  INV_X1 U30 ( .A(n291), .ZN(n12) );
  OAI21_X1 U31 ( .B1(n203), .B2(n20), .A(n19), .ZN(n372) );
  NAND2_X1 U32 ( .A1(n97), .A2(n345), .ZN(n19) );
  OAI22_X1 U33 ( .A1(n107), .A2(n248), .B1(n26), .B2(n55), .ZN(n139) );
  INV_X1 U34 ( .A(n251), .ZN(n248) );
  XNOR2_X1 U35 ( .A(n45), .B(\mult_x_1/a[2] ), .ZN(n251) );
  XNOR2_X1 U36 ( .A(n143), .B(n144), .ZN(n113) );
  XNOR2_X1 U37 ( .A(n65), .B(n64), .ZN(n84) );
  NAND2_X1 U38 ( .A1(n177), .A2(n176), .ZN(n228) );
  NAND2_X1 U39 ( .A1(n173), .A2(n172), .ZN(n177) );
  OR2_X1 U40 ( .A1(n98), .A2(n97), .ZN(n99) );
  XOR2_X1 U41 ( .A(n42), .B(n32), .Z(n21) );
  CLKBUF_X1 U42 ( .A(n560), .Z(n22) );
  OAI22_X1 U43 ( .A1(n164), .A2(n66), .B1(n238), .B2(n54), .ZN(n23) );
  XNOR2_X1 U44 ( .A(n24), .B(n560), .ZN(n53) );
  XNOR2_X1 U45 ( .A(n137), .B(n136), .ZN(n175) );
  XNOR2_X1 U46 ( .A(n135), .B(n134), .ZN(n137) );
  FA_X1 U47 ( .A(n140), .B(n27), .CI(n138), .CO(n25) );
  NAND2_X1 U48 ( .A1(n53), .A2(n52), .ZN(n26) );
  INV_X1 U49 ( .A(n109), .ZN(n27) );
  XNOR2_X1 U50 ( .A(n42), .B(n32), .ZN(n51) );
  INV_X1 U51 ( .A(n40), .ZN(n28) );
  XNOR2_X1 U52 ( .A(n146), .B(n113), .ZN(n131) );
  NAND2_X1 U53 ( .A1(n103), .A2(n102), .ZN(n104) );
  OR2_X1 U54 ( .A1(n61), .A2(n23), .ZN(n103) );
  AND2_X1 U55 ( .A1(n65), .A2(n63), .ZN(n30) );
  BUF_X1 U56 ( .A(en), .Z(n265) );
  INV_X1 U57 ( .A(n265), .ZN(n97) );
  OR2_X1 U58 ( .A1(n103), .A2(n102), .ZN(n43) );
  XOR2_X1 U59 ( .A(\mult_x_1/a[6] ), .B(n561), .Z(n46) );
  XNOR2_X1 U60 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n47) );
  XNOR2_X1 U61 ( .A(n561), .B(\mult_x_1/n287 ), .ZN(n70) );
  INV_X1 U62 ( .A(n47), .ZN(n48) );
  XNOR2_X1 U63 ( .A(n28), .B(\mult_x_1/n286 ), .ZN(n59) );
  OAI22_X1 U64 ( .A1(n7), .A2(n70), .B1(n184), .B2(n59), .ZN(n87) );
  NAND2_X1 U65 ( .A1(n559), .A2(n31), .ZN(n253) );
  XNOR2_X1 U66 ( .A(n559), .B(\mult_x_1/n281 ), .ZN(n89) );
  XNOR2_X1 U67 ( .A(n120), .B(n559), .ZN(n56) );
  OAI22_X1 U68 ( .A1(n253), .A2(n89), .B1(n56), .B2(n31), .ZN(n86) );
  INV_X1 U69 ( .A(n186), .ZN(n49) );
  AND2_X1 U70 ( .A1(\mult_x_1/n288 ), .A2(n49), .ZN(n85) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n311 ), .B(n42), .ZN(n50) );
  NAND2_X1 U72 ( .A1(n50), .A2(n51), .ZN(n164) );
  XNOR2_X1 U73 ( .A(n29), .B(\mult_x_1/n284 ), .ZN(n66) );
  INV_X2 U74 ( .A(n21), .ZN(n238) );
  XNOR2_X1 U75 ( .A(n29), .B(\mult_x_1/n283 ), .ZN(n54) );
  OAI22_X1 U76 ( .A1(n164), .A2(n66), .B1(n238), .B2(n54), .ZN(n60) );
  INV_X1 U77 ( .A(n251), .ZN(n52) );
  NAND2_X1 U78 ( .A1(n53), .A2(n52), .ZN(n67) );
  XNOR2_X1 U79 ( .A(n560), .B(\mult_x_1/n282 ), .ZN(n68) );
  XNOR2_X1 U80 ( .A(n560), .B(\mult_x_1/n281 ), .ZN(n55) );
  OAI22_X1 U81 ( .A1(n26), .A2(n68), .B1(n248), .B2(n55), .ZN(n61) );
  XNOR2_X1 U82 ( .A(n60), .B(n61), .ZN(n63) );
  XNOR2_X1 U83 ( .A(n28), .B(\mult_x_1/n285 ), .ZN(n58) );
  XNOR2_X1 U84 ( .A(n28), .B(\mult_x_1/n284 ), .ZN(n106) );
  OAI22_X1 U85 ( .A1(n7), .A2(n58), .B1(n184), .B2(n106), .ZN(n111) );
  XNOR2_X1 U86 ( .A(n29), .B(\mult_x_1/n282 ), .ZN(n112) );
  OAI22_X1 U87 ( .A1(n164), .A2(n54), .B1(n238), .B2(n112), .ZN(n110) );
  XNOR2_X1 U88 ( .A(n120), .B(n560), .ZN(n107) );
  INV_X1 U89 ( .A(n139), .ZN(n109) );
  AOI21_X1 U90 ( .B1(n253), .B2(n31), .A(n56), .ZN(n57) );
  INV_X1 U91 ( .A(n57), .ZN(n74) );
  NOR2_X1 U92 ( .A1(n34), .A2(n186), .ZN(n73) );
  OAI22_X1 U93 ( .A1(n6), .A2(n59), .B1(n184), .B2(n58), .ZN(n72) );
  NOR2_X1 U94 ( .A1(n35), .A2(n186), .ZN(n102) );
  XNOR2_X1 U95 ( .A(n103), .B(n102), .ZN(n62) );
  XNOR2_X1 U96 ( .A(n101), .B(n62), .ZN(n114) );
  INV_X1 U97 ( .A(n63), .ZN(n64) );
  XNOR2_X1 U98 ( .A(n29), .B(\mult_x_1/n285 ), .ZN(n88) );
  OAI22_X1 U99 ( .A1(n164), .A2(n88), .B1(n238), .B2(n66), .ZN(n93) );
  XNOR2_X1 U100 ( .A(n560), .B(\mult_x_1/n283 ), .ZN(n90) );
  OAI22_X1 U101 ( .A1(n67), .A2(n90), .B1(n248), .B2(n68), .ZN(n92) );
  OR2_X1 U102 ( .A1(\mult_x_1/n288 ), .A2(n40), .ZN(n69) );
  OAI22_X1 U103 ( .A1(n6), .A2(n40), .B1(n69), .B2(n184), .ZN(n156) );
  XNOR2_X1 U104 ( .A(n561), .B(\mult_x_1/n288 ), .ZN(n71) );
  OAI22_X1 U105 ( .A1(n5), .A2(n71), .B1(n184), .B2(n70), .ZN(n155) );
  NAND2_X1 U106 ( .A1(n84), .A2(n82), .ZN(n77) );
  FA_X1 U107 ( .A(n74), .B(n73), .CI(n72), .CO(n101), .S(n81) );
  NAND2_X1 U108 ( .A1(n84), .A2(n81), .ZN(n76) );
  NAND2_X1 U109 ( .A1(n82), .A2(n81), .ZN(n75) );
  NAND3_X1 U110 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n98) );
  OR2_X1 U111 ( .A1(n265), .A2(n337), .ZN(n78) );
  OAI21_X1 U112 ( .B1(n98), .B2(n97), .A(n78), .ZN(n79) );
  INV_X1 U113 ( .A(n79), .ZN(n80) );
  OAI21_X1 U114 ( .B1(n100), .B2(n97), .A(n80), .ZN(n390) );
  XOR2_X1 U115 ( .A(n82), .B(n81), .Z(n83) );
  XOR2_X1 U116 ( .A(n84), .B(n83), .Z(n232) );
  FA_X1 U117 ( .A(n87), .B(n86), .CI(n85), .CO(n65), .S(n206) );
  XNOR2_X1 U118 ( .A(n29), .B(\mult_x_1/n286 ), .ZN(n162) );
  OAI22_X1 U119 ( .A1(n164), .A2(n162), .B1(n238), .B2(n88), .ZN(n159) );
  XNOR2_X1 U120 ( .A(n559), .B(\mult_x_1/n282 ), .ZN(n152) );
  OAI22_X1 U121 ( .A1(n253), .A2(n152), .B1(n89), .B2(n31), .ZN(n158) );
  XNOR2_X1 U122 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n154) );
  OAI22_X1 U123 ( .A1(n67), .A2(n154), .B1(n248), .B2(n90), .ZN(n157) );
  FA_X1 U124 ( .A(n93), .B(n92), .CI(n91), .CO(n82), .S(n204) );
  NAND2_X1 U125 ( .A1(n232), .A2(n231), .ZN(n94) );
  NAND2_X1 U126 ( .A1(n94), .A2(en), .ZN(n96) );
  OR2_X1 U127 ( .A1(n265), .A2(n44), .ZN(n95) );
  NAND2_X1 U128 ( .A1(n96), .A2(n95), .ZN(n376) );
  OAI22_X1 U129 ( .A1(n100), .A2(n99), .B1(n265), .B2(n336), .ZN(n388) );
  NAND2_X1 U130 ( .A1(n101), .A2(n43), .ZN(n105) );
  NAND2_X1 U131 ( .A1(n105), .A2(n104), .ZN(n133) );
  XNOR2_X1 U132 ( .A(n561), .B(\mult_x_1/n283 ), .ZN(n124) );
  OAI22_X1 U133 ( .A1(n7), .A2(n106), .B1(n184), .B2(n124), .ZN(n140) );
  AOI21_X1 U134 ( .B1(n248), .B2(n67), .A(n107), .ZN(n108) );
  INV_X1 U135 ( .A(n108), .ZN(n138) );
  FA_X1 U136 ( .A(n110), .B(n111), .CI(n109), .CO(n146), .S(n115) );
  NOR2_X1 U137 ( .A1(n36), .A2(n186), .ZN(n143) );
  XNOR2_X1 U138 ( .A(n29), .B(\mult_x_1/n281 ), .ZN(n122) );
  OAI22_X1 U139 ( .A1(n164), .A2(n112), .B1(n238), .B2(n122), .ZN(n144) );
  FA_X1 U140 ( .A(n30), .B(n115), .CI(n114), .CO(n202), .S(n100) );
  NAND2_X1 U141 ( .A1(n203), .A2(n202), .ZN(n116) );
  NAND2_X1 U142 ( .A1(n116), .A2(en), .ZN(n118) );
  OR2_X1 U143 ( .A1(n265), .A2(n400), .ZN(n117) );
  NAND2_X1 U144 ( .A1(n118), .A2(n117), .ZN(n374) );
  NOR2_X1 U165 ( .A1(n37), .A2(n186), .ZN(n181) );
  XNOR2_X1 U166 ( .A(n28), .B(\mult_x_1/n281 ), .ZN(n119) );
  XNOR2_X1 U167 ( .A(n120), .B(n28), .ZN(n182) );
  OAI22_X1 U168 ( .A1(n6), .A2(n119), .B1(n182), .B2(n184), .ZN(n190) );
  INV_X1 U169 ( .A(n190), .ZN(n180) );
  XNOR2_X1 U170 ( .A(n561), .B(\mult_x_1/n282 ), .ZN(n123) );
  OAI22_X1 U171 ( .A1(n6), .A2(n123), .B1(n184), .B2(n119), .ZN(n129) );
  XNOR2_X1 U172 ( .A(n120), .B(n29), .ZN(n121) );
  OAI22_X1 U173 ( .A1(n164), .A2(n122), .B1(n121), .B2(n238), .ZN(n127) );
  INV_X1 U174 ( .A(n127), .ZN(n136) );
  OAI22_X1 U175 ( .A1(n5), .A2(n124), .B1(n184), .B2(n123), .ZN(n135) );
  NOR2_X1 U176 ( .A1(n38), .A2(n186), .ZN(n134) );
  OAI21_X1 U177 ( .B1(n136), .B2(n135), .A(n134), .ZN(n126) );
  NAND2_X1 U178 ( .A1(n136), .A2(n135), .ZN(n125) );
  NAND2_X1 U179 ( .A1(n126), .A2(n125), .ZN(n171) );
  NOR2_X1 U180 ( .A1(n39), .A2(n186), .ZN(n170) );
  FA_X1 U181 ( .A(n129), .B(n128), .CI(n127), .CO(n179), .S(n169) );
  OR2_X1 U182 ( .A1(n197), .A2(n196), .ZN(n130) );
  MUX2_X1 U183 ( .A(n338), .B(n130), .S(n334), .Z(n358) );
  FA_X1 U184 ( .A(n133), .B(n132), .CI(n131), .CO(n199), .S(n203) );
  INV_X1 U185 ( .A(n199), .ZN(n150) );
  FA_X1 U186 ( .A(n140), .B(n138), .CI(n27), .CO(n174), .S(n132) );
  XNOR2_X1 U187 ( .A(n175), .B(n25), .ZN(n148) );
  INV_X1 U188 ( .A(n144), .ZN(n142) );
  INV_X1 U189 ( .A(n143), .ZN(n141) );
  NAND2_X1 U190 ( .A1(n142), .A2(n141), .ZN(n145) );
  AOI22_X1 U191 ( .A1(n146), .A2(n145), .B1(n144), .B2(n143), .ZN(n147) );
  INV_X1 U192 ( .A(n147), .ZN(n172) );
  XNOR2_X1 U193 ( .A(n148), .B(n172), .ZN(n200) );
  INV_X1 U194 ( .A(n200), .ZN(n149) );
  NAND2_X1 U195 ( .A1(n150), .A2(n149), .ZN(n151) );
  MUX2_X1 U196 ( .A(n339), .B(n151), .S(n265), .Z(n360) );
  XNOR2_X1 U197 ( .A(n559), .B(\mult_x_1/n283 ), .ZN(n221) );
  OAI22_X1 U198 ( .A1(n253), .A2(n221), .B1(n152), .B2(n31), .ZN(n167) );
  INV_X1 U199 ( .A(n184), .ZN(n153) );
  AND2_X1 U200 ( .A1(\mult_x_1/n288 ), .A2(n153), .ZN(n166) );
  XNOR2_X1 U201 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n220) );
  OAI22_X1 U202 ( .A1(n67), .A2(n220), .B1(n248), .B2(n154), .ZN(n165) );
  HA_X1 U203 ( .A(n156), .B(n155), .CO(n91), .S(n208) );
  FA_X1 U204 ( .A(n159), .B(n158), .CI(n157), .CO(n205), .S(n207) );
  OR2_X1 U205 ( .A1(\mult_x_1/n288 ), .A2(n335), .ZN(n160) );
  OAI22_X1 U206 ( .A1(n164), .A2(n335), .B1(n160), .B2(n238), .ZN(n223) );
  XNOR2_X1 U207 ( .A(n29), .B(\mult_x_1/n288 ), .ZN(n161) );
  XNOR2_X1 U208 ( .A(n29), .B(\mult_x_1/n287 ), .ZN(n163) );
  OAI22_X1 U209 ( .A1(n164), .A2(n161), .B1(n238), .B2(n163), .ZN(n222) );
  OAI22_X1 U210 ( .A1(n164), .A2(n163), .B1(n238), .B2(n162), .ZN(n218) );
  FA_X1 U211 ( .A(n167), .B(n166), .CI(n165), .CO(n209), .S(n217) );
  OR2_X1 U212 ( .A1(n215), .A2(n214), .ZN(n168) );
  MUX2_X1 U213 ( .A(n340), .B(n168), .S(en), .Z(n362) );
  FA_X1 U214 ( .A(n171), .B(n170), .CI(n169), .CO(n196), .S(n229) );
  OR2_X1 U215 ( .A1(n174), .A2(n175), .ZN(n173) );
  NAND2_X1 U216 ( .A1(n175), .A2(n25), .ZN(n176) );
  OR2_X1 U217 ( .A1(n229), .A2(n228), .ZN(n178) );
  MUX2_X1 U218 ( .A(n341), .B(n178), .S(n334), .Z(n364) );
  FA_X1 U219 ( .A(n181), .B(n180), .CI(n179), .CO(n192), .S(n197) );
  AOI21_X1 U220 ( .B1(n184), .B2(n7), .A(n182), .ZN(n185) );
  INV_X1 U221 ( .A(n185), .ZN(n188) );
  NOR2_X1 U222 ( .A1(n33), .A2(n186), .ZN(n187) );
  XOR2_X1 U223 ( .A(n188), .B(n187), .Z(n189) );
  XOR2_X1 U224 ( .A(n190), .B(n189), .Z(n191) );
  OR2_X1 U225 ( .A1(n192), .A2(n191), .ZN(n194) );
  NAND2_X1 U226 ( .A1(n192), .A2(n191), .ZN(n193) );
  NAND2_X1 U227 ( .A1(n194), .A2(n193), .ZN(n195) );
  MUX2_X1 U228 ( .A(n342), .B(n195), .S(n334), .Z(n366) );
  NAND2_X1 U229 ( .A1(n197), .A2(n196), .ZN(n198) );
  MUX2_X1 U230 ( .A(n343), .B(n198), .S(en), .Z(n368) );
  NAND2_X1 U231 ( .A1(n200), .A2(n199), .ZN(n201) );
  MUX2_X1 U232 ( .A(n344), .B(n201), .S(en), .Z(n370) );
  FA_X1 U233 ( .A(n209), .B(n208), .CI(n207), .CO(n211), .S(n215) );
  NOR2_X1 U234 ( .A1(n212), .A2(n211), .ZN(n210) );
  MUX2_X1 U235 ( .A(n348), .B(n210), .S(en), .Z(n378) );
  NAND2_X1 U236 ( .A1(n212), .A2(n211), .ZN(n213) );
  MUX2_X1 U237 ( .A(n349), .B(n213), .S(en), .Z(n380) );
  NAND2_X1 U238 ( .A1(n215), .A2(n214), .ZN(n216) );
  MUX2_X1 U239 ( .A(n350), .B(n216), .S(n265), .Z(n382) );
  FA_X1 U240 ( .A(n219), .B(n218), .CI(n217), .CO(n214), .S(n226) );
  XNOR2_X1 U241 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n239) );
  OAI22_X1 U242 ( .A1(n67), .A2(n239), .B1(n248), .B2(n220), .ZN(n236) );
  XNOR2_X1 U243 ( .A(n559), .B(\mult_x_1/n284 ), .ZN(n237) );
  OAI22_X1 U244 ( .A1(n253), .A2(n237), .B1(n221), .B2(n31), .ZN(n235) );
  HA_X1 U245 ( .A(n223), .B(n222), .CO(n219), .S(n234) );
  NOR2_X1 U246 ( .A1(n226), .A2(n225), .ZN(n224) );
  MUX2_X1 U247 ( .A(n351), .B(n224), .S(n265), .Z(n384) );
  NAND2_X1 U248 ( .A1(n226), .A2(n225), .ZN(n227) );
  MUX2_X1 U249 ( .A(n352), .B(n227), .S(n265), .Z(n386) );
  NAND2_X1 U250 ( .A1(n229), .A2(n228), .ZN(n230) );
  MUX2_X1 U251 ( .A(n355), .B(n230), .S(n265), .Z(n392) );
  NOR2_X1 U252 ( .A1(n232), .A2(n231), .ZN(n233) );
  MUX2_X1 U253 ( .A(n356), .B(n233), .S(n265), .Z(n394) );
  FA_X1 U254 ( .A(n236), .B(n235), .CI(n234), .CO(n225), .S(n263) );
  XNOR2_X1 U255 ( .A(n559), .B(\mult_x_1/n285 ), .ZN(n245) );
  OAI22_X1 U256 ( .A1(n253), .A2(n245), .B1(n237), .B2(n31), .ZN(n242) );
  AND2_X1 U257 ( .A1(n21), .A2(\mult_x_1/n288 ), .ZN(n241) );
  XNOR2_X1 U258 ( .A(n560), .B(\mult_x_1/n287 ), .ZN(n243) );
  OAI22_X1 U259 ( .A1(n67), .A2(n243), .B1(n248), .B2(n239), .ZN(n240) );
  OR2_X1 U260 ( .A1(n263), .A2(n262), .ZN(n290) );
  FA_X1 U261 ( .A(n242), .B(n241), .CI(n240), .CO(n262), .S(n261) );
  XNOR2_X1 U262 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n244) );
  OAI22_X1 U263 ( .A1(n67), .A2(n244), .B1(n248), .B2(n243), .ZN(n247) );
  XNOR2_X1 U264 ( .A(n559), .B(\mult_x_1/n286 ), .ZN(n250) );
  OAI22_X1 U265 ( .A1(n253), .A2(n250), .B1(n245), .B2(n31), .ZN(n246) );
  NOR2_X1 U266 ( .A1(n261), .A2(n260), .ZN(n283) );
  HA_X1 U267 ( .A(n247), .B(n246), .CO(n260), .S(n258) );
  OR2_X1 U268 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n249) );
  OAI22_X1 U269 ( .A1(n67), .A2(n32), .B1(n249), .B2(n248), .ZN(n257) );
  OR2_X1 U270 ( .A1(n258), .A2(n257), .ZN(n279) );
  XNOR2_X1 U271 ( .A(n559), .B(\mult_x_1/n287 ), .ZN(n252) );
  OAI22_X1 U272 ( .A1(n253), .A2(n252), .B1(n250), .B2(n31), .ZN(n256) );
  AND2_X1 U273 ( .A1(\mult_x_1/n288 ), .A2(n251), .ZN(n255) );
  NOR2_X1 U274 ( .A1(n256), .A2(n255), .ZN(n272) );
  OAI22_X1 U275 ( .A1(n253), .A2(\mult_x_1/n288 ), .B1(n252), .B2(n31), .ZN(
        n269) );
  OR2_X1 U276 ( .A1(\mult_x_1/n288 ), .A2(n45), .ZN(n254) );
  NAND2_X1 U277 ( .A1(n254), .A2(n253), .ZN(n268) );
  NAND2_X1 U278 ( .A1(n269), .A2(n268), .ZN(n275) );
  NAND2_X1 U279 ( .A1(n256), .A2(n255), .ZN(n273) );
  OAI21_X1 U280 ( .B1(n272), .B2(n275), .A(n273), .ZN(n280) );
  NAND2_X1 U281 ( .A1(n258), .A2(n257), .ZN(n278) );
  INV_X1 U282 ( .A(n278), .ZN(n259) );
  AOI21_X1 U283 ( .B1(n279), .B2(n280), .A(n259), .ZN(n286) );
  NAND2_X1 U284 ( .A1(n261), .A2(n260), .ZN(n284) );
  OAI21_X1 U285 ( .B1(n283), .B2(n286), .A(n284), .ZN(n291) );
  NAND2_X1 U286 ( .A1(n263), .A2(n262), .ZN(n289) );
  INV_X1 U287 ( .A(n289), .ZN(n264) );
  AOI21_X1 U288 ( .B1(n290), .B2(n291), .A(n264), .ZN(n266) );
  MUX2_X1 U289 ( .A(n357), .B(n266), .S(n265), .Z(n396) );
  BUF_X4 U290 ( .A(en), .Z(n334) );
  MUX2_X1 U291 ( .A(product[0]), .B(n522), .S(n334), .Z(n412) );
  MUX2_X1 U292 ( .A(n522), .B(n523), .S(n334), .Z(n414) );
  AND2_X1 U293 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n267) );
  MUX2_X1 U294 ( .A(n523), .B(n267), .S(n334), .Z(n416) );
  MUX2_X1 U295 ( .A(product[1]), .B(n525), .S(n334), .Z(n418) );
  MUX2_X1 U296 ( .A(n525), .B(n526), .S(n334), .Z(n420) );
  OR2_X1 U297 ( .A1(n269), .A2(n268), .ZN(n270) );
  AND2_X1 U298 ( .A1(n270), .A2(n275), .ZN(n271) );
  MUX2_X1 U299 ( .A(n526), .B(n271), .S(n334), .Z(n422) );
  MUX2_X1 U300 ( .A(product[2]), .B(n528), .S(n334), .Z(n424) );
  MUX2_X1 U301 ( .A(n528), .B(n529), .S(n334), .Z(n426) );
  INV_X1 U302 ( .A(n272), .ZN(n274) );
  NAND2_X1 U303 ( .A1(n274), .A2(n273), .ZN(n276) );
  XOR2_X1 U304 ( .A(n276), .B(n275), .Z(n277) );
  MUX2_X1 U305 ( .A(n529), .B(n277), .S(n334), .Z(n428) );
  MUX2_X1 U306 ( .A(product[3]), .B(n531), .S(n334), .Z(n430) );
  MUX2_X1 U307 ( .A(n531), .B(n532), .S(n334), .Z(n432) );
  NAND2_X1 U308 ( .A1(n279), .A2(n278), .ZN(n281) );
  XNOR2_X1 U309 ( .A(n281), .B(n280), .ZN(n282) );
  MUX2_X1 U310 ( .A(n532), .B(n282), .S(n334), .Z(n434) );
  MUX2_X1 U311 ( .A(product[4]), .B(n534), .S(n334), .Z(n436) );
  MUX2_X1 U312 ( .A(n534), .B(n535), .S(n334), .Z(n438) );
  INV_X1 U313 ( .A(n283), .ZN(n285) );
  NAND2_X1 U314 ( .A1(n285), .A2(n284), .ZN(n287) );
  XOR2_X1 U315 ( .A(n287), .B(n286), .Z(n288) );
  MUX2_X1 U316 ( .A(n535), .B(n288), .S(n334), .Z(n440) );
  MUX2_X1 U317 ( .A(product[5]), .B(n537), .S(n334), .Z(n442) );
  MUX2_X1 U318 ( .A(n537), .B(n538), .S(n334), .Z(n444) );
  NAND2_X1 U319 ( .A1(n290), .A2(n289), .ZN(n292) );
  MUX2_X1 U320 ( .A(product[6]), .B(n540), .S(n334), .Z(n448) );
  NAND2_X1 U321 ( .A1(n401), .A2(n352), .ZN(n293) );
  XOR2_X1 U322 ( .A(n293), .B(n357), .Z(n294) );
  MUX2_X1 U323 ( .A(n540), .B(n294), .S(n334), .Z(n450) );
  MUX2_X1 U324 ( .A(product[7]), .B(n542), .S(n334), .Z(n452) );
  OAI21_X1 U325 ( .B1(n351), .B2(n357), .A(n352), .ZN(n297) );
  NAND2_X1 U326 ( .A1(n340), .A2(n350), .ZN(n295) );
  XNOR2_X1 U327 ( .A(n297), .B(n295), .ZN(n296) );
  MUX2_X1 U328 ( .A(n542), .B(n296), .S(n334), .Z(n454) );
  MUX2_X1 U329 ( .A(product[8]), .B(n544), .S(n334), .Z(n456) );
  AOI21_X1 U330 ( .B1(n297), .B2(n340), .A(n402), .ZN(n300) );
  NAND2_X1 U331 ( .A1(n403), .A2(n349), .ZN(n298) );
  XOR2_X1 U332 ( .A(n300), .B(n298), .Z(n299) );
  MUX2_X1 U333 ( .A(n544), .B(n299), .S(n334), .Z(n458) );
  MUX2_X1 U334 ( .A(product[9]), .B(n546), .S(n334), .Z(n460) );
  OAI21_X1 U335 ( .B1(n300), .B2(n348), .A(n349), .ZN(n308) );
  INV_X1 U336 ( .A(n308), .ZN(n303) );
  NAND2_X1 U337 ( .A1(n405), .A2(n347), .ZN(n301) );
  XOR2_X1 U338 ( .A(n303), .B(n301), .Z(n302) );
  MUX2_X1 U339 ( .A(n546), .B(n302), .S(n334), .Z(n462) );
  MUX2_X1 U340 ( .A(product[10]), .B(n548), .S(n334), .Z(n464) );
  OAI21_X1 U341 ( .B1(n303), .B2(n356), .A(n347), .ZN(n305) );
  NAND2_X1 U342 ( .A1(n336), .A2(n354), .ZN(n304) );
  XNOR2_X1 U343 ( .A(n305), .B(n304), .ZN(n306) );
  MUX2_X1 U344 ( .A(n548), .B(n306), .S(n334), .Z(n466) );
  MUX2_X1 U345 ( .A(product[11]), .B(n550), .S(n334), .Z(n468) );
  NOR2_X1 U346 ( .A1(n353), .A2(n356), .ZN(n309) );
  OAI21_X1 U347 ( .B1(n353), .B2(n347), .A(n354), .ZN(n307) );
  AOI21_X1 U348 ( .B1(n309), .B2(n308), .A(n307), .ZN(n331) );
  NAND2_X1 U349 ( .A1(n404), .A2(n346), .ZN(n310) );
  XOR2_X1 U350 ( .A(n331), .B(n310), .Z(n311) );
  MUX2_X1 U351 ( .A(n550), .B(n311), .S(n334), .Z(n470) );
  MUX2_X1 U352 ( .A(product[12]), .B(n552), .S(n334), .Z(n472) );
  OAI21_X1 U353 ( .B1(n331), .B2(n345), .A(n346), .ZN(n313) );
  NAND2_X1 U354 ( .A1(n339), .A2(n344), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n314) );
  MUX2_X1 U356 ( .A(n552), .B(n314), .S(n334), .Z(n474) );
  MUX2_X1 U357 ( .A(product[13]), .B(n554), .S(n334), .Z(n476) );
  NAND2_X1 U358 ( .A1(n404), .A2(n339), .ZN(n316) );
  AOI21_X1 U359 ( .B1(n400), .B2(n339), .A(n406), .ZN(n315) );
  OAI21_X1 U360 ( .B1(n331), .B2(n316), .A(n315), .ZN(n318) );
  NAND2_X1 U361 ( .A1(n341), .A2(n355), .ZN(n317) );
  XNOR2_X1 U362 ( .A(n318), .B(n317), .ZN(n319) );
  MUX2_X1 U363 ( .A(n554), .B(n319), .S(n334), .Z(n478) );
  MUX2_X1 U364 ( .A(product[14]), .B(n556), .S(n334), .Z(n480) );
  NAND2_X1 U365 ( .A1(n339), .A2(n341), .ZN(n321) );
  NOR2_X1 U366 ( .A1(n345), .A2(n321), .ZN(n327) );
  INV_X1 U367 ( .A(n327), .ZN(n323) );
  AOI21_X1 U368 ( .B1(n406), .B2(n341), .A(n399), .ZN(n320) );
  OAI21_X1 U369 ( .B1(n321), .B2(n346), .A(n320), .ZN(n328) );
  INV_X1 U370 ( .A(n328), .ZN(n322) );
  OAI21_X1 U371 ( .B1(n331), .B2(n323), .A(n322), .ZN(n325) );
  NAND2_X1 U372 ( .A1(n338), .A2(n343), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U374 ( .A(n556), .B(n326), .S(n334), .Z(n482) );
  MUX2_X1 U375 ( .A(product[15]), .B(n558), .S(n334), .Z(n484) );
  NAND2_X1 U376 ( .A1(n327), .A2(n338), .ZN(n330) );
  AOI21_X1 U377 ( .B1(n328), .B2(n338), .A(n398), .ZN(n329) );
  OAI21_X1 U378 ( .B1(n331), .B2(n330), .A(n329), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n332), .B(n342), .ZN(n333) );
  MUX2_X1 U380 ( .A(n558), .B(n333), .S(n334), .Z(n486) );
  MUX2_X1 U381 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n334), .Z(n488) );
  MUX2_X1 U382 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n334), .Z(n490) );
  MUX2_X1 U383 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n334), .Z(n492) );
  MUX2_X1 U384 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n334), .Z(n494) );
  MUX2_X1 U385 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n334), .Z(n496) );
  MUX2_X1 U386 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n334), .Z(n498) );
  MUX2_X1 U387 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n334), .Z(n500) );
  MUX2_X1 U388 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n334), .Z(n502) );
  MUX2_X1 U389 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n334), .Z(n504) );
  MUX2_X1 U390 ( .A(n559), .B(A_extended[1]), .S(n334), .Z(n506) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n334), .Z(n508) );
  MUX2_X1 U392 ( .A(n22), .B(A_extended[3]), .S(n334), .Z(n510) );
  MUX2_X1 U393 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n334), .Z(n512) );
  MUX2_X1 U394 ( .A(n29), .B(A_extended[5]), .S(n334), .Z(n514) );
  MUX2_X1 U395 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n334), .Z(n516) );
  MUX2_X1 U396 ( .A(n28), .B(A_extended[7]), .S(n334), .Z(n518) );
  OR2_X1 U397 ( .A1(n334), .A2(n562), .ZN(n520) );
endmodule


module conv_128_32_DW_mult_pipe_J1_16 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n352, n354, n356, n358, n360, n362, n364, n366, n368,
         n370, n372, n374, n376, n378, n380, n382, n384, n386, n388, n390,
         n392, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n405, n407, n409, n411, n413, n415, n417, n419, n421, n423, n425,
         n427, n429, n431, n433, n435, n437, n439, n441, n443, n445, n447,
         n449, n451, n453, n455, n457, n459, n461, n463, n465, n467, n469,
         n471, n473, n475, n477, n479, n481, n483, n485, n487, n489, n491,
         n493, n495, n497, n499, n501, n503, n505, n507, n509, n511, n513,
         n514, n516, n517, n519, n520, n522, n523, n525, n526, n528, n530,
         n532, n534, n536, n538, n540, n542, n544, n546, n548, n549, n550,
         n551;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n403), .SE(n511), .CK(clk), .Q(n550), 
        .QN(n326) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n403), .SE(n507), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n27) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n403), .SE(n503), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n28) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n403), .SE(n499), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n23) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n403), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n24) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n403), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n403), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n401), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n402), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n401), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n403), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n401), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n401), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n401), .SE(n477), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n401), .SE(n475), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n401), .SE(n473), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n401), .SE(n471), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n401), .SE(n469), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n402), .SE(n467), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n403), .SE(n465), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n401), .SE(n463), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n401), .SE(n461), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n401), .SE(n459), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n401), .SE(n457), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n401), .SE(n455), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n401), .SE(n453), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n401), .SE(n451), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n401), .SE(n449), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n402), .SE(n447), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n402), .SE(n445), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n402), .SE(n443), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n402), .SE(n441), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n402), .SE(n439), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n402), .SE(n437), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n402), .SE(n435), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n402), .SE(n433), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n402), .SE(n431), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n402), .SE(n429), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n402), .SE(n427), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n401), .SE(n425), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n401), .SE(n423), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n401), .SE(n421), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n401), .SE(n419), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n401), .SE(n417), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n401), .SE(n415), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n401), .SE(n413), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n401), .SE(n411), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n401), .SE(n409), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n401), .SE(n407), .CK(clk), .Q(n513)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n401), .SE(n405), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n551), .SE(n392), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2_IP  ( .D(1'b1), .SI(n551), .SE(n390), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n551), .SE(n388), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n551), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n551), .SE(n384), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n551), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n551), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n551), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n342), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n551), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n341), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n551), .SE(n374), .CK(
        clk), .Q(n327), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n551), .SE(n372), .CK(
        clk), .Q(n399), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n551), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n551), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n551), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n336), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n551), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n335), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n551), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n551), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n333), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n551), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n332), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n551), .SE(n356), .CK(
        clk), .QN(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n551), .SE(n354), .CK(
        clk), .QN(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n551), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n551), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n328) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n403), .SE(n505), .CK(clk), .Q(n549), 
        .QN(n26) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n403), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n25) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n403), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n29) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n403), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n325) );
  INV_X1 U2 ( .A(n26), .ZN(n22) );
  NAND2_X1 U3 ( .A1(n8), .A2(n5), .ZN(n378) );
  INV_X1 U4 ( .A(n6), .ZN(n5) );
  NOR2_X1 U5 ( .A1(n324), .A2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n342), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n9), .A2(n324), .ZN(n8) );
  NAND2_X1 U8 ( .A1(n206), .A2(n205), .ZN(n9) );
  CLKBUF_X2 U9 ( .A(n123), .Z(n15) );
  CLKBUF_X2 U10 ( .A(n123), .Z(n14) );
  BUF_X1 U11 ( .A(en), .Z(n123) );
  BUF_X1 U12 ( .A(n401), .Z(n403) );
  INV_X2 U13 ( .A(n551), .ZN(n401) );
  NAND2_X1 U14 ( .A1(n48), .A2(n49), .ZN(n66) );
  NAND2_X1 U15 ( .A1(n11), .A2(n10), .ZN(n109) );
  NAND2_X1 U16 ( .A1(n245), .A2(n12), .ZN(n11) );
  XNOR2_X1 U17 ( .A(n245), .B(n13), .ZN(n248) );
  XNOR2_X1 U18 ( .A(n247), .B(n246), .ZN(n13) );
  NAND2_X1 U19 ( .A1(n247), .A2(n246), .ZN(n10) );
  OR2_X1 U20 ( .A1(n247), .A2(n246), .ZN(n12) );
  BUF_X1 U21 ( .A(n401), .Z(n402) );
  INV_X1 U22 ( .A(rst_n), .ZN(n551) );
  OAI22_X1 U23 ( .A1(n146), .A2(n101), .B1(n145), .B2(n325), .ZN(n126) );
  BUF_X1 U24 ( .A(n49), .Z(n16) );
  INV_X1 U25 ( .A(n32), .ZN(n196) );
  OR2_X1 U26 ( .A1(n31), .A2(n32), .ZN(n136) );
  AND2_X2 U27 ( .A1(n550), .A2(\mult_x_1/n281 ), .ZN(n115) );
  OAI21_X1 U28 ( .B1(n46), .B2(n44), .A(n43), .ZN(n38) );
  NAND2_X1 U29 ( .A1(n46), .A2(n44), .ZN(n37) );
  NOR2_X2 U30 ( .A1(n325), .A2(n326), .ZN(n148) );
  OR2_X1 U31 ( .A1(n76), .A2(n75), .ZN(n56) );
  NAND2_X1 U32 ( .A1(n76), .A2(n75), .ZN(n57) );
  NAND2_X1 U33 ( .A1(n38), .A2(n37), .ZN(n122) );
  XNOR2_X1 U34 ( .A(n78), .B(n77), .ZN(n235) );
  XNOR2_X1 U35 ( .A(n76), .B(n75), .ZN(n77) );
  NAND2_X1 U36 ( .A1(n61), .A2(n60), .ZN(n352) );
  NAND2_X1 U37 ( .A1(n59), .A2(n329), .ZN(n60) );
  OAI21_X1 U38 ( .B1(n203), .B2(n202), .A(n14), .ZN(n61) );
  NAND2_X1 U39 ( .A1(n80), .A2(n79), .ZN(n380) );
  NAND2_X1 U40 ( .A1(n59), .A2(n343), .ZN(n79) );
  OAI21_X1 U41 ( .B1(n206), .B2(n205), .A(n15), .ZN(n80) );
  NAND2_X1 U42 ( .A1(n243), .A2(n242), .ZN(n244) );
  NAND2_X1 U43 ( .A1(n241), .A2(n240), .ZN(n242) );
  NAND2_X1 U44 ( .A1(n239), .A2(n30), .ZN(n243) );
  OAI22_X1 U45 ( .A1(n66), .A2(n67), .B1(n50), .B2(n16), .ZN(n17) );
  NAND2_X1 U46 ( .A1(n33), .A2(n34), .ZN(n18) );
  INV_X1 U47 ( .A(n325), .ZN(n19) );
  NAND2_X1 U48 ( .A1(n33), .A2(n34), .ZN(n145) );
  OAI22_X1 U49 ( .A1(n136), .A2(n99), .B1(n196), .B2(n65), .ZN(n20) );
  INV_X1 U50 ( .A(n25), .ZN(n21) );
  XNOR2_X1 U51 ( .A(n29), .B(n23), .ZN(n49) );
  INV_X1 U52 ( .A(n123), .ZN(n59) );
  OR2_X1 U53 ( .A1(n241), .A2(n240), .ZN(n30) );
  XNOR2_X1 U54 ( .A(\mult_x_1/a[4] ), .B(n549), .ZN(n31) );
  XNOR2_X1 U55 ( .A(\mult_x_1/n312 ), .B(n28), .ZN(n32) );
  XNOR2_X1 U56 ( .A(n22), .B(\mult_x_1/n281 ), .ZN(n53) );
  XNOR2_X1 U57 ( .A(n115), .B(n22), .ZN(n41) );
  OAI22_X1 U58 ( .A1(n136), .A2(n53), .B1(n41), .B2(n196), .ZN(n117) );
  INV_X1 U59 ( .A(n117), .ZN(n46) );
  XNOR2_X1 U60 ( .A(\mult_x_1/n310 ), .B(n27), .ZN(n33) );
  XNOR2_X1 U61 ( .A(n549), .B(\mult_x_1/a[6] ), .ZN(n34) );
  XNOR2_X1 U62 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n47) );
  INV_X1 U63 ( .A(n34), .ZN(n35) );
  INV_X2 U64 ( .A(n35), .ZN(n146) );
  XNOR2_X1 U65 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n40) );
  OAI22_X1 U66 ( .A1(n18), .A2(n47), .B1(n146), .B2(n40), .ZN(n44) );
  XNOR2_X1 U67 ( .A(n148), .B(\mult_x_1/n284 ), .ZN(n36) );
  NAND2_X1 U68 ( .A1(n326), .A2(\mult_x_1/n310 ), .ZN(n90) );
  NOR2_X1 U69 ( .A1(n36), .A2(n90), .ZN(n43) );
  XNOR2_X1 U70 ( .A(n148), .B(\mult_x_1/n283 ), .ZN(n39) );
  NOR2_X1 U71 ( .A1(n39), .A2(n90), .ZN(n121) );
  XNOR2_X1 U72 ( .A(n19), .B(\mult_x_1/n281 ), .ZN(n116) );
  OAI22_X1 U73 ( .A1(n18), .A2(n40), .B1(n146), .B2(n116), .ZN(n119) );
  AOI21_X1 U74 ( .B1(n196), .B2(n136), .A(n41), .ZN(n42) );
  INV_X1 U75 ( .A(n42), .ZN(n118) );
  XNOR2_X1 U76 ( .A(n44), .B(n43), .ZN(n45) );
  XNOR2_X1 U77 ( .A(n46), .B(n45), .ZN(n64) );
  XNOR2_X1 U78 ( .A(n19), .B(\mult_x_1/n284 ), .ZN(n52) );
  OAI22_X1 U79 ( .A1(n18), .A2(n52), .B1(n146), .B2(n47), .ZN(n74) );
  XOR2_X1 U80 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n48) );
  XNOR2_X1 U81 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n67) );
  XNOR2_X1 U82 ( .A(n115), .B(\mult_x_1/n312 ), .ZN(n50) );
  OAI22_X1 U83 ( .A1(n66), .A2(n67), .B1(n50), .B2(n16), .ZN(n73) );
  CLKBUF_X2 U84 ( .A(n66), .Z(n217) );
  AOI21_X1 U85 ( .B1(n16), .B2(n217), .A(n50), .ZN(n51) );
  INV_X1 U86 ( .A(n51), .ZN(n72) );
  XNOR2_X1 U87 ( .A(n19), .B(\mult_x_1/n285 ), .ZN(n71) );
  OAI22_X1 U88 ( .A1(n18), .A2(n71), .B1(n146), .B2(n52), .ZN(n94) );
  XNOR2_X1 U89 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n65) );
  XNOR2_X1 U90 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n54) );
  OAI22_X1 U91 ( .A1(n136), .A2(n65), .B1(n196), .B2(n54), .ZN(n93) );
  INV_X1 U92 ( .A(n73), .ZN(n92) );
  OAI22_X1 U93 ( .A1(n136), .A2(n54), .B1(n196), .B2(n53), .ZN(n76) );
  XNOR2_X1 U94 ( .A(n148), .B(\mult_x_1/n285 ), .ZN(n55) );
  NOR2_X1 U95 ( .A1(n55), .A2(n90), .ZN(n75) );
  NAND2_X1 U96 ( .A1(n78), .A2(n56), .ZN(n58) );
  NAND2_X1 U97 ( .A1(n58), .A2(n57), .ZN(n62) );
  FA_X1 U98 ( .A(n64), .B(n63), .CI(n62), .CO(n202), .S(n206) );
  XNOR2_X1 U99 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n99) );
  OAI22_X1 U100 ( .A1(n136), .A2(n99), .B1(n196), .B2(n65), .ZN(n85) );
  XNOR2_X1 U101 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n100) );
  OAI22_X1 U102 ( .A1(n66), .A2(n100), .B1(n16), .B2(n67), .ZN(n84) );
  OR2_X1 U103 ( .A1(n85), .A2(n84), .ZN(n83) );
  XNOR2_X1 U104 ( .A(n148), .B(\mult_x_1/n286 ), .ZN(n68) );
  NOR2_X1 U105 ( .A1(n68), .A2(n90), .ZN(n82) );
  NAND2_X1 U106 ( .A1(\mult_x_1/n313 ), .A2(n24), .ZN(n221) );
  XNOR2_X1 U107 ( .A(n115), .B(\mult_x_1/n313 ), .ZN(n89) );
  AOI21_X1 U108 ( .B1(n221), .B2(n24), .A(n89), .ZN(n69) );
  INV_X1 U109 ( .A(n69), .ZN(n98) );
  XNOR2_X1 U110 ( .A(n148), .B(\mult_x_1/n287 ), .ZN(n70) );
  NOR2_X1 U111 ( .A1(n70), .A2(n90), .ZN(n97) );
  XNOR2_X1 U112 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n88) );
  OAI22_X1 U113 ( .A1(n18), .A2(n88), .B1(n146), .B2(n71), .ZN(n96) );
  FA_X1 U114 ( .A(n74), .B(n17), .CI(n72), .CO(n63), .S(n236) );
  FA_X1 U115 ( .A(n83), .B(n82), .CI(n81), .CO(n237), .S(n239) );
  XNOR2_X1 U116 ( .A(n20), .B(n84), .ZN(n106) );
  INV_X1 U117 ( .A(n148), .ZN(n86) );
  OR2_X1 U118 ( .A1(\mult_x_1/n288 ), .A2(n86), .ZN(n87) );
  NOR2_X1 U119 ( .A1(n87), .A2(n90), .ZN(n105) );
  XNOR2_X1 U120 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n102) );
  OAI22_X1 U121 ( .A1(n145), .A2(n102), .B1(n146), .B2(n88), .ZN(n164) );
  XNOR2_X1 U122 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n128) );
  OAI22_X1 U123 ( .A1(n221), .A2(n128), .B1(n89), .B2(n24), .ZN(n163) );
  INV_X1 U124 ( .A(n90), .ZN(n91) );
  AND2_X1 U125 ( .A1(\mult_x_1/n288 ), .A2(n91), .ZN(n162) );
  FA_X1 U126 ( .A(n94), .B(n92), .CI(n93), .CO(n78), .S(n240) );
  XNOR2_X1 U127 ( .A(n241), .B(n240), .ZN(n95) );
  XNOR2_X1 U128 ( .A(n239), .B(n95), .ZN(n110) );
  FA_X1 U129 ( .A(n98), .B(n97), .CI(n96), .CO(n81), .S(n247) );
  XNOR2_X1 U130 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n127) );
  OAI22_X1 U131 ( .A1(n136), .A2(n127), .B1(n196), .B2(n99), .ZN(n170) );
  XNOR2_X1 U132 ( .A(n21), .B(\mult_x_1/n283 ), .ZN(n130) );
  OAI22_X1 U133 ( .A1(n217), .A2(n130), .B1(n16), .B2(n100), .ZN(n169) );
  OR2_X1 U134 ( .A1(\mult_x_1/n288 ), .A2(n325), .ZN(n101) );
  XNOR2_X1 U135 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n103) );
  OAI22_X1 U136 ( .A1(n145), .A2(n103), .B1(n146), .B2(n102), .ZN(n125) );
  FA_X1 U137 ( .A(n106), .B(n105), .CI(n104), .CO(n241), .S(n245) );
  INV_X1 U138 ( .A(n109), .ZN(n107) );
  NAND2_X1 U139 ( .A1(n107), .A2(n15), .ZN(n108) );
  OAI22_X1 U140 ( .A1(n110), .A2(n108), .B1(n324), .B2(n399), .ZN(n372) );
  NAND2_X1 U141 ( .A1(n110), .A2(n109), .ZN(n111) );
  NAND2_X1 U142 ( .A1(n111), .A2(n324), .ZN(n113) );
  OR2_X1 U143 ( .A1(n324), .A2(n327), .ZN(n112) );
  NAND2_X1 U144 ( .A1(n113), .A2(n112), .ZN(n374) );
  XNOR2_X1 U167 ( .A(n148), .B(\mult_x_1/n282 ), .ZN(n114) );
  NOR2_X1 U168 ( .A1(n114), .A2(n90), .ZN(n143) );
  XNOR2_X1 U169 ( .A(n115), .B(n19), .ZN(n144) );
  OAI22_X1 U170 ( .A1(n18), .A2(n116), .B1(n144), .B2(n146), .ZN(n153) );
  INV_X1 U171 ( .A(n153), .ZN(n142) );
  FA_X1 U172 ( .A(n119), .B(n118), .CI(n117), .CO(n141), .S(n120) );
  FA_X1 U173 ( .A(n122), .B(n121), .CI(n120), .CO(n159), .S(n203) );
  OR2_X1 U174 ( .A1(n160), .A2(n159), .ZN(n124) );
  MUX2_X1 U175 ( .A(n328), .B(n124), .S(n324), .Z(n350) );
  XNOR2_X1 U176 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n185) );
  XNOR2_X1 U177 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n129) );
  OAI22_X1 U178 ( .A1(n221), .A2(n185), .B1(n129), .B2(n24), .ZN(n139) );
  AND2_X1 U179 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n138) );
  XNOR2_X1 U180 ( .A(n21), .B(\mult_x_1/n285 ), .ZN(n184) );
  XNOR2_X1 U181 ( .A(n21), .B(\mult_x_1/n284 ), .ZN(n131) );
  OAI22_X1 U182 ( .A1(n217), .A2(n184), .B1(n16), .B2(n131), .ZN(n137) );
  HA_X1 U183 ( .A(n126), .B(n125), .CO(n168), .S(n172) );
  XNOR2_X1 U184 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n134) );
  OAI22_X1 U185 ( .A1(n136), .A2(n134), .B1(n196), .B2(n127), .ZN(n167) );
  OAI22_X1 U186 ( .A1(n221), .A2(n129), .B1(n128), .B2(n24), .ZN(n166) );
  OAI22_X1 U187 ( .A1(n217), .A2(n131), .B1(n16), .B2(n130), .ZN(n165) );
  OR2_X1 U188 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n132) );
  OAI22_X1 U189 ( .A1(n136), .A2(n26), .B1(n132), .B2(n196), .ZN(n187) );
  XNOR2_X1 U190 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n133) );
  XNOR2_X1 U191 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n135) );
  OAI22_X1 U192 ( .A1(n136), .A2(n133), .B1(n196), .B2(n135), .ZN(n186) );
  OAI22_X1 U193 ( .A1(n136), .A2(n135), .B1(n196), .B2(n134), .ZN(n182) );
  FA_X1 U194 ( .A(n139), .B(n138), .CI(n137), .CO(n173), .S(n181) );
  OR2_X1 U195 ( .A1(n179), .A2(n178), .ZN(n140) );
  MUX2_X1 U196 ( .A(n330), .B(n140), .S(n324), .Z(n354) );
  FA_X1 U197 ( .A(n143), .B(n142), .CI(n141), .CO(n155), .S(n160) );
  AOI21_X1 U198 ( .B1(n146), .B2(n18), .A(n144), .ZN(n147) );
  INV_X1 U199 ( .A(n147), .ZN(n151) );
  XNOR2_X1 U200 ( .A(n148), .B(\mult_x_1/n281 ), .ZN(n149) );
  NOR2_X1 U201 ( .A1(n149), .A2(n90), .ZN(n150) );
  XOR2_X1 U202 ( .A(n151), .B(n150), .Z(n152) );
  XOR2_X1 U203 ( .A(n153), .B(n152), .Z(n154) );
  OR2_X1 U204 ( .A1(n155), .A2(n154), .ZN(n157) );
  NAND2_X1 U205 ( .A1(n155), .A2(n154), .ZN(n156) );
  NAND2_X1 U206 ( .A1(n157), .A2(n156), .ZN(n158) );
  MUX2_X1 U207 ( .A(n331), .B(n158), .S(n324), .Z(n356) );
  NAND2_X1 U208 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2_X1 U209 ( .A(n332), .B(n161), .S(n15), .Z(n358) );
  FA_X1 U210 ( .A(n163), .B(n164), .CI(n162), .CO(n104), .S(n251) );
  FA_X1 U211 ( .A(n167), .B(n166), .CI(n165), .CO(n250), .S(n171) );
  FA_X1 U212 ( .A(n170), .B(n169), .CI(n168), .CO(n246), .S(n249) );
  FA_X1 U213 ( .A(n173), .B(n172), .CI(n171), .CO(n175), .S(n179) );
  NOR2_X1 U214 ( .A1(n176), .A2(n175), .ZN(n174) );
  MUX2_X1 U215 ( .A(n333), .B(n174), .S(n324), .Z(n360) );
  NAND2_X1 U216 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U217 ( .A(n334), .B(n177), .S(en), .Z(n362) );
  NAND2_X1 U218 ( .A1(n179), .A2(n178), .ZN(n180) );
  MUX2_X1 U219 ( .A(n335), .B(n180), .S(n14), .Z(n364) );
  FA_X1 U220 ( .A(n183), .B(n182), .CI(n181), .CO(n178), .S(n190) );
  XNOR2_X1 U221 ( .A(n21), .B(\mult_x_1/n286 ), .ZN(n198) );
  OAI22_X1 U222 ( .A1(n217), .A2(n198), .B1(n16), .B2(n184), .ZN(n194) );
  XNOR2_X1 U223 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n195) );
  OAI22_X1 U224 ( .A1(n221), .A2(n195), .B1(n185), .B2(n24), .ZN(n193) );
  HA_X1 U225 ( .A(n187), .B(n186), .CO(n183), .S(n192) );
  NOR2_X1 U226 ( .A1(n190), .A2(n189), .ZN(n188) );
  MUX2_X1 U227 ( .A(n336), .B(n188), .S(n324), .Z(n366) );
  NAND2_X1 U228 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U229 ( .A(n337), .B(n191), .S(n324), .Z(n368) );
  FA_X1 U230 ( .A(n194), .B(n193), .CI(n192), .CO(n189), .S(n200) );
  XNOR2_X1 U231 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n213) );
  OAI22_X1 U232 ( .A1(n221), .A2(n213), .B1(n195), .B2(n24), .ZN(n210) );
  INV_X1 U233 ( .A(n196), .ZN(n197) );
  AND2_X1 U234 ( .A1(\mult_x_1/n288 ), .A2(n197), .ZN(n209) );
  XNOR2_X1 U235 ( .A(n21), .B(\mult_x_1/n287 ), .ZN(n211) );
  OAI22_X1 U236 ( .A1(n217), .A2(n211), .B1(n16), .B2(n198), .ZN(n208) );
  OR2_X1 U237 ( .A1(n200), .A2(n199), .ZN(n232) );
  NAND2_X1 U238 ( .A1(n200), .A2(n199), .ZN(n230) );
  NAND2_X1 U239 ( .A1(n232), .A2(n230), .ZN(n201) );
  MUX2_X1 U240 ( .A(n338), .B(n201), .S(n324), .Z(n370) );
  NAND2_X1 U241 ( .A1(n203), .A2(n202), .ZN(n204) );
  MUX2_X1 U242 ( .A(n341), .B(n204), .S(n15), .Z(n376) );
  FA_X1 U243 ( .A(n210), .B(n209), .CI(n208), .CO(n199), .S(n229) );
  XNOR2_X1 U244 ( .A(n21), .B(\mult_x_1/n288 ), .ZN(n212) );
  OAI22_X1 U245 ( .A1(n217), .A2(n212), .B1(n16), .B2(n211), .ZN(n215) );
  XNOR2_X1 U246 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n218) );
  OAI22_X1 U247 ( .A1(n221), .A2(n218), .B1(n213), .B2(n24), .ZN(n214) );
  NOR2_X1 U248 ( .A1(n229), .A2(n228), .ZN(n269) );
  HA_X1 U249 ( .A(n215), .B(n214), .CO(n228), .S(n226) );
  OR2_X1 U250 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n216) );
  OAI22_X1 U251 ( .A1(n217), .A2(n25), .B1(n216), .B2(n16), .ZN(n225) );
  OR2_X1 U252 ( .A1(n226), .A2(n225), .ZN(n265) );
  XNOR2_X1 U253 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n220) );
  OAI22_X1 U254 ( .A1(n221), .A2(n220), .B1(n218), .B2(n24), .ZN(n224) );
  INV_X1 U255 ( .A(n16), .ZN(n219) );
  AND2_X1 U256 ( .A1(\mult_x_1/n288 ), .A2(n219), .ZN(n223) );
  NOR2_X1 U257 ( .A1(n224), .A2(n223), .ZN(n258) );
  OAI22_X1 U258 ( .A1(n221), .A2(\mult_x_1/n288 ), .B1(n220), .B2(n24), .ZN(
        n255) );
  OR2_X1 U259 ( .A1(\mult_x_1/n288 ), .A2(n29), .ZN(n222) );
  NAND2_X1 U260 ( .A1(n222), .A2(n221), .ZN(n254) );
  NAND2_X1 U261 ( .A1(n255), .A2(n254), .ZN(n261) );
  NAND2_X1 U262 ( .A1(n224), .A2(n223), .ZN(n259) );
  OAI21_X1 U263 ( .B1(n258), .B2(n261), .A(n259), .ZN(n266) );
  NAND2_X1 U264 ( .A1(n226), .A2(n225), .ZN(n264) );
  INV_X1 U265 ( .A(n264), .ZN(n227) );
  AOI21_X1 U266 ( .B1(n265), .B2(n266), .A(n227), .ZN(n272) );
  NAND2_X1 U267 ( .A1(n229), .A2(n228), .ZN(n270) );
  OAI21_X1 U268 ( .B1(n269), .B2(n272), .A(n270), .ZN(n234) );
  INV_X1 U269 ( .A(n230), .ZN(n231) );
  AOI21_X1 U270 ( .B1(n232), .B2(n234), .A(n231), .ZN(n233) );
  MUX2_X1 U271 ( .A(n344), .B(n233), .S(n324), .Z(n382) );
  MUX2_X1 U272 ( .A(n345), .B(n234), .S(n324), .Z(n384) );
  FA_X1 U273 ( .A(n237), .B(n236), .CI(n235), .CO(n205), .S(n238) );
  MUX2_X1 U274 ( .A(n346), .B(n238), .S(n324), .Z(n386) );
  MUX2_X1 U275 ( .A(n347), .B(n244), .S(n324), .Z(n388) );
  MUX2_X1 U276 ( .A(n348), .B(n248), .S(n324), .Z(n390) );
  FA_X1 U277 ( .A(n251), .B(n250), .CI(n249), .CO(n252), .S(n176) );
  MUX2_X1 U278 ( .A(n349), .B(n252), .S(n14), .Z(n392) );
  MUX2_X1 U279 ( .A(product[0]), .B(n513), .S(n324), .Z(n405) );
  MUX2_X1 U280 ( .A(n513), .B(n514), .S(n14), .Z(n407) );
  AND2_X1 U281 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n253) );
  MUX2_X1 U282 ( .A(n514), .B(n253), .S(n15), .Z(n409) );
  MUX2_X1 U283 ( .A(product[1]), .B(n516), .S(n14), .Z(n411) );
  MUX2_X1 U284 ( .A(n516), .B(n517), .S(n15), .Z(n413) );
  OR2_X1 U285 ( .A1(n255), .A2(n254), .ZN(n256) );
  AND2_X1 U286 ( .A1(n256), .A2(n261), .ZN(n257) );
  MUX2_X1 U287 ( .A(n517), .B(n257), .S(n324), .Z(n415) );
  MUX2_X1 U288 ( .A(product[2]), .B(n519), .S(n14), .Z(n417) );
  MUX2_X1 U289 ( .A(n519), .B(n520), .S(n324), .Z(n419) );
  INV_X1 U290 ( .A(n258), .ZN(n260) );
  NAND2_X1 U291 ( .A1(n260), .A2(n259), .ZN(n262) );
  XOR2_X1 U292 ( .A(n262), .B(n261), .Z(n263) );
  MUX2_X1 U293 ( .A(n520), .B(n263), .S(n324), .Z(n421) );
  MUX2_X1 U294 ( .A(product[3]), .B(n522), .S(n15), .Z(n423) );
  MUX2_X1 U295 ( .A(n522), .B(n523), .S(n324), .Z(n425) );
  NAND2_X1 U296 ( .A1(n265), .A2(n264), .ZN(n267) );
  XNOR2_X1 U297 ( .A(n267), .B(n266), .ZN(n268) );
  MUX2_X1 U298 ( .A(n523), .B(n268), .S(n324), .Z(n427) );
  MUX2_X1 U299 ( .A(product[4]), .B(n525), .S(n14), .Z(n429) );
  MUX2_X1 U300 ( .A(n525), .B(n526), .S(n324), .Z(n431) );
  INV_X1 U301 ( .A(n269), .ZN(n271) );
  NAND2_X1 U302 ( .A1(n271), .A2(n270), .ZN(n273) );
  XOR2_X1 U303 ( .A(n273), .B(n272), .Z(n274) );
  MUX2_X1 U304 ( .A(n526), .B(n274), .S(n324), .Z(n433) );
  MUX2_X1 U305 ( .A(product[5]), .B(n528), .S(n15), .Z(n435) );
  XNOR2_X1 U306 ( .A(n338), .B(n345), .ZN(n275) );
  MUX2_X1 U307 ( .A(n528), .B(n275), .S(n324), .Z(n437) );
  MUX2_X1 U308 ( .A(product[6]), .B(n530), .S(n324), .Z(n439) );
  NAND2_X1 U309 ( .A1(n395), .A2(n337), .ZN(n276) );
  XOR2_X1 U310 ( .A(n276), .B(n344), .Z(n277) );
  MUX2_X1 U311 ( .A(n530), .B(n277), .S(n324), .Z(n441) );
  MUX2_X1 U312 ( .A(product[7]), .B(n532), .S(n14), .Z(n443) );
  OAI21_X1 U313 ( .B1(n336), .B2(n344), .A(n337), .ZN(n280) );
  NAND2_X1 U314 ( .A1(n330), .A2(n335), .ZN(n278) );
  XNOR2_X1 U315 ( .A(n280), .B(n278), .ZN(n279) );
  BUF_X8 U316 ( .A(en), .Z(n324) );
  MUX2_X1 U317 ( .A(n532), .B(n279), .S(n324), .Z(n445) );
  MUX2_X1 U318 ( .A(product[8]), .B(n534), .S(n15), .Z(n447) );
  AOI21_X1 U319 ( .B1(n280), .B2(n330), .A(n397), .ZN(n283) );
  NAND2_X1 U320 ( .A1(n398), .A2(n334), .ZN(n281) );
  XOR2_X1 U321 ( .A(n283), .B(n281), .Z(n282) );
  MUX2_X1 U322 ( .A(n534), .B(n282), .S(n324), .Z(n449) );
  MUX2_X1 U323 ( .A(product[9]), .B(n536), .S(n14), .Z(n451) );
  OAI21_X1 U324 ( .B1(n283), .B2(n333), .A(n334), .ZN(n294) );
  INV_X1 U325 ( .A(n294), .ZN(n287) );
  NOR2_X1 U326 ( .A1(n348), .A2(n349), .ZN(n291) );
  INV_X1 U327 ( .A(n291), .ZN(n284) );
  NAND2_X1 U328 ( .A1(n348), .A2(n349), .ZN(n292) );
  NAND2_X1 U329 ( .A1(n284), .A2(n292), .ZN(n285) );
  XOR2_X1 U330 ( .A(n287), .B(n285), .Z(n286) );
  MUX2_X1 U331 ( .A(n536), .B(n286), .S(n324), .Z(n453) );
  MUX2_X1 U332 ( .A(product[10]), .B(n538), .S(n324), .Z(n455) );
  OAI21_X1 U333 ( .B1(n287), .B2(n291), .A(n292), .ZN(n289) );
  NAND2_X1 U334 ( .A1(n399), .A2(n340), .ZN(n288) );
  XNOR2_X1 U335 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U336 ( .A(n538), .B(n290), .S(n14), .Z(n457) );
  MUX2_X1 U337 ( .A(product[11]), .B(n540), .S(n324), .Z(n459) );
  NOR2_X1 U338 ( .A1(n339), .A2(n291), .ZN(n295) );
  OAI21_X1 U339 ( .B1(n339), .B2(n292), .A(n340), .ZN(n293) );
  AOI21_X1 U340 ( .B1(n295), .B2(n294), .A(n293), .ZN(n321) );
  NOR2_X1 U341 ( .A1(n346), .A2(n347), .ZN(n308) );
  INV_X1 U342 ( .A(n308), .ZN(n301) );
  NAND2_X1 U343 ( .A1(n346), .A2(n347), .ZN(n310) );
  NAND2_X1 U344 ( .A1(n301), .A2(n310), .ZN(n296) );
  XOR2_X1 U345 ( .A(n321), .B(n296), .Z(n297) );
  MUX2_X1 U346 ( .A(n540), .B(n297), .S(n14), .Z(n461) );
  MUX2_X1 U347 ( .A(product[12]), .B(n542), .S(n324), .Z(n463) );
  OAI21_X1 U348 ( .B1(n321), .B2(n308), .A(n310), .ZN(n299) );
  NAND2_X1 U349 ( .A1(n343), .A2(n342), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  MUX2_X1 U351 ( .A(n542), .B(n300), .S(n324), .Z(n465) );
  MUX2_X1 U352 ( .A(product[13]), .B(n544), .S(n14), .Z(n467) );
  NAND2_X1 U353 ( .A1(n301), .A2(n343), .ZN(n304) );
  INV_X1 U354 ( .A(n310), .ZN(n302) );
  AOI21_X1 U355 ( .B1(n302), .B2(n343), .A(n400), .ZN(n303) );
  OAI21_X1 U356 ( .B1(n321), .B2(n304), .A(n303), .ZN(n306) );
  NAND2_X1 U357 ( .A1(n329), .A2(n341), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  MUX2_X1 U359 ( .A(n544), .B(n307), .S(n324), .Z(n469) );
  MUX2_X1 U360 ( .A(product[14]), .B(n546), .S(n324), .Z(n471) );
  NAND2_X1 U361 ( .A1(n343), .A2(n329), .ZN(n311) );
  NOR2_X1 U362 ( .A1(n308), .A2(n311), .ZN(n317) );
  INV_X1 U363 ( .A(n317), .ZN(n313) );
  AOI21_X1 U364 ( .B1(n400), .B2(n329), .A(n396), .ZN(n309) );
  OAI21_X1 U365 ( .B1(n311), .B2(n310), .A(n309), .ZN(n318) );
  INV_X1 U366 ( .A(n318), .ZN(n312) );
  OAI21_X1 U367 ( .B1(n321), .B2(n313), .A(n312), .ZN(n315) );
  NAND2_X1 U368 ( .A1(n328), .A2(n332), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U370 ( .A(n546), .B(n316), .S(n15), .Z(n473) );
  MUX2_X1 U371 ( .A(product[15]), .B(n548), .S(n324), .Z(n475) );
  NAND2_X1 U372 ( .A1(n317), .A2(n328), .ZN(n320) );
  AOI21_X1 U373 ( .B1(n318), .B2(n328), .A(n394), .ZN(n319) );
  OAI21_X1 U374 ( .B1(n321), .B2(n320), .A(n319), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(n331), .ZN(n323) );
  MUX2_X1 U376 ( .A(n548), .B(n323), .S(n324), .Z(n477) );
  MUX2_X1 U377 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n324), .Z(n479) );
  MUX2_X1 U378 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n324), .Z(n481) );
  MUX2_X1 U379 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n15), .Z(n483) );
  MUX2_X1 U380 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n324), .Z(n485) );
  MUX2_X1 U381 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n14), .Z(n487) );
  MUX2_X1 U382 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n324), .Z(n489) );
  MUX2_X1 U383 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n15), .Z(n491) );
  MUX2_X1 U384 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n324), .Z(n493) );
  MUX2_X1 U385 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n15), .Z(n495) );
  MUX2_X1 U386 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n14), .Z(n497) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n324), .Z(n499) );
  MUX2_X1 U388 ( .A(n21), .B(A_extended[3]), .S(n324), .Z(n501) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n15), .Z(n503) );
  MUX2_X1 U390 ( .A(n22), .B(A_extended[5]), .S(n324), .Z(n505) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n324), .Z(n507) );
  MUX2_X1 U392 ( .A(n19), .B(A_extended[7]), .S(n324), .Z(n509) );
  OR2_X1 U393 ( .A1(n324), .A2(n550), .ZN(n511) );
endmodule


module conv_128_32_DW_mult_pipe_J1_17 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n378, n380, n382, n384, n386, n388, n390,
         n392, n394, n396, n398, n400, n402, n404, n406, n408, n410, n412,
         n414, n416, n418, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n432, n434, n436, n438, n440, n442, n444, n446,
         n448, n450, n452, n454, n456, n458, n460, n462, n464, n466, n468,
         n470, n472, n474, n476, n478, n480, n482, n484, n486, n488, n490,
         n492, n494, n496, n498, n500, n502, n504, n506, n508, n510, n512,
         n514, n516, n518, n520, n522, n524, n526, n528, n530, n532, n534,
         n536, n538, n540, n541, n543, n544, n546, n547, n549, n550, n552,
         n553, n555, n557, n559, n561, n563, n565, n567, n569, n571, n573,
         n575, n576, n577, n578, n579;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(rst_n), .SE(n538), .CK(clk), .Q(n578), 
        .QN(n429) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n534), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n23) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n530), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n15) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(rst_n), .SE(n526), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n13) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(rst_n), .SE(n524), .CK(clk), .Q(n576), 
        .QN(n24) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(rst_n), .SE(n522), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n18) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n520), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n518), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n516), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n512), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n510), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n508), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n504), .CK(clk), .Q(n575)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n502), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(rst_n), .SE(n500), .CK(clk), .Q(n573)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(rst_n), .SE(n498), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(rst_n), .SE(n496), .CK(clk), .Q(n571)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(rst_n), .SE(n492), .CK(clk), .Q(n569)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(rst_n), .SE(n490), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(rst_n), .SE(n488), .CK(clk), .Q(n567)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n486), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(rst_n), .SE(n484), .CK(clk), .Q(n565)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(rst_n), .SE(n482), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(rst_n), .SE(n480), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(rst_n), .SE(n478), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n476), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(rst_n), .SE(n474), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n470), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n468), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n466), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n464), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n462), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n460), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n458), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n456), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(rst_n), .SE(n454), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(rst_n), .SE(n452), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(rst_n), .SE(n450), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(rst_n), .SE(n448), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(rst_n), .SE(n446), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(rst_n), .SE(n444), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(rst_n), .SE(n442), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(rst_n), .SE(n440), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(rst_n), .SE(n438), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(rst_n), .SE(n436), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(rst_n), .SE(n434), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(rst_n), .SE(n432), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n536), .CK(clk), .Q(n577), 
        .QN(n430) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n579), .SI(1'b1), .SE(n412), .CK(clk), 
        .Q(n372), .QN(n25) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n579), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n361) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n579), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n364) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n579), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n579), .SE(n414), .CK(
        clk), .QN(n373) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n579), .SE(n418), .CK(
        clk), .QN(n375) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2_IP  ( .D(1'b1), .SI(n579), .SE(n416), .CK(
        clk), .QN(n374) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n579), .SE(n382), .CK(
        clk), .QN(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n579), .SE(n410), .CK(
        clk), .QN(n371) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n579), .SE(n402), .CK(
        clk), .Q(n353), .QN(n367) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n579), .SE(n384), .CK(
        clk), .QN(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n579), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n370), .QN(n428) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n579), .SE(n400), .CK(
        clk), .Q(n427), .QN(n366) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n579), .SE(n404), .CK(
        clk), .Q(n426), .QN(n368) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n579), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n365), .QN(n425) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n579), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n362), .QN(n424) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n579), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n360), .QN(n423) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n579), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n363), .QN(n422) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n579), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n369), .QN(n421) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n579), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n359), .QN(n420) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n579), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n579), .SE(n376), .CK(
        clk), .QN(n354) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(rst_n), .SE(n528), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n20) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n532), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n19) );
  INV_X1 U2 ( .A(rst_n), .ZN(n579) );
  XOR2_X1 U3 ( .A(n20), .B(n15), .Z(n5) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(n259) );
  NAND2_X1 U5 ( .A1(n52), .A2(n51), .ZN(n6) );
  XNOR2_X1 U6 ( .A(n52), .B(n51), .ZN(n8) );
  OR2_X1 U7 ( .A1(n30), .A2(n31), .ZN(n12) );
  NAND2_X1 U8 ( .A1(n27), .A2(n26), .ZN(n166) );
  CLKBUF_X2 U9 ( .A(n576), .Z(n351) );
  BUF_X1 U10 ( .A(\mult_x_1/n311 ), .Z(n17) );
  OAI21_X1 U11 ( .B1(n52), .B2(n51), .A(n50), .ZN(n7) );
  XNOR2_X1 U12 ( .A(n8), .B(n50), .ZN(n264) );
  NOR2_X1 U13 ( .A1(n101), .A2(n100), .ZN(n135) );
  INV_X1 U14 ( .A(n33), .ZN(n34) );
  NAND2_X1 U15 ( .A1(n126), .A2(n125), .ZN(n171) );
  NAND2_X1 U16 ( .A1(n136), .A2(n124), .ZN(n125) );
  OAI21_X1 U17 ( .B1(n136), .B2(n124), .A(n134), .ZN(n126) );
  INV_X1 U18 ( .A(n135), .ZN(n124) );
  XNOR2_X1 U19 ( .A(n137), .B(n136), .ZN(n143) );
  NAND2_X1 U20 ( .A1(n70), .A2(n69), .ZN(n71) );
  INV_X1 U21 ( .A(n73), .ZN(n69) );
  INV_X1 U22 ( .A(n74), .ZN(n70) );
  NAND2_X1 U23 ( .A1(n74), .A2(n73), .ZN(n75) );
  NAND2_X1 U24 ( .A1(n267), .A2(n266), .ZN(n268) );
  INV_X1 U25 ( .A(n270), .ZN(n266) );
  INV_X1 U26 ( .A(n271), .ZN(n267) );
  INV_X1 U27 ( .A(n5), .ZN(n164) );
  NAND2_X1 U28 ( .A1(n109), .A2(n108), .ZN(n145) );
  NAND2_X1 U29 ( .A1(n107), .A2(n106), .ZN(n108) );
  NAND2_X1 U30 ( .A1(n105), .A2(n21), .ZN(n109) );
  NAND2_X1 U31 ( .A1(n139), .A2(n138), .ZN(n191) );
  XNOR2_X1 U32 ( .A(n171), .B(n130), .ZN(n192) );
  XNOR2_X1 U33 ( .A(n173), .B(n172), .ZN(n130) );
  NAND2_X1 U34 ( .A1(n175), .A2(n174), .ZN(n187) );
  NAND2_X1 U35 ( .A1(n173), .A2(n172), .ZN(n174) );
  NAND2_X1 U36 ( .A1(n171), .A2(n22), .ZN(n175) );
  NAND2_X1 U37 ( .A1(n65), .A2(n64), .ZN(n89) );
  NAND2_X1 U38 ( .A1(n264), .A2(n63), .ZN(n65) );
  NAND2_X1 U39 ( .A1(n62), .A2(n61), .ZN(n63) );
  XNOR2_X1 U40 ( .A(n144), .B(n143), .ZN(n231) );
  XNOR2_X1 U41 ( .A(n269), .B(n203), .ZN(n209) );
  XNOR2_X1 U42 ( .A(n271), .B(n270), .ZN(n203) );
  XNOR2_X1 U43 ( .A(n105), .B(n85), .ZN(n94) );
  NAND2_X1 U44 ( .A1(n76), .A2(n75), .ZN(n96) );
  XNOR2_X1 U45 ( .A(n107), .B(n106), .ZN(n85) );
  XNOR2_X1 U46 ( .A(n264), .B(n263), .ZN(n265) );
  NAND2_X1 U47 ( .A1(n273), .A2(n272), .ZN(n274) );
  NAND2_X1 U48 ( .A1(n271), .A2(n270), .ZN(n272) );
  NAND2_X1 U49 ( .A1(n269), .A2(n268), .ZN(n273) );
  XOR2_X1 U50 ( .A(n13), .B(n20), .Z(n36) );
  INV_X1 U51 ( .A(n5), .ZN(n9) );
  OAI22_X1 U52 ( .A1(n166), .A2(n53), .B1(n164), .B2(n32), .ZN(n10) );
  NOR2_X2 U53 ( .A1(n429), .A2(n430), .ZN(n11) );
  NOR2_X1 U54 ( .A1(n429), .A2(n430), .ZN(n180) );
  OR2_X1 U55 ( .A1(n30), .A2(n31), .ZN(n177) );
  NAND2_X1 U56 ( .A1(n72), .A2(n71), .ZN(n76) );
  NAND2_X1 U57 ( .A1(n39), .A2(n38), .ZN(n103) );
  INV_X1 U58 ( .A(n78), .ZN(n37) );
  INV_X1 U59 ( .A(n262), .ZN(n62) );
  NAND2_X1 U60 ( .A1(n262), .A2(n261), .ZN(n64) );
  XNOR2_X1 U61 ( .A(n262), .B(n261), .ZN(n263) );
  INV_X1 U62 ( .A(n261), .ZN(n61) );
  OAI22_X1 U63 ( .A1(n250), .A2(n54), .B1(n248), .B2(n33), .ZN(n14) );
  INV_X1 U64 ( .A(n103), .ZN(n80) );
  XNOR2_X1 U65 ( .A(n20), .B(n15), .ZN(n27) );
  XOR2_X1 U66 ( .A(n180), .B(n352), .Z(n16) );
  BUF_X4 U67 ( .A(n577), .Z(n352) );
  OR2_X1 U68 ( .A1(n107), .A2(n106), .ZN(n21) );
  OR2_X1 U69 ( .A1(n173), .A2(n172), .ZN(n22) );
  XOR2_X1 U70 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n26) );
  XNOR2_X1 U71 ( .A(n17), .B(\mult_x_1/n284 ), .ZN(n53) );
  XNOR2_X1 U72 ( .A(n17), .B(\mult_x_1/n283 ), .ZN(n32) );
  OAI22_X1 U73 ( .A1(n166), .A2(n53), .B1(n164), .B2(n32), .ZN(n41) );
  XNOR2_X1 U74 ( .A(n576), .B(\mult_x_1/a[2] ), .ZN(n35) );
  NAND2_X2 U75 ( .A1(n36), .A2(n35), .ZN(n250) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n54) );
  INV_X1 U77 ( .A(n35), .ZN(n240) );
  INV_X2 U78 ( .A(n240), .ZN(n248) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n33) );
  OAI22_X1 U80 ( .A1(n250), .A2(n54), .B1(n248), .B2(n33), .ZN(n40) );
  XNOR2_X1 U81 ( .A(n40), .B(n41), .ZN(n52) );
  INV_X1 U82 ( .A(n11), .ZN(n28) );
  OR2_X1 U83 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n29) );
  XNOR2_X1 U84 ( .A(n180), .B(n352), .ZN(n47) );
  NOR2_X1 U85 ( .A1(n29), .A2(n47), .ZN(n51) );
  XNOR2_X1 U86 ( .A(\mult_x_1/a[6] ), .B(n352), .ZN(n30) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n311 ), .B(n23), .ZN(n31) );
  XNOR2_X1 U88 ( .A(n352), .B(\mult_x_1/n287 ), .ZN(n56) );
  INV_X1 U89 ( .A(n31), .ZN(n178) );
  XNOR2_X1 U90 ( .A(n352), .B(\mult_x_1/n286 ), .ZN(n46) );
  OAI22_X1 U91 ( .A1(n177), .A2(n56), .B1(n178), .B2(n46), .ZN(n199) );
  NAND2_X1 U92 ( .A1(n351), .A2(n18), .ZN(n242) );
  XNOR2_X1 U93 ( .A(n351), .B(\mult_x_1/n281 ), .ZN(n157) );
  AND2_X2 U94 ( .A1(n578), .A2(\mult_x_1/n281 ), .ZN(n127) );
  XNOR2_X1 U95 ( .A(n127), .B(n351), .ZN(n43) );
  OAI22_X1 U96 ( .A1(n242), .A2(n157), .B1(n43), .B2(n18), .ZN(n198) );
  AND2_X1 U97 ( .A1(\mult_x_1/n288 ), .A2(n16), .ZN(n197) );
  XNOR2_X1 U98 ( .A(n352), .B(\mult_x_1/n285 ), .ZN(n45) );
  XNOR2_X1 U99 ( .A(n352), .B(\mult_x_1/n284 ), .ZN(n77) );
  OAI22_X1 U100 ( .A1(n12), .A2(n45), .B1(n178), .B2(n77), .ZN(n82) );
  XNOR2_X1 U101 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n84) );
  OAI22_X1 U102 ( .A1(n166), .A2(n32), .B1(n164), .B2(n84), .ZN(n81) );
  NAND3_X1 U103 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n39) );
  XNOR2_X1 U104 ( .A(n127), .B(\mult_x_1/n312 ), .ZN(n78) );
  NAND2_X1 U105 ( .A1(n37), .A2(n240), .ZN(n38) );
  OR2_X2 U106 ( .A1(n10), .A2(n14), .ZN(n74) );
  XNOR2_X1 U107 ( .A(n11), .B(\mult_x_1/n286 ), .ZN(n42) );
  NOR2_X1 U108 ( .A1(n42), .A2(n47), .ZN(n73) );
  XNOR2_X1 U109 ( .A(n74), .B(n73), .ZN(n49) );
  AOI21_X1 U110 ( .B1(n242), .B2(n18), .A(n43), .ZN(n44) );
  INV_X1 U111 ( .A(n44), .ZN(n60) );
  OAI22_X1 U112 ( .A1(n177), .A2(n46), .B1(n178), .B2(n45), .ZN(n59) );
  XNOR2_X1 U113 ( .A(n11), .B(\mult_x_1/n287 ), .ZN(n48) );
  NOR2_X1 U114 ( .A1(n48), .A2(n47), .ZN(n58) );
  XNOR2_X1 U115 ( .A(n49), .B(n72), .ZN(n257) );
  XNOR2_X1 U116 ( .A(n17), .B(\mult_x_1/n285 ), .ZN(n156) );
  OAI22_X1 U117 ( .A1(n166), .A2(n156), .B1(n9), .B2(n53), .ZN(n196) );
  XNOR2_X1 U118 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n159) );
  OAI22_X1 U119 ( .A1(n250), .A2(n159), .B1(n248), .B2(n54), .ZN(n195) );
  OR2_X1 U120 ( .A1(\mult_x_1/n288 ), .A2(n430), .ZN(n55) );
  OAI22_X1 U121 ( .A1(n12), .A2(n430), .B1(n55), .B2(n178), .ZN(n155) );
  XNOR2_X1 U122 ( .A(n352), .B(\mult_x_1/n288 ), .ZN(n57) );
  OAI22_X1 U123 ( .A1(n177), .A2(n57), .B1(n178), .B2(n56), .ZN(n154) );
  FA_X1 U124 ( .A(n60), .B(n59), .CI(n58), .CO(n72), .S(n261) );
  INV_X1 U125 ( .A(n89), .ZN(n66) );
  INV_X1 U126 ( .A(en), .ZN(n120) );
  NAND2_X1 U127 ( .A1(n66), .A2(n299), .ZN(n68) );
  NAND2_X1 U128 ( .A1(n120), .A2(n366), .ZN(n67) );
  OAI21_X1 U129 ( .B1(n90), .B2(n68), .A(n67), .ZN(n400) );
  XNOR2_X1 U130 ( .A(n352), .B(\mult_x_1/n283 ), .ZN(n98) );
  OAI22_X1 U131 ( .A1(n12), .A2(n77), .B1(n178), .B2(n98), .ZN(n104) );
  AOI21_X1 U132 ( .B1(n248), .B2(n250), .A(n78), .ZN(n79) );
  INV_X1 U133 ( .A(n79), .ZN(n102) );
  FA_X1 U134 ( .A(n82), .B(n81), .CI(n80), .CO(n105), .S(n258) );
  XNOR2_X1 U135 ( .A(n11), .B(\mult_x_1/n285 ), .ZN(n83) );
  NOR2_X1 U136 ( .A1(n83), .A2(n47), .ZN(n107) );
  XNOR2_X1 U137 ( .A(n17), .B(\mult_x_1/n281 ), .ZN(n99) );
  OAI22_X1 U138 ( .A1(n166), .A2(n84), .B1(n9), .B2(n99), .ZN(n106) );
  NAND2_X1 U139 ( .A1(n86), .A2(n299), .ZN(n88) );
  OR2_X1 U140 ( .A1(n299), .A2(n25), .ZN(n87) );
  NAND2_X1 U141 ( .A1(n88), .A2(n87), .ZN(n412) );
  NAND2_X1 U142 ( .A1(n90), .A2(n89), .ZN(n91) );
  NAND2_X1 U143 ( .A1(n91), .A2(n299), .ZN(n93) );
  OR2_X1 U144 ( .A1(n299), .A2(n353), .ZN(n92) );
  NAND2_X1 U145 ( .A1(n93), .A2(n92), .ZN(n402) );
  FA_X1 U146 ( .A(n96), .B(n95), .CI(n94), .CO(n227), .S(n86) );
  XNOR2_X1 U147 ( .A(n11), .B(\mult_x_1/n284 ), .ZN(n97) );
  NOR2_X1 U148 ( .A1(n97), .A2(n47), .ZN(n133) );
  XNOR2_X1 U149 ( .A(n352), .B(\mult_x_1/n282 ), .ZN(n121) );
  OAI22_X1 U150 ( .A1(n12), .A2(n98), .B1(n178), .B2(n121), .ZN(n132) );
  XNOR2_X1 U151 ( .A(n127), .B(n17), .ZN(n122) );
  NOR2_X1 U152 ( .A1(n164), .A2(n122), .ZN(n101) );
  NOR2_X1 U153 ( .A1(n166), .A2(n99), .ZN(n100) );
  FA_X1 U154 ( .A(n104), .B(n102), .CI(n103), .CO(n146), .S(n95) );
  XNOR2_X1 U155 ( .A(n147), .B(n146), .ZN(n110) );
  XNOR2_X1 U156 ( .A(n110), .B(n145), .ZN(n228) );
  NAND2_X1 U157 ( .A1(n227), .A2(n228), .ZN(n111) );
  NAND2_X1 U158 ( .A1(n111), .A2(n299), .ZN(n113) );
  OR2_X1 U159 ( .A1(n299), .A2(n428), .ZN(n112) );
  NAND2_X1 U160 ( .A1(n113), .A2(n112), .ZN(n408) );
  XNOR2_X1 U183 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n117) );
  XNOR2_X1 U184 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n153) );
  OAI22_X1 U185 ( .A1(n250), .A2(n117), .B1(n248), .B2(n153), .ZN(n219) );
  XNOR2_X1 U186 ( .A(n351), .B(\mult_x_1/n284 ), .ZN(n116) );
  XNOR2_X1 U187 ( .A(n351), .B(\mult_x_1/n283 ), .ZN(n152) );
  OAI22_X1 U188 ( .A1(n242), .A2(n116), .B1(n152), .B2(n18), .ZN(n218) );
  OR2_X1 U189 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n114) );
  OAI22_X1 U190 ( .A1(n166), .A2(n19), .B1(n114), .B2(n9), .ZN(n162) );
  XNOR2_X1 U191 ( .A(n17), .B(\mult_x_1/n288 ), .ZN(n115) );
  XNOR2_X1 U192 ( .A(n17), .B(\mult_x_1/n287 ), .ZN(n165) );
  OAI22_X1 U193 ( .A1(n166), .A2(n115), .B1(n9), .B2(n165), .ZN(n161) );
  XNOR2_X1 U194 ( .A(n351), .B(\mult_x_1/n285 ), .ZN(n238) );
  OAI22_X1 U195 ( .A1(n242), .A2(n238), .B1(n116), .B2(n18), .ZN(n235) );
  AND2_X1 U196 ( .A1(\mult_x_1/n288 ), .A2(n5), .ZN(n234) );
  XNOR2_X1 U197 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n236) );
  OAI22_X1 U198 ( .A1(n250), .A2(n236), .B1(n248), .B2(n117), .ZN(n233) );
  NOR2_X1 U199 ( .A1(n225), .A2(n224), .ZN(n119) );
  NAND2_X1 U200 ( .A1(n120), .A2(n354), .ZN(n118) );
  OAI21_X1 U201 ( .B1(n120), .B2(n119), .A(n118), .ZN(n376) );
  XNOR2_X1 U202 ( .A(n352), .B(\mult_x_1/n281 ), .ZN(n128) );
  OAI22_X1 U203 ( .A1(n12), .A2(n121), .B1(n178), .B2(n128), .ZN(n136) );
  AOI21_X1 U204 ( .B1(n9), .B2(n166), .A(n122), .ZN(n123) );
  INV_X1 U205 ( .A(n123), .ZN(n134) );
  XNOR2_X1 U206 ( .A(n127), .B(n352), .ZN(n176) );
  OAI22_X1 U207 ( .A1(n12), .A2(n128), .B1(n176), .B2(n178), .ZN(n185) );
  INV_X1 U208 ( .A(n185), .ZN(n173) );
  XNOR2_X1 U209 ( .A(n11), .B(\mult_x_1/n282 ), .ZN(n129) );
  NOR2_X1 U210 ( .A1(n129), .A2(n47), .ZN(n172) );
  XNOR2_X1 U211 ( .A(n11), .B(\mult_x_1/n283 ), .ZN(n131) );
  NOR2_X1 U212 ( .A1(n131), .A2(n47), .ZN(n141) );
  FA_X1 U213 ( .A(n133), .B(n132), .CI(n135), .CO(n142), .S(n147) );
  XNOR2_X1 U214 ( .A(n135), .B(n123), .ZN(n137) );
  OAI21_X1 U215 ( .B1(n141), .B2(n142), .A(n143), .ZN(n139) );
  NAND2_X1 U216 ( .A1(n142), .A2(n141), .ZN(n138) );
  OR2_X1 U217 ( .A1(n192), .A2(n191), .ZN(n140) );
  MUX2_X1 U218 ( .A(n355), .B(n140), .S(n299), .Z(n378) );
  XNOR2_X1 U219 ( .A(n142), .B(n141), .ZN(n144) );
  NAND2_X1 U220 ( .A1(n145), .A2(n147), .ZN(n150) );
  NAND2_X1 U221 ( .A1(n145), .A2(n146), .ZN(n149) );
  NAND2_X1 U222 ( .A1(n147), .A2(n146), .ZN(n148) );
  NAND3_X1 U223 ( .A1(n150), .A2(n149), .A3(n148), .ZN(n230) );
  OR2_X1 U224 ( .A1(n231), .A2(n230), .ZN(n151) );
  MUX2_X1 U225 ( .A(n356), .B(n151), .S(n299), .Z(n380) );
  XNOR2_X1 U226 ( .A(n351), .B(\mult_x_1/n282 ), .ZN(n158) );
  OAI22_X1 U227 ( .A1(n242), .A2(n152), .B1(n158), .B2(n18), .ZN(n169) );
  AND2_X1 U228 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n168) );
  XNOR2_X1 U229 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n160) );
  OAI22_X1 U230 ( .A1(n250), .A2(n153), .B1(n248), .B2(n160), .ZN(n167) );
  HA_X1 U231 ( .A(n155), .B(n154), .CO(n194), .S(n205) );
  XNOR2_X1 U232 ( .A(n17), .B(\mult_x_1/n286 ), .ZN(n163) );
  OAI22_X1 U233 ( .A1(n166), .A2(n163), .B1(n9), .B2(n156), .ZN(n202) );
  OAI22_X1 U234 ( .A1(n242), .A2(n158), .B1(n157), .B2(n18), .ZN(n201) );
  OAI22_X1 U235 ( .A1(n250), .A2(n160), .B1(n248), .B2(n159), .ZN(n200) );
  HA_X1 U236 ( .A(n162), .B(n161), .CO(n216), .S(n217) );
  OAI22_X1 U237 ( .A1(n166), .A2(n165), .B1(n9), .B2(n163), .ZN(n215) );
  FA_X1 U238 ( .A(n169), .B(n168), .CI(n167), .CO(n206), .S(n214) );
  OR2_X1 U239 ( .A1(n212), .A2(n211), .ZN(n170) );
  MUX2_X1 U240 ( .A(n357), .B(n170), .S(n299), .Z(n382) );
  AOI21_X1 U241 ( .B1(n178), .B2(n12), .A(n176), .ZN(n179) );
  INV_X1 U242 ( .A(n179), .ZN(n183) );
  XNOR2_X1 U243 ( .A(\mult_x_1/n281 ), .B(n11), .ZN(n181) );
  NOR2_X1 U244 ( .A1(n181), .A2(n47), .ZN(n182) );
  XOR2_X1 U245 ( .A(n183), .B(n182), .Z(n184) );
  XOR2_X1 U246 ( .A(n185), .B(n184), .Z(n186) );
  OR2_X1 U247 ( .A1(n187), .A2(n186), .ZN(n189) );
  NAND2_X1 U248 ( .A1(n187), .A2(n186), .ZN(n188) );
  NAND2_X1 U249 ( .A1(n189), .A2(n188), .ZN(n190) );
  MUX2_X1 U250 ( .A(n358), .B(n190), .S(n299), .Z(n384) );
  NAND2_X1 U251 ( .A1(n192), .A2(n191), .ZN(n193) );
  MUX2_X1 U252 ( .A(n359), .B(n193), .S(n299), .Z(n386) );
  FA_X1 U253 ( .A(n196), .B(n195), .CI(n194), .CO(n262), .S(n269) );
  FA_X1 U254 ( .A(n197), .B(n198), .CI(n199), .CO(n50), .S(n271) );
  FA_X1 U255 ( .A(n202), .B(n201), .CI(n200), .CO(n270), .S(n204) );
  FA_X1 U256 ( .A(n206), .B(n205), .CI(n204), .CO(n208), .S(n212) );
  NOR2_X1 U257 ( .A1(n209), .A2(n208), .ZN(n207) );
  MUX2_X1 U258 ( .A(n360), .B(n207), .S(n299), .Z(n388) );
  NAND2_X1 U259 ( .A1(n209), .A2(n208), .ZN(n210) );
  MUX2_X1 U260 ( .A(n361), .B(n210), .S(n299), .Z(n390) );
  NAND2_X1 U261 ( .A1(n212), .A2(n211), .ZN(n213) );
  MUX2_X1 U262 ( .A(n362), .B(n213), .S(n299), .Z(n392) );
  FA_X1 U263 ( .A(n216), .B(n215), .CI(n214), .CO(n211), .S(n222) );
  FA_X1 U264 ( .A(n219), .B(n218), .CI(n217), .CO(n221), .S(n225) );
  NOR2_X1 U265 ( .A1(n222), .A2(n221), .ZN(n220) );
  MUX2_X1 U266 ( .A(n363), .B(n220), .S(n299), .Z(n394) );
  NAND2_X1 U267 ( .A1(n222), .A2(n221), .ZN(n223) );
  MUX2_X1 U268 ( .A(n364), .B(n223), .S(n299), .Z(n396) );
  NAND2_X1 U269 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U270 ( .A(n365), .B(n226), .S(n299), .Z(n398) );
  NOR2_X1 U271 ( .A1(n228), .A2(n227), .ZN(n229) );
  MUX2_X1 U272 ( .A(n368), .B(n229), .S(n299), .Z(n404) );
  NAND2_X1 U273 ( .A1(n231), .A2(n230), .ZN(n232) );
  MUX2_X1 U274 ( .A(n369), .B(n232), .S(n299), .Z(n406) );
  FA_X1 U275 ( .A(n235), .B(n234), .CI(n233), .CO(n224), .S(n255) );
  XNOR2_X1 U276 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n237) );
  OAI22_X1 U277 ( .A1(n250), .A2(n237), .B1(n248), .B2(n236), .ZN(n247) );
  XNOR2_X1 U278 ( .A(n351), .B(\mult_x_1/n286 ), .ZN(n239) );
  OAI22_X1 U279 ( .A1(n242), .A2(n239), .B1(n238), .B2(n18), .ZN(n246) );
  NOR2_X1 U280 ( .A1(n255), .A2(n254), .ZN(n291) );
  XNOR2_X1 U281 ( .A(n351), .B(\mult_x_1/n287 ), .ZN(n241) );
  OAI22_X1 U282 ( .A1(n242), .A2(n241), .B1(n239), .B2(n18), .ZN(n245) );
  AND2_X1 U283 ( .A1(\mult_x_1/n288 ), .A2(n240), .ZN(n244) );
  NOR2_X1 U284 ( .A1(n245), .A2(n244), .ZN(n280) );
  OAI22_X1 U285 ( .A1(n242), .A2(\mult_x_1/n288 ), .B1(n241), .B2(n18), .ZN(
        n277) );
  OR2_X1 U286 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n243) );
  NAND2_X1 U287 ( .A1(n243), .A2(n242), .ZN(n276) );
  NAND2_X1 U288 ( .A1(n277), .A2(n276), .ZN(n283) );
  NAND2_X1 U289 ( .A1(n245), .A2(n244), .ZN(n281) );
  OAI21_X1 U290 ( .B1(n280), .B2(n283), .A(n281), .ZN(n288) );
  HA_X1 U291 ( .A(n247), .B(n246), .CO(n254), .S(n252) );
  OR2_X1 U292 ( .A1(\mult_x_1/n288 ), .A2(n20), .ZN(n249) );
  OAI22_X1 U293 ( .A1(n250), .A2(n20), .B1(n249), .B2(n248), .ZN(n251) );
  OR2_X1 U294 ( .A1(n252), .A2(n251), .ZN(n287) );
  NAND2_X1 U295 ( .A1(n252), .A2(n251), .ZN(n286) );
  INV_X1 U296 ( .A(n286), .ZN(n253) );
  AOI21_X1 U297 ( .B1(n288), .B2(n287), .A(n253), .ZN(n294) );
  NAND2_X1 U298 ( .A1(n255), .A2(n254), .ZN(n293) );
  OAI21_X1 U299 ( .B1(n291), .B2(n294), .A(n293), .ZN(n256) );
  MUX2_X1 U300 ( .A(n371), .B(n256), .S(n299), .Z(n410) );
  FA_X1 U301 ( .A(n259), .B(n258), .CI(n257), .CO(n260), .S(n90) );
  MUX2_X1 U302 ( .A(n373), .B(n260), .S(n299), .Z(n414) );
  MUX2_X1 U303 ( .A(n374), .B(n265), .S(n299), .Z(n416) );
  MUX2_X1 U304 ( .A(n375), .B(n274), .S(n299), .Z(n418) );
  BUF_X4 U305 ( .A(en), .Z(n299) );
  MUX2_X1 U306 ( .A(product[0]), .B(n540), .S(n299), .Z(n432) );
  MUX2_X1 U307 ( .A(n540), .B(n541), .S(n299), .Z(n434) );
  AND2_X1 U308 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n275) );
  MUX2_X1 U309 ( .A(n541), .B(n275), .S(n299), .Z(n436) );
  MUX2_X1 U310 ( .A(product[1]), .B(n543), .S(n299), .Z(n438) );
  MUX2_X1 U311 ( .A(n543), .B(n544), .S(n299), .Z(n440) );
  OR2_X1 U312 ( .A1(n277), .A2(n276), .ZN(n278) );
  AND2_X1 U313 ( .A1(n278), .A2(n283), .ZN(n279) );
  MUX2_X1 U314 ( .A(n544), .B(n279), .S(n299), .Z(n442) );
  MUX2_X1 U315 ( .A(product[2]), .B(n546), .S(n299), .Z(n444) );
  MUX2_X1 U316 ( .A(n546), .B(n547), .S(n299), .Z(n446) );
  INV_X1 U317 ( .A(n280), .ZN(n282) );
  NAND2_X1 U318 ( .A1(n282), .A2(n281), .ZN(n284) );
  XOR2_X1 U319 ( .A(n284), .B(n283), .Z(n285) );
  MUX2_X1 U320 ( .A(n547), .B(n285), .S(n299), .Z(n448) );
  MUX2_X1 U321 ( .A(product[3]), .B(n549), .S(n299), .Z(n450) );
  MUX2_X1 U322 ( .A(n549), .B(n550), .S(n299), .Z(n452) );
  NAND2_X1 U323 ( .A1(n287), .A2(n286), .ZN(n289) );
  XNOR2_X1 U324 ( .A(n289), .B(n288), .ZN(n290) );
  MUX2_X1 U325 ( .A(n550), .B(n290), .S(n299), .Z(n454) );
  MUX2_X1 U326 ( .A(product[4]), .B(n552), .S(n299), .Z(n456) );
  MUX2_X1 U327 ( .A(n552), .B(n553), .S(n299), .Z(n458) );
  INV_X1 U328 ( .A(n291), .ZN(n292) );
  NAND2_X1 U329 ( .A1(n293), .A2(n292), .ZN(n296) );
  INV_X1 U330 ( .A(n294), .ZN(n295) );
  XNOR2_X1 U331 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U332 ( .A(n553), .B(n297), .S(n299), .Z(n460) );
  MUX2_X1 U333 ( .A(product[5]), .B(n555), .S(n299), .Z(n462) );
  NAND2_X1 U334 ( .A1(n354), .A2(n365), .ZN(n298) );
  XNOR2_X1 U335 ( .A(n298), .B(n371), .ZN(n300) );
  MUX2_X1 U336 ( .A(n555), .B(n300), .S(n299), .Z(n464) );
  CLKBUF_X1 U337 ( .A(en), .Z(n343) );
  MUX2_X1 U338 ( .A(product[6]), .B(n557), .S(n343), .Z(n466) );
  NAND2_X1 U339 ( .A1(n422), .A2(n364), .ZN(n301) );
  AOI21_X1 U340 ( .B1(n354), .B2(n371), .A(n425), .ZN(n303) );
  XOR2_X1 U341 ( .A(n301), .B(n303), .Z(n302) );
  MUX2_X1 U342 ( .A(n557), .B(n302), .S(n343), .Z(n468) );
  MUX2_X1 U343 ( .A(product[7]), .B(n559), .S(n343), .Z(n470) );
  OAI21_X1 U344 ( .B1(n363), .B2(n303), .A(n364), .ZN(n306) );
  NAND2_X1 U345 ( .A1(n357), .A2(n362), .ZN(n304) );
  XNOR2_X1 U346 ( .A(n306), .B(n304), .ZN(n305) );
  MUX2_X1 U347 ( .A(n559), .B(n305), .S(n343), .Z(n472) );
  MUX2_X1 U348 ( .A(product[8]), .B(n561), .S(n343), .Z(n474) );
  AOI21_X1 U349 ( .B1(n306), .B2(n357), .A(n424), .ZN(n309) );
  NAND2_X1 U350 ( .A1(n423), .A2(n361), .ZN(n307) );
  XOR2_X1 U351 ( .A(n309), .B(n307), .Z(n308) );
  MUX2_X1 U352 ( .A(n561), .B(n308), .S(n343), .Z(n476) );
  MUX2_X1 U353 ( .A(product[9]), .B(n563), .S(n343), .Z(n478) );
  OAI21_X1 U354 ( .B1(n309), .B2(n360), .A(n361), .ZN(n320) );
  INV_X1 U355 ( .A(n320), .ZN(n313) );
  NOR2_X1 U356 ( .A1(n374), .A2(n375), .ZN(n317) );
  INV_X1 U357 ( .A(n317), .ZN(n310) );
  NAND2_X1 U358 ( .A1(n374), .A2(n375), .ZN(n318) );
  NAND2_X1 U359 ( .A1(n310), .A2(n318), .ZN(n311) );
  XOR2_X1 U360 ( .A(n313), .B(n311), .Z(n312) );
  MUX2_X1 U361 ( .A(n563), .B(n312), .S(n343), .Z(n480) );
  MUX2_X1 U362 ( .A(product[10]), .B(n565), .S(n343), .Z(n482) );
  OAI21_X1 U363 ( .B1(n313), .B2(n317), .A(n318), .ZN(n315) );
  NAND2_X1 U364 ( .A1(n427), .A2(n367), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U366 ( .A(n565), .B(n316), .S(n343), .Z(n484) );
  MUX2_X1 U367 ( .A(product[11]), .B(n567), .S(n343), .Z(n486) );
  NOR2_X1 U368 ( .A1(n366), .A2(n317), .ZN(n321) );
  OAI21_X1 U369 ( .B1(n366), .B2(n318), .A(n367), .ZN(n319) );
  AOI21_X1 U370 ( .B1(n321), .B2(n320), .A(n319), .ZN(n348) );
  NOR2_X1 U371 ( .A1(n372), .A2(n373), .ZN(n334) );
  INV_X1 U372 ( .A(n334), .ZN(n327) );
  NAND2_X1 U373 ( .A1(n372), .A2(n373), .ZN(n336) );
  NAND2_X1 U374 ( .A1(n327), .A2(n336), .ZN(n322) );
  XOR2_X1 U375 ( .A(n348), .B(n322), .Z(n323) );
  MUX2_X1 U376 ( .A(n567), .B(n323), .S(n343), .Z(n488) );
  MUX2_X1 U377 ( .A(product[12]), .B(n569), .S(n343), .Z(n490) );
  OAI21_X1 U378 ( .B1(n348), .B2(n334), .A(n336), .ZN(n325) );
  NAND2_X1 U379 ( .A1(n426), .A2(n370), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U381 ( .A(n569), .B(n326), .S(n343), .Z(n492) );
  MUX2_X1 U382 ( .A(product[13]), .B(n571), .S(n343), .Z(n494) );
  NAND2_X1 U383 ( .A1(n327), .A2(n426), .ZN(n330) );
  INV_X1 U384 ( .A(n336), .ZN(n328) );
  AOI21_X1 U385 ( .B1(n328), .B2(n426), .A(n428), .ZN(n329) );
  OAI21_X1 U386 ( .B1(n348), .B2(n330), .A(n329), .ZN(n332) );
  NAND2_X1 U387 ( .A1(n356), .A2(n369), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  MUX2_X1 U389 ( .A(n571), .B(n333), .S(n343), .Z(n496) );
  MUX2_X1 U390 ( .A(product[14]), .B(n573), .S(n343), .Z(n498) );
  NAND2_X1 U391 ( .A1(n426), .A2(n356), .ZN(n337) );
  NOR2_X1 U392 ( .A1(n334), .A2(n337), .ZN(n344) );
  INV_X1 U393 ( .A(n344), .ZN(n339) );
  AOI21_X1 U394 ( .B1(n428), .B2(n356), .A(n421), .ZN(n335) );
  OAI21_X1 U395 ( .B1(n337), .B2(n336), .A(n335), .ZN(n345) );
  INV_X1 U396 ( .A(n345), .ZN(n338) );
  OAI21_X1 U397 ( .B1(n348), .B2(n339), .A(n338), .ZN(n341) );
  NAND2_X1 U398 ( .A1(n355), .A2(n359), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  MUX2_X1 U400 ( .A(n573), .B(n342), .S(n343), .Z(n500) );
  MUX2_X1 U401 ( .A(product[15]), .B(n575), .S(n343), .Z(n502) );
  NAND2_X1 U402 ( .A1(n344), .A2(n355), .ZN(n347) );
  AOI21_X1 U403 ( .B1(n345), .B2(n355), .A(n420), .ZN(n346) );
  OAI21_X1 U404 ( .B1(n348), .B2(n347), .A(n346), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n349), .B(n358), .ZN(n350) );
  MUX2_X1 U406 ( .A(n575), .B(n350), .S(n299), .Z(n504) );
  MUX2_X1 U407 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n299), .Z(n506) );
  MUX2_X1 U408 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n299), .Z(n508) );
  MUX2_X1 U409 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n299), .Z(n510) );
  MUX2_X1 U410 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n299), .Z(n512) );
  MUX2_X1 U411 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n299), .Z(n514) );
  MUX2_X1 U412 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n299), .Z(n516) );
  MUX2_X1 U413 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n299), .Z(n518) );
  MUX2_X1 U414 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n299), .Z(n520) );
  MUX2_X1 U415 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n299), .Z(n522) );
  MUX2_X1 U416 ( .A(n351), .B(A_extended[1]), .S(n299), .Z(n524) );
  MUX2_X1 U417 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n299), .Z(n526) );
  MUX2_X1 U418 ( .A(\mult_x_1/n312 ), .B(A_extended[3]), .S(n299), .Z(n528) );
  MUX2_X1 U419 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n299), .Z(n530) );
  MUX2_X1 U420 ( .A(n17), .B(A_extended[5]), .S(n299), .Z(n532) );
  MUX2_X1 U421 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n299), .Z(n534) );
  MUX2_X1 U422 ( .A(n352), .B(A_extended[7]), .S(n299), .Z(n536) );
  OR2_X1 U423 ( .A1(n299), .A2(n578), .ZN(n538) );
endmodule


module conv_128_32_DW_mult_pipe_J1_18 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n310 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n361, n363, n365, n367, n369,
         n371, n373, n375, n377, n379, n381, n383, n385, n387, n389, n391,
         n393, n395, n397, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n414, n416, n418, n420, n422,
         n424, n426, n428, n430, n432, n434, n436, n438, n440, n442, n444,
         n446, n448, n450, n452, n454, n456, n458, n460, n462, n464, n466,
         n468, n470, n472, n474, n476, n478, n480, n482, n484, n486, n488,
         n490, n492, n494, n496, n498, n500, n502, n504, n506, n508, n510,
         n512, n514, n516, n518, n520, n522, n524, n525, n527, n528, n530,
         n531, n533, n534, n536, n537, n539, n540, n542, n544, n546, n548,
         n550, n552, n554, n556, n558, n560, n561, n562, n563, n564, n565;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n412), .SE(n522), .CK(clk), .Q(n564)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n412), .SE(n518), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n338) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n412), .SE(n516), .CK(clk), .Q(n563), 
        .QN(n337) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n412), .SE(n514), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n37) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n412), .SE(n512), .CK(clk), .Q(n562), 
        .QN(n38) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n412), .SE(n510), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n412), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n36) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n412), .SE(n504), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n27) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n412), .SE(n502), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n410), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n411), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n409), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n412), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n409), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n409), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n6) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n409), .SE(n488), .CK(clk), .Q(n560)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n409), .SE(n486), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n409), .SE(n484), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n409), .SE(n482), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n409), .SE(n480), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n411), .SE(n478), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n410), .SE(n476), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n412), .SE(n474), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n409), .SE(n472), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n409), .SE(n470), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n409), .SE(n468), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n409), .SE(n466), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n409), .SE(n464), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n409), .SE(n462), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n409), .SE(n460), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n409), .SE(n458), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n411), .SE(n456), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n411), .SE(n454), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n411), .SE(n452), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n411), .SE(n450), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n411), .SE(n448), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n411), .SE(n446), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n411), .SE(n444), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n411), .SE(n442), .CK(clk), .Q(n537)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n411), .SE(n440), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n411), .SE(n438), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n411), .SE(n436), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n410), .SE(n434), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n410), .SE(n432), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n410), .SE(n430), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n410), .SE(n428), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n410), .SE(n426), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n410), .SE(n424), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n410), .SE(n422), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n410), .SE(n420), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n410), .SE(n418), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n410), .SE(n416), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n410), .SE(n414), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n565), .SI(1'b1), .SE(n397), .CK(clk), 
        .Q(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n565), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n565), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n565), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n355), .QN(n39) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n565), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n354), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n565), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n352), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n565), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n565), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n350), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n565), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n349), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n565), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n565), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n347), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n565), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n346), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n565), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n345), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n565), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n344), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n565), .SE(n367), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n565), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n565), .SE(n363), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n565), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n565), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n339), .QN(n401) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n412), .SE(n520), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n7) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n412), .SE(n508), .CK(clk), .Q(n561), 
        .QN(n40) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n565), .SE(n387), .CK(
        clk), .Q(n407), .QN(n353) );
  NAND2_X1 U2 ( .A1(n5), .A2(n216), .ZN(n218) );
  XNOR2_X1 U3 ( .A(n159), .B(n160), .ZN(n5) );
  BUF_X2 U4 ( .A(\mult_x_1/n310 ), .Z(n8) );
  XNOR2_X2 U5 ( .A(n175), .B(n8), .ZN(n56) );
  BUF_X1 U6 ( .A(n409), .Z(n412) );
  BUF_X1 U7 ( .A(n409), .Z(n411) );
  BUF_X1 U8 ( .A(n409), .Z(n410) );
  INV_X1 U9 ( .A(n565), .ZN(n409) );
  CLKBUF_X1 U10 ( .A(n83), .Z(n34) );
  OR2_X1 U11 ( .A1(n43), .A2(n29), .ZN(n83) );
  NAND2_X1 U12 ( .A1(n36), .A2(n561), .ZN(n237) );
  NAND2_X1 U13 ( .A1(n19), .A2(n18), .ZN(n71) );
  XNOR2_X1 U14 ( .A(n14), .B(n93), .ZN(n257) );
  OAI21_X1 U15 ( .B1(n24), .B2(n23), .A(n22), .ZN(n163) );
  NAND2_X1 U16 ( .A1(n189), .A2(n20), .ZN(n19) );
  XNOR2_X1 U17 ( .A(n95), .B(n94), .ZN(n14) );
  NAND2_X1 U18 ( .A1(n191), .A2(n190), .ZN(n18) );
  OR2_X1 U19 ( .A1(n191), .A2(n190), .ZN(n20) );
  NOR2_X1 U20 ( .A1(n101), .A2(n100), .ZN(n23) );
  NAND2_X1 U21 ( .A1(n101), .A2(n100), .ZN(n22) );
  INV_X1 U22 ( .A(n99), .ZN(n24) );
  OR2_X1 U23 ( .A1(n128), .A2(n127), .ZN(n17) );
  INV_X1 U24 ( .A(rst_n), .ZN(n565) );
  CLKBUF_X1 U25 ( .A(n83), .Z(n35) );
  INV_X1 U26 ( .A(n48), .ZN(n173) );
  INV_X1 U27 ( .A(n42), .ZN(n223) );
  INV_X1 U28 ( .A(n43), .ZN(n9) );
  AND2_X1 U29 ( .A1(n564), .A2(\mult_x_1/n281 ), .ZN(n111) );
  NAND2_X1 U30 ( .A1(n166), .A2(n10), .ZN(n167) );
  XNOR2_X1 U31 ( .A(n159), .B(n11), .ZN(n10) );
  INV_X1 U32 ( .A(n160), .ZN(n11) );
  NAND2_X1 U33 ( .A1(n13), .A2(n12), .ZN(n252) );
  NAND2_X1 U34 ( .A1(n95), .A2(n94), .ZN(n12) );
  OAI21_X1 U35 ( .B1(n94), .B2(n95), .A(n93), .ZN(n13) );
  NAND2_X1 U36 ( .A1(n16), .A2(n15), .ZN(n140) );
  INV_X1 U37 ( .A(n214), .ZN(n15) );
  INV_X1 U38 ( .A(n213), .ZN(n16) );
  NAND2_X1 U39 ( .A1(n126), .A2(n17), .ZN(n130) );
  NOR2_X1 U40 ( .A1(n56), .A2(n6), .ZN(n60) );
  NAND2_X1 U41 ( .A1(n197), .A2(n196), .ZN(n198) );
  XNOR2_X1 U42 ( .A(n189), .B(n21), .ZN(n197) );
  XNOR2_X1 U43 ( .A(n191), .B(n190), .ZN(n21) );
  NAND2_X1 U44 ( .A1(n46), .A2(n47), .ZN(n172) );
  XNOR2_X1 U45 ( .A(n337), .B(n338), .ZN(n47) );
  XNOR2_X1 U46 ( .A(n25), .B(n99), .ZN(n250) );
  XNOR2_X1 U47 ( .A(n101), .B(n100), .ZN(n25) );
  XNOR2_X1 U48 ( .A(n257), .B(n59), .ZN(n72) );
  XNOR2_X1 U49 ( .A(n258), .B(n259), .ZN(n59) );
  NAND2_X1 U50 ( .A1(n255), .A2(n254), .ZN(n256) );
  INV_X1 U51 ( .A(n259), .ZN(n255) );
  INV_X1 U52 ( .A(n258), .ZN(n254) );
  NAND2_X1 U53 ( .A1(n128), .A2(n127), .ZN(n129) );
  NAND2_X1 U54 ( .A1(n69), .A2(n336), .ZN(n70) );
  INV_X1 U55 ( .A(n71), .ZN(n69) );
  NAND2_X1 U56 ( .A1(n261), .A2(n260), .ZN(n262) );
  NAND2_X1 U57 ( .A1(n259), .A2(n258), .ZN(n260) );
  NAND2_X1 U58 ( .A1(n257), .A2(n256), .ZN(n261) );
  XNOR2_X1 U59 ( .A(n111), .B(n561), .ZN(n26) );
  INV_X1 U60 ( .A(n27), .ZN(n28) );
  XNOR2_X1 U61 ( .A(\mult_x_1/a[2] ), .B(n562), .ZN(n29) );
  OAI22_X1 U62 ( .A1(n152), .A2(n112), .B1(n113), .B2(n223), .ZN(n30) );
  NAND2_X1 U63 ( .A1(n130), .A2(n129), .ZN(n160) );
  INV_X1 U64 ( .A(n31), .ZN(n33) );
  AND2_X2 U65 ( .A1(n564), .A2(\mult_x_1/n310 ), .ZN(n175) );
  INV_X1 U66 ( .A(n563), .ZN(n31) );
  INV_X1 U67 ( .A(n31), .ZN(n32) );
  NAND2_X1 U68 ( .A1(n163), .A2(n162), .ZN(n164) );
  OAI21_X1 U69 ( .B1(n163), .B2(n162), .A(n161), .ZN(n165) );
  OAI22_X1 U70 ( .A1(n83), .A2(n82), .B1(n84), .B2(n9), .ZN(n135) );
  XNOR2_X1 U71 ( .A(n40), .B(\mult_x_1/a[2] ), .ZN(n43) );
  BUF_X2 U72 ( .A(en), .Z(n293) );
  BUF_X2 U73 ( .A(n562), .Z(n335) );
  XNOR2_X1 U74 ( .A(\mult_x_1/a[4] ), .B(n32), .ZN(n41) );
  XNOR2_X1 U75 ( .A(n562), .B(n37), .ZN(n42) );
  OR2_X2 U76 ( .A1(n41), .A2(n42), .ZN(n152) );
  XNOR2_X1 U77 ( .A(n33), .B(\mult_x_1/n284 ), .ZN(n49) );
  XNOR2_X1 U78 ( .A(n33), .B(\mult_x_1/n283 ), .ZN(n87) );
  OAI22_X1 U79 ( .A1(n152), .A2(n49), .B1(n223), .B2(n87), .ZN(n77) );
  XNOR2_X1 U80 ( .A(n335), .B(\mult_x_1/n282 ), .ZN(n50) );
  XNOR2_X1 U81 ( .A(n335), .B(\mult_x_1/n281 ), .ZN(n82) );
  OAI22_X1 U82 ( .A1(n83), .A2(n50), .B1(n9), .B2(n82), .ZN(n76) );
  XNOR2_X1 U83 ( .A(n77), .B(n76), .ZN(n95) );
  INV_X1 U84 ( .A(n175), .ZN(n44) );
  OR2_X1 U85 ( .A1(\mult_x_1/n288 ), .A2(n44), .ZN(n45) );
  NOR2_X1 U86 ( .A1(n45), .A2(n56), .ZN(n94) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n310 ), .B(n338), .ZN(n46) );
  XNOR2_X1 U88 ( .A(n8), .B(\mult_x_1/n287 ), .ZN(n52) );
  INV_X1 U89 ( .A(n47), .ZN(n48) );
  XNOR2_X1 U90 ( .A(n8), .B(\mult_x_1/n286 ), .ZN(n58) );
  OAI22_X1 U91 ( .A1(n172), .A2(n52), .B1(n173), .B2(n58), .ZN(n62) );
  XNOR2_X1 U92 ( .A(n561), .B(n28), .ZN(n64) );
  XNOR2_X1 U93 ( .A(n111), .B(n561), .ZN(n54) );
  OAI22_X1 U94 ( .A1(n237), .A2(n64), .B1(n54), .B2(n36), .ZN(n61) );
  XNOR2_X1 U95 ( .A(n33), .B(\mult_x_1/n285 ), .ZN(n63) );
  OAI22_X1 U96 ( .A1(n152), .A2(n63), .B1(n223), .B2(n49), .ZN(n68) );
  XNOR2_X1 U97 ( .A(n335), .B(\mult_x_1/n283 ), .ZN(n65) );
  OAI22_X1 U98 ( .A1(n35), .A2(n65), .B1(n9), .B2(n50), .ZN(n67) );
  OR2_X1 U99 ( .A1(\mult_x_1/n288 ), .A2(n7), .ZN(n51) );
  OAI22_X1 U100 ( .A1(n172), .A2(n7), .B1(n51), .B2(n173), .ZN(n144) );
  XNOR2_X1 U101 ( .A(n8), .B(\mult_x_1/n288 ), .ZN(n53) );
  OAI22_X1 U102 ( .A1(n172), .A2(n53), .B1(n173), .B2(n52), .ZN(n143) );
  AOI21_X1 U103 ( .B1(n237), .B2(n36), .A(n26), .ZN(n55) );
  INV_X1 U104 ( .A(n55), .ZN(n81) );
  XNOR2_X1 U105 ( .A(n175), .B(\mult_x_1/n287 ), .ZN(n57) );
  NOR2_X1 U106 ( .A1(n57), .A2(n56), .ZN(n80) );
  XNOR2_X1 U107 ( .A(n8), .B(\mult_x_1/n285 ), .ZN(n90) );
  OAI22_X1 U108 ( .A1(n172), .A2(n58), .B1(n173), .B2(n90), .ZN(n79) );
  FA_X1 U109 ( .A(n60), .B(n61), .CI(n62), .CO(n93), .S(n191) );
  XNOR2_X1 U110 ( .A(n33), .B(\mult_x_1/n286 ), .ZN(n150) );
  OAI22_X1 U111 ( .A1(n152), .A2(n150), .B1(n223), .B2(n63), .ZN(n147) );
  XNOR2_X1 U112 ( .A(n561), .B(\mult_x_1/n282 ), .ZN(n141) );
  OAI22_X1 U113 ( .A1(n237), .A2(n141), .B1(n64), .B2(n36), .ZN(n146) );
  XNOR2_X1 U114 ( .A(n335), .B(\mult_x_1/n284 ), .ZN(n142) );
  OAI22_X1 U115 ( .A1(n34), .A2(n142), .B1(n9), .B2(n65), .ZN(n145) );
  FA_X1 U116 ( .A(n68), .B(n67), .CI(n66), .CO(n258), .S(n189) );
  OAI22_X1 U117 ( .A1(n72), .A2(n70), .B1(n336), .B2(n406), .ZN(n373) );
  NAND2_X1 U118 ( .A1(n72), .A2(n71), .ZN(n73) );
  NAND2_X1 U119 ( .A1(n73), .A2(n293), .ZN(n75) );
  OR2_X1 U120 ( .A1(n293), .A2(n39), .ZN(n74) );
  NAND2_X1 U121 ( .A1(n75), .A2(n74), .ZN(n391) );
  OR2_X1 U122 ( .A1(n77), .A2(n76), .ZN(n101) );
  XNOR2_X1 U123 ( .A(n175), .B(\mult_x_1/n286 ), .ZN(n78) );
  NOR2_X1 U124 ( .A1(n78), .A2(n56), .ZN(n100) );
  FA_X1 U125 ( .A(n81), .B(n80), .CI(n79), .CO(n99), .S(n259) );
  XNOR2_X1 U126 ( .A(n8), .B(\mult_x_1/n284 ), .ZN(n89) );
  XNOR2_X1 U127 ( .A(n8), .B(\mult_x_1/n283 ), .ZN(n116) );
  OAI22_X1 U128 ( .A1(n172), .A2(n89), .B1(n173), .B2(n116), .ZN(n136) );
  XNOR2_X1 U129 ( .A(n111), .B(n335), .ZN(n84) );
  AOI21_X1 U130 ( .B1(n9), .B2(n35), .A(n84), .ZN(n85) );
  INV_X1 U131 ( .A(n85), .ZN(n134) );
  XNOR2_X1 U132 ( .A(n163), .B(n162), .ZN(n92) );
  XNOR2_X1 U133 ( .A(n175), .B(\mult_x_1/n285 ), .ZN(n86) );
  NOR2_X1 U134 ( .A1(n86), .A2(n56), .ZN(n128) );
  XNOR2_X1 U135 ( .A(n33), .B(\mult_x_1/n282 ), .ZN(n88) );
  XNOR2_X1 U136 ( .A(n33), .B(\mult_x_1/n281 ), .ZN(n112) );
  OAI22_X1 U137 ( .A1(n152), .A2(n88), .B1(n223), .B2(n112), .ZN(n127) );
  XNOR2_X1 U138 ( .A(n128), .B(n127), .ZN(n91) );
  INV_X1 U139 ( .A(n135), .ZN(n98) );
  OAI22_X1 U140 ( .A1(n223), .A2(n88), .B1(n152), .B2(n87), .ZN(n97) );
  OAI22_X1 U141 ( .A1(n172), .A2(n90), .B1(n173), .B2(n89), .ZN(n96) );
  XNOR2_X1 U142 ( .A(n91), .B(n126), .ZN(n161) );
  XNOR2_X1 U143 ( .A(n92), .B(n161), .ZN(n105) );
  FA_X1 U144 ( .A(n98), .B(n97), .CI(n96), .CO(n126), .S(n251) );
  INV_X1 U145 ( .A(n104), .ZN(n102) );
  NAND2_X1 U146 ( .A1(n102), .A2(n293), .ZN(n103) );
  OAI22_X1 U147 ( .A1(n105), .A2(n103), .B1(n293), .B2(n407), .ZN(n387) );
  NAND2_X1 U148 ( .A1(n105), .A2(n104), .ZN(n106) );
  NAND2_X1 U149 ( .A1(n106), .A2(n336), .ZN(n108) );
  OR2_X1 U150 ( .A1(n336), .A2(n400), .ZN(n107) );
  NAND2_X1 U151 ( .A1(n108), .A2(n107), .ZN(n371) );
  XNOR2_X1 U172 ( .A(n175), .B(\mult_x_1/n282 ), .ZN(n109) );
  NOR2_X1 U173 ( .A1(n109), .A2(n56), .ZN(n170) );
  XNOR2_X1 U174 ( .A(n8), .B(n28), .ZN(n110) );
  XNOR2_X1 U175 ( .A(n111), .B(n8), .ZN(n171) );
  OAI22_X1 U176 ( .A1(n172), .A2(n110), .B1(n171), .B2(n173), .ZN(n180) );
  INV_X1 U177 ( .A(n180), .ZN(n169) );
  XNOR2_X1 U178 ( .A(n8), .B(\mult_x_1/n282 ), .ZN(n115) );
  OAI22_X1 U179 ( .A1(n172), .A2(n115), .B1(n173), .B2(n110), .ZN(n121) );
  XNOR2_X1 U180 ( .A(n111), .B(n33), .ZN(n113) );
  OAI22_X1 U181 ( .A1(n152), .A2(n112), .B1(n113), .B2(n223), .ZN(n120) );
  AOI21_X1 U182 ( .B1(n223), .B2(n152), .A(n113), .ZN(n114) );
  INV_X1 U183 ( .A(n114), .ZN(n119) );
  INV_X1 U184 ( .A(n120), .ZN(n133) );
  OAI22_X1 U185 ( .A1(n172), .A2(n116), .B1(n173), .B2(n115), .ZN(n132) );
  XNOR2_X1 U186 ( .A(n175), .B(\mult_x_1/n284 ), .ZN(n117) );
  NOR2_X1 U187 ( .A1(n117), .A2(n56), .ZN(n131) );
  XNOR2_X1 U188 ( .A(n175), .B(\mult_x_1/n283 ), .ZN(n118) );
  NOR2_X1 U189 ( .A1(n118), .A2(n56), .ZN(n124) );
  FA_X1 U190 ( .A(n121), .B(n30), .CI(n119), .CO(n168), .S(n123) );
  OR2_X1 U191 ( .A1(n187), .A2(n186), .ZN(n122) );
  MUX2_X1 U192 ( .A(n339), .B(n122), .S(n336), .Z(n359) );
  FA_X1 U193 ( .A(n125), .B(n124), .CI(n123), .CO(n186), .S(n214) );
  FA_X1 U194 ( .A(n133), .B(n131), .CI(n132), .CO(n125), .S(n158) );
  NAND2_X1 U195 ( .A1(n160), .A2(n158), .ZN(n139) );
  FA_X1 U196 ( .A(n136), .B(n135), .CI(n134), .CO(n157), .S(n162) );
  NAND2_X1 U197 ( .A1(n160), .A2(n157), .ZN(n138) );
  NAND2_X1 U198 ( .A1(n158), .A2(n157), .ZN(n137) );
  NAND3_X1 U199 ( .A1(n139), .A2(n138), .A3(n137), .ZN(n213) );
  MUX2_X1 U200 ( .A(n340), .B(n140), .S(n336), .Z(n361) );
  XNOR2_X1 U201 ( .A(n561), .B(\mult_x_1/n283 ), .ZN(n206) );
  OAI22_X1 U202 ( .A1(n237), .A2(n206), .B1(n141), .B2(n36), .ZN(n155) );
  AND2_X1 U203 ( .A1(\mult_x_1/n288 ), .A2(n48), .ZN(n154) );
  XNOR2_X1 U204 ( .A(n335), .B(\mult_x_1/n285 ), .ZN(n205) );
  OAI22_X1 U205 ( .A1(n35), .A2(n205), .B1(n9), .B2(n142), .ZN(n153) );
  HA_X1 U206 ( .A(n144), .B(n143), .CO(n66), .S(n193) );
  FA_X1 U207 ( .A(n147), .B(n146), .CI(n145), .CO(n190), .S(n192) );
  OR2_X1 U208 ( .A1(\mult_x_1/n288 ), .A2(n337), .ZN(n148) );
  OAI22_X1 U209 ( .A1(n152), .A2(n337), .B1(n148), .B2(n223), .ZN(n208) );
  XNOR2_X1 U210 ( .A(n33), .B(\mult_x_1/n288 ), .ZN(n149) );
  XNOR2_X1 U211 ( .A(n33), .B(\mult_x_1/n287 ), .ZN(n151) );
  OAI22_X1 U212 ( .A1(n152), .A2(n149), .B1(n223), .B2(n151), .ZN(n207) );
  OAI22_X1 U213 ( .A1(n152), .A2(n151), .B1(n223), .B2(n150), .ZN(n203) );
  FA_X1 U214 ( .A(n155), .B(n154), .CI(n153), .CO(n194), .S(n202) );
  OR2_X1 U215 ( .A1(n200), .A2(n199), .ZN(n156) );
  MUX2_X1 U216 ( .A(n341), .B(n156), .S(n336), .Z(n363) );
  XNOR2_X1 U217 ( .A(n158), .B(n157), .ZN(n159) );
  NAND2_X1 U218 ( .A1(n165), .A2(n164), .ZN(n216) );
  INV_X1 U219 ( .A(n216), .ZN(n166) );
  MUX2_X1 U220 ( .A(n342), .B(n167), .S(n336), .Z(n365) );
  FA_X1 U221 ( .A(n170), .B(n169), .CI(n168), .CO(n182), .S(n187) );
  AOI21_X1 U222 ( .B1(n173), .B2(n172), .A(n171), .ZN(n174) );
  INV_X1 U223 ( .A(n174), .ZN(n178) );
  XNOR2_X1 U224 ( .A(n175), .B(n28), .ZN(n176) );
  NOR2_X1 U225 ( .A1(n176), .A2(n56), .ZN(n177) );
  XOR2_X1 U226 ( .A(n178), .B(n177), .Z(n179) );
  XOR2_X1 U227 ( .A(n180), .B(n179), .Z(n181) );
  OR2_X1 U228 ( .A1(n182), .A2(n181), .ZN(n184) );
  NAND2_X1 U229 ( .A1(n182), .A2(n181), .ZN(n183) );
  NAND2_X1 U230 ( .A1(n184), .A2(n183), .ZN(n185) );
  MUX2_X1 U231 ( .A(n343), .B(n185), .S(n336), .Z(n367) );
  NAND2_X1 U232 ( .A1(n187), .A2(n186), .ZN(n188) );
  MUX2_X1 U233 ( .A(n344), .B(n188), .S(n336), .Z(n369) );
  FA_X1 U234 ( .A(n194), .B(n193), .CI(n192), .CO(n196), .S(n200) );
  NOR2_X1 U235 ( .A1(n197), .A2(n196), .ZN(n195) );
  MUX2_X1 U236 ( .A(n347), .B(n195), .S(n336), .Z(n375) );
  MUX2_X1 U237 ( .A(n348), .B(n198), .S(n336), .Z(n377) );
  NAND2_X1 U238 ( .A1(n200), .A2(n199), .ZN(n201) );
  MUX2_X1 U239 ( .A(n349), .B(n201), .S(n336), .Z(n379) );
  FA_X1 U240 ( .A(n204), .B(n203), .CI(n202), .CO(n199), .S(n211) );
  XNOR2_X1 U241 ( .A(n335), .B(\mult_x_1/n286 ), .ZN(n224) );
  OAI22_X1 U242 ( .A1(n35), .A2(n224), .B1(n9), .B2(n205), .ZN(n221) );
  XNOR2_X1 U243 ( .A(n561), .B(\mult_x_1/n284 ), .ZN(n222) );
  OAI22_X1 U244 ( .A1(n237), .A2(n222), .B1(n206), .B2(n36), .ZN(n220) );
  HA_X1 U245 ( .A(n208), .B(n207), .CO(n204), .S(n219) );
  NOR2_X1 U246 ( .A1(n211), .A2(n210), .ZN(n209) );
  MUX2_X1 U247 ( .A(n350), .B(n209), .S(n336), .Z(n381) );
  NAND2_X1 U248 ( .A1(n211), .A2(n210), .ZN(n212) );
  MUX2_X1 U249 ( .A(n351), .B(n212), .S(n293), .Z(n383) );
  NAND2_X1 U250 ( .A1(n214), .A2(n213), .ZN(n215) );
  MUX2_X1 U251 ( .A(n352), .B(n215), .S(n293), .Z(n385) );
  MUX2_X1 U252 ( .A(n354), .B(n218), .S(n293), .Z(n389) );
  FA_X1 U253 ( .A(n221), .B(n220), .CI(n219), .CO(n210), .S(n247) );
  XNOR2_X1 U254 ( .A(n561), .B(\mult_x_1/n285 ), .ZN(n230) );
  OAI22_X1 U255 ( .A1(n237), .A2(n230), .B1(n222), .B2(n36), .ZN(n227) );
  AND2_X1 U256 ( .A1(\mult_x_1/n288 ), .A2(n42), .ZN(n226) );
  XNOR2_X1 U257 ( .A(n335), .B(\mult_x_1/n287 ), .ZN(n228) );
  OAI22_X1 U258 ( .A1(n34), .A2(n228), .B1(n9), .B2(n224), .ZN(n225) );
  OR2_X1 U259 ( .A1(n247), .A2(n246), .ZN(n286) );
  FA_X1 U260 ( .A(n227), .B(n226), .CI(n225), .CO(n246), .S(n245) );
  XNOR2_X1 U261 ( .A(n335), .B(\mult_x_1/n288 ), .ZN(n229) );
  OAI22_X1 U262 ( .A1(n34), .A2(n229), .B1(n9), .B2(n228), .ZN(n232) );
  XNOR2_X1 U263 ( .A(n561), .B(\mult_x_1/n286 ), .ZN(n234) );
  OAI22_X1 U264 ( .A1(n237), .A2(n234), .B1(n230), .B2(n36), .ZN(n231) );
  NOR2_X1 U265 ( .A1(n245), .A2(n244), .ZN(n279) );
  HA_X1 U266 ( .A(n232), .B(n231), .CO(n244), .S(n242) );
  OR2_X1 U267 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n233) );
  OAI22_X1 U268 ( .A1(n34), .A2(n38), .B1(n233), .B2(n9), .ZN(n241) );
  OR2_X1 U269 ( .A1(n242), .A2(n241), .ZN(n275) );
  XNOR2_X1 U270 ( .A(n561), .B(\mult_x_1/n287 ), .ZN(n236) );
  OAI22_X1 U271 ( .A1(n237), .A2(n236), .B1(n234), .B2(n36), .ZN(n240) );
  INV_X1 U272 ( .A(n9), .ZN(n235) );
  AND2_X1 U273 ( .A1(\mult_x_1/n288 ), .A2(n235), .ZN(n239) );
  NOR2_X1 U274 ( .A1(n240), .A2(n239), .ZN(n268) );
  OAI22_X1 U275 ( .A1(n237), .A2(\mult_x_1/n288 ), .B1(n236), .B2(n36), .ZN(
        n265) );
  OR2_X1 U276 ( .A1(\mult_x_1/n288 ), .A2(n40), .ZN(n238) );
  NAND2_X1 U277 ( .A1(n238), .A2(n237), .ZN(n264) );
  NAND2_X1 U278 ( .A1(n265), .A2(n264), .ZN(n271) );
  NAND2_X1 U279 ( .A1(n240), .A2(n239), .ZN(n269) );
  OAI21_X1 U280 ( .B1(n268), .B2(n271), .A(n269), .ZN(n276) );
  NAND2_X1 U281 ( .A1(n242), .A2(n241), .ZN(n274) );
  INV_X1 U282 ( .A(n274), .ZN(n243) );
  AOI21_X1 U283 ( .B1(n275), .B2(n276), .A(n243), .ZN(n282) );
  NAND2_X1 U284 ( .A1(n245), .A2(n244), .ZN(n280) );
  OAI21_X1 U285 ( .B1(n279), .B2(n282), .A(n280), .ZN(n287) );
  NAND2_X1 U286 ( .A1(n247), .A2(n246), .ZN(n285) );
  INV_X1 U287 ( .A(n285), .ZN(n248) );
  AOI21_X1 U288 ( .B1(n286), .B2(n287), .A(n248), .ZN(n249) );
  MUX2_X1 U289 ( .A(n356), .B(n249), .S(n293), .Z(n393) );
  FA_X1 U290 ( .A(n252), .B(n251), .CI(n250), .CO(n104), .S(n253) );
  MUX2_X1 U291 ( .A(n357), .B(n253), .S(n293), .Z(n395) );
  MUX2_X1 U292 ( .A(n358), .B(n262), .S(n293), .Z(n397) );
  MUX2_X1 U293 ( .A(product[0]), .B(n524), .S(n293), .Z(n414) );
  MUX2_X1 U294 ( .A(n524), .B(n525), .S(n293), .Z(n416) );
  AND2_X1 U295 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n263) );
  MUX2_X1 U296 ( .A(n525), .B(n263), .S(n293), .Z(n418) );
  MUX2_X1 U297 ( .A(product[1]), .B(n527), .S(n293), .Z(n420) );
  MUX2_X1 U298 ( .A(n527), .B(n528), .S(n293), .Z(n422) );
  OR2_X1 U299 ( .A1(n265), .A2(n264), .ZN(n266) );
  AND2_X1 U300 ( .A1(n266), .A2(n271), .ZN(n267) );
  MUX2_X1 U301 ( .A(n528), .B(n267), .S(n293), .Z(n424) );
  MUX2_X1 U302 ( .A(product[2]), .B(n530), .S(n293), .Z(n426) );
  MUX2_X1 U303 ( .A(n530), .B(n531), .S(n293), .Z(n428) );
  INV_X1 U304 ( .A(n268), .ZN(n270) );
  NAND2_X1 U305 ( .A1(n270), .A2(n269), .ZN(n272) );
  XOR2_X1 U306 ( .A(n272), .B(n271), .Z(n273) );
  MUX2_X1 U307 ( .A(n531), .B(n273), .S(n293), .Z(n430) );
  MUX2_X1 U308 ( .A(product[3]), .B(n533), .S(n293), .Z(n432) );
  MUX2_X1 U309 ( .A(n533), .B(n534), .S(n293), .Z(n434) );
  NAND2_X1 U310 ( .A1(n275), .A2(n274), .ZN(n277) );
  XNOR2_X1 U311 ( .A(n277), .B(n276), .ZN(n278) );
  MUX2_X1 U312 ( .A(n534), .B(n278), .S(n293), .Z(n436) );
  MUX2_X1 U313 ( .A(product[4]), .B(n536), .S(n293), .Z(n438) );
  MUX2_X1 U314 ( .A(n536), .B(n537), .S(n293), .Z(n440) );
  INV_X1 U315 ( .A(n279), .ZN(n281) );
  NAND2_X1 U316 ( .A1(n281), .A2(n280), .ZN(n283) );
  XOR2_X1 U317 ( .A(n283), .B(n282), .Z(n284) );
  MUX2_X1 U318 ( .A(n537), .B(n284), .S(n293), .Z(n442) );
  MUX2_X1 U319 ( .A(product[5]), .B(n539), .S(n293), .Z(n444) );
  MUX2_X1 U320 ( .A(n539), .B(n540), .S(n293), .Z(n446) );
  NAND2_X1 U321 ( .A1(n286), .A2(n285), .ZN(n288) );
  XNOR2_X1 U322 ( .A(n288), .B(n287), .ZN(n289) );
  MUX2_X1 U323 ( .A(n540), .B(n289), .S(n293), .Z(n448) );
  MUX2_X1 U324 ( .A(product[6]), .B(n542), .S(n293), .Z(n450) );
  NAND2_X1 U325 ( .A1(n402), .A2(n351), .ZN(n290) );
  XOR2_X1 U326 ( .A(n290), .B(n356), .Z(n291) );
  MUX2_X1 U327 ( .A(n542), .B(n291), .S(n293), .Z(n452) );
  MUX2_X1 U328 ( .A(product[7]), .B(n544), .S(n293), .Z(n454) );
  OAI21_X1 U329 ( .B1(n350), .B2(n356), .A(n351), .ZN(n295) );
  NAND2_X1 U330 ( .A1(n341), .A2(n349), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n295), .B(n292), .ZN(n294) );
  MUX2_X1 U332 ( .A(n544), .B(n294), .S(n293), .Z(n456) );
  BUF_X4 U333 ( .A(en), .Z(n336) );
  MUX2_X1 U334 ( .A(product[8]), .B(n546), .S(n336), .Z(n458) );
  AOI21_X1 U335 ( .B1(n295), .B2(n341), .A(n404), .ZN(n298) );
  NAND2_X1 U336 ( .A1(n405), .A2(n348), .ZN(n296) );
  XOR2_X1 U337 ( .A(n298), .B(n296), .Z(n297) );
  MUX2_X1 U338 ( .A(n546), .B(n297), .S(n336), .Z(n460) );
  MUX2_X1 U339 ( .A(product[9]), .B(n548), .S(n336), .Z(n462) );
  OAI21_X1 U340 ( .B1(n298), .B2(n347), .A(n348), .ZN(n309) );
  INV_X1 U341 ( .A(n309), .ZN(n301) );
  NAND2_X1 U342 ( .A1(n406), .A2(n355), .ZN(n299) );
  XOR2_X1 U343 ( .A(n301), .B(n299), .Z(n300) );
  MUX2_X1 U344 ( .A(n548), .B(n300), .S(n336), .Z(n464) );
  MUX2_X1 U345 ( .A(product[10]), .B(n550), .S(n336), .Z(n466) );
  OAI21_X1 U346 ( .B1(n301), .B2(n346), .A(n355), .ZN(n304) );
  NOR2_X1 U347 ( .A1(n357), .A2(n358), .ZN(n307) );
  INV_X1 U348 ( .A(n307), .ZN(n302) );
  NAND2_X1 U349 ( .A1(n357), .A2(n358), .ZN(n306) );
  NAND2_X1 U350 ( .A1(n302), .A2(n306), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  MUX2_X1 U352 ( .A(n550), .B(n305), .S(n336), .Z(n468) );
  MUX2_X1 U353 ( .A(product[11]), .B(n552), .S(n336), .Z(n470) );
  NOR2_X1 U354 ( .A1(n307), .A2(n346), .ZN(n310) );
  OAI21_X1 U355 ( .B1(n307), .B2(n355), .A(n306), .ZN(n308) );
  AOI21_X1 U356 ( .B1(n310), .B2(n309), .A(n308), .ZN(n332) );
  NAND2_X1 U357 ( .A1(n407), .A2(n345), .ZN(n311) );
  XOR2_X1 U358 ( .A(n332), .B(n311), .Z(n312) );
  MUX2_X1 U359 ( .A(n552), .B(n312), .S(n336), .Z(n472) );
  MUX2_X1 U360 ( .A(product[12]), .B(n554), .S(n336), .Z(n474) );
  OAI21_X1 U361 ( .B1(n332), .B2(n353), .A(n345), .ZN(n314) );
  NAND2_X1 U362 ( .A1(n342), .A2(n354), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U364 ( .A(n554), .B(n315), .S(n336), .Z(n476) );
  MUX2_X1 U365 ( .A(product[13]), .B(n556), .S(n336), .Z(n478) );
  NAND2_X1 U366 ( .A1(n407), .A2(n342), .ZN(n317) );
  AOI21_X1 U367 ( .B1(n400), .B2(n342), .A(n408), .ZN(n316) );
  OAI21_X1 U368 ( .B1(n332), .B2(n317), .A(n316), .ZN(n319) );
  NAND2_X1 U369 ( .A1(n340), .A2(n352), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  MUX2_X1 U371 ( .A(n556), .B(n320), .S(n336), .Z(n480) );
  MUX2_X1 U372 ( .A(product[14]), .B(n558), .S(n336), .Z(n482) );
  NAND2_X1 U373 ( .A1(n342), .A2(n340), .ZN(n327) );
  OR2_X1 U374 ( .A1(n353), .A2(n327), .ZN(n323) );
  AOI21_X1 U375 ( .B1(n408), .B2(n340), .A(n403), .ZN(n321) );
  OAI21_X1 U376 ( .B1(n327), .B2(n345), .A(n321), .ZN(n329) );
  INV_X1 U377 ( .A(n329), .ZN(n322) );
  OAI21_X1 U378 ( .B1(n332), .B2(n323), .A(n322), .ZN(n325) );
  NAND2_X1 U379 ( .A1(n339), .A2(n344), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U381 ( .A(n558), .B(n326), .S(n336), .Z(n484) );
  MUX2_X1 U382 ( .A(product[15]), .B(n560), .S(n336), .Z(n486) );
  NOR2_X1 U383 ( .A1(n327), .A2(n401), .ZN(n328) );
  NAND2_X1 U384 ( .A1(n407), .A2(n328), .ZN(n331) );
  AOI21_X1 U385 ( .B1(n329), .B2(n339), .A(n399), .ZN(n330) );
  OAI21_X1 U386 ( .B1(n332), .B2(n331), .A(n330), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n333), .B(n343), .ZN(n334) );
  MUX2_X1 U388 ( .A(n560), .B(n334), .S(n336), .Z(n488) );
  MUX2_X1 U389 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n336), .Z(n490) );
  MUX2_X1 U390 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n336), .Z(n492) );
  MUX2_X1 U391 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n336), .Z(n494) );
  MUX2_X1 U392 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n336), .Z(n496) );
  MUX2_X1 U393 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n336), .Z(n498) );
  MUX2_X1 U394 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n336), .Z(n500) );
  MUX2_X1 U395 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n336), .Z(n502) );
  MUX2_X1 U396 ( .A(n28), .B(B_extended[7]), .S(n336), .Z(n504) );
  MUX2_X1 U397 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n336), .Z(n506) );
  MUX2_X1 U398 ( .A(n561), .B(A_extended[1]), .S(n336), .Z(n508) );
  MUX2_X1 U399 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n336), .Z(n510) );
  MUX2_X1 U400 ( .A(n335), .B(A_extended[3]), .S(n336), .Z(n512) );
  MUX2_X1 U401 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n336), .Z(n514) );
  MUX2_X1 U402 ( .A(n32), .B(A_extended[5]), .S(n336), .Z(n516) );
  MUX2_X1 U403 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n336), .Z(n518) );
  MUX2_X1 U404 ( .A(n8), .B(A_extended[7]), .S(n336), .Z(n520) );
  OR2_X1 U405 ( .A1(n336), .A2(n564), .ZN(n522) );
endmodule


module conv_128_32_DW_mult_pipe_J1_19 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n350, n352, n354, n356, n358,
         n360, n362, n364, n366, n368, n370, n372, n374, n376, n378, n380,
         n382, n384, n386, n388, n390, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n403, n405, n407, n409, n411, n413, n415,
         n417, n419, n421, n423, n425, n427, n429, n431, n433, n435, n437,
         n439, n441, n443, n445, n447, n449, n451, n453, n455, n457, n459,
         n461, n463, n465, n467, n469, n471, n473, n475, n477, n479, n481,
         n483, n485, n487, n489, n491, n493, n495, n497, n499, n501, n503,
         n505, n507, n509, n511, n512, n514, n515, n517, n518, n520, n521,
         n523, n524, n526, n528, n530, n532, n534, n536, n538, n540, n542,
         n544, n546, n547, n548, n549, n550, n551;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(rst_n), .SE(n509), .CK(clk), .Q(n550), 
        .QN(n400) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n507), .CK(clk), .Q(n549), 
        .QN(n401) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n505), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n501), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(rst_n), .SE(n497), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(rst_n), .SE(n495), .CK(clk), .Q(n547), 
        .QN(n26) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n399), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n399), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n20), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n399), .SE(n479), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n20), .SE(n477), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n325) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n399), .SE(n475), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n20), .SE(n473), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n399), .SE(n471), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n20), .SE(n469), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n20), .SE(n467), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n20), .SE(n465), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(rst_n), .SE(n463), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n20), .SE(n461), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n399), .SE(n459), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n20), .SE(n457), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n399), .SE(n455), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n20), .SE(n453), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n399), .SE(n451), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n20), .SE(n449), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n399), .SE(n447), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n20), .SE(n445), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n399), .SE(n443), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n20), .SE(n441), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n399), .SE(n439), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n20), .SE(n437), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n399), .SE(n435), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n20), .SE(n433), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n399), .SE(n431), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n399), .SE(n429), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n20), .SE(n427), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n399), .SE(n425), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n20), .SE(n423), .CK(clk), .Q(n520)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n399), .SE(n421), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n20), .SE(n419), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n399), .SE(n417), .CK(clk), .Q(n517)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(rst_n), .SE(n415), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(rst_n), .SE(n413), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(rst_n), .SE(n411), .CK(clk), .Q(n514)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n20), .SE(n409), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n399), .SE(n407), .CK(clk), .Q(n512)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(rst_n), .SE(n405), .CK(clk), .Q(n511)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(rst_n), .SE(n403), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n551), .SE(n390), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n551), .SE(n388), .CK(
        clk), .QN(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2_IP  ( .D(1'b1), .SI(n551), .SE(n386), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n551), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2_IP  ( .D(1'b1), .SI(n551), .SE(n382), .CK(
        clk), .QN(n343) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n551), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n551), .SE(n378), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n551), .SE(n376), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2_IP  ( .D(1'b1), .SI(n551), .SE(n374), .CK(
        clk), .Q(n392), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n551), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n338), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n551), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n337), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n551), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n551), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n335), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n551), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n334), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n551), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n333) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n551), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n332), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n551), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n331), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n551), .SE(n356), .CK(
        clk), .QN(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n551), .SE(n354), .CK(
        clk), .QN(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n551), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n328) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n551), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n327) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2_IP  ( .D(1'b1), .SI(n551), .SE(n348), .CK(
        clk), .QN(n326) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(rst_n), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n25) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n503), .CK(clk), .Q(n548), 
        .QN(n24) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(rst_n), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n23) );
  NAND2_X1 U2 ( .A1(n35), .A2(n36), .ZN(n130) );
  NAND2_X2 U3 ( .A1(n28), .A2(n29), .ZN(n66) );
  INV_X1 U4 ( .A(n551), .ZN(n20) );
  INV_X1 U5 ( .A(n551), .ZN(n399) );
  BUF_X4 U6 ( .A(en), .Z(n324) );
  CLKBUF_X2 U7 ( .A(n195), .Z(n5) );
  CLKBUF_X2 U8 ( .A(n549), .Z(n21) );
  INV_X1 U9 ( .A(n73), .ZN(n242) );
  XNOR2_X1 U10 ( .A(n21), .B(\mult_x_1/n287 ), .ZN(n57) );
  OAI22_X1 U11 ( .A1(n44), .A2(n23), .B1(n200), .B2(n114), .ZN(n148) );
  XNOR2_X1 U12 ( .A(n76), .B(n547), .ZN(n44) );
  OAI22_X1 U13 ( .A1(n195), .A2(n40), .B1(n197), .B2(n95), .ZN(n218) );
  NAND2_X1 U14 ( .A1(n221), .A2(n220), .ZN(n106) );
  NAND2_X1 U15 ( .A1(n104), .A2(n103), .ZN(n105) );
  INV_X1 U16 ( .A(n221), .ZN(n103) );
  INV_X1 U17 ( .A(n220), .ZN(n104) );
  XNOR2_X1 U18 ( .A(n221), .B(n220), .ZN(n222) );
  NAND2_X1 U19 ( .A1(n233), .A2(n232), .ZN(n234) );
  INV_X1 U20 ( .A(n26), .ZN(n7) );
  INV_X1 U21 ( .A(n73), .ZN(n8) );
  INV_X1 U22 ( .A(n73), .ZN(n9) );
  INV_X1 U23 ( .A(n73), .ZN(n10) );
  XOR2_X1 U24 ( .A(n241), .B(n240), .Z(n11) );
  XOR2_X1 U25 ( .A(n239), .B(n11), .Z(n161) );
  NAND2_X1 U26 ( .A1(n239), .A2(n241), .ZN(n12) );
  NAND2_X1 U27 ( .A1(n239), .A2(n240), .ZN(n13) );
  NAND2_X1 U28 ( .A1(n241), .A2(n240), .ZN(n14) );
  NAND3_X1 U29 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n243) );
  BUF_X2 U30 ( .A(n29), .Z(n15) );
  INV_X1 U31 ( .A(n25), .ZN(n16) );
  NAND2_X1 U32 ( .A1(n30), .A2(n31), .ZN(n195) );
  INV_X1 U33 ( .A(n32), .ZN(n17) );
  INV_X1 U34 ( .A(n32), .ZN(n197) );
  XNOR2_X1 U35 ( .A(n133), .B(n21), .ZN(n18) );
  XNOR2_X1 U36 ( .A(n133), .B(n21), .ZN(n19) );
  NAND2_X1 U37 ( .A1(n107), .A2(n106), .ZN(n210) );
  INV_X1 U38 ( .A(n24), .ZN(n22) );
  INV_X1 U39 ( .A(n73), .ZN(n172) );
  BUF_X1 U40 ( .A(en), .Z(n253) );
  OR2_X1 U41 ( .A1(n231), .A2(n230), .ZN(n27) );
  XOR2_X1 U42 ( .A(\mult_x_1/a[4] ), .B(n548), .Z(n28) );
  XNOR2_X1 U43 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n29) );
  XNOR2_X1 U44 ( .A(n22), .B(\mult_x_1/n284 ), .ZN(n53) );
  XNOR2_X1 U45 ( .A(n22), .B(\mult_x_1/n283 ), .ZN(n39) );
  OAI22_X1 U46 ( .A1(n66), .A2(n53), .B1(n15), .B2(n39), .ZN(n42) );
  XOR2_X1 U47 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n30) );
  XNOR2_X1 U48 ( .A(\mult_x_1/a[2] ), .B(n547), .ZN(n31) );
  XNOR2_X1 U49 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n54) );
  INV_X1 U50 ( .A(n31), .ZN(n32) );
  XNOR2_X1 U51 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n40) );
  OAI22_X1 U52 ( .A1(n195), .A2(n54), .B1(n197), .B2(n40), .ZN(n41) );
  XNOR2_X1 U53 ( .A(n42), .B(n41), .ZN(n61) );
  NOR2_X4 U54 ( .A1(n400), .A2(n401), .ZN(n133) );
  INV_X1 U55 ( .A(n133), .ZN(n33) );
  OR2_X1 U56 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n34) );
  XNOR2_X1 U57 ( .A(n133), .B(n21), .ZN(n38) );
  NOR2_X1 U58 ( .A1(n34), .A2(n18), .ZN(n60) );
  XOR2_X1 U59 ( .A(\mult_x_1/a[6] ), .B(n549), .Z(n35) );
  XNOR2_X1 U60 ( .A(n548), .B(\mult_x_1/a[6] ), .ZN(n36) );
  INV_X1 U61 ( .A(n36), .ZN(n37) );
  INV_X2 U62 ( .A(n37), .ZN(n131) );
  XNOR2_X1 U63 ( .A(n21), .B(\mult_x_1/n286 ), .ZN(n47) );
  OAI22_X1 U64 ( .A1(n130), .A2(n57), .B1(n131), .B2(n47), .ZN(n149) );
  NAND2_X1 U65 ( .A1(n547), .A2(n23), .ZN(n200) );
  XNOR2_X1 U66 ( .A(n547), .B(\mult_x_1/n281 ), .ZN(n114) );
  AND2_X2 U67 ( .A1(n550), .A2(\mult_x_1/n281 ), .ZN(n76) );
  NOR2_X1 U68 ( .A1(n325), .A2(n38), .ZN(n147) );
  XNOR2_X1 U69 ( .A(n21), .B(\mult_x_1/n285 ), .ZN(n46) );
  XNOR2_X1 U70 ( .A(n21), .B(\mult_x_1/n284 ), .ZN(n94) );
  OAI22_X1 U71 ( .A1(n130), .A2(n46), .B1(n131), .B2(n94), .ZN(n99) );
  XNOR2_X1 U72 ( .A(n22), .B(\mult_x_1/n282 ), .ZN(n101) );
  OAI22_X1 U73 ( .A1(n66), .A2(n39), .B1(n15), .B2(n101), .ZN(n98) );
  XNOR2_X1 U74 ( .A(n76), .B(\mult_x_1/n312 ), .ZN(n95) );
  INV_X1 U75 ( .A(n218), .ZN(n97) );
  XNOR2_X1 U76 ( .A(n231), .B(n230), .ZN(n49) );
  OR2_X1 U77 ( .A1(n42), .A2(n41), .ZN(n216) );
  XNOR2_X1 U78 ( .A(n133), .B(\mult_x_1/n286 ), .ZN(n43) );
  NOR2_X1 U79 ( .A1(n43), .A2(n19), .ZN(n215) );
  AOI21_X1 U80 ( .B1(n200), .B2(n23), .A(n44), .ZN(n45) );
  INV_X1 U81 ( .A(n45), .ZN(n52) );
  OAI22_X1 U82 ( .A1(n130), .A2(n47), .B1(n131), .B2(n46), .ZN(n51) );
  XNOR2_X1 U83 ( .A(n133), .B(\mult_x_1/n287 ), .ZN(n48) );
  NOR2_X1 U84 ( .A1(n48), .A2(n18), .ZN(n50) );
  XNOR2_X1 U85 ( .A(n229), .B(n49), .ZN(n184) );
  FA_X1 U86 ( .A(n52), .B(n51), .CI(n50), .CO(n214), .S(n237) );
  XNOR2_X1 U87 ( .A(n22), .B(\mult_x_1/n285 ), .ZN(n113) );
  OAI22_X1 U88 ( .A1(n66), .A2(n113), .B1(n15), .B2(n53), .ZN(n155) );
  XNOR2_X1 U89 ( .A(n16), .B(\mult_x_1/n283 ), .ZN(n116) );
  OAI22_X1 U90 ( .A1(n5), .A2(n116), .B1(n17), .B2(n54), .ZN(n154) );
  INV_X1 U91 ( .A(n21), .ZN(n56) );
  OR2_X1 U92 ( .A1(\mult_x_1/n288 ), .A2(n56), .ZN(n55) );
  OAI22_X1 U93 ( .A1(n130), .A2(n56), .B1(n55), .B2(n131), .ZN(n112) );
  XNOR2_X1 U94 ( .A(n21), .B(\mult_x_1/n288 ), .ZN(n58) );
  OAI22_X1 U95 ( .A1(n130), .A2(n58), .B1(n131), .B2(n57), .ZN(n111) );
  FA_X1 U96 ( .A(n61), .B(n60), .CI(n59), .CO(n231), .S(n235) );
  NAND2_X1 U97 ( .A1(n184), .A2(n183), .ZN(n62) );
  INV_X2 U98 ( .A(n253), .ZN(n73) );
  NAND2_X1 U99 ( .A1(n62), .A2(n10), .ZN(n64) );
  NAND2_X1 U100 ( .A1(n73), .A2(n340), .ZN(n63) );
  NAND2_X1 U101 ( .A1(n64), .A2(n63), .ZN(n376) );
  XNOR2_X1 U124 ( .A(n16), .B(\mult_x_1/n286 ), .ZN(n70) );
  XNOR2_X1 U125 ( .A(n16), .B(\mult_x_1/n285 ), .ZN(n110) );
  OAI22_X1 U126 ( .A1(n5), .A2(n70), .B1(n17), .B2(n110), .ZN(n171) );
  XNOR2_X1 U127 ( .A(n547), .B(\mult_x_1/n284 ), .ZN(n68) );
  XNOR2_X1 U128 ( .A(n7), .B(\mult_x_1/n283 ), .ZN(n109) );
  OAI22_X1 U129 ( .A1(n200), .A2(n68), .B1(n109), .B2(n23), .ZN(n170) );
  OR2_X1 U130 ( .A1(\mult_x_1/n288 ), .A2(n24), .ZN(n65) );
  OAI22_X1 U131 ( .A1(n66), .A2(n24), .B1(n65), .B2(n15), .ZN(n119) );
  XNOR2_X1 U132 ( .A(n22), .B(\mult_x_1/n288 ), .ZN(n67) );
  XNOR2_X1 U133 ( .A(n22), .B(\mult_x_1/n287 ), .ZN(n121) );
  OAI22_X1 U134 ( .A1(n66), .A2(n67), .B1(n15), .B2(n121), .ZN(n118) );
  XNOR2_X1 U135 ( .A(n7), .B(\mult_x_1/n285 ), .ZN(n191) );
  OAI22_X1 U136 ( .A1(n200), .A2(n191), .B1(n68), .B2(n23), .ZN(n188) );
  INV_X1 U137 ( .A(n15), .ZN(n69) );
  AND2_X1 U138 ( .A1(\mult_x_1/n288 ), .A2(n69), .ZN(n187) );
  XNOR2_X1 U139 ( .A(n16), .B(\mult_x_1/n287 ), .ZN(n189) );
  OAI22_X1 U140 ( .A1(n5), .A2(n189), .B1(n17), .B2(n70), .ZN(n186) );
  NOR2_X1 U141 ( .A1(n178), .A2(n177), .ZN(n72) );
  NAND2_X1 U142 ( .A1(n73), .A2(n326), .ZN(n71) );
  OAI21_X1 U143 ( .B1(n73), .B2(n72), .A(n71), .ZN(n348) );
  XNOR2_X1 U144 ( .A(n133), .B(\mult_x_1/n282 ), .ZN(n74) );
  NOR2_X1 U145 ( .A1(n74), .A2(n18), .ZN(n128) );
  XNOR2_X1 U146 ( .A(n21), .B(\mult_x_1/n281 ), .ZN(n75) );
  XNOR2_X1 U147 ( .A(n76), .B(n21), .ZN(n129) );
  OAI22_X1 U148 ( .A1(n130), .A2(n75), .B1(n129), .B2(n131), .ZN(n138) );
  INV_X1 U149 ( .A(n138), .ZN(n127) );
  XNOR2_X1 U150 ( .A(n21), .B(\mult_x_1/n282 ), .ZN(n80) );
  OAI22_X1 U151 ( .A1(n130), .A2(n80), .B1(n131), .B2(n75), .ZN(n85) );
  XNOR2_X1 U152 ( .A(n548), .B(\mult_x_1/n281 ), .ZN(n100) );
  XNOR2_X1 U153 ( .A(n76), .B(n548), .ZN(n78) );
  OAI22_X1 U154 ( .A1(n66), .A2(n100), .B1(n78), .B2(n15), .ZN(n84) );
  AOI21_X1 U155 ( .B1(n15), .B2(n66), .A(n78), .ZN(n77) );
  INV_X1 U156 ( .A(n77), .ZN(n83) );
  OAI22_X1 U157 ( .A1(n66), .A2(n100), .B1(n78), .B2(n15), .ZN(n79) );
  INV_X1 U158 ( .A(n79), .ZN(n92) );
  XNOR2_X1 U159 ( .A(n21), .B(\mult_x_1/n283 ), .ZN(n93) );
  OAI22_X1 U160 ( .A1(n130), .A2(n93), .B1(n131), .B2(n80), .ZN(n91) );
  XNOR2_X1 U161 ( .A(n133), .B(\mult_x_1/n284 ), .ZN(n81) );
  NOR2_X1 U162 ( .A1(n81), .A2(n19), .ZN(n90) );
  XNOR2_X1 U163 ( .A(n133), .B(\mult_x_1/n283 ), .ZN(n82) );
  NOR2_X1 U164 ( .A1(n82), .A2(n19), .ZN(n88) );
  FA_X1 U165 ( .A(n85), .B(n84), .CI(n83), .CO(n126), .S(n87) );
  OR2_X1 U166 ( .A1(n145), .A2(n144), .ZN(n86) );
  MUX2_X1 U167 ( .A(n327), .B(n86), .S(n242), .Z(n350) );
  FA_X1 U168 ( .A(n89), .B(n88), .CI(n87), .CO(n144), .S(n181) );
  FA_X1 U169 ( .A(n92), .B(n91), .CI(n90), .CO(n89), .S(n212) );
  OAI22_X1 U170 ( .A1(n130), .A2(n94), .B1(n131), .B2(n93), .ZN(n219) );
  AOI21_X1 U171 ( .B1(n17), .B2(n5), .A(n95), .ZN(n96) );
  INV_X1 U172 ( .A(n96), .ZN(n217) );
  FA_X1 U173 ( .A(n99), .B(n98), .CI(n97), .CO(n223), .S(n230) );
  OAI22_X1 U174 ( .A1(n66), .A2(n101), .B1(n15), .B2(n100), .ZN(n220) );
  XNOR2_X1 U175 ( .A(n133), .B(\mult_x_1/n285 ), .ZN(n102) );
  NOR2_X1 U176 ( .A1(n102), .A2(n19), .ZN(n221) );
  NAND2_X1 U177 ( .A1(n223), .A2(n105), .ZN(n107) );
  OR2_X1 U178 ( .A1(n180), .A2(n181), .ZN(n108) );
  MUX2_X1 U179 ( .A(n328), .B(n108), .S(n9), .Z(n352) );
  XNOR2_X1 U180 ( .A(n547), .B(\mult_x_1/n282 ), .ZN(n115) );
  OAI22_X1 U181 ( .A1(n200), .A2(n109), .B1(n115), .B2(n23), .ZN(n124) );
  AND2_X1 U182 ( .A1(\mult_x_1/n288 ), .A2(n37), .ZN(n123) );
  XNOR2_X1 U183 ( .A(n16), .B(\mult_x_1/n284 ), .ZN(n117) );
  OAI22_X1 U184 ( .A1(n5), .A2(n110), .B1(n17), .B2(n117), .ZN(n122) );
  HA_X1 U185 ( .A(n112), .B(n111), .CO(n153), .S(n157) );
  XNOR2_X1 U186 ( .A(n22), .B(\mult_x_1/n286 ), .ZN(n120) );
  OAI22_X1 U187 ( .A1(n66), .A2(n120), .B1(n15), .B2(n113), .ZN(n152) );
  OAI22_X1 U188 ( .A1(n200), .A2(n115), .B1(n114), .B2(n23), .ZN(n151) );
  OAI22_X1 U189 ( .A1(n5), .A2(n117), .B1(n17), .B2(n116), .ZN(n150) );
  HA_X1 U190 ( .A(n119), .B(n118), .CO(n168), .S(n169) );
  OAI22_X1 U191 ( .A1(n66), .A2(n121), .B1(n15), .B2(n120), .ZN(n167) );
  FA_X1 U192 ( .A(n124), .B(n123), .CI(n122), .CO(n158), .S(n166) );
  OR2_X1 U193 ( .A1(n164), .A2(n163), .ZN(n125) );
  MUX2_X1 U194 ( .A(n329), .B(n125), .S(n172), .Z(n354) );
  FA_X1 U195 ( .A(n128), .B(n127), .CI(n126), .CO(n140), .S(n145) );
  AOI21_X1 U196 ( .B1(n131), .B2(n130), .A(n129), .ZN(n132) );
  INV_X1 U197 ( .A(n132), .ZN(n136) );
  XNOR2_X1 U198 ( .A(n133), .B(\mult_x_1/n281 ), .ZN(n134) );
  NOR2_X1 U199 ( .A1(n134), .A2(n18), .ZN(n135) );
  XOR2_X1 U200 ( .A(n136), .B(n135), .Z(n137) );
  XOR2_X1 U201 ( .A(n138), .B(n137), .Z(n139) );
  OR2_X1 U202 ( .A1(n140), .A2(n139), .ZN(n142) );
  NAND2_X1 U203 ( .A1(n140), .A2(n139), .ZN(n141) );
  NAND2_X1 U204 ( .A1(n142), .A2(n141), .ZN(n143) );
  MUX2_X1 U205 ( .A(n330), .B(n143), .S(n242), .Z(n356) );
  NAND2_X1 U206 ( .A1(n145), .A2(n144), .ZN(n146) );
  MUX2_X1 U207 ( .A(n331), .B(n146), .S(n9), .Z(n358) );
  FA_X1 U208 ( .A(n147), .B(n148), .CI(n149), .CO(n59), .S(n241) );
  FA_X1 U209 ( .A(n152), .B(n151), .CI(n150), .CO(n240), .S(n156) );
  FA_X1 U210 ( .A(n155), .B(n154), .CI(n153), .CO(n236), .S(n239) );
  FA_X1 U211 ( .A(n158), .B(n157), .CI(n156), .CO(n160), .S(n164) );
  NOR2_X1 U212 ( .A1(n161), .A2(n160), .ZN(n159) );
  MUX2_X1 U213 ( .A(n332), .B(n159), .S(n10), .Z(n360) );
  NAND2_X1 U214 ( .A1(n161), .A2(n160), .ZN(n162) );
  MUX2_X1 U215 ( .A(n333), .B(n162), .S(n172), .Z(n362) );
  NAND2_X1 U216 ( .A1(n164), .A2(n163), .ZN(n165) );
  MUX2_X1 U217 ( .A(n334), .B(n165), .S(n242), .Z(n364) );
  FA_X1 U218 ( .A(n168), .B(n167), .CI(n166), .CO(n163), .S(n175) );
  FA_X1 U219 ( .A(n171), .B(n170), .CI(n169), .CO(n174), .S(n178) );
  NOR2_X1 U220 ( .A1(n175), .A2(n174), .ZN(n173) );
  MUX2_X1 U221 ( .A(n335), .B(n173), .S(n9), .Z(n366) );
  NAND2_X1 U222 ( .A1(n175), .A2(n174), .ZN(n176) );
  MUX2_X1 U223 ( .A(n336), .B(n176), .S(n242), .Z(n368) );
  NAND2_X1 U224 ( .A1(n178), .A2(n177), .ZN(n179) );
  MUX2_X1 U225 ( .A(n337), .B(n179), .S(n9), .Z(n370) );
  NAND2_X1 U226 ( .A1(n181), .A2(n180), .ZN(n182) );
  MUX2_X1 U227 ( .A(n338), .B(n182), .S(n10), .Z(n372) );
  NOR2_X1 U228 ( .A1(n184), .A2(n183), .ZN(n185) );
  MUX2_X1 U229 ( .A(n339), .B(n185), .S(n172), .Z(n374) );
  FA_X1 U230 ( .A(n188), .B(n187), .CI(n186), .CO(n177), .S(n208) );
  XNOR2_X1 U231 ( .A(n16), .B(\mult_x_1/n288 ), .ZN(n190) );
  OAI22_X1 U232 ( .A1(n5), .A2(n190), .B1(n17), .B2(n189), .ZN(n193) );
  XNOR2_X1 U233 ( .A(n7), .B(\mult_x_1/n286 ), .ZN(n196) );
  OAI22_X1 U234 ( .A1(n200), .A2(n196), .B1(n191), .B2(n23), .ZN(n192) );
  NOR2_X1 U235 ( .A1(n208), .A2(n207), .ZN(n244) );
  HA_X1 U236 ( .A(n193), .B(n192), .CO(n207), .S(n205) );
  OR2_X1 U237 ( .A1(\mult_x_1/n288 ), .A2(n25), .ZN(n194) );
  OAI22_X1 U238 ( .A1(n5), .A2(n25), .B1(n194), .B2(n17), .ZN(n204) );
  OR2_X1 U239 ( .A1(n205), .A2(n204), .ZN(n266) );
  XNOR2_X1 U240 ( .A(n7), .B(\mult_x_1/n287 ), .ZN(n199) );
  OAI22_X1 U241 ( .A1(n200), .A2(n199), .B1(n196), .B2(n23), .ZN(n203) );
  INV_X1 U242 ( .A(n17), .ZN(n198) );
  AND2_X1 U243 ( .A1(\mult_x_1/n288 ), .A2(n198), .ZN(n202) );
  NOR2_X1 U244 ( .A1(n203), .A2(n202), .ZN(n259) );
  OAI22_X1 U245 ( .A1(n200), .A2(\mult_x_1/n288 ), .B1(n199), .B2(n23), .ZN(
        n256) );
  OR2_X1 U246 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n201) );
  NAND2_X1 U247 ( .A1(n201), .A2(n200), .ZN(n255) );
  NAND2_X1 U248 ( .A1(n256), .A2(n255), .ZN(n262) );
  NAND2_X1 U249 ( .A1(n203), .A2(n202), .ZN(n260) );
  OAI21_X1 U250 ( .B1(n259), .B2(n262), .A(n260), .ZN(n267) );
  NAND2_X1 U251 ( .A1(n205), .A2(n204), .ZN(n265) );
  INV_X1 U252 ( .A(n265), .ZN(n206) );
  AOI21_X1 U253 ( .B1(n266), .B2(n267), .A(n206), .ZN(n247) );
  NAND2_X1 U254 ( .A1(n208), .A2(n207), .ZN(n246) );
  OAI21_X1 U255 ( .B1(n244), .B2(n247), .A(n246), .ZN(n209) );
  MUX2_X1 U256 ( .A(n341), .B(n209), .S(n242), .Z(n378) );
  FA_X1 U257 ( .A(n212), .B(n211), .CI(n210), .CO(n180), .S(n213) );
  MUX2_X1 U258 ( .A(n342), .B(n213), .S(n9), .Z(n380) );
  FA_X1 U259 ( .A(n216), .B(n215), .CI(n214), .CO(n227), .S(n229) );
  FA_X1 U260 ( .A(n219), .B(n218), .CI(n217), .CO(n211), .S(n226) );
  XNOR2_X1 U261 ( .A(n223), .B(n222), .ZN(n225) );
  MUX2_X1 U262 ( .A(n343), .B(n224), .S(n10), .Z(n382) );
  FA_X1 U263 ( .A(n227), .B(n226), .CI(n225), .CO(n224), .S(n228) );
  MUX2_X1 U264 ( .A(n344), .B(n228), .S(n10), .Z(n384) );
  NAND2_X1 U265 ( .A1(n229), .A2(n27), .ZN(n233) );
  NAND2_X1 U266 ( .A1(n231), .A2(n230), .ZN(n232) );
  MUX2_X1 U267 ( .A(n345), .B(n234), .S(n172), .Z(n386) );
  FA_X1 U268 ( .A(n237), .B(n236), .CI(n235), .CO(n183), .S(n238) );
  MUX2_X1 U269 ( .A(n346), .B(n238), .S(n242), .Z(n388) );
  MUX2_X1 U270 ( .A(n347), .B(n243), .S(n9), .Z(n390) );
  INV_X2 U271 ( .A(rst_n), .ZN(n551) );
  INV_X1 U272 ( .A(n244), .ZN(n245) );
  NAND2_X1 U273 ( .A1(n246), .A2(n245), .ZN(n248) );
  XOR2_X1 U274 ( .A(n248), .B(n247), .Z(n249) );
  NAND2_X1 U275 ( .A1(n249), .A2(n8), .ZN(n252) );
  INV_X1 U276 ( .A(n324), .ZN(n250) );
  NAND2_X1 U277 ( .A1(n250), .A2(n524), .ZN(n251) );
  NAND2_X1 U278 ( .A1(n252), .A2(n251), .ZN(n431) );
  MUX2_X1 U279 ( .A(product[0]), .B(n511), .S(n324), .Z(n403) );
  MUX2_X1 U280 ( .A(n511), .B(n512), .S(n324), .Z(n405) );
  AND2_X1 U281 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n254) );
  MUX2_X1 U282 ( .A(n512), .B(n254), .S(n324), .Z(n407) );
  MUX2_X1 U283 ( .A(product[1]), .B(n514), .S(n324), .Z(n409) );
  MUX2_X1 U284 ( .A(n514), .B(n515), .S(n324), .Z(n411) );
  OR2_X1 U285 ( .A1(n256), .A2(n255), .ZN(n257) );
  AND2_X1 U286 ( .A1(n257), .A2(n262), .ZN(n258) );
  MUX2_X1 U287 ( .A(n515), .B(n258), .S(n324), .Z(n413) );
  MUX2_X1 U288 ( .A(product[2]), .B(n517), .S(n324), .Z(n415) );
  MUX2_X1 U289 ( .A(n517), .B(n518), .S(n324), .Z(n417) );
  INV_X1 U290 ( .A(n259), .ZN(n261) );
  NAND2_X1 U291 ( .A1(n261), .A2(n260), .ZN(n263) );
  XOR2_X1 U292 ( .A(n263), .B(n262), .Z(n264) );
  MUX2_X1 U293 ( .A(n518), .B(n264), .S(n324), .Z(n419) );
  MUX2_X1 U294 ( .A(product[3]), .B(n520), .S(n324), .Z(n421) );
  MUX2_X1 U295 ( .A(n520), .B(n521), .S(n324), .Z(n423) );
  NAND2_X1 U296 ( .A1(n266), .A2(n265), .ZN(n268) );
  XNOR2_X1 U297 ( .A(n268), .B(n267), .ZN(n269) );
  MUX2_X1 U298 ( .A(n521), .B(n269), .S(n324), .Z(n425) );
  MUX2_X1 U299 ( .A(product[4]), .B(n523), .S(n324), .Z(n427) );
  MUX2_X1 U300 ( .A(n523), .B(n524), .S(n324), .Z(n429) );
  MUX2_X1 U301 ( .A(product[5]), .B(n526), .S(n324), .Z(n433) );
  NAND2_X1 U302 ( .A1(n326), .A2(n337), .ZN(n270) );
  XNOR2_X1 U303 ( .A(n270), .B(n341), .ZN(n271) );
  MUX2_X1 U304 ( .A(n526), .B(n271), .S(n324), .Z(n435) );
  MUX2_X1 U305 ( .A(product[6]), .B(n528), .S(n324), .Z(n437) );
  NAND2_X1 U306 ( .A1(n395), .A2(n336), .ZN(n272) );
  AOI21_X1 U307 ( .B1(n326), .B2(n341), .A(n397), .ZN(n274) );
  XOR2_X1 U308 ( .A(n272), .B(n274), .Z(n273) );
  MUX2_X1 U309 ( .A(n528), .B(n273), .S(n324), .Z(n439) );
  MUX2_X1 U310 ( .A(product[7]), .B(n530), .S(n324), .Z(n441) );
  OAI21_X1 U311 ( .B1(n335), .B2(n274), .A(n336), .ZN(n277) );
  NAND2_X1 U312 ( .A1(n329), .A2(n334), .ZN(n275) );
  XNOR2_X1 U313 ( .A(n277), .B(n275), .ZN(n276) );
  MUX2_X1 U314 ( .A(n530), .B(n276), .S(n324), .Z(n443) );
  MUX2_X1 U315 ( .A(product[8]), .B(n532), .S(n324), .Z(n445) );
  AOI21_X1 U316 ( .B1(n277), .B2(n329), .A(n396), .ZN(n280) );
  NAND2_X1 U317 ( .A1(n398), .A2(n333), .ZN(n278) );
  XOR2_X1 U318 ( .A(n280), .B(n278), .Z(n279) );
  MUX2_X1 U319 ( .A(n532), .B(n279), .S(n324), .Z(n447) );
  MUX2_X1 U320 ( .A(product[9]), .B(n534), .S(n324), .Z(n449) );
  OAI21_X1 U321 ( .B1(n280), .B2(n332), .A(n333), .ZN(n291) );
  INV_X1 U322 ( .A(n291), .ZN(n284) );
  NOR2_X1 U323 ( .A1(n346), .A2(n347), .ZN(n288) );
  INV_X1 U324 ( .A(n288), .ZN(n281) );
  NAND2_X1 U325 ( .A1(n346), .A2(n347), .ZN(n289) );
  NAND2_X1 U326 ( .A1(n281), .A2(n289), .ZN(n282) );
  XOR2_X1 U327 ( .A(n284), .B(n282), .Z(n283) );
  MUX2_X1 U328 ( .A(n534), .B(n283), .S(n324), .Z(n451) );
  MUX2_X1 U329 ( .A(product[10]), .B(n536), .S(n324), .Z(n453) );
  OAI21_X1 U330 ( .B1(n284), .B2(n288), .A(n289), .ZN(n286) );
  NAND2_X1 U331 ( .A1(n392), .A2(n340), .ZN(n285) );
  XNOR2_X1 U332 ( .A(n286), .B(n285), .ZN(n287) );
  MUX2_X1 U333 ( .A(n536), .B(n287), .S(n324), .Z(n455) );
  MUX2_X1 U334 ( .A(product[11]), .B(n538), .S(n324), .Z(n457) );
  NOR2_X1 U335 ( .A1(n339), .A2(n288), .ZN(n292) );
  OAI21_X1 U336 ( .B1(n339), .B2(n289), .A(n340), .ZN(n290) );
  AOI21_X1 U337 ( .B1(n292), .B2(n291), .A(n290), .ZN(n321) );
  NOR2_X1 U338 ( .A1(n344), .A2(n345), .ZN(n307) );
  INV_X1 U339 ( .A(n307), .ZN(n298) );
  NAND2_X1 U340 ( .A1(n344), .A2(n345), .ZN(n310) );
  NAND2_X1 U341 ( .A1(n298), .A2(n310), .ZN(n293) );
  XOR2_X1 U342 ( .A(n321), .B(n293), .Z(n294) );
  MUX2_X1 U343 ( .A(n538), .B(n294), .S(n324), .Z(n459) );
  MUX2_X1 U344 ( .A(product[12]), .B(n540), .S(n324), .Z(n461) );
  OAI21_X1 U345 ( .B1(n321), .B2(n307), .A(n310), .ZN(n296) );
  OR2_X1 U346 ( .A1(n342), .A2(n343), .ZN(n306) );
  NAND2_X1 U347 ( .A1(n342), .A2(n343), .ZN(n299) );
  NAND2_X1 U348 ( .A1(n306), .A2(n299), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  MUX2_X1 U350 ( .A(n540), .B(n297), .S(n324), .Z(n463) );
  MUX2_X1 U351 ( .A(product[13]), .B(n542), .S(n324), .Z(n465) );
  NAND2_X1 U352 ( .A1(n298), .A2(n306), .ZN(n302) );
  INV_X1 U353 ( .A(n310), .ZN(n300) );
  INV_X1 U354 ( .A(n299), .ZN(n308) );
  AOI21_X1 U355 ( .B1(n300), .B2(n306), .A(n308), .ZN(n301) );
  OAI21_X1 U356 ( .B1(n321), .B2(n302), .A(n301), .ZN(n304) );
  NAND2_X1 U357 ( .A1(n328), .A2(n338), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  MUX2_X1 U359 ( .A(n542), .B(n305), .S(n10), .Z(n467) );
  MUX2_X1 U360 ( .A(product[14]), .B(n544), .S(n324), .Z(n469) );
  NAND2_X1 U361 ( .A1(n306), .A2(n328), .ZN(n311) );
  NOR2_X1 U362 ( .A1(n307), .A2(n311), .ZN(n317) );
  INV_X1 U363 ( .A(n317), .ZN(n313) );
  AOI21_X1 U364 ( .B1(n308), .B2(n328), .A(n393), .ZN(n309) );
  OAI21_X1 U365 ( .B1(n311), .B2(n310), .A(n309), .ZN(n318) );
  INV_X1 U366 ( .A(n318), .ZN(n312) );
  OAI21_X1 U367 ( .B1(n321), .B2(n313), .A(n312), .ZN(n315) );
  NAND2_X1 U368 ( .A1(n327), .A2(n331), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U370 ( .A(n544), .B(n316), .S(n172), .Z(n471) );
  MUX2_X1 U371 ( .A(product[15]), .B(n546), .S(en), .Z(n473) );
  NAND2_X1 U372 ( .A1(n317), .A2(n327), .ZN(n320) );
  AOI21_X1 U373 ( .B1(n318), .B2(n327), .A(n394), .ZN(n319) );
  OAI21_X1 U374 ( .B1(n321), .B2(n320), .A(n319), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(n330), .ZN(n323) );
  MUX2_X1 U376 ( .A(n546), .B(n323), .S(n324), .Z(n475) );
  MUX2_X1 U377 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n324), .Z(n477) );
  MUX2_X1 U378 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n324), .Z(n479) );
  MUX2_X1 U379 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n324), .Z(n481) );
  MUX2_X1 U380 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n324), .Z(n483) );
  MUX2_X1 U381 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n324), .Z(n485) );
  MUX2_X1 U382 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n324), .Z(n487) );
  MUX2_X1 U383 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n324), .Z(n489) );
  MUX2_X1 U384 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n324), .Z(n491) );
  MUX2_X1 U385 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n324), .Z(n493) );
  MUX2_X1 U386 ( .A(n7), .B(A_extended[1]), .S(n324), .Z(n495) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n324), .Z(n497) );
  MUX2_X1 U388 ( .A(n16), .B(A_extended[3]), .S(n8), .Z(n499) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n324), .Z(n501) );
  MUX2_X1 U390 ( .A(n22), .B(A_extended[5]), .S(n8), .Z(n503) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n8), .Z(n505) );
  MUX2_X1 U392 ( .A(n21), .B(A_extended[7]), .S(n324), .Z(n507) );
  OR2_X1 U393 ( .A1(n8), .A2(n550), .ZN(n509) );
endmodule


module conv_128_32_DW_mult_pipe_J1_20 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n368, n370, n372, n374,
         n376, n378, n380, n382, n384, n386, n388, n390, n392, n394, n396,
         n398, n400, n402, n404, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n419, n421, n423, n425, n427, n429,
         n431, n433, n435, n437, n439, n441, n443, n445, n447, n449, n451,
         n453, n455, n457, n459, n461, n463, n465, n467, n469, n471, n473,
         n475, n477, n479, n481, n483, n485, n487, n489, n491, n493, n495,
         n497, n499, n501, n503, n505, n507, n509, n511, n513, n515, n517,
         n519, n521, n523, n525, n527, n529, n530, n532, n533, n535, n536,
         n538, n539, n541, n542, n544, n545, n547, n549, n551, n553, n555,
         n557, n559, n561, n563, n565, n566, n567, n568;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n415), .SE(n527), .CK(clk), .Q(n567), 
        .QN(n28) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n415), .SE(n523), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n35) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n415), .SE(n519), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n34) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n415), .SE(n515), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n18) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n415), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n29) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n415), .SE(n509), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n20) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n415), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n27) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n416), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n26) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n417), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n25) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n415), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n24) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n415), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n22) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n415), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n23) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n415), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n415), .SE(n493), .CK(clk), .Q(n565)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n415), .SE(n491), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n415), .SE(n489), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n415), .SE(n487), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n415), .SE(n485), .CK(clk), .Q(n561)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n417), .SE(n483), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n416), .SE(n481), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n415), .SE(n479), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG18_S3 ( .D(1'b0), .SI(n415), .SE(n477), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG19_S4 ( .D(1'b0), .SI(n415), .SE(n475), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n415), .SE(n473), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n415), .SE(n471), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n415), .SE(n469), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n415), .SE(n467), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n415), .SE(n465), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n415), .SE(n463), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n417), .SE(n461), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n417), .SE(n459), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n417), .SE(n457), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n417), .SE(n455), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n417), .SE(n453), .CK(clk), .Q(n545), 
        .QN(n40) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n417), .SE(n451), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n417), .SE(n449), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n417), .SE(n447), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n417), .SE(n445), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n417), .SE(n443), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n417), .SE(n441), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n416), .SE(n439), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n416), .SE(n437), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n416), .SE(n435), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n416), .SE(n433), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n416), .SE(n431), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n416), .SE(n429), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n416), .SE(n427), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n416), .SE(n425), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n416), .SE(n423), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n416), .SE(n421), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n416), .SE(n419), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n415), .SE(n517), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n21) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n568), .SI(1'b1), .SE(n404), .CK(clk), 
        .Q(n365) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n568), .SI(1'b1), .SE(n402), .CK(clk), 
        .Q(n364) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n568), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n363) );
  SDFF_X1 \mult_x_1/clk_r_REG13_S2  ( .D(n568), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n362), .QN(n412) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n568), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n361), .QN(n39) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n568), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n360), .QN(n414) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n568), .SE(n392), .CK(
        clk), .Q(n413), .QN(n359) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n568), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n358), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n568), .SI(1'b1), .SE(n388), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n568), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n356), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n568), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n355), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n568), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n568), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n353), .QN(n411) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n568), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n352), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n568), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n351), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n568), .SE(n374), .CK(
        clk), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n568), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n349), .QN(n36) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n568), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n348), .QN(n38) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n568), .SE(n368), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n568), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n346) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n415), .SE(n521), .CK(clk), .Q(n566), 
        .QN(n31) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n415), .SE(n525), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n30) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n415), .SE(n513), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n33) );
  INV_X2 U2 ( .A(n53), .ZN(n213) );
  XNOR2_X1 U3 ( .A(n227), .B(n5), .ZN(n235) );
  XNOR2_X1 U4 ( .A(n229), .B(n228), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n43), .A2(n12), .ZN(n193) );
  INV_X2 U6 ( .A(n568), .ZN(n415) );
  BUF_X1 U7 ( .A(n67), .Z(n7) );
  INV_X1 U8 ( .A(n301), .ZN(n6) );
  BUF_X1 U9 ( .A(n415), .Z(n416) );
  BUF_X1 U10 ( .A(n415), .Z(n417) );
  INV_X1 U11 ( .A(rst_n), .ZN(n568) );
  OR2_X1 U12 ( .A1(n139), .A2(n140), .ZN(n145) );
  BUF_X1 U13 ( .A(\mult_x_1/n312 ), .Z(n344) );
  NOR2_X1 U14 ( .A1(n254), .A2(n255), .ZN(n256) );
  XNOR2_X1 U15 ( .A(n133), .B(n134), .ZN(n254) );
  NAND2_X1 U16 ( .A1(n9), .A2(n8), .ZN(n382) );
  NAND2_X1 U17 ( .A1(n6), .A2(n354), .ZN(n8) );
  NAND2_X1 U18 ( .A1(n10), .A2(n301), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n235), .A2(n234), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n257), .A2(n37), .ZN(n258) );
  XNOR2_X1 U21 ( .A(n81), .B(n11), .ZN(n37) );
  INV_X1 U22 ( .A(n90), .ZN(n11) );
  NAND2_X1 U23 ( .A1(n268), .A2(n267), .ZN(n269) );
  INV_X1 U24 ( .A(n272), .ZN(n268) );
  INV_X1 U25 ( .A(n271), .ZN(n267) );
  OAI22_X1 U26 ( .A1(n203), .A2(n60), .B1(n7), .B2(n65), .ZN(n78) );
  OAI21_X1 U27 ( .B1(n7), .B2(n59), .A(n42), .ZN(n139) );
  INV_X1 U28 ( .A(n154), .ZN(n41) );
  OAI22_X1 U29 ( .A1(n203), .A2(n99), .B1(n7), .B2(n202), .ZN(n199) );
  OAI22_X1 U30 ( .A1(n203), .A2(n31), .B1(n7), .B2(n98), .ZN(n200) );
  OAI22_X1 U31 ( .A1(n203), .A2(n59), .B1(n7), .B2(n60), .ZN(n142) );
  OAI22_X1 U32 ( .A1(n203), .A2(n166), .B1(n7), .B2(n154), .ZN(n171) );
  OAI21_X1 U33 ( .B1(n88), .B2(n7), .A(n69), .ZN(n182) );
  INV_X1 U34 ( .A(n65), .ZN(n66) );
  XNOR2_X1 U35 ( .A(n200), .B(n199), .ZN(n246) );
  NAND2_X1 U36 ( .A1(n78), .A2(n77), .ZN(n79) );
  OR2_X1 U37 ( .A1(n78), .A2(n77), .ZN(n75) );
  NAND2_X1 U38 ( .A1(n145), .A2(n144), .ZN(n50) );
  XNOR2_X1 U39 ( .A(n76), .B(n61), .ZN(n134) );
  XNOR2_X1 U40 ( .A(n78), .B(n77), .ZN(n61) );
  OAI22_X1 U41 ( .A1(n203), .A2(n201), .B1(n7), .B2(n166), .ZN(n198) );
  XNOR2_X1 U42 ( .A(n246), .B(n101), .ZN(n106) );
  XNOR2_X1 U43 ( .A(n243), .B(n100), .ZN(n101) );
  INV_X1 U44 ( .A(n242), .ZN(n100) );
  OAI22_X1 U45 ( .A1(n203), .A2(n202), .B1(n7), .B2(n201), .ZN(n240) );
  OAI21_X1 U46 ( .B1(n246), .B2(n245), .A(n244), .ZN(n248) );
  NAND2_X1 U47 ( .A1(n243), .A2(n242), .ZN(n244) );
  NOR2_X1 U48 ( .A1(n243), .A2(n242), .ZN(n245) );
  XNOR2_X1 U49 ( .A(n147), .B(n146), .ZN(n264) );
  XNOR2_X1 U50 ( .A(n145), .B(n144), .ZN(n146) );
  NAND2_X1 U51 ( .A1(n97), .A2(n96), .ZN(n370) );
  OR2_X1 U52 ( .A1(n301), .A2(n38), .ZN(n96) );
  OAI21_X1 U53 ( .B1(n252), .B2(n251), .A(n301), .ZN(n97) );
  NAND2_X1 U54 ( .A1(n274), .A2(n273), .ZN(n275) );
  NAND2_X1 U55 ( .A1(n272), .A2(n271), .ZN(n273) );
  NAND2_X1 U56 ( .A1(n270), .A2(n269), .ZN(n274) );
  NAND2_X1 U57 ( .A1(n67), .A2(n68), .ZN(n203) );
  XNOR2_X1 U58 ( .A(n33), .B(n18), .ZN(n12) );
  NAND2_X1 U59 ( .A1(n227), .A2(n229), .ZN(n14) );
  NAND2_X1 U60 ( .A1(n227), .A2(n228), .ZN(n15) );
  NAND2_X1 U61 ( .A1(n229), .A2(n228), .ZN(n16) );
  NAND3_X1 U62 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n175) );
  INV_X1 U63 ( .A(n175), .ZN(n172) );
  INV_X1 U64 ( .A(n30), .ZN(n17) );
  XNOR2_X1 U65 ( .A(n33), .B(n18), .ZN(n44) );
  INV_X1 U66 ( .A(n31), .ZN(n19) );
  NAND2_X1 U67 ( .A1(n48), .A2(n52), .ZN(n212) );
  XNOR2_X1 U68 ( .A(n566), .B(n34), .ZN(n68) );
  AND2_X1 U69 ( .A1(n152), .A2(n151), .ZN(n32) );
  XNOR2_X1 U70 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n67) );
  XNOR2_X1 U71 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n59) );
  XNOR2_X1 U72 ( .A(n566), .B(\mult_x_1/n284 ), .ZN(n154) );
  NAND3_X1 U73 ( .A1(n68), .A2(n67), .A3(n41), .ZN(n42) );
  XOR2_X1 U74 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n43) );
  XNOR2_X1 U75 ( .A(n344), .B(\mult_x_1/n282 ), .ZN(n155) );
  INV_X1 U76 ( .A(n44), .ZN(n117) );
  XNOR2_X1 U77 ( .A(n344), .B(\mult_x_1/n281 ), .ZN(n55) );
  OAI22_X1 U78 ( .A1(n193), .A2(n155), .B1(n44), .B2(n55), .ZN(n140) );
  INV_X1 U79 ( .A(n145), .ZN(n46) );
  NAND2_X1 U80 ( .A1(n28), .A2(\mult_x_1/n310 ), .ZN(n137) );
  NOR2_X1 U81 ( .A1(n22), .A2(n137), .ZN(n144) );
  INV_X1 U82 ( .A(n144), .ZN(n45) );
  NAND2_X1 U83 ( .A1(n46), .A2(n45), .ZN(n49) );
  NAND2_X1 U84 ( .A1(\mult_x_1/n313 ), .A2(n29), .ZN(n190) );
  AND2_X1 U85 ( .A1(n567), .A2(\mult_x_1/n281 ), .ZN(n179) );
  XNOR2_X1 U86 ( .A(n179), .B(\mult_x_1/n313 ), .ZN(n136) );
  AOI21_X1 U87 ( .B1(n190), .B2(n29), .A(n136), .ZN(n47) );
  INV_X1 U88 ( .A(n47), .ZN(n161) );
  XNOR2_X1 U89 ( .A(\mult_x_1/a[6] ), .B(n566), .ZN(n52) );
  XNOR2_X1 U90 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n58) );
  XNOR2_X1 U91 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n135) );
  XNOR2_X1 U92 ( .A(n35), .B(\mult_x_1/n310 ), .ZN(n48) );
  OAI22_X1 U93 ( .A1(n52), .A2(n58), .B1(n135), .B2(n212), .ZN(n160) );
  NOR2_X1 U94 ( .A1(n23), .A2(n137), .ZN(n159) );
  NAND2_X1 U95 ( .A1(n49), .A2(n147), .ZN(n51) );
  NAND2_X1 U96 ( .A1(n51), .A2(n50), .ZN(n132) );
  XNOR2_X1 U97 ( .A(n17), .B(\mult_x_1/n284 ), .ZN(n57) );
  INV_X1 U98 ( .A(n52), .ZN(n53) );
  XNOR2_X1 U99 ( .A(n17), .B(\mult_x_1/n283 ), .ZN(n70) );
  OAI22_X1 U100 ( .A1(n212), .A2(n57), .B1(n213), .B2(n70), .ZN(n73) );
  XNOR2_X1 U101 ( .A(n179), .B(n344), .ZN(n56) );
  AOI21_X1 U102 ( .B1(n193), .B2(n44), .A(n56), .ZN(n54) );
  INV_X1 U103 ( .A(n54), .ZN(n72) );
  OAI22_X1 U104 ( .A1(n44), .A2(n56), .B1(n193), .B2(n55), .ZN(n71) );
  OR2_X1 U105 ( .A1(n132), .A2(n131), .ZN(n62) );
  OAI22_X1 U106 ( .A1(n212), .A2(n58), .B1(n213), .B2(n57), .ZN(n143) );
  XNOR2_X1 U107 ( .A(n19), .B(\mult_x_1/n282 ), .ZN(n60) );
  INV_X1 U108 ( .A(n71), .ZN(n141) );
  XNOR2_X1 U109 ( .A(n566), .B(\mult_x_1/n281 ), .ZN(n65) );
  NOR2_X1 U110 ( .A1(n24), .A2(n137), .ZN(n77) );
  NAND2_X1 U111 ( .A1(n62), .A2(n134), .ZN(n64) );
  NAND2_X1 U112 ( .A1(n132), .A2(n131), .ZN(n63) );
  NAND2_X1 U113 ( .A1(n64), .A2(n63), .ZN(n257) );
  XNOR2_X1 U114 ( .A(n179), .B(n19), .ZN(n88) );
  NAND3_X1 U115 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n69) );
  INV_X1 U116 ( .A(n182), .ZN(n86) );
  XNOR2_X1 U117 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n87) );
  OAI22_X1 U118 ( .A1(n212), .A2(n70), .B1(n213), .B2(n87), .ZN(n85) );
  NOR2_X1 U119 ( .A1(n25), .A2(n137), .ZN(n84) );
  FA_X1 U120 ( .A(n73), .B(n72), .CI(n71), .CO(n91), .S(n131) );
  INV_X1 U121 ( .A(n91), .ZN(n74) );
  XNOR2_X1 U122 ( .A(n92), .B(n74), .ZN(n81) );
  NAND2_X1 U123 ( .A1(n76), .A2(n75), .ZN(n80) );
  NAND2_X1 U124 ( .A1(n80), .A2(n79), .ZN(n90) );
  BUF_X4 U125 ( .A(en), .Z(n301) );
  OAI21_X1 U126 ( .B1(n257), .B2(n37), .A(n301), .ZN(n83) );
  OR2_X1 U127 ( .A1(n301), .A2(n36), .ZN(n82) );
  NAND2_X1 U128 ( .A1(n83), .A2(n82), .ZN(n372) );
  FA_X1 U129 ( .A(n86), .B(n85), .CI(n84), .CO(n186), .S(n92) );
  NOR2_X1 U130 ( .A1(n26), .A2(n137), .ZN(n185) );
  XNOR2_X1 U131 ( .A(n17), .B(\mult_x_1/n281 ), .ZN(n180) );
  OAI22_X1 U132 ( .A1(n212), .A2(n87), .B1(n213), .B2(n180), .ZN(n183) );
  AOI21_X1 U133 ( .B1(n7), .B2(n203), .A(n88), .ZN(n89) );
  INV_X1 U134 ( .A(n89), .ZN(n181) );
  NAND2_X1 U135 ( .A1(n90), .A2(n92), .ZN(n95) );
  NAND2_X1 U136 ( .A1(n90), .A2(n91), .ZN(n94) );
  NAND2_X1 U137 ( .A1(n92), .A2(n91), .ZN(n93) );
  NAND3_X1 U138 ( .A1(n95), .A2(n94), .A3(n93), .ZN(n251) );
  OR2_X1 U139 ( .A1(\mult_x_1/n288 ), .A2(n31), .ZN(n98) );
  XNOR2_X1 U140 ( .A(n19), .B(\mult_x_1/n288 ), .ZN(n99) );
  XNOR2_X1 U141 ( .A(n19), .B(\mult_x_1/n287 ), .ZN(n202) );
  XNOR2_X1 U142 ( .A(n344), .B(\mult_x_1/n286 ), .ZN(n104) );
  XNOR2_X1 U143 ( .A(n344), .B(\mult_x_1/n285 ), .ZN(n192) );
  OAI22_X1 U144 ( .A1(n193), .A2(n104), .B1(n44), .B2(n192), .ZN(n243) );
  XNOR2_X1 U145 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n102) );
  XNOR2_X1 U146 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n189) );
  OAI22_X1 U147 ( .A1(n190), .A2(n102), .B1(n189), .B2(n29), .ZN(n242) );
  XNOR2_X1 U148 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n112) );
  OAI22_X1 U149 ( .A1(n190), .A2(n112), .B1(n102), .B2(n29), .ZN(n109) );
  INV_X1 U150 ( .A(n7), .ZN(n103) );
  AND2_X1 U151 ( .A1(\mult_x_1/n288 ), .A2(n103), .ZN(n108) );
  XNOR2_X1 U152 ( .A(n344), .B(\mult_x_1/n287 ), .ZN(n110) );
  OAI22_X1 U153 ( .A1(n193), .A2(n110), .B1(n44), .B2(n104), .ZN(n107) );
  OR2_X1 U154 ( .A1(n106), .A2(n105), .ZN(n262) );
  NAND2_X1 U155 ( .A1(n106), .A2(n105), .ZN(n259) );
  NAND2_X1 U156 ( .A1(n262), .A2(n259), .ZN(n128) );
  FA_X1 U157 ( .A(n109), .B(n108), .CI(n107), .CO(n105), .S(n126) );
  XNOR2_X1 U158 ( .A(n344), .B(\mult_x_1/n288 ), .ZN(n111) );
  OAI22_X1 U159 ( .A1(n193), .A2(n111), .B1(n44), .B2(n110), .ZN(n114) );
  XNOR2_X1 U160 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n116) );
  OAI22_X1 U161 ( .A1(n190), .A2(n116), .B1(n112), .B2(n29), .ZN(n113) );
  NOR2_X1 U162 ( .A1(n126), .A2(n125), .ZN(n292) );
  HA_X1 U163 ( .A(n114), .B(n113), .CO(n125), .S(n123) );
  OR2_X1 U164 ( .A1(\mult_x_1/n288 ), .A2(n21), .ZN(n115) );
  OAI22_X1 U165 ( .A1(n193), .A2(n21), .B1(n115), .B2(n44), .ZN(n122) );
  OR2_X1 U166 ( .A1(n123), .A2(n122), .ZN(n288) );
  XNOR2_X1 U167 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n118) );
  OAI22_X1 U168 ( .A1(n190), .A2(n118), .B1(n116), .B2(n29), .ZN(n121) );
  AND2_X1 U169 ( .A1(n117), .A2(\mult_x_1/n288 ), .ZN(n120) );
  NOR2_X1 U170 ( .A1(n121), .A2(n120), .ZN(n281) );
  OAI22_X1 U171 ( .A1(n190), .A2(\mult_x_1/n288 ), .B1(n118), .B2(n29), .ZN(
        n278) );
  OR2_X1 U172 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n119) );
  NAND2_X1 U173 ( .A1(n119), .A2(n190), .ZN(n277) );
  NAND2_X1 U174 ( .A1(n278), .A2(n277), .ZN(n284) );
  NAND2_X1 U175 ( .A1(n121), .A2(n120), .ZN(n282) );
  OAI21_X1 U176 ( .B1(n281), .B2(n284), .A(n282), .ZN(n289) );
  NAND2_X1 U177 ( .A1(n123), .A2(n122), .ZN(n287) );
  INV_X1 U178 ( .A(n287), .ZN(n124) );
  AOI21_X1 U179 ( .B1(n288), .B2(n289), .A(n124), .ZN(n295) );
  NAND2_X1 U180 ( .A1(n126), .A2(n125), .ZN(n293) );
  OAI21_X1 U181 ( .B1(n292), .B2(n295), .A(n293), .ZN(n261) );
  INV_X1 U182 ( .A(n261), .ZN(n127) );
  XNOR2_X1 U183 ( .A(n128), .B(n127), .ZN(n130) );
  OR2_X1 U184 ( .A1(n301), .A2(n40), .ZN(n129) );
  OAI21_X1 U185 ( .B1(n130), .B2(n6), .A(n129), .ZN(n453) );
  XNOR2_X1 U186 ( .A(n132), .B(n131), .ZN(n133) );
  XNOR2_X1 U187 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n157) );
  OAI22_X1 U188 ( .A1(n212), .A2(n157), .B1(n213), .B2(n135), .ZN(n165) );
  XNOR2_X1 U189 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n167) );
  OAI22_X1 U190 ( .A1(n190), .A2(n167), .B1(n136), .B2(n29), .ZN(n164) );
  INV_X1 U191 ( .A(n137), .ZN(n138) );
  AND2_X1 U192 ( .A1(\mult_x_1/n288 ), .A2(n138), .ZN(n163) );
  XNOR2_X1 U193 ( .A(n140), .B(n139), .ZN(n151) );
  FA_X1 U194 ( .A(n143), .B(n142), .CI(n141), .CO(n76), .S(n265) );
  NAND2_X1 U195 ( .A1(n254), .A2(n255), .ZN(n148) );
  NAND2_X1 U196 ( .A1(n148), .A2(n301), .ZN(n150) );
  OR2_X1 U197 ( .A1(n301), .A2(n408), .ZN(n149) );
  NAND2_X1 U198 ( .A1(n150), .A2(n149), .ZN(n378) );
  INV_X1 U199 ( .A(n151), .ZN(n153) );
  XNOR2_X1 U200 ( .A(n153), .B(n152), .ZN(n270) );
  XNOR2_X1 U201 ( .A(n19), .B(\mult_x_1/n285 ), .ZN(n166) );
  XNOR2_X1 U202 ( .A(n344), .B(\mult_x_1/n283 ), .ZN(n168) );
  OAI22_X1 U203 ( .A1(n193), .A2(n168), .B1(n44), .B2(n155), .ZN(n170) );
  OR2_X1 U204 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n156) );
  OAI22_X1 U205 ( .A1(n212), .A2(n30), .B1(n156), .B2(n213), .ZN(n195) );
  XNOR2_X1 U206 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n158) );
  OAI22_X1 U207 ( .A1(n212), .A2(n158), .B1(n213), .B2(n157), .ZN(n194) );
  FA_X1 U208 ( .A(n161), .B(n160), .CI(n159), .CO(n147), .S(n272) );
  XNOR2_X1 U209 ( .A(n271), .B(n272), .ZN(n162) );
  XNOR2_X1 U210 ( .A(n270), .B(n162), .ZN(n174) );
  FA_X1 U211 ( .A(n163), .B(n164), .CI(n165), .CO(n152), .S(n229) );
  XNOR2_X1 U212 ( .A(n19), .B(\mult_x_1/n286 ), .ZN(n201) );
  XNOR2_X1 U213 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n188) );
  OAI22_X1 U214 ( .A1(n190), .A2(n188), .B1(n167), .B2(n29), .ZN(n197) );
  XNOR2_X1 U215 ( .A(n344), .B(\mult_x_1/n284 ), .ZN(n191) );
  OAI22_X1 U216 ( .A1(n193), .A2(n191), .B1(n44), .B2(n168), .ZN(n196) );
  FA_X1 U217 ( .A(n171), .B(n170), .CI(n169), .CO(n271), .S(n227) );
  NAND2_X1 U218 ( .A1(n301), .A2(n172), .ZN(n173) );
  OAI22_X1 U219 ( .A1(n174), .A2(n173), .B1(n345), .B2(n412), .ZN(n398) );
  NAND2_X1 U220 ( .A1(n175), .A2(n174), .ZN(n176) );
  NAND2_X1 U221 ( .A1(n301), .A2(n176), .ZN(n178) );
  OR2_X1 U222 ( .A1(n301), .A2(n39), .ZN(n177) );
  NAND2_X1 U223 ( .A1(n178), .A2(n177), .ZN(n396) );
  NOR2_X1 U244 ( .A1(n27), .A2(n137), .ZN(n210) );
  XNOR2_X1 U245 ( .A(n179), .B(n17), .ZN(n211) );
  OAI22_X1 U246 ( .A1(n212), .A2(n180), .B1(n211), .B2(n213), .ZN(n218) );
  INV_X1 U247 ( .A(n218), .ZN(n209) );
  FA_X1 U248 ( .A(n183), .B(n181), .CI(n182), .CO(n208), .S(n184) );
  FA_X1 U249 ( .A(n186), .B(n185), .CI(n184), .CO(n224), .S(n252) );
  OR2_X1 U250 ( .A1(n225), .A2(n224), .ZN(n187) );
  MUX2_X1 U251 ( .A(n346), .B(n187), .S(n301), .Z(n366) );
  OAI22_X1 U252 ( .A1(n190), .A2(n189), .B1(n188), .B2(n29), .ZN(n206) );
  AND2_X1 U253 ( .A1(\mult_x_1/n288 ), .A2(n53), .ZN(n205) );
  OAI22_X1 U254 ( .A1(n193), .A2(n192), .B1(n44), .B2(n191), .ZN(n204) );
  HA_X1 U255 ( .A(n194), .B(n195), .CO(n169), .S(n231) );
  FA_X1 U256 ( .A(n198), .B(n197), .CI(n196), .CO(n228), .S(n230) );
  AND2_X1 U257 ( .A1(n200), .A2(n199), .ZN(n241) );
  FA_X1 U258 ( .A(n206), .B(n205), .CI(n204), .CO(n232), .S(n239) );
  OR2_X1 U259 ( .A1(n237), .A2(n236), .ZN(n207) );
  MUX2_X1 U260 ( .A(n347), .B(n207), .S(n301), .Z(n368) );
  FA_X1 U261 ( .A(n210), .B(n209), .CI(n208), .CO(n220), .S(n225) );
  AOI21_X1 U262 ( .B1(n213), .B2(n212), .A(n211), .ZN(n214) );
  INV_X1 U263 ( .A(n214), .ZN(n216) );
  NOR2_X1 U264 ( .A1(n20), .A2(n137), .ZN(n215) );
  XOR2_X1 U265 ( .A(n216), .B(n215), .Z(n217) );
  XOR2_X1 U266 ( .A(n218), .B(n217), .Z(n219) );
  OR2_X1 U267 ( .A1(n220), .A2(n219), .ZN(n222) );
  NAND2_X1 U268 ( .A1(n220), .A2(n219), .ZN(n221) );
  NAND2_X1 U269 ( .A1(n222), .A2(n221), .ZN(n223) );
  MUX2_X1 U270 ( .A(n350), .B(n223), .S(n301), .Z(n374) );
  NAND2_X1 U271 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U272 ( .A(n351), .B(n226), .S(n301), .Z(n376) );
  FA_X1 U273 ( .A(n232), .B(n231), .CI(n230), .CO(n234), .S(n237) );
  NOR2_X1 U274 ( .A1(n235), .A2(n234), .ZN(n233) );
  MUX2_X1 U275 ( .A(n353), .B(n233), .S(n301), .Z(n380) );
  NAND2_X1 U276 ( .A1(n237), .A2(n236), .ZN(n238) );
  MUX2_X1 U277 ( .A(n355), .B(n238), .S(n301), .Z(n384) );
  FA_X1 U278 ( .A(n241), .B(n240), .CI(n239), .CO(n236), .S(n249) );
  NOR2_X1 U279 ( .A1(n249), .A2(n248), .ZN(n247) );
  MUX2_X1 U280 ( .A(n356), .B(n247), .S(n301), .Z(n386) );
  NAND2_X1 U281 ( .A1(n249), .A2(n248), .ZN(n250) );
  MUX2_X1 U282 ( .A(n357), .B(n250), .S(n301), .Z(n388) );
  NAND2_X1 U283 ( .A1(n252), .A2(n251), .ZN(n253) );
  MUX2_X1 U284 ( .A(n358), .B(n253), .S(n301), .Z(n390) );
  MUX2_X1 U285 ( .A(n359), .B(n256), .S(n301), .Z(n392) );
  MUX2_X1 U286 ( .A(n360), .B(n258), .S(n301), .Z(n394) );
  INV_X1 U287 ( .A(n259), .ZN(n260) );
  AOI21_X1 U288 ( .B1(n262), .B2(n261), .A(n260), .ZN(n263) );
  MUX2_X1 U289 ( .A(n363), .B(n263), .S(n301), .Z(n400) );
  FA_X1 U290 ( .A(n32), .B(n265), .CI(n264), .CO(n255), .S(n266) );
  MUX2_X1 U291 ( .A(n364), .B(n266), .S(n301), .Z(n402) );
  MUX2_X1 U292 ( .A(n365), .B(n275), .S(n301), .Z(n404) );
  MUX2_X1 U293 ( .A(product[0]), .B(n529), .S(n301), .Z(n419) );
  MUX2_X1 U294 ( .A(n529), .B(n530), .S(n301), .Z(n421) );
  AND2_X1 U295 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n276) );
  MUX2_X1 U296 ( .A(n530), .B(n276), .S(n301), .Z(n423) );
  MUX2_X1 U297 ( .A(product[1]), .B(n532), .S(n301), .Z(n425) );
  MUX2_X1 U298 ( .A(n532), .B(n533), .S(n301), .Z(n427) );
  OR2_X1 U299 ( .A1(n278), .A2(n277), .ZN(n279) );
  AND2_X1 U300 ( .A1(n279), .A2(n284), .ZN(n280) );
  MUX2_X1 U301 ( .A(n533), .B(n280), .S(n301), .Z(n429) );
  MUX2_X1 U302 ( .A(product[2]), .B(n535), .S(n301), .Z(n431) );
  MUX2_X1 U303 ( .A(n535), .B(n536), .S(n301), .Z(n433) );
  INV_X1 U304 ( .A(n281), .ZN(n283) );
  NAND2_X1 U305 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U306 ( .A(n285), .B(n284), .Z(n286) );
  MUX2_X1 U307 ( .A(n536), .B(n286), .S(n301), .Z(n435) );
  MUX2_X1 U308 ( .A(product[3]), .B(n538), .S(n301), .Z(n437) );
  MUX2_X1 U309 ( .A(n538), .B(n539), .S(n301), .Z(n439) );
  NAND2_X1 U310 ( .A1(n288), .A2(n287), .ZN(n290) );
  XNOR2_X1 U311 ( .A(n290), .B(n289), .ZN(n291) );
  MUX2_X1 U312 ( .A(n539), .B(n291), .S(n301), .Z(n441) );
  MUX2_X1 U313 ( .A(product[4]), .B(n541), .S(n301), .Z(n443) );
  MUX2_X1 U314 ( .A(n541), .B(n542), .S(n301), .Z(n445) );
  INV_X1 U315 ( .A(n292), .ZN(n294) );
  NAND2_X1 U316 ( .A1(n294), .A2(n293), .ZN(n296) );
  XOR2_X1 U317 ( .A(n296), .B(n295), .Z(n297) );
  MUX2_X1 U318 ( .A(n542), .B(n297), .S(n301), .Z(n447) );
  MUX2_X1 U319 ( .A(product[5]), .B(n544), .S(n301), .Z(n449) );
  MUX2_X1 U320 ( .A(n544), .B(n545), .S(n301), .Z(n451) );
  MUX2_X1 U321 ( .A(product[6]), .B(n547), .S(n301), .Z(n455) );
  NAND2_X1 U322 ( .A1(n409), .A2(n357), .ZN(n298) );
  XOR2_X1 U323 ( .A(n298), .B(n363), .Z(n299) );
  MUX2_X1 U324 ( .A(n547), .B(n299), .S(n301), .Z(n457) );
  MUX2_X1 U325 ( .A(product[7]), .B(n549), .S(n301), .Z(n459) );
  OAI21_X1 U326 ( .B1(n356), .B2(n363), .A(n357), .ZN(n303) );
  NAND2_X1 U327 ( .A1(n347), .A2(n355), .ZN(n300) );
  XNOR2_X1 U328 ( .A(n303), .B(n300), .ZN(n302) );
  MUX2_X1 U329 ( .A(n549), .B(n302), .S(n301), .Z(n461) );
  BUF_X2 U330 ( .A(en), .Z(n345) );
  MUX2_X1 U331 ( .A(product[8]), .B(n551), .S(n345), .Z(n463) );
  AOI21_X1 U332 ( .B1(n303), .B2(n347), .A(n410), .ZN(n306) );
  NAND2_X1 U333 ( .A1(n411), .A2(n354), .ZN(n304) );
  XOR2_X1 U334 ( .A(n306), .B(n304), .Z(n305) );
  MUX2_X1 U335 ( .A(n551), .B(n305), .S(n345), .Z(n465) );
  MUX2_X1 U336 ( .A(product[9]), .B(n553), .S(n345), .Z(n467) );
  OAI21_X1 U337 ( .B1(n306), .B2(n353), .A(n354), .ZN(n317) );
  INV_X1 U338 ( .A(n317), .ZN(n309) );
  NAND2_X1 U339 ( .A1(n412), .A2(n361), .ZN(n307) );
  XOR2_X1 U340 ( .A(n309), .B(n307), .Z(n308) );
  MUX2_X1 U341 ( .A(n553), .B(n308), .S(n345), .Z(n469) );
  MUX2_X1 U342 ( .A(product[10]), .B(n555), .S(n345), .Z(n471) );
  OAI21_X1 U343 ( .B1(n309), .B2(n362), .A(n361), .ZN(n312) );
  NOR2_X1 U344 ( .A1(n364), .A2(n365), .ZN(n315) );
  INV_X1 U345 ( .A(n315), .ZN(n310) );
  NAND2_X1 U346 ( .A1(n364), .A2(n365), .ZN(n314) );
  NAND2_X1 U347 ( .A1(n310), .A2(n314), .ZN(n311) );
  XNOR2_X1 U348 ( .A(n312), .B(n311), .ZN(n313) );
  MUX2_X1 U349 ( .A(n555), .B(n313), .S(n345), .Z(n473) );
  MUX2_X1 U350 ( .A(product[11]), .B(n557), .S(n345), .Z(n475) );
  NOR2_X1 U351 ( .A1(n315), .A2(n362), .ZN(n318) );
  OAI21_X1 U352 ( .B1(n315), .B2(n361), .A(n314), .ZN(n316) );
  AOI21_X1 U353 ( .B1(n318), .B2(n317), .A(n316), .ZN(n341) );
  NAND2_X1 U354 ( .A1(n413), .A2(n352), .ZN(n319) );
  XOR2_X1 U355 ( .A(n341), .B(n319), .Z(n320) );
  MUX2_X1 U356 ( .A(n557), .B(n320), .S(n345), .Z(n477) );
  MUX2_X1 U357 ( .A(product[12]), .B(n559), .S(n345), .Z(n479) );
  OAI21_X1 U358 ( .B1(n341), .B2(n359), .A(n352), .ZN(n322) );
  NAND2_X1 U359 ( .A1(n349), .A2(n360), .ZN(n321) );
  XNOR2_X1 U360 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U361 ( .A(n559), .B(n323), .S(n345), .Z(n481) );
  MUX2_X1 U362 ( .A(product[13]), .B(n561), .S(n345), .Z(n483) );
  NAND2_X1 U363 ( .A1(n413), .A2(n349), .ZN(n325) );
  AOI21_X1 U364 ( .B1(n408), .B2(n349), .A(n414), .ZN(n324) );
  OAI21_X1 U365 ( .B1(n341), .B2(n325), .A(n324), .ZN(n327) );
  NAND2_X1 U366 ( .A1(n348), .A2(n358), .ZN(n326) );
  XNOR2_X1 U367 ( .A(n327), .B(n326), .ZN(n328) );
  MUX2_X1 U368 ( .A(n561), .B(n328), .S(n345), .Z(n485) );
  MUX2_X1 U369 ( .A(product[14]), .B(n563), .S(n345), .Z(n487) );
  AND2_X1 U370 ( .A1(n349), .A2(n348), .ZN(n336) );
  NAND2_X1 U371 ( .A1(n413), .A2(n336), .ZN(n332) );
  NAND2_X1 U372 ( .A1(n349), .A2(n348), .ZN(n330) );
  AOI21_X1 U373 ( .B1(n414), .B2(n348), .A(n407), .ZN(n329) );
  OAI21_X1 U374 ( .B1(n330), .B2(n352), .A(n329), .ZN(n338) );
  INV_X1 U375 ( .A(n338), .ZN(n331) );
  OAI21_X1 U376 ( .B1(n341), .B2(n332), .A(n331), .ZN(n334) );
  NAND2_X1 U377 ( .A1(n346), .A2(n351), .ZN(n333) );
  XNOR2_X1 U378 ( .A(n334), .B(n333), .ZN(n335) );
  MUX2_X1 U379 ( .A(n563), .B(n335), .S(n345), .Z(n489) );
  MUX2_X1 U380 ( .A(product[15]), .B(n565), .S(n345), .Z(n491) );
  AND2_X1 U381 ( .A1(n413), .A2(n346), .ZN(n337) );
  NAND2_X1 U382 ( .A1(n337), .A2(n336), .ZN(n340) );
  AOI21_X1 U383 ( .B1(n338), .B2(n346), .A(n406), .ZN(n339) );
  OAI21_X1 U384 ( .B1(n341), .B2(n340), .A(n339), .ZN(n342) );
  XNOR2_X1 U385 ( .A(n342), .B(n350), .ZN(n343) );
  MUX2_X1 U386 ( .A(n565), .B(n343), .S(n345), .Z(n493) );
  MUX2_X1 U387 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n345), .Z(n495) );
  MUX2_X1 U388 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n345), .Z(n497) );
  MUX2_X1 U389 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n345), .Z(n499) );
  MUX2_X1 U390 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n345), .Z(n501) );
  MUX2_X1 U391 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n345), .Z(n503) );
  MUX2_X1 U392 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n345), .Z(n505) );
  MUX2_X1 U393 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n345), .Z(n507) );
  MUX2_X1 U394 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n345), .Z(n509) );
  MUX2_X1 U395 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n345), .Z(n511) );
  MUX2_X1 U396 ( .A(\mult_x_1/n313 ), .B(A_extended[1]), .S(n345), .Z(n513) );
  MUX2_X1 U397 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n345), .Z(n515) );
  MUX2_X1 U398 ( .A(n344), .B(A_extended[3]), .S(n345), .Z(n517) );
  MUX2_X1 U399 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n345), .Z(n519) );
  MUX2_X1 U400 ( .A(n19), .B(A_extended[5]), .S(n345), .Z(n521) );
  MUX2_X1 U401 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n345), .Z(n523) );
  MUX2_X1 U402 ( .A(n17), .B(A_extended[7]), .S(n345), .Z(n525) );
  OR2_X1 U403 ( .A1(n345), .A2(n567), .ZN(n527) );
endmodule


module conv_128_32_DW_mult_pipe_J1_21 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n310 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n355, n357, n359, n361, n363, n365, n367, n369, n371, n373,
         n375, n377, n379, n381, n383, n385, n387, n389, n391, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n408, n410, n412, n414, n416, n418, n420, n422, n424, n426,
         n428, n430, n432, n434, n436, n438, n440, n442, n444, n446, n448,
         n450, n452, n454, n456, n458, n460, n462, n464, n466, n468, n470,
         n472, n474, n476, n478, n480, n482, n484, n486, n488, n490, n492,
         n494, n496, n498, n500, n502, n504, n506, n508, n510, n512, n514,
         n516, n518, n519, n521, n522, n524, n525, n527, n528, n530, n531,
         n533, n534, n536, n538, n540, n542, n544, n546, n548, n550, n552,
         n554, n555, n556, n557, n558, n559;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n516), .CK(clk), .Q(n558), 
        .QN(n405) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n514), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n406) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n506), .CK(clk), .Q(n556), 
        .QN(n12) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(rst_n), .SE(n504), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n8) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n10) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n404), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n9), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n404), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n9), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n404), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n9), .SE(n482), .CK(clk), .Q(n554) );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n404), .SE(n480), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n9), .SE(n478), .CK(clk), .Q(n552) );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n404), .SE(n476), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n9), .SE(n474), .CK(clk), .Q(n550) );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(rst_n), .SE(n472), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n404), .SE(n470), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n9), .SE(n468), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n404), .SE(n466), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n9), .SE(n464), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG23_S3 ( .D(1'b0), .SI(n404), .SE(n462), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG24_S4 ( .D(1'b0), .SI(n9), .SE(n460), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG21_S3 ( .D(1'b0), .SI(n404), .SE(n458), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG22_S4 ( .D(1'b0), .SI(n9), .SE(n456), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n404), .SE(n454), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n9), .SE(n452), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n404), .SE(n450), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n9), .SE(n448), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n404), .SE(n446), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n9), .SE(n444), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n404), .SE(n442), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n9), .SE(n440), .CK(clk), .Q(n533) );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n404), .SE(n438), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n9), .SE(n436), .CK(clk), .Q(n531) );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n404), .SE(n434), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n9), .SE(n432), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n404), .SE(n430), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n9), .SE(n428), .CK(clk), .Q(n527) );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n404), .SE(n426), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n424), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n422), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n420), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n9), .SE(n418), .CK(clk), .Q(n522) );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n416), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n414), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n412), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n404), .SE(n410), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n9), .SE(n408), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n559), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n559), .SE(n389), .CK(
        clk), .Q(n402), .QN(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n559), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n350), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n559), .SE(n385), .CK(
        clk), .Q(n332), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n559), .SE(n383), .CK(
        clk), .Q(n401), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n559), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n559), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n346), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n559), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n345), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n559), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n559), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n343), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n559), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n342), .QN(n16) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n559), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n341), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n559), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n340), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n559), .SI(1'b1), .SE(n365), .CK(clk), 
        .Q(n339), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n559), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n338), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n559), .SE(n361), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n559), .SE(n359), .CK(
        clk), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n559), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n559), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n559), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n333), .QN(n396) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(rst_n), .SE(n502), .CK(clk), .Q(n555), 
        .QN(n15) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n510), .CK(clk), .Q(n557), 
        .QN(n11) );
  INV_X1 U2 ( .A(rst_n), .ZN(n559) );
  INV_X2 U3 ( .A(n233), .ZN(n162) );
  BUF_X1 U4 ( .A(n25), .Z(n178) );
  CLKBUF_X2 U5 ( .A(n24), .Z(n174) );
  NAND2_X1 U6 ( .A1(n17), .A2(n18), .ZN(n164) );
  NAND2_X1 U7 ( .A1(n19), .A2(n20), .ZN(n244) );
  INV_X1 U8 ( .A(n11), .ZN(n6) );
  BUF_X1 U9 ( .A(n556), .Z(n330) );
  OR2_X1 U10 ( .A1(n191), .A2(n190), .ZN(n150) );
  XNOR2_X1 U11 ( .A(n149), .B(n148), .ZN(n191) );
  INV_X1 U12 ( .A(n117), .ZN(n126) );
  OAI22_X1 U13 ( .A1(n110), .A2(n162), .B1(n164), .B2(n111), .ZN(n117) );
  INV_X1 U14 ( .A(n88), .ZN(n53) );
  NAND2_X1 U15 ( .A1(n125), .A2(n124), .ZN(n148) );
  NAND2_X1 U16 ( .A1(n123), .A2(n122), .ZN(n124) );
  NAND2_X1 U17 ( .A1(n121), .A2(n13), .ZN(n125) );
  XNOR2_X1 U18 ( .A(n121), .B(n69), .ZN(n140) );
  XNOR2_X1 U19 ( .A(n123), .B(n122), .ZN(n69) );
  XNOR2_X1 U20 ( .A(n70), .B(n38), .ZN(n80) );
  XNOR2_X1 U21 ( .A(n72), .B(n71), .ZN(n38) );
  XNOR2_X1 U22 ( .A(n91), .B(n90), .ZN(n194) );
  XNOR2_X1 U23 ( .A(n101), .B(n100), .ZN(n196) );
  NAND2_X1 U24 ( .A1(n54), .A2(n53), .ZN(n58) );
  NAND2_X1 U25 ( .A1(n147), .A2(n146), .ZN(n132) );
  OR2_X1 U26 ( .A1(n147), .A2(n146), .ZN(n131) );
  NAND2_X1 U27 ( .A1(n84), .A2(n83), .ZN(n226) );
  NAND2_X1 U28 ( .A1(n82), .A2(n81), .ZN(n83) );
  OAI21_X1 U29 ( .B1(n82), .B2(n81), .A(n80), .ZN(n84) );
  BUF_X8 U30 ( .A(en), .Z(n331) );
  INV_X1 U31 ( .A(n36), .ZN(n5) );
  NOR2_X1 U32 ( .A1(n405), .A2(n406), .ZN(n112) );
  INV_X1 U33 ( .A(n36), .ZN(n177) );
  BUF_X1 U34 ( .A(\mult_x_1/n310 ), .Z(n7) );
  XNOR2_X1 U35 ( .A(\mult_x_1/a[2] ), .B(n12), .ZN(n19) );
  XNOR2_X1 U36 ( .A(n15), .B(n8), .ZN(n20) );
  INV_X1 U37 ( .A(n559), .ZN(n9) );
  OR2_X1 U38 ( .A1(n35), .A2(n34), .ZN(n72) );
  INV_X1 U39 ( .A(n559), .ZN(n404) );
  OR2_X1 U40 ( .A1(n123), .A2(n122), .ZN(n13) );
  OR2_X1 U41 ( .A1(n72), .A2(n71), .ZN(n14) );
  XOR2_X1 U42 ( .A(\mult_x_1/a[4] ), .B(n557), .Z(n17) );
  XNOR2_X1 U43 ( .A(n556), .B(\mult_x_1/a[4] ), .ZN(n18) );
  XNOR2_X1 U44 ( .A(n6), .B(\mult_x_1/n284 ), .ZN(n44) );
  INV_X1 U45 ( .A(n18), .ZN(n233) );
  XNOR2_X1 U46 ( .A(n6), .B(\mult_x_1/n283 ), .ZN(n27) );
  OAI22_X1 U47 ( .A1(n164), .A2(n44), .B1(n162), .B2(n27), .ZN(n35) );
  XNOR2_X1 U48 ( .A(n330), .B(\mult_x_1/n282 ), .ZN(n43) );
  INV_X1 U49 ( .A(n20), .ZN(n21) );
  INV_X2 U50 ( .A(n21), .ZN(n246) );
  XNOR2_X1 U51 ( .A(n330), .B(\mult_x_1/n281 ), .ZN(n28) );
  OAI22_X1 U52 ( .A1(n244), .A2(n43), .B1(n246), .B2(n28), .ZN(n34) );
  XNOR2_X1 U53 ( .A(n35), .B(n34), .ZN(n57) );
  INV_X1 U54 ( .A(n112), .ZN(n36) );
  OR2_X1 U55 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n22) );
  XNOR2_X1 U56 ( .A(n112), .B(\mult_x_1/n310 ), .ZN(n25) );
  NOR2_X1 U57 ( .A1(n22), .A2(n178), .ZN(n56) );
  XOR2_X1 U58 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n23) );
  XNOR2_X1 U59 ( .A(n557), .B(\mult_x_1/a[6] ), .ZN(n24) );
  NAND2_X2 U60 ( .A1(n23), .A2(n24), .ZN(n173) );
  XNOR2_X1 U61 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n41) );
  XNOR2_X1 U62 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n32) );
  OAI22_X1 U63 ( .A1(n173), .A2(n41), .B1(n174), .B2(n32), .ZN(n94) );
  NAND2_X1 U64 ( .A1(n555), .A2(n10), .ZN(n249) );
  XNOR2_X1 U65 ( .A(n555), .B(\mult_x_1/n281 ), .ZN(n96) );
  AND2_X1 U66 ( .A1(n558), .A2(\mult_x_1/n281 ), .ZN(n107) );
  XNOR2_X1 U67 ( .A(n107), .B(n555), .ZN(n29) );
  OAI22_X1 U68 ( .A1(n249), .A2(n96), .B1(n29), .B2(n10), .ZN(n93) );
  INV_X1 U69 ( .A(n25), .ZN(n26) );
  AND2_X1 U70 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n92) );
  XNOR2_X1 U71 ( .A(n7), .B(\mult_x_1/n285 ), .ZN(n31) );
  XNOR2_X1 U72 ( .A(n7), .B(\mult_x_1/n284 ), .ZN(n75) );
  OAI22_X1 U73 ( .A1(n173), .A2(n31), .B1(n174), .B2(n75), .ZN(n66) );
  XNOR2_X1 U74 ( .A(n6), .B(\mult_x_1/n282 ), .ZN(n68) );
  OAI22_X1 U75 ( .A1(n164), .A2(n27), .B1(n162), .B2(n68), .ZN(n65) );
  XNOR2_X1 U76 ( .A(n107), .B(n330), .ZN(n76) );
  OAI22_X1 U77 ( .A1(n244), .A2(n28), .B1(n76), .B2(n246), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n64) );
  XNOR2_X1 U79 ( .A(n82), .B(n81), .ZN(n39) );
  AOI21_X1 U80 ( .B1(n249), .B2(n10), .A(n29), .ZN(n30) );
  INV_X1 U81 ( .A(n30), .ZN(n52) );
  OAI22_X1 U82 ( .A1(n173), .A2(n32), .B1(n174), .B2(n31), .ZN(n51) );
  XNOR2_X1 U83 ( .A(n5), .B(\mult_x_1/n287 ), .ZN(n33) );
  NOR2_X1 U84 ( .A1(n33), .A2(n178), .ZN(n50) );
  XNOR2_X1 U85 ( .A(n177), .B(\mult_x_1/n286 ), .ZN(n37) );
  NOR2_X1 U86 ( .A1(n37), .A2(n178), .ZN(n71) );
  XNOR2_X1 U87 ( .A(n39), .B(n80), .ZN(n221) );
  OR2_X1 U88 ( .A1(\mult_x_1/n288 ), .A2(n406), .ZN(n40) );
  OAI22_X1 U89 ( .A1(n173), .A2(n406), .B1(n40), .B2(n174), .ZN(n155) );
  XNOR2_X1 U90 ( .A(n7), .B(\mult_x_1/n288 ), .ZN(n42) );
  OAI22_X1 U91 ( .A1(n173), .A2(n42), .B1(n174), .B2(n41), .ZN(n154) );
  XNOR2_X1 U92 ( .A(n330), .B(\mult_x_1/n283 ), .ZN(n97) );
  OAI22_X1 U93 ( .A1(n244), .A2(n97), .B1(n246), .B2(n43), .ZN(n98) );
  INV_X1 U94 ( .A(n98), .ZN(n46) );
  XNOR2_X1 U95 ( .A(n6), .B(\mult_x_1/n285 ), .ZN(n95) );
  OAI22_X1 U96 ( .A1(n164), .A2(n95), .B1(n162), .B2(n44), .ZN(n99) );
  INV_X1 U97 ( .A(n99), .ZN(n45) );
  NAND2_X1 U98 ( .A1(n46), .A2(n45), .ZN(n47) );
  NAND2_X1 U99 ( .A1(n101), .A2(n47), .ZN(n49) );
  NAND2_X1 U100 ( .A1(n98), .A2(n99), .ZN(n48) );
  NAND2_X1 U101 ( .A1(n49), .A2(n48), .ZN(n89) );
  INV_X1 U102 ( .A(n89), .ZN(n54) );
  FA_X1 U103 ( .A(n52), .B(n51), .CI(n50), .CO(n70), .S(n88) );
  FA_X1 U104 ( .A(n57), .B(n56), .CI(n55), .CO(n82), .S(n91) );
  NAND2_X1 U105 ( .A1(n58), .A2(n91), .ZN(n60) );
  NAND2_X1 U106 ( .A1(n89), .A2(n88), .ZN(n59) );
  NAND2_X1 U107 ( .A1(n60), .A2(n59), .ZN(n220) );
  NAND2_X1 U108 ( .A1(n221), .A2(n220), .ZN(n61) );
  NAND2_X1 U109 ( .A1(n61), .A2(n331), .ZN(n63) );
  OR2_X1 U110 ( .A1(n331), .A2(n332), .ZN(n62) );
  NAND2_X1 U111 ( .A1(n63), .A2(n62), .ZN(n385) );
  FA_X1 U112 ( .A(n66), .B(n65), .CI(n64), .CO(n121), .S(n81) );
  XNOR2_X1 U113 ( .A(n177), .B(\mult_x_1/n285 ), .ZN(n67) );
  NOR2_X1 U114 ( .A1(n67), .A2(n178), .ZN(n123) );
  XNOR2_X1 U115 ( .A(n557), .B(\mult_x_1/n281 ), .ZN(n111) );
  OAI22_X1 U116 ( .A1(n164), .A2(n68), .B1(n162), .B2(n111), .ZN(n122) );
  NAND2_X1 U117 ( .A1(n70), .A2(n14), .ZN(n74) );
  NAND2_X1 U118 ( .A1(n72), .A2(n71), .ZN(n73) );
  NAND2_X1 U119 ( .A1(n74), .A2(n73), .ZN(n142) );
  XNOR2_X1 U120 ( .A(n7), .B(\mult_x_1/n283 ), .ZN(n115) );
  OAI22_X1 U121 ( .A1(n173), .A2(n75), .B1(n174), .B2(n115), .ZN(n130) );
  AOI21_X1 U122 ( .B1(n246), .B2(n244), .A(n76), .ZN(n77) );
  INV_X1 U123 ( .A(n77), .ZN(n129) );
  XNOR2_X1 U124 ( .A(n142), .B(n141), .ZN(n79) );
  XNOR2_X1 U125 ( .A(n140), .B(n79), .ZN(n227) );
  NAND2_X1 U126 ( .A1(n227), .A2(n226), .ZN(n85) );
  NAND2_X1 U127 ( .A1(n85), .A2(n331), .ZN(n87) );
  OR2_X1 U128 ( .A1(n331), .A2(n395), .ZN(n86) );
  NAND2_X1 U129 ( .A1(n87), .A2(n86), .ZN(n367) );
  XNOR2_X1 U130 ( .A(n89), .B(n88), .ZN(n90) );
  FA_X1 U131 ( .A(n92), .B(n94), .CI(n93), .CO(n55), .S(n198) );
  XNOR2_X1 U132 ( .A(n6), .B(\mult_x_1/n286 ), .ZN(n161) );
  OAI22_X1 U133 ( .A1(n164), .A2(n161), .B1(n162), .B2(n95), .ZN(n158) );
  XNOR2_X1 U134 ( .A(n555), .B(\mult_x_1/n282 ), .ZN(n151) );
  OAI22_X1 U135 ( .A1(n249), .A2(n151), .B1(n96), .B2(n10), .ZN(n157) );
  XNOR2_X1 U136 ( .A(n330), .B(\mult_x_1/n284 ), .ZN(n153) );
  OAI22_X1 U137 ( .A1(n244), .A2(n153), .B1(n246), .B2(n97), .ZN(n156) );
  XNOR2_X1 U138 ( .A(n99), .B(n98), .ZN(n100) );
  NAND2_X1 U139 ( .A1(n194), .A2(n193), .ZN(n102) );
  NAND2_X1 U140 ( .A1(n102), .A2(n331), .ZN(n104) );
  OR2_X1 U141 ( .A1(n331), .A2(n16), .ZN(n103) );
  NAND2_X1 U142 ( .A1(n104), .A2(n103), .ZN(n371) );
  XNOR2_X1 U163 ( .A(n177), .B(\mult_x_1/n282 ), .ZN(n105) );
  NOR2_X1 U164 ( .A1(n105), .A2(n178), .ZN(n171) );
  XNOR2_X1 U165 ( .A(n7), .B(\mult_x_1/n281 ), .ZN(n106) );
  XNOR2_X1 U166 ( .A(n107), .B(n7), .ZN(n172) );
  OAI22_X1 U167 ( .A1(n173), .A2(n106), .B1(n172), .B2(n174), .ZN(n175) );
  INV_X1 U168 ( .A(n175), .ZN(n170) );
  XNOR2_X1 U169 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n114) );
  OAI22_X1 U170 ( .A1(n173), .A2(n114), .B1(n174), .B2(n106), .ZN(n119) );
  NAND2_X1 U171 ( .A1(n162), .A2(n164), .ZN(n109) );
  XNOR2_X1 U172 ( .A(n107), .B(n557), .ZN(n110) );
  INV_X1 U173 ( .A(n110), .ZN(n108) );
  NAND2_X1 U174 ( .A1(n109), .A2(n108), .ZN(n118) );
  XNOR2_X1 U175 ( .A(n5), .B(\mult_x_1/n284 ), .ZN(n113) );
  NOR2_X1 U176 ( .A1(n113), .A2(n178), .ZN(n128) );
  OAI22_X1 U177 ( .A1(n173), .A2(n115), .B1(n174), .B2(n114), .ZN(n127) );
  XNOR2_X1 U178 ( .A(n177), .B(\mult_x_1/n283 ), .ZN(n116) );
  NOR2_X1 U179 ( .A1(n116), .A2(n178), .ZN(n135) );
  FA_X1 U180 ( .A(n119), .B(n118), .CI(n117), .CO(n169), .S(n134) );
  OR2_X1 U181 ( .A1(n188), .A2(n187), .ZN(n120) );
  MUX2_X1 U182 ( .A(n333), .B(n120), .S(n331), .Z(n353) );
  FA_X1 U183 ( .A(n128), .B(n127), .CI(n126), .CO(n136), .S(n147) );
  FA_X1 U184 ( .A(n130), .B(n129), .CI(n78), .CO(n146), .S(n141) );
  NAND2_X1 U185 ( .A1(n148), .A2(n131), .ZN(n133) );
  NAND2_X1 U186 ( .A1(n133), .A2(n132), .ZN(n223) );
  INV_X1 U187 ( .A(n223), .ZN(n138) );
  FA_X1 U188 ( .A(n136), .B(n135), .CI(n134), .CO(n187), .S(n224) );
  INV_X1 U189 ( .A(n224), .ZN(n137) );
  NAND2_X1 U190 ( .A1(n138), .A2(n137), .ZN(n139) );
  MUX2_X1 U191 ( .A(n334), .B(n139), .S(n331), .Z(n355) );
  NAND2_X1 U192 ( .A1(n140), .A2(n142), .ZN(n145) );
  NAND2_X1 U193 ( .A1(n140), .A2(n141), .ZN(n144) );
  NAND2_X1 U194 ( .A1(n142), .A2(n141), .ZN(n143) );
  NAND3_X1 U195 ( .A1(n145), .A2(n144), .A3(n143), .ZN(n190) );
  XNOR2_X1 U196 ( .A(n147), .B(n146), .ZN(n149) );
  MUX2_X1 U197 ( .A(n335), .B(n150), .S(n331), .Z(n357) );
  XNOR2_X1 U198 ( .A(n555), .B(\mult_x_1/n283 ), .ZN(n213) );
  OAI22_X1 U199 ( .A1(n249), .A2(n213), .B1(n151), .B2(n10), .ZN(n167) );
  INV_X1 U200 ( .A(n174), .ZN(n152) );
  AND2_X1 U201 ( .A1(\mult_x_1/n288 ), .A2(n152), .ZN(n166) );
  XNOR2_X1 U202 ( .A(n330), .B(\mult_x_1/n285 ), .ZN(n212) );
  OAI22_X1 U203 ( .A1(n244), .A2(n212), .B1(n246), .B2(n153), .ZN(n165) );
  HA_X1 U204 ( .A(n155), .B(n154), .CO(n101), .S(n200) );
  FA_X1 U205 ( .A(n158), .B(n157), .CI(n156), .CO(n197), .S(n199) );
  OR2_X1 U206 ( .A1(\mult_x_1/n288 ), .A2(n11), .ZN(n159) );
  OAI22_X1 U207 ( .A1(n164), .A2(n11), .B1(n159), .B2(n162), .ZN(n215) );
  XNOR2_X1 U208 ( .A(n6), .B(\mult_x_1/n288 ), .ZN(n160) );
  XNOR2_X1 U209 ( .A(n6), .B(\mult_x_1/n287 ), .ZN(n163) );
  OAI22_X1 U210 ( .A1(n164), .A2(n160), .B1(n162), .B2(n163), .ZN(n214) );
  OAI22_X1 U211 ( .A1(n164), .A2(n163), .B1(n162), .B2(n161), .ZN(n210) );
  FA_X1 U212 ( .A(n167), .B(n166), .CI(n165), .CO(n201), .S(n209) );
  OR2_X1 U213 ( .A1(n207), .A2(n206), .ZN(n168) );
  MUX2_X1 U214 ( .A(n336), .B(n168), .S(n331), .Z(n359) );
  FA_X1 U215 ( .A(n171), .B(n170), .CI(n169), .CO(n183), .S(n188) );
  AOI21_X1 U216 ( .B1(n174), .B2(n173), .A(n172), .ZN(n176) );
  XNOR2_X1 U217 ( .A(n176), .B(n175), .ZN(n181) );
  XNOR2_X1 U218 ( .A(n177), .B(\mult_x_1/n281 ), .ZN(n179) );
  OR2_X1 U219 ( .A1(n179), .A2(n178), .ZN(n180) );
  XNOR2_X1 U220 ( .A(n181), .B(n180), .ZN(n182) );
  OR2_X1 U221 ( .A1(n183), .A2(n182), .ZN(n185) );
  NAND2_X1 U222 ( .A1(n183), .A2(n182), .ZN(n184) );
  NAND2_X1 U223 ( .A1(n185), .A2(n184), .ZN(n186) );
  MUX2_X1 U224 ( .A(n337), .B(n186), .S(n331), .Z(n361) );
  NAND2_X1 U225 ( .A1(n188), .A2(n187), .ZN(n189) );
  MUX2_X1 U226 ( .A(n338), .B(n189), .S(n331), .Z(n363) );
  NAND2_X1 U227 ( .A1(n191), .A2(n190), .ZN(n192) );
  MUX2_X1 U228 ( .A(n339), .B(n192), .S(n331), .Z(n365) );
  NOR2_X1 U229 ( .A1(n194), .A2(n193), .ZN(n195) );
  MUX2_X1 U230 ( .A(n341), .B(n195), .S(n331), .Z(n369) );
  FA_X1 U231 ( .A(n198), .B(n197), .CI(n196), .CO(n193), .S(n204) );
  FA_X1 U232 ( .A(n201), .B(n200), .CI(n199), .CO(n203), .S(n207) );
  NOR2_X1 U233 ( .A1(n204), .A2(n203), .ZN(n202) );
  MUX2_X1 U234 ( .A(n343), .B(n202), .S(n331), .Z(n373) );
  NAND2_X1 U235 ( .A1(n204), .A2(n203), .ZN(n205) );
  MUX2_X1 U236 ( .A(n344), .B(n205), .S(n331), .Z(n375) );
  NAND2_X1 U237 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U238 ( .A(n345), .B(n208), .S(n331), .Z(n377) );
  FA_X1 U239 ( .A(n211), .B(n210), .CI(n209), .CO(n206), .S(n218) );
  XNOR2_X1 U240 ( .A(n330), .B(\mult_x_1/n286 ), .ZN(n234) );
  OAI22_X1 U241 ( .A1(n244), .A2(n234), .B1(n246), .B2(n212), .ZN(n231) );
  XNOR2_X1 U242 ( .A(n555), .B(\mult_x_1/n284 ), .ZN(n232) );
  OAI22_X1 U243 ( .A1(n249), .A2(n232), .B1(n213), .B2(n10), .ZN(n230) );
  HA_X1 U244 ( .A(n215), .B(n214), .CO(n211), .S(n229) );
  NOR2_X1 U245 ( .A1(n218), .A2(n217), .ZN(n216) );
  MUX2_X1 U246 ( .A(n346), .B(n216), .S(n331), .Z(n379) );
  NAND2_X1 U247 ( .A1(n218), .A2(n217), .ZN(n219) );
  MUX2_X1 U248 ( .A(n347), .B(n219), .S(n331), .Z(n381) );
  NOR2_X1 U249 ( .A1(n221), .A2(n220), .ZN(n222) );
  MUX2_X1 U250 ( .A(n348), .B(n222), .S(n331), .Z(n383) );
  NAND2_X1 U251 ( .A1(n224), .A2(n223), .ZN(n225) );
  MUX2_X1 U252 ( .A(n350), .B(n225), .S(n331), .Z(n387) );
  NOR2_X1 U253 ( .A1(n227), .A2(n226), .ZN(n228) );
  MUX2_X1 U254 ( .A(n351), .B(n228), .S(n331), .Z(n389) );
  FA_X1 U255 ( .A(n231), .B(n230), .CI(n229), .CO(n217), .S(n259) );
  XNOR2_X1 U256 ( .A(n555), .B(\mult_x_1/n285 ), .ZN(n240) );
  OAI22_X1 U257 ( .A1(n249), .A2(n240), .B1(n232), .B2(n10), .ZN(n237) );
  AND2_X1 U258 ( .A1(\mult_x_1/n288 ), .A2(n233), .ZN(n236) );
  XNOR2_X1 U259 ( .A(n330), .B(\mult_x_1/n287 ), .ZN(n238) );
  OAI22_X1 U260 ( .A1(n244), .A2(n238), .B1(n246), .B2(n234), .ZN(n235) );
  OR2_X1 U261 ( .A1(n259), .A2(n258), .ZN(n285) );
  FA_X1 U262 ( .A(n237), .B(n236), .CI(n235), .CO(n258), .S(n257) );
  XNOR2_X1 U263 ( .A(n330), .B(\mult_x_1/n288 ), .ZN(n239) );
  OAI22_X1 U264 ( .A1(n244), .A2(n239), .B1(n246), .B2(n238), .ZN(n242) );
  XNOR2_X1 U265 ( .A(n555), .B(\mult_x_1/n286 ), .ZN(n245) );
  OAI22_X1 U266 ( .A1(n249), .A2(n245), .B1(n240), .B2(n10), .ZN(n241) );
  NOR2_X1 U267 ( .A1(n257), .A2(n256), .ZN(n278) );
  HA_X1 U268 ( .A(n242), .B(n241), .CO(n256), .S(n254) );
  OR2_X1 U269 ( .A1(\mult_x_1/n288 ), .A2(n12), .ZN(n243) );
  OAI22_X1 U270 ( .A1(n244), .A2(n12), .B1(n243), .B2(n246), .ZN(n253) );
  OR2_X1 U271 ( .A1(n254), .A2(n253), .ZN(n274) );
  XNOR2_X1 U272 ( .A(n555), .B(\mult_x_1/n287 ), .ZN(n248) );
  OAI22_X1 U273 ( .A1(n249), .A2(n248), .B1(n245), .B2(n10), .ZN(n252) );
  INV_X1 U274 ( .A(n246), .ZN(n247) );
  AND2_X1 U275 ( .A1(\mult_x_1/n288 ), .A2(n247), .ZN(n251) );
  NOR2_X1 U276 ( .A1(n252), .A2(n251), .ZN(n267) );
  OAI22_X1 U277 ( .A1(n249), .A2(\mult_x_1/n288 ), .B1(n248), .B2(n10), .ZN(
        n264) );
  OR2_X1 U278 ( .A1(\mult_x_1/n288 ), .A2(n15), .ZN(n250) );
  NAND2_X1 U279 ( .A1(n250), .A2(n249), .ZN(n263) );
  NAND2_X1 U280 ( .A1(n264), .A2(n263), .ZN(n270) );
  NAND2_X1 U281 ( .A1(n252), .A2(n251), .ZN(n268) );
  OAI21_X1 U282 ( .B1(n267), .B2(n270), .A(n268), .ZN(n275) );
  NAND2_X1 U283 ( .A1(n254), .A2(n253), .ZN(n273) );
  INV_X1 U284 ( .A(n273), .ZN(n255) );
  AOI21_X1 U285 ( .B1(n274), .B2(n275), .A(n255), .ZN(n281) );
  NAND2_X1 U286 ( .A1(n257), .A2(n256), .ZN(n279) );
  OAI21_X1 U287 ( .B1(n278), .B2(n281), .A(n279), .ZN(n286) );
  NAND2_X1 U288 ( .A1(n259), .A2(n258), .ZN(n284) );
  INV_X1 U289 ( .A(n284), .ZN(n260) );
  AOI21_X1 U290 ( .B1(n285), .B2(n286), .A(n260), .ZN(n261) );
  MUX2_X1 U291 ( .A(n352), .B(n261), .S(n331), .Z(n391) );
  MUX2_X1 U292 ( .A(product[0]), .B(n518), .S(n331), .Z(n408) );
  MUX2_X1 U293 ( .A(n518), .B(n519), .S(n331), .Z(n410) );
  AND2_X1 U294 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n262) );
  MUX2_X1 U295 ( .A(n519), .B(n262), .S(n331), .Z(n412) );
  MUX2_X1 U296 ( .A(product[1]), .B(n521), .S(n331), .Z(n414) );
  MUX2_X1 U297 ( .A(n521), .B(n522), .S(n331), .Z(n416) );
  OR2_X1 U298 ( .A1(n264), .A2(n263), .ZN(n265) );
  AND2_X1 U299 ( .A1(n265), .A2(n270), .ZN(n266) );
  MUX2_X1 U300 ( .A(n522), .B(n266), .S(n331), .Z(n418) );
  MUX2_X1 U301 ( .A(product[2]), .B(n524), .S(n331), .Z(n420) );
  MUX2_X1 U302 ( .A(n524), .B(n525), .S(n331), .Z(n422) );
  INV_X1 U303 ( .A(n267), .ZN(n269) );
  NAND2_X1 U304 ( .A1(n269), .A2(n268), .ZN(n271) );
  XOR2_X1 U305 ( .A(n271), .B(n270), .Z(n272) );
  MUX2_X1 U306 ( .A(n525), .B(n272), .S(n331), .Z(n424) );
  MUX2_X1 U307 ( .A(product[3]), .B(n527), .S(n331), .Z(n426) );
  MUX2_X1 U308 ( .A(n527), .B(n528), .S(n331), .Z(n428) );
  NAND2_X1 U309 ( .A1(n274), .A2(n273), .ZN(n276) );
  XNOR2_X1 U310 ( .A(n276), .B(n275), .ZN(n277) );
  MUX2_X1 U311 ( .A(n528), .B(n277), .S(n331), .Z(n430) );
  MUX2_X1 U312 ( .A(product[4]), .B(n530), .S(n331), .Z(n432) );
  MUX2_X1 U313 ( .A(n530), .B(n531), .S(n331), .Z(n434) );
  INV_X1 U314 ( .A(n278), .ZN(n280) );
  NAND2_X1 U315 ( .A1(n280), .A2(n279), .ZN(n282) );
  XOR2_X1 U316 ( .A(n282), .B(n281), .Z(n283) );
  MUX2_X1 U317 ( .A(n531), .B(n283), .S(n331), .Z(n436) );
  MUX2_X1 U318 ( .A(product[5]), .B(n533), .S(n331), .Z(n438) );
  MUX2_X1 U319 ( .A(n533), .B(n534), .S(n331), .Z(n440) );
  NAND2_X1 U320 ( .A1(n285), .A2(n284), .ZN(n287) );
  XNOR2_X1 U321 ( .A(n287), .B(n286), .ZN(n288) );
  MUX2_X1 U322 ( .A(n534), .B(n288), .S(n331), .Z(n442) );
  MUX2_X1 U323 ( .A(product[6]), .B(n536), .S(n331), .Z(n444) );
  NAND2_X1 U324 ( .A1(n397), .A2(n347), .ZN(n289) );
  XOR2_X1 U325 ( .A(n289), .B(n352), .Z(n290) );
  MUX2_X1 U326 ( .A(n536), .B(n290), .S(n331), .Z(n446) );
  MUX2_X1 U327 ( .A(product[7]), .B(n538), .S(n331), .Z(n448) );
  OAI21_X1 U328 ( .B1(n346), .B2(n352), .A(n347), .ZN(n293) );
  NAND2_X1 U329 ( .A1(n336), .A2(n345), .ZN(n291) );
  XNOR2_X1 U330 ( .A(n293), .B(n291), .ZN(n292) );
  MUX2_X1 U331 ( .A(n538), .B(n292), .S(n331), .Z(n450) );
  MUX2_X1 U332 ( .A(product[8]), .B(n540), .S(n331), .Z(n452) );
  AOI21_X1 U333 ( .B1(n293), .B2(n336), .A(n398), .ZN(n296) );
  NAND2_X1 U334 ( .A1(n399), .A2(n344), .ZN(n294) );
  XOR2_X1 U335 ( .A(n296), .B(n294), .Z(n295) );
  MUX2_X1 U336 ( .A(n540), .B(n295), .S(n331), .Z(n454) );
  MUX2_X1 U337 ( .A(product[9]), .B(n542), .S(n331), .Z(n456) );
  OAI21_X1 U338 ( .B1(n296), .B2(n343), .A(n344), .ZN(n304) );
  INV_X1 U339 ( .A(n304), .ZN(n299) );
  NAND2_X1 U340 ( .A1(n400), .A2(n342), .ZN(n297) );
  XOR2_X1 U341 ( .A(n299), .B(n297), .Z(n298) );
  MUX2_X1 U342 ( .A(n542), .B(n298), .S(n331), .Z(n458) );
  MUX2_X1 U343 ( .A(product[10]), .B(n544), .S(n331), .Z(n460) );
  OAI21_X1 U344 ( .B1(n299), .B2(n341), .A(n342), .ZN(n301) );
  NAND2_X1 U345 ( .A1(n401), .A2(n349), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  MUX2_X1 U347 ( .A(n544), .B(n302), .S(n331), .Z(n462) );
  MUX2_X1 U348 ( .A(product[11]), .B(n546), .S(n331), .Z(n464) );
  NOR2_X1 U349 ( .A1(n348), .A2(n341), .ZN(n305) );
  OAI21_X1 U350 ( .B1(n348), .B2(n342), .A(n349), .ZN(n303) );
  AOI21_X1 U351 ( .B1(n305), .B2(n304), .A(n303), .ZN(n327) );
  NAND2_X1 U352 ( .A1(n402), .A2(n340), .ZN(n306) );
  XOR2_X1 U353 ( .A(n327), .B(n306), .Z(n307) );
  MUX2_X1 U354 ( .A(n546), .B(n307), .S(n331), .Z(n466) );
  MUX2_X1 U355 ( .A(product[12]), .B(n548), .S(n331), .Z(n468) );
  OAI21_X1 U356 ( .B1(n327), .B2(n351), .A(n340), .ZN(n309) );
  NAND2_X1 U357 ( .A1(n335), .A2(n339), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U359 ( .A(n548), .B(n310), .S(n331), .Z(n470) );
  MUX2_X1 U360 ( .A(product[13]), .B(n550), .S(n331), .Z(n472) );
  NAND2_X1 U361 ( .A1(n402), .A2(n335), .ZN(n312) );
  AOI21_X1 U362 ( .B1(n395), .B2(n335), .A(n403), .ZN(n311) );
  OAI21_X1 U363 ( .B1(n327), .B2(n312), .A(n311), .ZN(n314) );
  NAND2_X1 U364 ( .A1(n334), .A2(n350), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  MUX2_X1 U366 ( .A(n550), .B(n315), .S(n331), .Z(n474) );
  MUX2_X1 U367 ( .A(product[14]), .B(n552), .S(n331), .Z(n476) );
  NAND2_X1 U368 ( .A1(n335), .A2(n334), .ZN(n322) );
  OR2_X1 U369 ( .A1(n351), .A2(n322), .ZN(n318) );
  AOI21_X1 U370 ( .B1(n403), .B2(n334), .A(n394), .ZN(n316) );
  OAI21_X1 U371 ( .B1(n322), .B2(n340), .A(n316), .ZN(n324) );
  INV_X1 U372 ( .A(n324), .ZN(n317) );
  OAI21_X1 U373 ( .B1(n327), .B2(n318), .A(n317), .ZN(n320) );
  NAND2_X1 U374 ( .A1(n333), .A2(n338), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U376 ( .A(n552), .B(n321), .S(n331), .Z(n478) );
  MUX2_X1 U377 ( .A(product[15]), .B(n554), .S(n331), .Z(n480) );
  NOR2_X1 U378 ( .A1(n322), .A2(n396), .ZN(n323) );
  NAND2_X1 U379 ( .A1(n402), .A2(n323), .ZN(n326) );
  AOI21_X1 U380 ( .B1(n324), .B2(n333), .A(n393), .ZN(n325) );
  OAI21_X1 U381 ( .B1(n327), .B2(n326), .A(n325), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n328), .B(n337), .ZN(n329) );
  MUX2_X1 U383 ( .A(n554), .B(n329), .S(n331), .Z(n482) );
  MUX2_X1 U384 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n331), .Z(n484) );
  MUX2_X1 U385 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n331), .Z(n486) );
  MUX2_X1 U386 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n331), .Z(n488) );
  MUX2_X1 U387 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n331), .Z(n490) );
  MUX2_X1 U388 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n331), .Z(n492) );
  MUX2_X1 U389 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n331), .Z(n494) );
  MUX2_X1 U390 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n331), .Z(n496) );
  MUX2_X1 U391 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n331), .Z(n498) );
  MUX2_X1 U392 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n331), .Z(n500) );
  MUX2_X1 U393 ( .A(n555), .B(A_extended[1]), .S(n331), .Z(n502) );
  MUX2_X1 U394 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n331), .Z(n504) );
  MUX2_X1 U395 ( .A(n330), .B(A_extended[3]), .S(n331), .Z(n506) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n331), .Z(n508) );
  MUX2_X1 U397 ( .A(n6), .B(A_extended[5]), .S(n331), .Z(n510) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n331), .Z(n512) );
  MUX2_X1 U399 ( .A(n7), .B(A_extended[7]), .S(n331), .Z(n514) );
  OR2_X1 U400 ( .A1(n331), .A2(n558), .ZN(n516) );
endmodule


module conv_128_32_DW_mult_pipe_J1_22 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n361, n363, n365, n367, n369, n371, n373,
         n375, n377, n379, n381, n383, n385, n387, n389, n391, n393, n395,
         n397, n399, n401, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n415, n417, n419, n421, n423, n425, n427, n429,
         n431, n433, n435, n437, n439, n441, n443, n445, n447, n449, n451,
         n453, n455, n457, n459, n461, n463, n465, n467, n469, n471, n473,
         n475, n477, n479, n481, n483, n485, n487, n489, n491, n493, n495,
         n497, n499, n501, n503, n505, n507, n509, n511, n513, n515, n517,
         n519, n521, n523, n524, n526, n527, n529, n530, n532, n533, n535,
         n536, n538, n540, n542, n544, n546, n548, n550, n552, n554, n556,
         n558, n559, n560;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n411), .SE(n521), .CK(clk), .Q(n559), 
        .QN(n41) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n411), .SE(n517), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n28) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n411), .SE(n513), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n24) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n411), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n45) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n411), .SE(n509), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n46) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n411), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n43) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n411), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n34) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n411), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n39) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n412), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n40) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n413), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n35) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n411), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n36) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n411), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n38) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n411), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n37) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n411), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n411), .SE(n487), .CK(clk), .Q(n558)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n411), .SE(n485), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n411), .SE(n483), .CK(clk), .Q(n556)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n411), .SE(n481), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n411), .SE(n479), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n413), .SE(n477), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n411), .SE(n475), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n412), .SE(n473), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n411), .SE(n471), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n411), .SE(n469), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n411), .SE(n467), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n411), .SE(n465), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n411), .SE(n463), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n411), .SE(n461), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n411), .SE(n459), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n413), .SE(n457), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n413), .SE(n455), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n413), .SE(n453), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n413), .SE(n451), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n413), .SE(n449), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n413), .SE(n447), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n413), .SE(n445), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n413), .SE(n443), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n413), .SE(n441), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n413), .SE(n439), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n413), .SE(n437), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n412), .SE(n435), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n412), .SE(n433), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n412), .SE(n431), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n412), .SE(n429), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n412), .SE(n427), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n412), .SE(n425), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n412), .SE(n423), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n412), .SE(n421), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n412), .SE(n419), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n412), .SE(n417), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n412), .SE(n415), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2_IP  ( .D(1'b1), .SI(n560), .SE(n401), .CK(
        clk), .QN(n358) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n560), .SI(1'b1), .SE(n399), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n560), .SE(n397), .CK(
        clk), .QN(n356) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n560), .SI(1'b1), .SE(n395), .CK(clk), 
        .Q(n355) );
  SDFF_X1 \mult_x_1/clk_r_REG16_S2  ( .D(n560), .SI(1'b1), .SE(n393), .CK(clk), 
        .Q(n354) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2_IP  ( .D(1'b1), .SI(n560), .SE(n391), .CK(
        clk), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n560), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n352), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n560), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2_IP  ( .D(1'b1), .SI(n560), .SE(n385), .CK(
        clk), .Q(n403), .QN(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n560), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n560), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n560), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n347), .QN(n406) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n560), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n346), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n560), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n560), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n344), .QN(n408) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n560), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n343), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n560), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n342), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n560), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n341), .QN(n405) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n560), .SE(n365), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n560), .SE(n363), .CK(
        clk), .QN(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n560), .SI(1'b1), .SE(n361), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n560), .SI(1'b1), .SE(n359), .CK(clk), 
        .Q(n337) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n411), .SE(n519), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n335) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n411), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n48) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n411), .SE(n515), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n336) );
  INV_X1 U2 ( .A(n53), .ZN(n183) );
  XOR2_X1 U3 ( .A(n148), .B(n25), .Z(n5) );
  BUF_X1 U4 ( .A(n411), .Z(n412) );
  INV_X2 U5 ( .A(n560), .ZN(n411) );
  INV_X1 U6 ( .A(n6), .ZN(n240) );
  NAND2_X1 U7 ( .A1(n52), .A2(n92), .ZN(n182) );
  BUF_X1 U8 ( .A(\mult_x_1/n313 ), .Z(n23) );
  NAND2_X1 U9 ( .A1(n8), .A2(n7), .ZN(n226) );
  NAND2_X1 U10 ( .A1(n17), .A2(n16), .ZN(n194) );
  OAI21_X1 U11 ( .B1(n163), .B2(n162), .A(n10), .ZN(n8) );
  NAND2_X1 U12 ( .A1(n159), .A2(n18), .ZN(n17) );
  OR2_X1 U13 ( .A1(n161), .A2(n160), .ZN(n18) );
  NAND2_X1 U14 ( .A1(n161), .A2(n160), .ZN(n16) );
  NAND2_X1 U15 ( .A1(n163), .A2(n162), .ZN(n7) );
  BUF_X1 U16 ( .A(n411), .Z(n413) );
  OR2_X1 U17 ( .A1(n76), .A2(n75), .ZN(n60) );
  INV_X1 U18 ( .A(rst_n), .ZN(n560) );
  INV_X1 U19 ( .A(n218), .ZN(n172) );
  NAND2_X2 U20 ( .A1(n50), .A2(n51), .ZN(n174) );
  INV_X1 U21 ( .A(n68), .ZN(n6) );
  BUF_X2 U22 ( .A(\mult_x_1/n312 ), .Z(n25) );
  XNOR2_X1 U23 ( .A(\mult_x_1/n311 ), .B(n24), .ZN(n50) );
  XNOR2_X1 U24 ( .A(n9), .B(n163), .ZN(n145) );
  XNOR2_X1 U25 ( .A(n10), .B(n162), .ZN(n9) );
  NAND2_X1 U26 ( .A1(n11), .A2(n49), .ZN(n10) );
  NAND2_X1 U27 ( .A1(n78), .A2(n60), .ZN(n11) );
  NAND2_X1 U28 ( .A1(n154), .A2(n152), .ZN(n32) );
  NOR2_X1 U29 ( .A1(n13), .A2(n12), .ZN(n154) );
  NOR2_X1 U30 ( .A1(n172), .A2(n151), .ZN(n12) );
  NOR2_X1 U31 ( .A1(n174), .A2(n58), .ZN(n13) );
  XNOR2_X1 U32 ( .A(n161), .B(n160), .ZN(n19) );
  XNOR2_X1 U33 ( .A(n159), .B(n19), .ZN(n227) );
  NAND2_X1 U34 ( .A1(n15), .A2(n14), .ZN(n155) );
  INV_X1 U35 ( .A(n151), .ZN(n14) );
  NAND2_X1 U36 ( .A1(n174), .A2(n172), .ZN(n15) );
  NAND2_X1 U37 ( .A1(n21), .A2(n20), .ZN(n363) );
  NAND2_X1 U38 ( .A1(n97), .A2(n339), .ZN(n20) );
  OAI21_X1 U39 ( .B1(n201), .B2(n200), .A(n290), .ZN(n21) );
  XNOR2_X1 U40 ( .A(n153), .B(n22), .ZN(n30) );
  INV_X1 U41 ( .A(n152), .ZN(n22) );
  OAI22_X1 U42 ( .A1(n183), .A2(n150), .B1(n182), .B2(n54), .ZN(n153) );
  NAND2_X1 U43 ( .A1(n5), .A2(n6), .ZN(n29) );
  INV_X1 U44 ( .A(n136), .ZN(n71) );
  NOR2_X1 U45 ( .A1(n135), .A2(n134), .ZN(n70) );
  NAND2_X1 U46 ( .A1(n135), .A2(n134), .ZN(n69) );
  NAND2_X1 U47 ( .A1(n113), .A2(n112), .ZN(n108) );
  NAND2_X1 U48 ( .A1(n115), .A2(n107), .ZN(n109) );
  OR2_X1 U49 ( .A1(n113), .A2(n112), .ZN(n107) );
  XNOR2_X1 U50 ( .A(n336), .B(n28), .ZN(n92) );
  INV_X1 U51 ( .A(n27), .ZN(n67) );
  INV_X1 U52 ( .A(n86), .ZN(n64) );
  XNOR2_X1 U53 ( .A(n115), .B(n114), .ZN(n198) );
  XNOR2_X1 U54 ( .A(n113), .B(n112), .ZN(n114) );
  XNOR2_X1 U55 ( .A(n120), .B(n119), .ZN(n166) );
  INV_X1 U56 ( .A(n118), .ZN(n119) );
  OAI21_X1 U57 ( .B1(n71), .B2(n70), .A(n69), .ZN(n258) );
  OAI211_X1 U58 ( .C1(n128), .C2(n97), .A(n111), .B(n110), .ZN(n393) );
  NAND2_X1 U59 ( .A1(n263), .A2(n262), .ZN(n264) );
  NAND2_X1 U60 ( .A1(n44), .A2(n261), .ZN(n262) );
  OAI21_X1 U61 ( .B1(n44), .B2(n261), .A(n260), .ZN(n263) );
  XNOR2_X1 U62 ( .A(n24), .B(n45), .ZN(n51) );
  INV_X1 U63 ( .A(n335), .ZN(n26) );
  XNOR2_X1 U64 ( .A(n25), .B(n34), .ZN(n27) );
  NAND2_X1 U65 ( .A1(n29), .A2(n55), .ZN(n73) );
  XOR2_X1 U66 ( .A(n154), .B(n30), .Z(n163) );
  NAND2_X1 U67 ( .A1(n154), .A2(n153), .ZN(n31) );
  NAND2_X1 U68 ( .A1(n153), .A2(n152), .ZN(n33) );
  NAND3_X1 U69 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n161) );
  XNOR2_X1 U70 ( .A(n25), .B(n46), .ZN(n65) );
  BUF_X4 U71 ( .A(en), .Z(n334) );
  AND2_X1 U72 ( .A1(n109), .A2(n108), .ZN(n42) );
  AND2_X1 U73 ( .A1(n129), .A2(n130), .ZN(n44) );
  XOR2_X1 U74 ( .A(n130), .B(n129), .Z(n47) );
  NAND2_X1 U75 ( .A1(n76), .A2(n75), .ZN(n49) );
  XNOR2_X1 U76 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n58) );
  AND2_X1 U77 ( .A1(n559), .A2(\mult_x_1/n281 ), .ZN(n148) );
  XNOR2_X1 U78 ( .A(n148), .B(\mult_x_1/n311 ), .ZN(n151) );
  INV_X1 U79 ( .A(n51), .ZN(n218) );
  OAI22_X1 U80 ( .A1(n174), .A2(n58), .B1(n151), .B2(n172), .ZN(n156) );
  XOR2_X1 U81 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n52) );
  XNOR2_X1 U82 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n54) );
  INV_X1 U83 ( .A(n92), .ZN(n53) );
  XNOR2_X1 U84 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n150) );
  NAND2_X1 U85 ( .A1(n41), .A2(\mult_x_1/n310 ), .ZN(n95) );
  NOR2_X1 U86 ( .A1(n35), .A2(n95), .ZN(n152) );
  XNOR2_X1 U87 ( .A(n26), .B(\mult_x_1/n284 ), .ZN(n57) );
  OAI22_X1 U88 ( .A1(n182), .A2(n57), .B1(n183), .B2(n54), .ZN(n74) );
  XNOR2_X1 U89 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/a[2] ), .ZN(n68) );
  NAND3_X1 U90 ( .A1(n65), .A2(n68), .A3(n27), .ZN(n55) );
  NAND2_X1 U91 ( .A1(n65), .A2(n68), .ZN(n237) );
  NAND2_X1 U92 ( .A1(n240), .A2(n237), .ZN(n56) );
  NAND2_X1 U93 ( .A1(n56), .A2(n5), .ZN(n72) );
  INV_X1 U94 ( .A(n73), .ZN(n133) );
  XNOR2_X1 U95 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n63) );
  XNOR2_X1 U96 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n59) );
  OAI22_X1 U97 ( .A1(n174), .A2(n63), .B1(n51), .B2(n59), .ZN(n132) );
  XNOR2_X1 U98 ( .A(n26), .B(\mult_x_1/n285 ), .ZN(n62) );
  OAI22_X1 U99 ( .A1(n182), .A2(n62), .B1(n92), .B2(n57), .ZN(n131) );
  OAI22_X1 U100 ( .A1(n174), .A2(n59), .B1(n172), .B2(n58), .ZN(n76) );
  NOR2_X1 U101 ( .A1(n36), .A2(n95), .ZN(n75) );
  NAND2_X1 U102 ( .A1(n23), .A2(n43), .ZN(n242) );
  XNOR2_X1 U103 ( .A(n148), .B(n23), .ZN(n94) );
  AOI21_X1 U104 ( .B1(n242), .B2(n43), .A(n94), .ZN(n61) );
  INV_X1 U105 ( .A(n61), .ZN(n84) );
  XNOR2_X1 U106 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n91) );
  OAI22_X1 U107 ( .A1(n182), .A2(n91), .B1(n183), .B2(n62), .ZN(n83) );
  NOR2_X1 U108 ( .A1(n37), .A2(n95), .ZN(n82) );
  XNOR2_X1 U109 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n85) );
  OAI22_X1 U110 ( .A1(n174), .A2(n85), .B1(n172), .B2(n63), .ZN(n90) );
  XNOR2_X1 U111 ( .A(n25), .B(\mult_x_1/n282 ), .ZN(n86) );
  NAND3_X1 U112 ( .A1(n65), .A2(n68), .A3(n64), .ZN(n66) );
  OAI21_X1 U113 ( .B1(n68), .B2(n67), .A(n66), .ZN(n89) );
  OR2_X1 U114 ( .A1(n90), .A2(n89), .ZN(n135) );
  NOR2_X1 U115 ( .A1(n38), .A2(n95), .ZN(n134) );
  FA_X1 U116 ( .A(n74), .B(n73), .CI(n72), .CO(n162), .S(n257) );
  XOR2_X1 U117 ( .A(n76), .B(n75), .Z(n77) );
  XOR2_X1 U118 ( .A(n78), .B(n77), .Z(n256) );
  NAND2_X1 U119 ( .A1(n145), .A2(n144), .ZN(n79) );
  NAND2_X1 U120 ( .A1(n79), .A2(n334), .ZN(n81) );
  NAND2_X1 U121 ( .A1(n97), .A2(n342), .ZN(n80) );
  NAND2_X1 U122 ( .A1(n81), .A2(n80), .ZN(n369) );
  FA_X1 U123 ( .A(n84), .B(n83), .CI(n82), .CO(n136), .S(n140) );
  XNOR2_X1 U124 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n285 ), .ZN(n101) );
  OAI22_X1 U125 ( .A1(n174), .A2(n101), .B1(n172), .B2(n85), .ZN(n100) );
  XNOR2_X1 U126 ( .A(n25), .B(\mult_x_1/n283 ), .ZN(n103) );
  OAI22_X1 U127 ( .A1(n240), .A2(n86), .B1(n237), .B2(n103), .ZN(n99) );
  XNOR2_X1 U128 ( .A(n26), .B(\mult_x_1/n288 ), .ZN(n87) );
  XNOR2_X1 U129 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n93) );
  OAI22_X1 U130 ( .A1(n182), .A2(n87), .B1(n183), .B2(n93), .ZN(n120) );
  OR2_X1 U131 ( .A1(\mult_x_1/n288 ), .A2(n335), .ZN(n88) );
  OAI22_X1 U132 ( .A1(n183), .A2(n88), .B1(n182), .B2(n335), .ZN(n118) );
  AND2_X1 U133 ( .A1(n120), .A2(n118), .ZN(n98) );
  XNOR2_X1 U134 ( .A(n90), .B(n89), .ZN(n130) );
  OAI22_X1 U135 ( .A1(n182), .A2(n93), .B1(n183), .B2(n91), .ZN(n106) );
  XNOR2_X1 U136 ( .A(n23), .B(\mult_x_1/n281 ), .ZN(n102) );
  OAI22_X1 U137 ( .A1(n242), .A2(n102), .B1(n94), .B2(n43), .ZN(n105) );
  INV_X1 U138 ( .A(n95), .ZN(n96) );
  AND2_X1 U139 ( .A1(\mult_x_1/n288 ), .A2(n96), .ZN(n104) );
  INV_X1 U140 ( .A(en), .ZN(n97) );
  NAND2_X1 U141 ( .A1(n97), .A2(n354), .ZN(n111) );
  FA_X1 U142 ( .A(n100), .B(n99), .CI(n98), .CO(n139), .S(n115) );
  XNOR2_X1 U143 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n286 ), .ZN(n171) );
  OAI22_X1 U144 ( .A1(n174), .A2(n171), .B1(n172), .B2(n101), .ZN(n123) );
  XNOR2_X1 U145 ( .A(n23), .B(\mult_x_1/n282 ), .ZN(n116) );
  OAI22_X1 U146 ( .A1(n242), .A2(n116), .B1(n102), .B2(n43), .ZN(n122) );
  XNOR2_X1 U147 ( .A(n25), .B(\mult_x_1/n284 ), .ZN(n117) );
  OAI22_X1 U148 ( .A1(n240), .A2(n103), .B1(n237), .B2(n117), .ZN(n121) );
  FA_X1 U149 ( .A(n106), .B(n105), .CI(n104), .CO(n129), .S(n112) );
  NAND2_X1 U150 ( .A1(n42), .A2(n290), .ZN(n110) );
  XNOR2_X1 U151 ( .A(n23), .B(\mult_x_1/n283 ), .ZN(n207) );
  OAI22_X1 U152 ( .A1(n242), .A2(n207), .B1(n116), .B2(n43), .ZN(n177) );
  AND2_X1 U153 ( .A1(\mult_x_1/n288 ), .A2(n53), .ZN(n176) );
  XNOR2_X1 U154 ( .A(n25), .B(\mult_x_1/n285 ), .ZN(n206) );
  OAI22_X1 U155 ( .A1(n240), .A2(n117), .B1(n237), .B2(n206), .ZN(n175) );
  FA_X1 U156 ( .A(n123), .B(n122), .CI(n121), .CO(n113), .S(n165) );
  NAND2_X1 U157 ( .A1(n198), .A2(n197), .ZN(n124) );
  NAND2_X1 U158 ( .A1(n124), .A2(n290), .ZN(n126) );
  NAND2_X1 U159 ( .A1(n97), .A2(n345), .ZN(n125) );
  NAND2_X1 U160 ( .A1(n126), .A2(n125), .ZN(n375) );
  NAND2_X1 U161 ( .A1(n290), .A2(n42), .ZN(n127) );
  OAI22_X1 U162 ( .A1(n128), .A2(n127), .B1(n290), .B2(n409), .ZN(n371) );
  FA_X1 U163 ( .A(n131), .B(n132), .CI(n133), .CO(n78), .S(n261) );
  XNOR2_X1 U164 ( .A(n44), .B(n261), .ZN(n138) );
  XNOR2_X1 U165 ( .A(n135), .B(n134), .ZN(n137) );
  XNOR2_X1 U166 ( .A(n137), .B(n136), .ZN(n260) );
  XNOR2_X1 U167 ( .A(n138), .B(n260), .ZN(n224) );
  FA_X1 U168 ( .A(n140), .B(n139), .CI(n47), .CO(n223), .S(n128) );
  NAND2_X1 U169 ( .A1(n224), .A2(n223), .ZN(n141) );
  NAND2_X1 U170 ( .A1(n141), .A2(n290), .ZN(n143) );
  NAND2_X1 U171 ( .A1(n97), .A2(n353), .ZN(n142) );
  NAND2_X1 U172 ( .A1(n143), .A2(n142), .ZN(n391) );
  OAI21_X1 U173 ( .B1(n145), .B2(n144), .A(n290), .ZN(n147) );
  NAND2_X1 U174 ( .A1(n97), .A2(n351), .ZN(n146) );
  NAND2_X1 U175 ( .A1(n147), .A2(n146), .ZN(n387) );
  NOR2_X1 U198 ( .A1(n39), .A2(n95), .ZN(n180) );
  XNOR2_X1 U199 ( .A(n26), .B(\mult_x_1/n281 ), .ZN(n149) );
  XNOR2_X1 U200 ( .A(n148), .B(n26), .ZN(n181) );
  OAI22_X1 U201 ( .A1(n182), .A2(n149), .B1(n181), .B2(n183), .ZN(n188) );
  INV_X1 U202 ( .A(n188), .ZN(n179) );
  OAI22_X1 U203 ( .A1(n182), .A2(n150), .B1(n183), .B2(n149), .ZN(n157) );
  NOR2_X1 U204 ( .A1(n40), .A2(n95), .ZN(n160) );
  FA_X1 U205 ( .A(n157), .B(n156), .CI(n155), .CO(n178), .S(n159) );
  OR2_X1 U206 ( .A1(n195), .A2(n194), .ZN(n158) );
  MUX2_X1 U207 ( .A(n337), .B(n158), .S(n290), .Z(n359) );
  OR2_X1 U208 ( .A1(n226), .A2(n227), .ZN(n164) );
  MUX2_X1 U209 ( .A(n338), .B(n164), .S(en), .Z(n361) );
  FA_X1 U210 ( .A(n167), .B(n166), .CI(n165), .CO(n197), .S(n201) );
  INV_X1 U211 ( .A(\mult_x_1/n311 ), .ZN(n169) );
  OR2_X1 U212 ( .A1(\mult_x_1/n288 ), .A2(n169), .ZN(n168) );
  OAI22_X1 U213 ( .A1(n174), .A2(n169), .B1(n168), .B2(n172), .ZN(n209) );
  XNOR2_X1 U214 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n288 ), .ZN(n170) );
  XNOR2_X1 U215 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n173) );
  OAI22_X1 U216 ( .A1(n174), .A2(n170), .B1(n172), .B2(n173), .ZN(n208) );
  OAI22_X1 U217 ( .A1(n174), .A2(n173), .B1(n172), .B2(n171), .ZN(n204) );
  FA_X1 U218 ( .A(n177), .B(n176), .CI(n175), .CO(n167), .S(n203) );
  FA_X1 U219 ( .A(n180), .B(n179), .CI(n178), .CO(n190), .S(n195) );
  AOI21_X1 U220 ( .B1(n183), .B2(n182), .A(n181), .ZN(n184) );
  INV_X1 U221 ( .A(n184), .ZN(n186) );
  NOR2_X1 U222 ( .A1(n34), .A2(n95), .ZN(n185) );
  XOR2_X1 U223 ( .A(n186), .B(n185), .Z(n187) );
  XOR2_X1 U224 ( .A(n188), .B(n187), .Z(n189) );
  OR2_X1 U225 ( .A1(n190), .A2(n189), .ZN(n192) );
  NAND2_X1 U226 ( .A1(n190), .A2(n189), .ZN(n191) );
  NAND2_X1 U227 ( .A1(n192), .A2(n191), .ZN(n193) );
  MUX2_X1 U228 ( .A(n340), .B(n193), .S(en), .Z(n365) );
  NAND2_X1 U229 ( .A1(n195), .A2(n194), .ZN(n196) );
  MUX2_X1 U230 ( .A(n341), .B(n196), .S(n290), .Z(n367) );
  NOR2_X1 U231 ( .A1(n198), .A2(n197), .ZN(n199) );
  MUX2_X1 U232 ( .A(n344), .B(n199), .S(n290), .Z(n373) );
  NAND2_X1 U233 ( .A1(n201), .A2(n200), .ZN(n202) );
  MUX2_X1 U234 ( .A(n346), .B(n202), .S(n334), .Z(n377) );
  FA_X1 U235 ( .A(n205), .B(n204), .CI(n203), .CO(n200), .S(n212) );
  XNOR2_X1 U236 ( .A(n25), .B(\mult_x_1/n286 ), .ZN(n219) );
  OAI22_X1 U237 ( .A1(n240), .A2(n206), .B1(n237), .B2(n219), .ZN(n216) );
  XNOR2_X1 U238 ( .A(n23), .B(\mult_x_1/n284 ), .ZN(n217) );
  OAI22_X1 U239 ( .A1(n242), .A2(n217), .B1(n207), .B2(n43), .ZN(n215) );
  HA_X1 U240 ( .A(n209), .B(n208), .CO(n205), .S(n214) );
  NOR2_X1 U241 ( .A1(n212), .A2(n211), .ZN(n210) );
  MUX2_X1 U242 ( .A(n347), .B(n210), .S(n290), .Z(n379) );
  NAND2_X1 U243 ( .A1(n212), .A2(n211), .ZN(n213) );
  MUX2_X1 U244 ( .A(n348), .B(n213), .S(n334), .Z(n381) );
  FA_X1 U245 ( .A(n216), .B(n215), .CI(n214), .CO(n211), .S(n221) );
  XNOR2_X1 U246 ( .A(n23), .B(\mult_x_1/n285 ), .ZN(n234) );
  OAI22_X1 U247 ( .A1(n242), .A2(n234), .B1(n217), .B2(n43), .ZN(n231) );
  AND2_X1 U248 ( .A1(\mult_x_1/n288 ), .A2(n218), .ZN(n230) );
  XNOR2_X1 U249 ( .A(n25), .B(\mult_x_1/n287 ), .ZN(n233) );
  OAI22_X1 U250 ( .A1(n240), .A2(n219), .B1(n237), .B2(n233), .ZN(n229) );
  OR2_X1 U251 ( .A1(n221), .A2(n220), .ZN(n253) );
  NAND2_X1 U252 ( .A1(n221), .A2(n220), .ZN(n251) );
  NAND2_X1 U253 ( .A1(n253), .A2(n251), .ZN(n222) );
  MUX2_X1 U254 ( .A(n349), .B(n222), .S(n290), .Z(n383) );
  NOR2_X1 U255 ( .A1(n224), .A2(n223), .ZN(n225) );
  MUX2_X1 U256 ( .A(n350), .B(n225), .S(n290), .Z(n385) );
  NAND2_X1 U257 ( .A1(n227), .A2(n226), .ZN(n228) );
  MUX2_X1 U258 ( .A(n352), .B(n228), .S(n334), .Z(n389) );
  FA_X1 U259 ( .A(n231), .B(n230), .CI(n229), .CO(n220), .S(n250) );
  XNOR2_X1 U260 ( .A(n25), .B(\mult_x_1/n288 ), .ZN(n232) );
  OAI22_X1 U261 ( .A1(n240), .A2(n233), .B1(n237), .B2(n232), .ZN(n236) );
  XNOR2_X1 U262 ( .A(n23), .B(\mult_x_1/n286 ), .ZN(n239) );
  OAI22_X1 U263 ( .A1(n242), .A2(n239), .B1(n234), .B2(n43), .ZN(n235) );
  NOR2_X1 U264 ( .A1(n250), .A2(n249), .ZN(n281) );
  HA_X1 U265 ( .A(n236), .B(n235), .CO(n249), .S(n247) );
  OR2_X1 U266 ( .A1(\mult_x_1/n288 ), .A2(n45), .ZN(n238) );
  OAI22_X1 U267 ( .A1(n240), .A2(n238), .B1(n237), .B2(n45), .ZN(n246) );
  OR2_X1 U268 ( .A1(n247), .A2(n246), .ZN(n277) );
  XNOR2_X1 U269 ( .A(n23), .B(\mult_x_1/n287 ), .ZN(n241) );
  OAI22_X1 U270 ( .A1(n242), .A2(n241), .B1(n239), .B2(n43), .ZN(n245) );
  AND2_X1 U271 ( .A1(\mult_x_1/n288 ), .A2(n6), .ZN(n244) );
  NOR2_X1 U272 ( .A1(n245), .A2(n244), .ZN(n270) );
  OAI22_X1 U273 ( .A1(n242), .A2(\mult_x_1/n288 ), .B1(n241), .B2(n43), .ZN(
        n267) );
  OR2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(n48), .ZN(n243) );
  NAND2_X1 U275 ( .A1(n243), .A2(n242), .ZN(n266) );
  NAND2_X1 U276 ( .A1(n267), .A2(n266), .ZN(n273) );
  NAND2_X1 U277 ( .A1(n245), .A2(n244), .ZN(n271) );
  OAI21_X1 U278 ( .B1(n270), .B2(n273), .A(n271), .ZN(n278) );
  NAND2_X1 U279 ( .A1(n247), .A2(n246), .ZN(n276) );
  INV_X1 U280 ( .A(n276), .ZN(n248) );
  AOI21_X1 U281 ( .B1(n277), .B2(n278), .A(n248), .ZN(n284) );
  NAND2_X1 U282 ( .A1(n250), .A2(n249), .ZN(n282) );
  OAI21_X1 U283 ( .B1(n281), .B2(n284), .A(n282), .ZN(n255) );
  INV_X1 U284 ( .A(n251), .ZN(n252) );
  AOI21_X1 U285 ( .B1(n253), .B2(n255), .A(n252), .ZN(n254) );
  MUX2_X1 U286 ( .A(n355), .B(n254), .S(n290), .Z(n395) );
  MUX2_X1 U287 ( .A(n356), .B(n255), .S(n334), .Z(n397) );
  FA_X1 U288 ( .A(n258), .B(n257), .CI(n256), .CO(n144), .S(n259) );
  MUX2_X1 U289 ( .A(n357), .B(n259), .S(n290), .Z(n399) );
  MUX2_X1 U290 ( .A(n358), .B(n264), .S(n290), .Z(n401) );
  BUF_X4 U291 ( .A(en), .Z(n290) );
  MUX2_X1 U292 ( .A(product[0]), .B(n523), .S(n290), .Z(n415) );
  MUX2_X1 U293 ( .A(n523), .B(n524), .S(n290), .Z(n417) );
  AND2_X1 U294 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n265) );
  MUX2_X1 U295 ( .A(n524), .B(n265), .S(n290), .Z(n419) );
  MUX2_X1 U296 ( .A(product[1]), .B(n526), .S(n290), .Z(n421) );
  MUX2_X1 U297 ( .A(n526), .B(n527), .S(n290), .Z(n423) );
  OR2_X1 U298 ( .A1(n267), .A2(n266), .ZN(n268) );
  AND2_X1 U299 ( .A1(n268), .A2(n273), .ZN(n269) );
  MUX2_X1 U300 ( .A(n527), .B(n269), .S(n290), .Z(n425) );
  MUX2_X1 U301 ( .A(product[2]), .B(n529), .S(n290), .Z(n427) );
  MUX2_X1 U302 ( .A(n529), .B(n530), .S(n290), .Z(n429) );
  INV_X1 U303 ( .A(n270), .ZN(n272) );
  NAND2_X1 U304 ( .A1(n272), .A2(n271), .ZN(n274) );
  XOR2_X1 U305 ( .A(n274), .B(n273), .Z(n275) );
  MUX2_X1 U306 ( .A(n530), .B(n275), .S(n290), .Z(n431) );
  MUX2_X1 U307 ( .A(product[3]), .B(n532), .S(n290), .Z(n433) );
  MUX2_X1 U308 ( .A(n532), .B(n533), .S(n290), .Z(n435) );
  NAND2_X1 U309 ( .A1(n277), .A2(n276), .ZN(n279) );
  XNOR2_X1 U310 ( .A(n279), .B(n278), .ZN(n280) );
  MUX2_X1 U311 ( .A(n533), .B(n280), .S(n290), .Z(n437) );
  MUX2_X1 U312 ( .A(product[4]), .B(n535), .S(n290), .Z(n439) );
  MUX2_X1 U313 ( .A(n535), .B(n536), .S(n290), .Z(n441) );
  INV_X1 U314 ( .A(n281), .ZN(n283) );
  NAND2_X1 U315 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U316 ( .A(n285), .B(n284), .Z(n286) );
  MUX2_X1 U317 ( .A(n536), .B(n286), .S(n290), .Z(n443) );
  MUX2_X1 U318 ( .A(product[5]), .B(n538), .S(n290), .Z(n445) );
  XNOR2_X1 U319 ( .A(n349), .B(n356), .ZN(n287) );
  MUX2_X1 U320 ( .A(n538), .B(n287), .S(n290), .Z(n447) );
  MUX2_X1 U321 ( .A(product[6]), .B(n540), .S(n290), .Z(n449) );
  NAND2_X1 U322 ( .A1(n406), .A2(n348), .ZN(n288) );
  XOR2_X1 U323 ( .A(n288), .B(n355), .Z(n289) );
  MUX2_X1 U324 ( .A(n540), .B(n289), .S(n290), .Z(n451) );
  MUX2_X1 U325 ( .A(product[7]), .B(n542), .S(n290), .Z(n453) );
  OAI21_X1 U326 ( .B1(n347), .B2(n355), .A(n348), .ZN(n293) );
  NAND2_X1 U327 ( .A1(n339), .A2(n346), .ZN(n291) );
  XNOR2_X1 U328 ( .A(n293), .B(n291), .ZN(n292) );
  MUX2_X1 U329 ( .A(n542), .B(n292), .S(n334), .Z(n455) );
  MUX2_X1 U330 ( .A(product[8]), .B(n544), .S(n334), .Z(n457) );
  AOI21_X1 U331 ( .B1(n293), .B2(n339), .A(n407), .ZN(n296) );
  NAND2_X1 U332 ( .A1(n408), .A2(n345), .ZN(n294) );
  XOR2_X1 U333 ( .A(n296), .B(n294), .Z(n295) );
  MUX2_X1 U334 ( .A(n544), .B(n295), .S(n334), .Z(n459) );
  MUX2_X1 U335 ( .A(product[9]), .B(n546), .S(n334), .Z(n461) );
  OAI21_X1 U336 ( .B1(n296), .B2(n344), .A(n345), .ZN(n304) );
  INV_X1 U337 ( .A(n304), .ZN(n299) );
  NAND2_X1 U338 ( .A1(n409), .A2(n354), .ZN(n297) );
  XOR2_X1 U339 ( .A(n299), .B(n297), .Z(n298) );
  MUX2_X1 U340 ( .A(n546), .B(n298), .S(n334), .Z(n463) );
  MUX2_X1 U341 ( .A(product[10]), .B(n548), .S(n334), .Z(n465) );
  OAI21_X1 U342 ( .B1(n299), .B2(n343), .A(n354), .ZN(n301) );
  NAND2_X1 U343 ( .A1(n403), .A2(n353), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n302) );
  MUX2_X1 U345 ( .A(n548), .B(n302), .S(n334), .Z(n467) );
  MUX2_X1 U346 ( .A(product[11]), .B(n550), .S(n334), .Z(n469) );
  NOR2_X1 U347 ( .A1(n350), .A2(n343), .ZN(n305) );
  OAI21_X1 U348 ( .B1(n350), .B2(n354), .A(n353), .ZN(n303) );
  AOI21_X1 U349 ( .B1(n305), .B2(n304), .A(n303), .ZN(n331) );
  NOR2_X1 U350 ( .A1(n357), .A2(n358), .ZN(n318) );
  INV_X1 U351 ( .A(n318), .ZN(n311) );
  NAND2_X1 U352 ( .A1(n357), .A2(n358), .ZN(n320) );
  NAND2_X1 U353 ( .A1(n311), .A2(n320), .ZN(n306) );
  XOR2_X1 U354 ( .A(n331), .B(n306), .Z(n307) );
  MUX2_X1 U355 ( .A(n550), .B(n307), .S(n334), .Z(n471) );
  MUX2_X1 U356 ( .A(product[12]), .B(n552), .S(n334), .Z(n473) );
  OAI21_X1 U357 ( .B1(n331), .B2(n318), .A(n320), .ZN(n309) );
  NAND2_X1 U358 ( .A1(n351), .A2(n342), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  MUX2_X1 U360 ( .A(n552), .B(n310), .S(n334), .Z(n475) );
  MUX2_X1 U361 ( .A(product[13]), .B(n554), .S(n334), .Z(n477) );
  NAND2_X1 U362 ( .A1(n311), .A2(n351), .ZN(n314) );
  INV_X1 U363 ( .A(n320), .ZN(n312) );
  AOI21_X1 U364 ( .B1(n312), .B2(n351), .A(n410), .ZN(n313) );
  OAI21_X1 U365 ( .B1(n331), .B2(n314), .A(n313), .ZN(n316) );
  NAND2_X1 U366 ( .A1(n338), .A2(n352), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  MUX2_X1 U368 ( .A(n554), .B(n317), .S(n334), .Z(n479) );
  MUX2_X1 U369 ( .A(product[14]), .B(n556), .S(n334), .Z(n481) );
  NAND2_X1 U370 ( .A1(n351), .A2(n338), .ZN(n321) );
  NOR2_X1 U371 ( .A1(n318), .A2(n321), .ZN(n327) );
  INV_X1 U372 ( .A(n327), .ZN(n323) );
  AOI21_X1 U373 ( .B1(n410), .B2(n338), .A(n404), .ZN(n319) );
  OAI21_X1 U374 ( .B1(n321), .B2(n320), .A(n319), .ZN(n328) );
  INV_X1 U375 ( .A(n328), .ZN(n322) );
  OAI21_X1 U376 ( .B1(n331), .B2(n323), .A(n322), .ZN(n325) );
  NAND2_X1 U377 ( .A1(n337), .A2(n341), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  MUX2_X1 U379 ( .A(n556), .B(n326), .S(n334), .Z(n483) );
  MUX2_X1 U380 ( .A(product[15]), .B(n558), .S(n334), .Z(n485) );
  NAND2_X1 U381 ( .A1(n327), .A2(n337), .ZN(n330) );
  AOI21_X1 U382 ( .B1(n328), .B2(n337), .A(n405), .ZN(n329) );
  OAI21_X1 U383 ( .B1(n331), .B2(n330), .A(n329), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(n340), .ZN(n333) );
  MUX2_X1 U385 ( .A(n558), .B(n333), .S(n334), .Z(n487) );
  MUX2_X1 U386 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n334), .Z(n489) );
  MUX2_X1 U387 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n334), .Z(n491) );
  MUX2_X1 U388 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n334), .Z(n493) );
  MUX2_X1 U389 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n334), .Z(n495) );
  MUX2_X1 U390 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n334), .Z(n497) );
  MUX2_X1 U391 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n334), .Z(n499) );
  MUX2_X1 U392 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n334), .Z(n501) );
  MUX2_X1 U393 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n334), .Z(n503) );
  MUX2_X1 U394 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n334), .Z(n505) );
  MUX2_X1 U395 ( .A(n23), .B(A_extended[1]), .S(n334), .Z(n507) );
  MUX2_X1 U396 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n334), .Z(n509) );
  MUX2_X1 U397 ( .A(n25), .B(A_extended[3]), .S(n334), .Z(n511) );
  MUX2_X1 U398 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n334), .Z(n513) );
  MUX2_X1 U399 ( .A(\mult_x_1/n311 ), .B(A_extended[5]), .S(n334), .Z(n515) );
  MUX2_X1 U400 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n334), .Z(n517) );
  MUX2_X1 U401 ( .A(n26), .B(A_extended[7]), .S(n334), .Z(n519) );
  OR2_X1 U402 ( .A1(n334), .A2(n559), .ZN(n521) );
endmodule


module conv_128_32_DW_mult_pipe_J1_23 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n355,
         n357, n359, n361, n363, n365, n367, n369, n371, n373, n375, n377,
         n379, n381, n383, n385, n387, n389, n391, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n408,
         n410, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n442, n444, n446, n448, n450, n452,
         n454, n456, n458, n460, n462, n464, n466, n468, n470, n472, n474,
         n476, n478, n480, n482, n484, n486, n488, n490, n492, n494, n496,
         n498, n500, n502, n504, n506, n508, n510, n512, n514, n516, n518,
         n519, n521, n522, n524, n525, n527, n528, n530, n531, n533, n534,
         n536, n538, n540, n542, n544, n546, n548, n550, n552, n554, n555,
         n556, n557, n558, n559;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n406), .SE(n516), .CK(clk), .Q(n558), 
        .QN(n402) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n406), .SE(n514), .CK(clk), .Q(n557), 
        .QN(n403) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n406), .SE(n512), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n406), .SE(n510), .CK(clk), .Q(n556), 
        .QN(n35) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n406), .SE(n508), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n36) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n406), .SE(n504), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n37) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n406), .SE(n500), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n34) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n406), .SE(n498), .CK(clk), .Q(
        \mult_x_1/n281 ) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n406), .SE(n496), .CK(clk), .Q(
        \mult_x_1/n282 ) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n404), .SE(n494), .CK(clk), .Q(
        \mult_x_1/n283 ) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n405), .SE(n492), .CK(clk), .Q(
        \mult_x_1/n284 ) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n401), .SE(n490), .CK(clk), .Q(
        \mult_x_1/n285 ) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n406), .SE(n488), .CK(clk), .Q(
        \mult_x_1/n286 ) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n401), .SE(n486), .CK(clk), .Q(
        \mult_x_1/n287 ) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n401), .SE(n484), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n401), .SE(n482), .CK(clk), .Q(n554)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n401), .SE(n480), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n401), .SE(n478), .CK(clk), .Q(n552)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n401), .SE(n476), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n401), .SE(n474), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n405), .SE(n472), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n404), .SE(n470), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n406), .SE(n468), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n401), .SE(n466), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n401), .SE(n464), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n401), .SE(n462), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n401), .SE(n460), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n401), .SE(n458), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n401), .SE(n456), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n401), .SE(n454), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n401), .SE(n452), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n405), .SE(n450), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n405), .SE(n448), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n405), .SE(n446), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n405), .SE(n444), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n405), .SE(n442), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n405), .SE(n440), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n405), .SE(n438), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n405), .SE(n436), .CK(clk), .Q(n531)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n405), .SE(n434), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n405), .SE(n432), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n405), .SE(n430), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n404), .SE(n428), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n404), .SE(n426), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n404), .SE(n424), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n404), .SE(n422), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n404), .SE(n420), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n404), .SE(n418), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n404), .SE(n416), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n404), .SE(n414), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n404), .SE(n412), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n404), .SE(n410), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n404), .SE(n408), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n559), .SI(1'b1), .SE(n391), .CK(clk), 
        .Q(n352) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2  ( .D(n559), .SI(1'b1), .SE(n389), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n559), .SI(1'b1), .SE(n387), .CK(clk), 
        .Q(n350) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n559), .SI(1'b1), .SE(n385), .CK(clk), 
        .Q(n349), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n559), .SI(1'b1), .SE(n383), .CK(clk), 
        .Q(n348), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n559), .SI(1'b1), .SE(n381), .CK(clk), 
        .Q(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n559), .SI(1'b1), .SE(n379), .CK(clk), 
        .Q(n346), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n559), .SI(1'b1), .SE(n377), .CK(clk), 
        .Q(n345), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n559), .SI(1'b1), .SE(n375), .CK(clk), 
        .Q(n344), .QN(n39) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n559), .SI(1'b1), .SE(n373), .CK(clk), 
        .Q(n343), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n559), .SI(1'b1), .SE(n371), .CK(clk), 
        .Q(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n559), .SI(1'b1), .SE(n369), .CK(clk), 
        .Q(n341), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n559), .SI(1'b1), .SE(n367), .CK(clk), 
        .Q(n340), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n559), .SI(1'b1), .SE(n363), .CK(clk), 
        .Q(n338), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n559), .SE(n361), .CK(
        clk), .QN(n337) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n559), .SE(n359), .CK(
        clk), .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n559), .SI(1'b1), .SE(n357), .CK(clk), 
        .Q(n335), .QN(n38) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n559), .SI(1'b1), .SE(n355), .CK(clk), 
        .Q(n334) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n559), .SI(1'b1), .SE(n353), .CK(clk), 
        .Q(n333) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n406), .SE(n506), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n331) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n406), .SE(n502), .CK(clk), .Q(n555), 
        .QN(n40) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n559), .SE(n365), .CK(
        clk), .Q(n332), .QN(n339) );
  NAND2_X1 U2 ( .A1(n6), .A2(n5), .ZN(n212) );
  OAI21_X1 U3 ( .B1(n140), .B2(n139), .A(n138), .ZN(n6) );
  NAND2_X2 U4 ( .A1(n140), .A2(n139), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n209), .A2(n210), .ZN(n211) );
  XNOR2_X1 U6 ( .A(n7), .B(n140), .ZN(n210) );
  XNOR2_X1 U7 ( .A(n138), .B(n139), .ZN(n7) );
  AND2_X2 U8 ( .A1(n558), .A2(\mult_x_1/n281 ), .ZN(n121) );
  INV_X1 U9 ( .A(n330), .ZN(n8) );
  BUF_X1 U10 ( .A(n401), .Z(n405) );
  BUF_X1 U11 ( .A(n401), .Z(n404) );
  BUF_X1 U12 ( .A(n401), .Z(n406) );
  INV_X1 U13 ( .A(n559), .ZN(n401) );
  BUF_X4 U14 ( .A(en), .Z(n28) );
  BUF_X4 U15 ( .A(en), .Z(n330) );
  INV_X1 U16 ( .A(rst_n), .ZN(n559) );
  BUF_X1 U17 ( .A(n87), .Z(n161) );
  CLKBUF_X2 U18 ( .A(n70), .Z(n230) );
  INV_X1 U19 ( .A(n331), .ZN(n31) );
  INV_X1 U20 ( .A(n50), .ZN(n232) );
  INV_X2 U21 ( .A(n43), .ZN(n11) );
  INV_X1 U22 ( .A(n35), .ZN(n33) );
  BUF_X1 U23 ( .A(n555), .Z(n29) );
  NAND2_X1 U24 ( .A1(n34), .A2(n555), .ZN(n235) );
  OAI21_X1 U25 ( .B1(n13), .B2(n8), .A(n12), .ZN(n442) );
  NAND2_X1 U26 ( .A1(n8), .A2(n534), .ZN(n12) );
  XNOR2_X1 U27 ( .A(n284), .B(n14), .ZN(n13) );
  INV_X1 U28 ( .A(n283), .ZN(n14) );
  NAND2_X1 U29 ( .A1(n16), .A2(n15), .ZN(n183) );
  NAND2_X1 U30 ( .A1(n235), .A2(n34), .ZN(n15) );
  INV_X1 U31 ( .A(n84), .ZN(n16) );
  NAND2_X1 U32 ( .A1(n18), .A2(n17), .ZN(n389) );
  NAND2_X1 U33 ( .A1(n8), .A2(n351), .ZN(n17) );
  NAND2_X1 U34 ( .A1(n251), .A2(n330), .ZN(n18) );
  OAI22_X1 U35 ( .A1(n19), .A2(n119), .B1(n28), .B2(n332), .ZN(n365) );
  NAND2_X1 U36 ( .A1(n118), .A2(n28), .ZN(n19) );
  OR2_X1 U37 ( .A1(n255), .A2(n254), .ZN(n252) );
  XNOR2_X1 U38 ( .A(n109), .B(n110), .ZN(n249) );
  NAND2_X1 U39 ( .A1(n96), .A2(n95), .ZN(n357) );
  OR2_X1 U40 ( .A1(n28), .A2(n38), .ZN(n95) );
  OAI21_X1 U41 ( .B1(n210), .B2(n209), .A(n28), .ZN(n96) );
  NAND2_X1 U42 ( .A1(n255), .A2(n254), .ZN(n256) );
  NAND2_X1 U43 ( .A1(n253), .A2(n252), .ZN(n257) );
  XNOR2_X1 U44 ( .A(\mult_x_1/a[6] ), .B(n403), .ZN(n41) );
  INV_X1 U45 ( .A(n557), .ZN(n54) );
  XOR2_X1 U46 ( .A(n187), .B(n186), .Z(n20) );
  XOR2_X1 U47 ( .A(n185), .B(n20), .Z(n193) );
  NAND2_X1 U48 ( .A1(n185), .A2(n187), .ZN(n21) );
  NAND2_X1 U49 ( .A1(n185), .A2(n186), .ZN(n22) );
  NAND2_X1 U50 ( .A1(n187), .A2(n186), .ZN(n23) );
  NAND3_X1 U51 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n189) );
  OR2_X1 U52 ( .A1(n158), .A2(n56), .ZN(n24) );
  OR2_X1 U53 ( .A1(n11), .A2(n55), .ZN(n25) );
  NAND2_X1 U54 ( .A1(n24), .A2(n25), .ZN(n59) );
  INV_X1 U55 ( .A(n102), .ZN(n26) );
  NOR2_X2 U56 ( .A1(n403), .A2(n402), .ZN(n160) );
  NAND2_X1 U57 ( .A1(n41), .A2(n42), .ZN(n27) );
  NAND2_X1 U58 ( .A1(n41), .A2(n42), .ZN(n158) );
  OAI22_X1 U59 ( .A1(n230), .A2(n82), .B1(n232), .B2(n81), .ZN(n30) );
  INV_X1 U60 ( .A(n109), .ZN(n32) );
  XNOR2_X1 U61 ( .A(\mult_x_1/a[6] ), .B(n556), .ZN(n42) );
  XNOR2_X1 U62 ( .A(n557), .B(\mult_x_1/n287 ), .ZN(n55) );
  INV_X1 U63 ( .A(n42), .ZN(n43) );
  XNOR2_X1 U64 ( .A(n557), .B(\mult_x_1/n286 ), .ZN(n86) );
  OAI22_X1 U65 ( .A1(n27), .A2(n55), .B1(n11), .B2(n86), .ZN(n106) );
  XNOR2_X1 U66 ( .A(n29), .B(\mult_x_1/n281 ), .ZN(n47) );
  XNOR2_X1 U67 ( .A(n121), .B(n29), .ZN(n84) );
  OAI22_X1 U68 ( .A1(n235), .A2(n47), .B1(n84), .B2(n34), .ZN(n105) );
  XNOR2_X1 U69 ( .A(n54), .B(n160), .ZN(n67) );
  AND2_X1 U70 ( .A1(\mult_x_1/n288 ), .A2(n67), .ZN(n104) );
  XNOR2_X1 U71 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n45) );
  XNOR2_X1 U72 ( .A(n556), .B(n36), .ZN(n44) );
  NAND2_X1 U73 ( .A1(n45), .A2(n44), .ZN(n149) );
  XNOR2_X1 U74 ( .A(n33), .B(\mult_x_1/n286 ), .ZN(n147) );
  INV_X1 U75 ( .A(n45), .ZN(n46) );
  INV_X2 U76 ( .A(n46), .ZN(n219) );
  XNOR2_X1 U77 ( .A(n33), .B(\mult_x_1/n285 ), .ZN(n51) );
  OAI22_X1 U78 ( .A1(n149), .A2(n147), .B1(n219), .B2(n51), .ZN(n63) );
  XNOR2_X1 U79 ( .A(n29), .B(\mult_x_1/n282 ), .ZN(n57) );
  OAI22_X1 U80 ( .A1(n235), .A2(n57), .B1(n47), .B2(n34), .ZN(n62) );
  XOR2_X1 U81 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .Z(n49) );
  XNOR2_X1 U82 ( .A(n555), .B(n37), .ZN(n50) );
  INV_X1 U83 ( .A(n50), .ZN(n48) );
  NAND2_X1 U84 ( .A1(n49), .A2(n48), .ZN(n70) );
  XNOR2_X1 U85 ( .A(n31), .B(\mult_x_1/n284 ), .ZN(n58) );
  XNOR2_X1 U86 ( .A(n31), .B(\mult_x_1/n283 ), .ZN(n52) );
  OAI22_X1 U87 ( .A1(n230), .A2(n58), .B1(n232), .B2(n52), .ZN(n61) );
  XNOR2_X1 U88 ( .A(n33), .B(\mult_x_1/n284 ), .ZN(n80) );
  OAI22_X1 U89 ( .A1(n149), .A2(n51), .B1(n219), .B2(n80), .ZN(n180) );
  XNOR2_X1 U90 ( .A(n31), .B(\mult_x_1/n282 ), .ZN(n82) );
  OAI22_X1 U91 ( .A1(n230), .A2(n52), .B1(n232), .B2(n82), .ZN(n179) );
  OR2_X1 U92 ( .A1(\mult_x_1/n288 ), .A2(n54), .ZN(n53) );
  OAI22_X1 U93 ( .A1(n158), .A2(n54), .B1(n53), .B2(n11), .ZN(n60) );
  XNOR2_X1 U94 ( .A(n557), .B(\mult_x_1/n288 ), .ZN(n56) );
  XNOR2_X1 U95 ( .A(n29), .B(\mult_x_1/n283 ), .ZN(n202) );
  OAI22_X1 U96 ( .A1(n235), .A2(n202), .B1(n57), .B2(n34), .ZN(n152) );
  AND2_X1 U97 ( .A1(\mult_x_1/n288 ), .A2(n43), .ZN(n151) );
  XNOR2_X1 U98 ( .A(n31), .B(\mult_x_1/n285 ), .ZN(n201) );
  OAI22_X1 U99 ( .A1(n230), .A2(n201), .B1(n232), .B2(n58), .ZN(n150) );
  HA_X1 U100 ( .A(n60), .B(n59), .CO(n178), .S(n143) );
  FA_X1 U101 ( .A(n63), .B(n62), .CI(n61), .CO(n186), .S(n142) );
  NAND2_X1 U102 ( .A1(n193), .A2(n192), .ZN(n64) );
  NAND2_X1 U103 ( .A1(n64), .A2(n28), .ZN(n66) );
  OR2_X1 U104 ( .A1(n28), .A2(n39), .ZN(n65) );
  NAND2_X1 U105 ( .A1(n66), .A2(n65), .ZN(n375) );
  XNOR2_X1 U106 ( .A(n26), .B(\mult_x_1/n284 ), .ZN(n68) );
  INV_X1 U107 ( .A(n67), .ZN(n87) );
  NOR2_X1 U108 ( .A1(n68), .A2(n87), .ZN(n129) );
  XNOR2_X1 U109 ( .A(n557), .B(\mult_x_1/n283 ), .ZN(n69) );
  XNOR2_X1 U110 ( .A(n557), .B(\mult_x_1/n282 ), .ZN(n123) );
  OAI22_X1 U111 ( .A1(n27), .A2(n69), .B1(n11), .B2(n123), .ZN(n128) );
  XNOR2_X1 U112 ( .A(n33), .B(\mult_x_1/n281 ), .ZN(n74) );
  XNOR2_X1 U113 ( .A(n121), .B(n33), .ZN(n124) );
  OAI22_X1 U114 ( .A1(n149), .A2(n74), .B1(n124), .B2(n219), .ZN(n131) );
  INV_X1 U115 ( .A(n131), .ZN(n127) );
  XNOR2_X1 U116 ( .A(n557), .B(\mult_x_1/n284 ), .ZN(n76) );
  OAI22_X1 U117 ( .A1(n27), .A2(n76), .B1(n11), .B2(n69), .ZN(n91) );
  XNOR2_X1 U118 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n81) );
  XNOR2_X1 U119 ( .A(n121), .B(\mult_x_1/n312 ), .ZN(n71) );
  OAI22_X1 U120 ( .A1(n70), .A2(n81), .B1(n71), .B2(n232), .ZN(n90) );
  AOI21_X1 U121 ( .B1(n232), .B2(n230), .A(n71), .ZN(n72) );
  INV_X1 U122 ( .A(n72), .ZN(n89) );
  XNOR2_X1 U123 ( .A(n160), .B(\mult_x_1/n285 ), .ZN(n73) );
  NOR2_X1 U124 ( .A1(n73), .A2(n161), .ZN(n94) );
  XNOR2_X1 U125 ( .A(n33), .B(\mult_x_1/n282 ), .ZN(n75) );
  OAI22_X1 U126 ( .A1(n149), .A2(n75), .B1(n219), .B2(n74), .ZN(n93) );
  XNOR2_X1 U127 ( .A(n33), .B(\mult_x_1/n283 ), .ZN(n79) );
  OAI22_X1 U128 ( .A1(n149), .A2(n79), .B1(n219), .B2(n75), .ZN(n108) );
  XNOR2_X1 U129 ( .A(n557), .B(\mult_x_1/n285 ), .ZN(n85) );
  OAI22_X1 U130 ( .A1(n158), .A2(n85), .B1(n11), .B2(n76), .ZN(n107) );
  INV_X1 U131 ( .A(n90), .ZN(n109) );
  OAI21_X1 U132 ( .B1(n108), .B2(n107), .A(n109), .ZN(n78) );
  NAND2_X1 U133 ( .A1(n108), .A2(n107), .ZN(n77) );
  NAND2_X1 U134 ( .A1(n78), .A2(n77), .ZN(n92) );
  OAI22_X1 U135 ( .A1(n149), .A2(n80), .B1(n219), .B2(n79), .ZN(n101) );
  OAI22_X1 U136 ( .A1(n230), .A2(n82), .B1(n232), .B2(n81), .ZN(n100) );
  OR2_X1 U137 ( .A1(n101), .A2(n30), .ZN(n113) );
  XNOR2_X1 U138 ( .A(n26), .B(\mult_x_1/n286 ), .ZN(n83) );
  NOR2_X1 U139 ( .A1(n83), .A2(n161), .ZN(n112) );
  OAI22_X1 U140 ( .A1(n158), .A2(n86), .B1(n11), .B2(n85), .ZN(n182) );
  XNOR2_X1 U141 ( .A(n160), .B(\mult_x_1/n287 ), .ZN(n88) );
  NOR2_X1 U142 ( .A1(n88), .A2(n87), .ZN(n181) );
  FA_X1 U143 ( .A(n91), .B(n32), .CI(n89), .CO(n139), .S(n98) );
  FA_X1 U144 ( .A(n94), .B(n93), .CI(n92), .CO(n138), .S(n97) );
  FA_X1 U145 ( .A(n99), .B(n98), .CI(n97), .CO(n209), .S(n119) );
  INV_X1 U146 ( .A(n28), .ZN(n117) );
  OR2_X1 U147 ( .A1(n28), .A2(n394), .ZN(n116) );
  XNOR2_X1 U148 ( .A(n101), .B(n100), .ZN(n177) );
  INV_X1 U149 ( .A(n160), .ZN(n102) );
  OR2_X1 U150 ( .A1(\mult_x_1/n288 ), .A2(n102), .ZN(n103) );
  NOR2_X1 U151 ( .A1(n103), .A2(n161), .ZN(n176) );
  FA_X1 U152 ( .A(n106), .B(n105), .CI(n104), .CO(n175), .S(n187) );
  XNOR2_X1 U153 ( .A(n108), .B(n107), .ZN(n110) );
  FA_X1 U154 ( .A(n113), .B(n112), .CI(n111), .CO(n99), .S(n248) );
  INV_X1 U155 ( .A(n114), .ZN(n118) );
  NAND2_X1 U156 ( .A1(n118), .A2(n28), .ZN(n115) );
  OAI211_X1 U157 ( .C1(n119), .C2(n117), .A(n116), .B(n115), .ZN(n367) );
  XNOR2_X1 U178 ( .A(n26), .B(\mult_x_1/n282 ), .ZN(n120) );
  NOR2_X1 U179 ( .A1(n120), .A2(n161), .ZN(n156) );
  XNOR2_X1 U180 ( .A(n557), .B(\mult_x_1/n281 ), .ZN(n122) );
  XNOR2_X1 U181 ( .A(n121), .B(n557), .ZN(n157) );
  OAI22_X1 U182 ( .A1(n27), .A2(n122), .B1(n157), .B2(n11), .ZN(n166) );
  INV_X1 U183 ( .A(n166), .ZN(n155) );
  OAI22_X1 U184 ( .A1(n27), .A2(n123), .B1(n11), .B2(n122), .ZN(n133) );
  INV_X1 U185 ( .A(n124), .ZN(n126) );
  NAND2_X1 U186 ( .A1(n219), .A2(n149), .ZN(n125) );
  NAND2_X1 U187 ( .A1(n126), .A2(n125), .ZN(n132) );
  FA_X1 U188 ( .A(n129), .B(n128), .CI(n127), .CO(n137), .S(n140) );
  XNOR2_X1 U189 ( .A(n26), .B(\mult_x_1/n283 ), .ZN(n130) );
  NOR2_X1 U190 ( .A1(n130), .A2(n161), .ZN(n136) );
  FA_X1 U191 ( .A(n133), .B(n132), .CI(n131), .CO(n154), .S(n135) );
  OR2_X1 U192 ( .A1(n173), .A2(n172), .ZN(n134) );
  MUX2_X1 U193 ( .A(n333), .B(n134), .S(n28), .Z(n353) );
  FA_X1 U194 ( .A(n137), .B(n136), .CI(n135), .CO(n172), .S(n213) );
  OR2_X1 U195 ( .A1(n213), .A2(n212), .ZN(n141) );
  MUX2_X1 U196 ( .A(n334), .B(n141), .S(n28), .Z(n355) );
  FA_X1 U197 ( .A(n144), .B(n143), .CI(n142), .CO(n192), .S(n196) );
  OR2_X1 U198 ( .A1(\mult_x_1/n288 ), .A2(n35), .ZN(n145) );
  OAI22_X1 U199 ( .A1(n149), .A2(n35), .B1(n145), .B2(n219), .ZN(n204) );
  XNOR2_X1 U200 ( .A(n33), .B(\mult_x_1/n288 ), .ZN(n146) );
  XNOR2_X1 U201 ( .A(n33), .B(\mult_x_1/n287 ), .ZN(n148) );
  OAI22_X1 U202 ( .A1(n149), .A2(n146), .B1(n219), .B2(n148), .ZN(n203) );
  OAI22_X1 U203 ( .A1(n149), .A2(n148), .B1(n219), .B2(n147), .ZN(n199) );
  FA_X1 U204 ( .A(n152), .B(n151), .CI(n150), .CO(n144), .S(n198) );
  OR2_X1 U205 ( .A1(n196), .A2(n195), .ZN(n153) );
  MUX2_X1 U206 ( .A(n336), .B(n153), .S(n28), .Z(n359) );
  FA_X1 U207 ( .A(n156), .B(n155), .CI(n154), .CO(n168), .S(n173) );
  AOI21_X1 U208 ( .B1(n11), .B2(n27), .A(n157), .ZN(n159) );
  INV_X1 U209 ( .A(n159), .ZN(n164) );
  XNOR2_X1 U210 ( .A(n26), .B(\mult_x_1/n281 ), .ZN(n162) );
  NOR2_X1 U211 ( .A1(n162), .A2(n161), .ZN(n163) );
  XOR2_X1 U212 ( .A(n164), .B(n163), .Z(n165) );
  XOR2_X1 U213 ( .A(n166), .B(n165), .Z(n167) );
  OR2_X1 U214 ( .A1(n168), .A2(n167), .ZN(n170) );
  NAND2_X1 U215 ( .A1(n168), .A2(n167), .ZN(n169) );
  NAND2_X1 U216 ( .A1(n170), .A2(n169), .ZN(n171) );
  MUX2_X1 U217 ( .A(n337), .B(n171), .S(n28), .Z(n361) );
  NAND2_X1 U218 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2_X1 U219 ( .A(n338), .B(n174), .S(n28), .Z(n363) );
  FA_X1 U220 ( .A(n177), .B(n176), .CI(n175), .CO(n250), .S(n253) );
  FA_X1 U221 ( .A(n180), .B(n179), .CI(n178), .CO(n254), .S(n185) );
  FA_X1 U222 ( .A(n183), .B(n182), .CI(n181), .CO(n111), .S(n255) );
  XNOR2_X1 U223 ( .A(n254), .B(n255), .ZN(n184) );
  XNOR2_X1 U224 ( .A(n253), .B(n184), .ZN(n190) );
  NOR2_X1 U225 ( .A1(n190), .A2(n189), .ZN(n188) );
  MUX2_X1 U226 ( .A(n341), .B(n188), .S(n28), .Z(n369) );
  NAND2_X1 U227 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U228 ( .A(n342), .B(n191), .S(n28), .Z(n371) );
  NOR2_X1 U229 ( .A1(n193), .A2(n192), .ZN(n194) );
  MUX2_X1 U230 ( .A(n343), .B(n194), .S(n28), .Z(n373) );
  NAND2_X1 U231 ( .A1(n196), .A2(n195), .ZN(n197) );
  MUX2_X1 U232 ( .A(n345), .B(n197), .S(n28), .Z(n377) );
  FA_X1 U233 ( .A(n200), .B(n199), .CI(n198), .CO(n195), .S(n207) );
  XNOR2_X1 U234 ( .A(n31), .B(\mult_x_1/n286 ), .ZN(n220) );
  OAI22_X1 U235 ( .A1(n230), .A2(n220), .B1(n232), .B2(n201), .ZN(n217) );
  XNOR2_X1 U236 ( .A(n29), .B(\mult_x_1/n284 ), .ZN(n218) );
  OAI22_X1 U237 ( .A1(n235), .A2(n218), .B1(n202), .B2(n34), .ZN(n216) );
  HA_X1 U238 ( .A(n204), .B(n203), .CO(n200), .S(n215) );
  NOR2_X1 U239 ( .A1(n207), .A2(n206), .ZN(n205) );
  MUX2_X1 U240 ( .A(n346), .B(n205), .S(n330), .Z(n379) );
  NAND2_X1 U241 ( .A1(n207), .A2(n206), .ZN(n208) );
  MUX2_X1 U242 ( .A(n347), .B(n208), .S(n28), .Z(n381) );
  MUX2_X1 U243 ( .A(n348), .B(n211), .S(n330), .Z(n383) );
  NAND2_X1 U244 ( .A1(n213), .A2(n212), .ZN(n214) );
  MUX2_X1 U245 ( .A(n349), .B(n214), .S(n330), .Z(n385) );
  FA_X1 U246 ( .A(n217), .B(n216), .CI(n215), .CO(n206), .S(n245) );
  XNOR2_X1 U247 ( .A(n29), .B(\mult_x_1/n285 ), .ZN(n226) );
  OAI22_X1 U248 ( .A1(n235), .A2(n226), .B1(n218), .B2(n34), .ZN(n223) );
  AND2_X1 U249 ( .A1(\mult_x_1/n288 ), .A2(n46), .ZN(n222) );
  XNOR2_X1 U250 ( .A(n31), .B(\mult_x_1/n287 ), .ZN(n224) );
  OAI22_X1 U251 ( .A1(n230), .A2(n224), .B1(n232), .B2(n220), .ZN(n221) );
  OR2_X1 U252 ( .A1(n245), .A2(n244), .ZN(n282) );
  FA_X1 U253 ( .A(n223), .B(n222), .CI(n221), .CO(n244), .S(n243) );
  XNOR2_X1 U254 ( .A(n31), .B(\mult_x_1/n288 ), .ZN(n225) );
  OAI22_X1 U255 ( .A1(n230), .A2(n225), .B1(n232), .B2(n224), .ZN(n228) );
  XNOR2_X1 U256 ( .A(n29), .B(\mult_x_1/n286 ), .ZN(n231) );
  OAI22_X1 U257 ( .A1(n235), .A2(n231), .B1(n226), .B2(n34), .ZN(n227) );
  NOR2_X1 U258 ( .A1(n243), .A2(n242), .ZN(n275) );
  HA_X1 U259 ( .A(n228), .B(n227), .CO(n242), .S(n240) );
  OR2_X1 U260 ( .A1(\mult_x_1/n288 ), .A2(n331), .ZN(n229) );
  OAI22_X1 U261 ( .A1(n230), .A2(n331), .B1(n229), .B2(n232), .ZN(n239) );
  OR2_X1 U262 ( .A1(n240), .A2(n239), .ZN(n271) );
  XNOR2_X1 U263 ( .A(n29), .B(\mult_x_1/n287 ), .ZN(n234) );
  OAI22_X1 U264 ( .A1(n235), .A2(n234), .B1(n231), .B2(n34), .ZN(n238) );
  INV_X1 U265 ( .A(n232), .ZN(n233) );
  AND2_X1 U266 ( .A1(\mult_x_1/n288 ), .A2(n233), .ZN(n237) );
  NOR2_X1 U267 ( .A1(n238), .A2(n237), .ZN(n264) );
  OAI22_X1 U268 ( .A1(n235), .A2(\mult_x_1/n288 ), .B1(n234), .B2(n34), .ZN(
        n261) );
  OR2_X1 U269 ( .A1(\mult_x_1/n288 ), .A2(n40), .ZN(n236) );
  NAND2_X1 U270 ( .A1(n236), .A2(n235), .ZN(n260) );
  NAND2_X1 U271 ( .A1(n261), .A2(n260), .ZN(n267) );
  NAND2_X1 U272 ( .A1(n238), .A2(n237), .ZN(n265) );
  OAI21_X1 U273 ( .B1(n264), .B2(n267), .A(n265), .ZN(n272) );
  NAND2_X1 U274 ( .A1(n240), .A2(n239), .ZN(n270) );
  INV_X1 U275 ( .A(n270), .ZN(n241) );
  AOI21_X1 U276 ( .B1(n271), .B2(n272), .A(n241), .ZN(n278) );
  NAND2_X1 U277 ( .A1(n243), .A2(n242), .ZN(n276) );
  OAI21_X1 U278 ( .B1(n275), .B2(n278), .A(n276), .ZN(n283) );
  NAND2_X1 U279 ( .A1(n245), .A2(n244), .ZN(n281) );
  INV_X1 U280 ( .A(n281), .ZN(n246) );
  AOI21_X1 U281 ( .B1(n282), .B2(n283), .A(n246), .ZN(n247) );
  MUX2_X1 U282 ( .A(n350), .B(n247), .S(n28), .Z(n387) );
  FA_X1 U283 ( .A(n250), .B(n249), .CI(n248), .CO(n114), .S(n251) );
  NAND2_X1 U284 ( .A1(n257), .A2(n256), .ZN(n258) );
  MUX2_X1 U285 ( .A(n352), .B(n258), .S(n330), .Z(n391) );
  MUX2_X1 U286 ( .A(product[0]), .B(n518), .S(n330), .Z(n408) );
  MUX2_X1 U287 ( .A(n518), .B(n519), .S(n330), .Z(n410) );
  AND2_X1 U288 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n259) );
  MUX2_X1 U289 ( .A(n519), .B(n259), .S(n28), .Z(n412) );
  MUX2_X1 U290 ( .A(product[1]), .B(n521), .S(n330), .Z(n414) );
  MUX2_X1 U291 ( .A(n521), .B(n522), .S(n330), .Z(n416) );
  OR2_X1 U292 ( .A1(n261), .A2(n260), .ZN(n262) );
  AND2_X1 U293 ( .A1(n262), .A2(n267), .ZN(n263) );
  MUX2_X1 U294 ( .A(n522), .B(n263), .S(n28), .Z(n418) );
  MUX2_X1 U295 ( .A(product[2]), .B(n524), .S(n330), .Z(n420) );
  MUX2_X1 U296 ( .A(n524), .B(n525), .S(n330), .Z(n422) );
  INV_X1 U297 ( .A(n264), .ZN(n266) );
  NAND2_X1 U298 ( .A1(n266), .A2(n265), .ZN(n268) );
  XOR2_X1 U299 ( .A(n268), .B(n267), .Z(n269) );
  MUX2_X1 U300 ( .A(n525), .B(n269), .S(n28), .Z(n424) );
  MUX2_X1 U301 ( .A(product[3]), .B(n527), .S(n330), .Z(n426) );
  MUX2_X1 U302 ( .A(n527), .B(n528), .S(n330), .Z(n428) );
  NAND2_X1 U303 ( .A1(n271), .A2(n270), .ZN(n273) );
  XNOR2_X1 U304 ( .A(n273), .B(n272), .ZN(n274) );
  MUX2_X1 U305 ( .A(n528), .B(n274), .S(n28), .Z(n430) );
  MUX2_X1 U306 ( .A(product[4]), .B(n530), .S(n330), .Z(n432) );
  MUX2_X1 U307 ( .A(n530), .B(n531), .S(n28), .Z(n434) );
  INV_X1 U308 ( .A(n275), .ZN(n277) );
  NAND2_X1 U309 ( .A1(n277), .A2(n276), .ZN(n279) );
  XOR2_X1 U310 ( .A(n279), .B(n278), .Z(n280) );
  MUX2_X1 U311 ( .A(n531), .B(n280), .S(n330), .Z(n436) );
  MUX2_X1 U312 ( .A(product[5]), .B(n533), .S(n330), .Z(n438) );
  MUX2_X1 U313 ( .A(n533), .B(n534), .S(n28), .Z(n440) );
  NAND2_X1 U314 ( .A1(n282), .A2(n281), .ZN(n284) );
  MUX2_X1 U315 ( .A(product[6]), .B(n536), .S(n330), .Z(n444) );
  NAND2_X1 U316 ( .A1(n395), .A2(n347), .ZN(n285) );
  XOR2_X1 U317 ( .A(n285), .B(n350), .Z(n286) );
  MUX2_X1 U318 ( .A(n536), .B(n286), .S(n28), .Z(n446) );
  MUX2_X1 U319 ( .A(product[7]), .B(n538), .S(n330), .Z(n448) );
  OAI21_X1 U320 ( .B1(n346), .B2(n350), .A(n347), .ZN(n289) );
  NAND2_X1 U321 ( .A1(n336), .A2(n345), .ZN(n287) );
  XNOR2_X1 U322 ( .A(n289), .B(n287), .ZN(n288) );
  MUX2_X1 U323 ( .A(n538), .B(n288), .S(n330), .Z(n450) );
  MUX2_X1 U324 ( .A(product[8]), .B(n540), .S(n28), .Z(n452) );
  AOI21_X1 U325 ( .B1(n289), .B2(n336), .A(n397), .ZN(n292) );
  NAND2_X1 U326 ( .A1(n398), .A2(n344), .ZN(n290) );
  XOR2_X1 U327 ( .A(n292), .B(n290), .Z(n291) );
  MUX2_X1 U328 ( .A(n540), .B(n291), .S(n330), .Z(n454) );
  MUX2_X1 U329 ( .A(product[9]), .B(n542), .S(n330), .Z(n456) );
  OAI21_X1 U330 ( .B1(n292), .B2(n343), .A(n344), .ZN(n303) );
  INV_X1 U331 ( .A(n303), .ZN(n295) );
  NAND2_X1 U332 ( .A1(n399), .A2(n342), .ZN(n293) );
  XOR2_X1 U333 ( .A(n295), .B(n293), .Z(n294) );
  MUX2_X1 U334 ( .A(n542), .B(n294), .S(n330), .Z(n458) );
  MUX2_X1 U335 ( .A(product[10]), .B(n544), .S(n330), .Z(n460) );
  OAI21_X1 U336 ( .B1(n295), .B2(n341), .A(n342), .ZN(n298) );
  NOR2_X1 U337 ( .A1(n351), .A2(n352), .ZN(n301) );
  INV_X1 U338 ( .A(n301), .ZN(n296) );
  NAND2_X1 U339 ( .A1(n351), .A2(n352), .ZN(n300) );
  NAND2_X1 U340 ( .A1(n296), .A2(n300), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  MUX2_X1 U342 ( .A(n544), .B(n299), .S(n28), .Z(n462) );
  MUX2_X1 U343 ( .A(product[11]), .B(n546), .S(n28), .Z(n464) );
  NOR2_X1 U344 ( .A1(n301), .A2(n341), .ZN(n304) );
  OAI21_X1 U345 ( .B1(n301), .B2(n342), .A(n300), .ZN(n302) );
  AOI21_X1 U346 ( .B1(n304), .B2(n303), .A(n302), .ZN(n326) );
  NAND2_X1 U347 ( .A1(n332), .A2(n340), .ZN(n305) );
  XOR2_X1 U348 ( .A(n326), .B(n305), .Z(n306) );
  MUX2_X1 U349 ( .A(n546), .B(n306), .S(n28), .Z(n466) );
  MUX2_X1 U350 ( .A(product[12]), .B(n548), .S(n330), .Z(n468) );
  OAI21_X1 U351 ( .B1(n326), .B2(n339), .A(n340), .ZN(n308) );
  NAND2_X1 U352 ( .A1(n335), .A2(n348), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  MUX2_X1 U354 ( .A(n548), .B(n309), .S(n330), .Z(n470) );
  MUX2_X1 U355 ( .A(product[13]), .B(n550), .S(n28), .Z(n472) );
  NAND2_X1 U356 ( .A1(n332), .A2(n335), .ZN(n311) );
  AOI21_X1 U357 ( .B1(n394), .B2(n335), .A(n400), .ZN(n310) );
  OAI21_X1 U358 ( .B1(n326), .B2(n311), .A(n310), .ZN(n313) );
  NAND2_X1 U359 ( .A1(n334), .A2(n349), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  MUX2_X1 U361 ( .A(n550), .B(n314), .S(n330), .Z(n474) );
  MUX2_X1 U362 ( .A(product[14]), .B(n552), .S(n330), .Z(n476) );
  NAND2_X1 U363 ( .A1(n335), .A2(n334), .ZN(n316) );
  NOR2_X1 U364 ( .A1(n339), .A2(n316), .ZN(n322) );
  INV_X1 U365 ( .A(n322), .ZN(n318) );
  AOI21_X1 U366 ( .B1(n400), .B2(n334), .A(n396), .ZN(n315) );
  OAI21_X1 U367 ( .B1(n316), .B2(n340), .A(n315), .ZN(n323) );
  INV_X1 U368 ( .A(n323), .ZN(n317) );
  OAI21_X1 U369 ( .B1(n326), .B2(n318), .A(n317), .ZN(n320) );
  NAND2_X1 U370 ( .A1(n333), .A2(n338), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  MUX2_X1 U372 ( .A(n552), .B(n321), .S(n28), .Z(n478) );
  MUX2_X1 U373 ( .A(product[15]), .B(n554), .S(n330), .Z(n480) );
  NAND2_X1 U374 ( .A1(n322), .A2(n333), .ZN(n325) );
  AOI21_X1 U375 ( .B1(n323), .B2(n333), .A(n393), .ZN(n324) );
  OAI21_X1 U376 ( .B1(n326), .B2(n325), .A(n324), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n327), .B(n337), .ZN(n328) );
  MUX2_X1 U378 ( .A(n554), .B(n328), .S(n330), .Z(n482) );
  MUX2_X1 U379 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n28), .Z(n484) );
  MUX2_X1 U380 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n330), .Z(n486) );
  MUX2_X1 U381 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n28), .Z(n488) );
  MUX2_X1 U382 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n330), .Z(n490) );
  MUX2_X1 U383 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n330), .Z(n492) );
  MUX2_X1 U384 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n28), .Z(n494) );
  MUX2_X1 U385 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n330), .Z(n496) );
  MUX2_X1 U386 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n330), .Z(n498) );
  MUX2_X1 U387 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n28), .Z(n500) );
  MUX2_X1 U388 ( .A(n29), .B(A_extended[1]), .S(n330), .Z(n502) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n28), .Z(n504) );
  MUX2_X1 U390 ( .A(n31), .B(A_extended[3]), .S(n330), .Z(n506) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n28), .Z(n508) );
  MUX2_X1 U392 ( .A(n33), .B(A_extended[5]), .S(n28), .Z(n510) );
  MUX2_X1 U393 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n28), .Z(n512) );
  MUX2_X1 U394 ( .A(n557), .B(A_extended[7]), .S(n330), .Z(n514) );
  OR2_X1 U395 ( .A1(n28), .A2(n558), .ZN(n516) );
endmodule


module conv_128_32_DW_mult_pipe_J1_24 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n310 ,
         \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 ,
         \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 ,
         \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n360, n362, n364, n366, n368, n370,
         n372, n374, n376, n378, n380, n382, n384, n386, n388, n390, n392,
         n394, n396, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n415, n417, n419, n421, n423,
         n425, n427, n429, n431, n433, n435, n437, n439, n441, n443, n445,
         n447, n449, n451, n453, n455, n457, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n515, n517, n519, n521, n523, n524, n526, n527, n529, n530,
         n532, n533, n535, n536, n538, n539, n541, n543, n545, n547, n549,
         n551, n553, n555, n557, n559, n560, n561, n562, n563, n564;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n411), .SE(n521), .CK(clk), .Q(n563)
         );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n411), .SE(n517), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n411), .SE(n515), .CK(clk), .Q(n562), 
        .QN(n30) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n411), .SE(n513), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n335) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n411), .SE(n509), .CK(clk), .Q(
        \mult_x_1/a[2] ) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n411), .SE(n507), .CK(clk), .Q(n560), 
        .QN(n38) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n411), .SE(n505), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n27) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n411), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n29) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n411), .SE(n501), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n35) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n409), .SE(n499), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n36) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n410), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n32) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n408), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n33) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n411), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n34) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n408), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n31) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n408), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n288 ) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n408), .SE(n487), .CK(clk), .Q(n559)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n408), .SE(n485), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n408), .SE(n483), .CK(clk), .Q(n557)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n408), .SE(n481), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n408), .SE(n479), .CK(clk), .Q(n555)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n410), .SE(n477), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n409), .SE(n475), .CK(clk), .Q(n553)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n411), .SE(n473), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n408), .SE(n471), .CK(clk), .Q(n551)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n408), .SE(n469), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n408), .SE(n467), .CK(clk), .Q(n549)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n408), .SE(n465), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n408), .SE(n463), .CK(clk), .Q(n547)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n408), .SE(n461), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n408), .SE(n459), .CK(clk), .Q(n545)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n408), .SE(n457), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n410), .SE(n455), .CK(clk), .Q(n543)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n410), .SE(n453), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n410), .SE(n451), .CK(clk), .Q(n541)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n410), .SE(n449), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n410), .SE(n447), .CK(clk), .Q(n539)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n410), .SE(n445), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n410), .SE(n443), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n410), .SE(n441), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n410), .SE(n439), .CK(clk), .Q(n535)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n410), .SE(n437), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n410), .SE(n435), .CK(clk), .Q(n533)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n409), .SE(n433), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n409), .SE(n431), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n409), .SE(n429), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n409), .SE(n427), .CK(clk), .Q(n529)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n409), .SE(n425), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n409), .SE(n423), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n409), .SE(n421), .CK(clk), .Q(n526)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n409), .SE(n419), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n409), .SE(n417), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n409), .SE(n415), .CK(clk), .Q(n523)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n409), .SE(n413), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n411), .SE(n511), .CK(clk), .Q(n561), 
        .QN(n336) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n564), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n357) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n564), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n356), .QN(n39) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n564), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n355), .QN(n407) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n564), .SI(1'b1), .SE(n390), .CK(clk), 
        .Q(n354), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n564), .SE(n388), .CK(
        clk), .Q(n337), .QN(n353) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n564), .SI(1'b1), .SE(n384), .CK(clk), 
        .Q(n351) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n564), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n350), .QN(n400) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n564), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n349), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n564), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n564), .SI(1'b1), .SE(n376), .CK(clk), 
        .Q(n347), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n564), .SI(1'b1), .SE(n374), .CK(clk), 
        .Q(n346), .QN(n403) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n564), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n345), .QN(n404) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n564), .SE(n370), .CK(
        clk), .Q(n406), .QN(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n564), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n343), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2_IP  ( .D(1'b1), .SI(n564), .SE(n366), .CK(
        clk), .QN(n342) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n564), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n564), .SE(n362), .CK(
        clk), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n564), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n339), .QN(n37) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n564), .SI(1'b1), .SE(n358), .CK(clk), 
        .Q(n338) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n411), .SE(n519), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n28) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n564), .SE(n386), .CK(
        clk), .Q(n405), .QN(n352) );
  BUF_X1 U2 ( .A(n408), .Z(n411) );
  BUF_X1 U3 ( .A(n408), .Z(n409) );
  BUF_X1 U4 ( .A(n408), .Z(n410) );
  INV_X1 U5 ( .A(n564), .ZN(n408) );
  BUF_X1 U6 ( .A(n562), .Z(n333) );
  OR2_X1 U7 ( .A1(n260), .A2(n259), .ZN(n286) );
  AND2_X1 U8 ( .A1(n563), .A2(\mult_x_1/n281 ), .ZN(n150) );
  CLKBUF_X2 U9 ( .A(n560), .Z(n331) );
  FA_X1 U10 ( .A(n123), .B(1'b0), .CI(n121), .CO(n136), .S(n137) );
  OAI21_X1 U11 ( .B1(n209), .B2(n7), .A(n5), .ZN(n376) );
  NAND2_X1 U12 ( .A1(n6), .A2(n347), .ZN(n5) );
  INV_X1 U13 ( .A(n334), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n334), .A2(n8), .ZN(n7) );
  INV_X1 U15 ( .A(n208), .ZN(n8) );
  INV_X2 U16 ( .A(n25), .ZN(n234) );
  OAI21_X1 U17 ( .B1(n11), .B2(n10), .A(n9), .ZN(n447) );
  NAND2_X1 U18 ( .A1(n10), .A2(n539), .ZN(n9) );
  INV_X1 U19 ( .A(n292), .ZN(n10) );
  XNOR2_X1 U20 ( .A(n288), .B(n12), .ZN(n11) );
  INV_X1 U21 ( .A(n287), .ZN(n12) );
  OAI21_X1 U22 ( .B1(n204), .B2(n15), .A(n13), .ZN(n370) );
  NAND2_X1 U23 ( .A1(n14), .A2(n344), .ZN(n13) );
  INV_X1 U24 ( .A(n334), .ZN(n14) );
  NAND2_X1 U25 ( .A1(n16), .A2(n334), .ZN(n15) );
  INV_X1 U26 ( .A(n203), .ZN(n16) );
  INV_X1 U27 ( .A(n41), .ZN(n188) );
  XNOR2_X1 U28 ( .A(n155), .B(n156), .ZN(n87) );
  AND2_X1 U29 ( .A1(n43), .A2(\mult_x_1/n288 ), .ZN(n68) );
  NAND2_X1 U30 ( .A1(n70), .A2(n69), .ZN(n71) );
  AND2_X1 U31 ( .A1(n563), .A2(\mult_x_1/n310 ), .ZN(n42) );
  NAND2_X1 U32 ( .A1(n130), .A2(n106), .ZN(n108) );
  XNOR2_X1 U33 ( .A(n87), .B(n157), .ZN(n181) );
  XNOR2_X1 U34 ( .A(n44), .B(n68), .ZN(n82) );
  XNOR2_X1 U35 ( .A(n70), .B(n69), .ZN(n44) );
  INV_X1 U36 ( .A(rst_n), .ZN(n564) );
  CLKBUF_X1 U37 ( .A(n561), .Z(n332) );
  NAND2_X1 U38 ( .A1(n128), .A2(n127), .ZN(n107) );
  OR2_X1 U39 ( .A1(n128), .A2(n127), .ZN(n106) );
  CLKBUF_X1 U40 ( .A(n245), .Z(n17) );
  NAND2_X1 U41 ( .A1(n45), .A2(n46), .ZN(n18) );
  INV_X1 U42 ( .A(n234), .ZN(n19) );
  XOR2_X1 U43 ( .A(n126), .B(n125), .Z(n20) );
  XOR2_X1 U44 ( .A(n124), .B(n20), .Z(n135) );
  NAND2_X1 U45 ( .A1(n124), .A2(n126), .ZN(n21) );
  NAND2_X1 U46 ( .A1(n124), .A2(n125), .ZN(n22) );
  NAND2_X1 U47 ( .A1(n126), .A2(n125), .ZN(n23) );
  NAND3_X1 U48 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n115) );
  INV_X1 U49 ( .A(n124), .ZN(n24) );
  OAI22_X1 U50 ( .A1(n90), .A2(n89), .B1(n247), .B2(n91), .ZN(n110) );
  XOR2_X1 U51 ( .A(n335), .B(n336), .Z(n25) );
  NAND2_X1 U52 ( .A1(n108), .A2(n107), .ZN(n120) );
  INV_X1 U53 ( .A(n28), .ZN(n26) );
  OR2_X1 U54 ( .A1(n105), .A2(n104), .ZN(n127) );
  XNOR2_X1 U55 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n40) );
  XOR2_X1 U56 ( .A(\mult_x_1/a[6] ), .B(n562), .Z(n41) );
  OR2_X2 U57 ( .A1(n40), .A2(n41), .ZN(n187) );
  XNOR2_X1 U58 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n54) );
  XNOR2_X1 U59 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n78) );
  OAI22_X1 U60 ( .A1(n187), .A2(n54), .B1(n188), .B2(n78), .ZN(n70) );
  NAND2_X1 U61 ( .A1(n331), .A2(n27), .ZN(n250) );
  XNOR2_X1 U62 ( .A(n331), .B(\mult_x_1/n281 ), .ZN(n47) );
  XNOR2_X1 U63 ( .A(n150), .B(n331), .ZN(n76) );
  OAI22_X1 U64 ( .A1(n250), .A2(n47), .B1(n76), .B2(n27), .ZN(n69) );
  XNOR2_X1 U65 ( .A(n42), .B(\mult_x_1/n310 ), .ZN(n86) );
  INV_X1 U66 ( .A(n86), .ZN(n43) );
  XOR2_X1 U67 ( .A(\mult_x_1/a[4] ), .B(n562), .Z(n45) );
  XNOR2_X1 U68 ( .A(n335), .B(n336), .ZN(n46) );
  NAND2_X1 U69 ( .A1(n45), .A2(n46), .ZN(n167) );
  XNOR2_X1 U70 ( .A(n333), .B(\mult_x_1/n286 ), .ZN(n170) );
  XNOR2_X1 U71 ( .A(n333), .B(\mult_x_1/n285 ), .ZN(n51) );
  OAI22_X1 U72 ( .A1(n18), .A2(n170), .B1(n234), .B2(n51), .ZN(n62) );
  XNOR2_X1 U73 ( .A(n331), .B(\mult_x_1/n282 ), .ZN(n56) );
  OAI22_X1 U74 ( .A1(n250), .A2(n56), .B1(n47), .B2(n27), .ZN(n61) );
  XOR2_X1 U75 ( .A(\mult_x_1/a[2] ), .B(n561), .Z(n48) );
  XNOR2_X1 U76 ( .A(\mult_x_1/a[2] ), .B(n560), .ZN(n49) );
  NAND2_X1 U77 ( .A1(n48), .A2(n49), .ZN(n90) );
  BUF_X2 U78 ( .A(n90), .Z(n245) );
  XNOR2_X1 U79 ( .A(n332), .B(\mult_x_1/n284 ), .ZN(n57) );
  INV_X1 U80 ( .A(n49), .ZN(n50) );
  INV_X2 U81 ( .A(n50), .ZN(n247) );
  XNOR2_X1 U82 ( .A(n561), .B(\mult_x_1/n283 ), .ZN(n52) );
  OAI22_X1 U83 ( .A1(n245), .A2(n57), .B1(n247), .B2(n52), .ZN(n60) );
  XNOR2_X1 U84 ( .A(n333), .B(\mult_x_1/n284 ), .ZN(n66) );
  OAI22_X1 U85 ( .A1(n18), .A2(n51), .B1(n234), .B2(n66), .ZN(n75) );
  XNOR2_X1 U86 ( .A(n561), .B(\mult_x_1/n282 ), .ZN(n67) );
  OAI22_X1 U87 ( .A1(n245), .A2(n52), .B1(n247), .B2(n67), .ZN(n74) );
  OR2_X1 U88 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n53) );
  OAI22_X1 U89 ( .A1(n187), .A2(n28), .B1(n53), .B2(n188), .ZN(n59) );
  XNOR2_X1 U90 ( .A(n26), .B(\mult_x_1/n288 ), .ZN(n55) );
  OAI22_X1 U91 ( .A1(n187), .A2(n55), .B1(n188), .B2(n54), .ZN(n58) );
  XNOR2_X1 U92 ( .A(n331), .B(\mult_x_1/n283 ), .ZN(n217) );
  OAI22_X1 U93 ( .A1(n250), .A2(n217), .B1(n56), .B2(n27), .ZN(n174) );
  AND2_X1 U94 ( .A1(\mult_x_1/n288 ), .A2(n41), .ZN(n173) );
  XNOR2_X1 U95 ( .A(n332), .B(\mult_x_1/n285 ), .ZN(n216) );
  OAI22_X1 U96 ( .A1(n216), .A2(n245), .B1(n247), .B2(n57), .ZN(n172) );
  HA_X1 U97 ( .A(n58), .B(n59), .CO(n73), .S(n165) );
  FA_X1 U98 ( .A(n62), .B(n61), .CI(n60), .CO(n81), .S(n164) );
  NAND2_X1 U99 ( .A1(n209), .A2(n208), .ZN(n63) );
  BUF_X8 U100 ( .A(en), .Z(n334) );
  NAND2_X1 U101 ( .A1(n63), .A2(n334), .ZN(n65) );
  NAND2_X1 U102 ( .A1(n10), .A2(n348), .ZN(n64) );
  NAND2_X1 U103 ( .A1(n65), .A2(n64), .ZN(n378) );
  XNOR2_X1 U104 ( .A(n333), .B(\mult_x_1/n283 ), .ZN(n95) );
  OAI22_X1 U105 ( .A1(n167), .A2(n66), .B1(n234), .B2(n95), .ZN(n105) );
  XNOR2_X1 U106 ( .A(n561), .B(\mult_x_1/n281 ), .ZN(n89) );
  OAI22_X1 U107 ( .A1(n67), .A2(n90), .B1(n247), .B2(n89), .ZN(n104) );
  XNOR2_X1 U108 ( .A(n105), .B(n104), .ZN(n123) );
  OAI21_X1 U110 ( .B1(n70), .B2(n69), .A(n68), .ZN(n72) );
  NAND2_X1 U111 ( .A1(n72), .A2(n71), .ZN(n121) );
  FA_X1 U112 ( .A(n75), .B(n74), .CI(n73), .CO(n139), .S(n80) );
  AOI21_X1 U113 ( .B1(n250), .B2(n27), .A(n76), .ZN(n77) );
  INV_X1 U114 ( .A(n77), .ZN(n103) );
  XNOR2_X1 U115 ( .A(n26), .B(\mult_x_1/n285 ), .ZN(n94) );
  OAI22_X1 U116 ( .A1(n187), .A2(n78), .B1(n188), .B2(n94), .ZN(n102) );
  NOR2_X1 U117 ( .A1(n31), .A2(n86), .ZN(n101) );
  XOR2_X1 U118 ( .A(n139), .B(n138), .Z(n79) );
  XOR2_X1 U119 ( .A(n137), .B(n79), .Z(n206) );
  FA_X1 U120 ( .A(n82), .B(n81), .CI(n80), .CO(n205), .S(n209) );
  NAND2_X1 U121 ( .A1(n206), .A2(n205), .ZN(n83) );
  BUF_X4 U122 ( .A(en), .Z(n292) );
  NAND2_X1 U123 ( .A1(n83), .A2(n292), .ZN(n85) );
  OR2_X1 U124 ( .A1(n292), .A2(n39), .ZN(n84) );
  NAND2_X1 U125 ( .A1(n85), .A2(n84), .ZN(n394) );
  CLKBUF_X1 U126 ( .A(n86), .Z(n190) );
  NOR2_X1 U127 ( .A1(n32), .A2(n190), .ZN(n155) );
  XNOR2_X1 U128 ( .A(n26), .B(\mult_x_1/n283 ), .ZN(n88) );
  XNOR2_X1 U129 ( .A(n26), .B(\mult_x_1/n282 ), .ZN(n152) );
  OAI22_X1 U130 ( .A1(n187), .A2(n88), .B1(n188), .B2(n152), .ZN(n156) );
  XNOR2_X1 U131 ( .A(n333), .B(\mult_x_1/n281 ), .ZN(n96) );
  XNOR2_X1 U132 ( .A(n150), .B(n333), .ZN(n153) );
  OAI22_X1 U133 ( .A1(n167), .A2(n96), .B1(n153), .B2(n234), .ZN(n161) );
  INV_X1 U134 ( .A(n161), .ZN(n157) );
  XNOR2_X1 U135 ( .A(n26), .B(\mult_x_1/n284 ), .ZN(n93) );
  OAI22_X1 U136 ( .A1(n187), .A2(n93), .B1(n188), .B2(n88), .ZN(n111) );
  XNOR2_X1 U137 ( .A(n150), .B(n561), .ZN(n91) );
  AOI21_X1 U138 ( .B1(n245), .B2(n247), .A(n91), .ZN(n92) );
  INV_X1 U139 ( .A(n92), .ZN(n109) );
  OAI22_X1 U140 ( .A1(n187), .A2(n94), .B1(n188), .B2(n93), .ZN(n126) );
  XNOR2_X1 U141 ( .A(n333), .B(\mult_x_1/n282 ), .ZN(n97) );
  OAI22_X1 U142 ( .A1(n167), .A2(n95), .B1(n234), .B2(n97), .ZN(n125) );
  INV_X1 U143 ( .A(n110), .ZN(n124) );
  NOR2_X1 U144 ( .A1(n33), .A2(n190), .ZN(n113) );
  NAND2_X1 U145 ( .A1(n115), .A2(n113), .ZN(n100) );
  OAI22_X1 U146 ( .A1(n167), .A2(n97), .B1(n234), .B2(n96), .ZN(n112) );
  NAND2_X1 U147 ( .A1(n115), .A2(n112), .ZN(n99) );
  NAND2_X1 U148 ( .A1(n113), .A2(n112), .ZN(n98) );
  NAND3_X1 U149 ( .A1(n100), .A2(n99), .A3(n98), .ZN(n179) );
  FA_X1 U150 ( .A(n103), .B(n102), .CI(n101), .CO(n130), .S(n138) );
  NOR2_X1 U151 ( .A1(n34), .A2(n190), .ZN(n128) );
  FA_X1 U152 ( .A(n111), .B(n109), .CI(n24), .CO(n180), .S(n119) );
  XNOR2_X1 U153 ( .A(n113), .B(n112), .ZN(n114) );
  XNOR2_X1 U154 ( .A(n115), .B(n114), .ZN(n118) );
  OAI21_X1 U155 ( .B1(n228), .B2(n227), .A(n334), .ZN(n117) );
  OR2_X1 U156 ( .A1(n334), .A2(n37), .ZN(n116) );
  NAND2_X1 U157 ( .A1(n117), .A2(n116), .ZN(n360) );
  FA_X1 U158 ( .A(n120), .B(n119), .CI(n118), .CO(n227), .S(n204) );
  XNOR2_X1 U159 ( .A(n128), .B(n127), .ZN(n129) );
  XNOR2_X1 U160 ( .A(n130), .B(n129), .ZN(n134) );
  NAND2_X1 U161 ( .A1(n204), .A2(n203), .ZN(n131) );
  NAND2_X1 U162 ( .A1(n131), .A2(n334), .ZN(n133) );
  OR2_X1 U163 ( .A1(n334), .A2(n404), .ZN(n132) );
  NAND2_X1 U164 ( .A1(n133), .A2(n132), .ZN(n372) );
  FA_X1 U165 ( .A(n136), .B(n135), .CI(n134), .CO(n203), .S(n146) );
  NAND2_X1 U166 ( .A1(n137), .A2(n139), .ZN(n142) );
  NAND2_X1 U167 ( .A1(n137), .A2(n138), .ZN(n141) );
  NAND2_X1 U168 ( .A1(n139), .A2(n138), .ZN(n140) );
  NAND3_X1 U169 ( .A1(n142), .A2(n141), .A3(n140), .ZN(n145) );
  INV_X1 U170 ( .A(n145), .ZN(n143) );
  NAND2_X1 U171 ( .A1(n143), .A2(n292), .ZN(n144) );
  OAI22_X1 U172 ( .A1(n146), .A2(n144), .B1(n292), .B2(n405), .ZN(n386) );
  NAND2_X1 U173 ( .A1(n146), .A2(n145), .ZN(n147) );
  NAND2_X1 U174 ( .A1(n147), .A2(n292), .ZN(n149) );
  OR2_X1 U175 ( .A1(n292), .A2(n337), .ZN(n148) );
  NAND2_X1 U176 ( .A1(n149), .A2(n148), .ZN(n388) );
  NOR2_X1 U197 ( .A1(n35), .A2(n190), .ZN(n185) );
  XNOR2_X1 U198 ( .A(n26), .B(\mult_x_1/n281 ), .ZN(n151) );
  XNOR2_X1 U199 ( .A(n150), .B(n26), .ZN(n186) );
  OAI22_X1 U200 ( .A1(n187), .A2(n151), .B1(n186), .B2(n188), .ZN(n194) );
  INV_X1 U201 ( .A(n194), .ZN(n184) );
  OAI22_X1 U202 ( .A1(n187), .A2(n152), .B1(n188), .B2(n151), .ZN(n162) );
  AOI21_X1 U203 ( .B1(n234), .B2(n167), .A(n153), .ZN(n154) );
  INV_X1 U204 ( .A(n154), .ZN(n160) );
  OAI21_X1 U205 ( .B1(n157), .B2(n156), .A(n155), .ZN(n159) );
  NAND2_X1 U206 ( .A1(n157), .A2(n156), .ZN(n158) );
  NAND2_X1 U207 ( .A1(n159), .A2(n158), .ZN(n178) );
  NOR2_X1 U208 ( .A1(n36), .A2(n190), .ZN(n177) );
  FA_X1 U209 ( .A(n162), .B(n161), .CI(n160), .CO(n183), .S(n176) );
  OR2_X1 U210 ( .A1(n201), .A2(n200), .ZN(n163) );
  MUX2_X1 U211 ( .A(n338), .B(n163), .S(n334), .Z(n358) );
  FA_X1 U212 ( .A(n166), .B(n165), .CI(n164), .CO(n208), .S(n211) );
  OR2_X1 U213 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n168) );
  OAI22_X1 U214 ( .A1(n18), .A2(n30), .B1(n168), .B2(n234), .ZN(n219) );
  XNOR2_X1 U215 ( .A(n333), .B(\mult_x_1/n288 ), .ZN(n169) );
  XNOR2_X1 U216 ( .A(n333), .B(\mult_x_1/n287 ), .ZN(n171) );
  OAI22_X1 U217 ( .A1(n18), .A2(n169), .B1(n234), .B2(n171), .ZN(n218) );
  AND2_X1 U218 ( .A1(n219), .A2(n218), .ZN(n215) );
  OAI22_X1 U219 ( .A1(n18), .A2(n171), .B1(n234), .B2(n170), .ZN(n214) );
  FA_X1 U220 ( .A(n174), .B(n173), .CI(n172), .CO(n166), .S(n213) );
  OR2_X1 U221 ( .A1(n211), .A2(n210), .ZN(n175) );
  MUX2_X1 U222 ( .A(n340), .B(n175), .S(n334), .Z(n362) );
  FA_X1 U223 ( .A(n178), .B(n177), .CI(n176), .CO(n200), .S(n225) );
  FA_X1 U224 ( .A(n181), .B(n180), .CI(n179), .CO(n224), .S(n228) );
  OR2_X1 U225 ( .A1(n225), .A2(n224), .ZN(n182) );
  MUX2_X1 U226 ( .A(n341), .B(n182), .S(n334), .Z(n364) );
  FA_X1 U227 ( .A(n185), .B(n184), .CI(n183), .CO(n196), .S(n201) );
  AOI21_X1 U228 ( .B1(n188), .B2(n187), .A(n186), .ZN(n189) );
  INV_X1 U229 ( .A(n189), .ZN(n192) );
  NOR2_X1 U230 ( .A1(n29), .A2(n190), .ZN(n191) );
  XOR2_X1 U231 ( .A(n192), .B(n191), .Z(n193) );
  XOR2_X1 U232 ( .A(n194), .B(n193), .Z(n195) );
  OR2_X1 U233 ( .A1(n196), .A2(n195), .ZN(n198) );
  NAND2_X1 U234 ( .A1(n196), .A2(n195), .ZN(n197) );
  NAND2_X1 U235 ( .A1(n198), .A2(n197), .ZN(n199) );
  MUX2_X1 U236 ( .A(n342), .B(n199), .S(n334), .Z(n366) );
  NAND2_X1 U237 ( .A1(n201), .A2(n200), .ZN(n202) );
  MUX2_X1 U238 ( .A(n343), .B(n202), .S(n334), .Z(n368) );
  NOR2_X1 U239 ( .A1(n206), .A2(n205), .ZN(n207) );
  MUX2_X1 U240 ( .A(n346), .B(n207), .S(n334), .Z(n374) );
  NAND2_X1 U241 ( .A1(n211), .A2(n210), .ZN(n212) );
  MUX2_X1 U242 ( .A(n349), .B(n212), .S(n334), .Z(n380) );
  FA_X1 U243 ( .A(n215), .B(n214), .CI(n213), .CO(n210), .S(n222) );
  XNOR2_X1 U244 ( .A(n332), .B(\mult_x_1/n286 ), .ZN(n235) );
  OAI22_X1 U245 ( .A1(n17), .A2(n235), .B1(n247), .B2(n216), .ZN(n232) );
  XNOR2_X1 U246 ( .A(n331), .B(\mult_x_1/n284 ), .ZN(n233) );
  OAI22_X1 U247 ( .A1(n250), .A2(n233), .B1(n217), .B2(n27), .ZN(n231) );
  XOR2_X1 U248 ( .A(n218), .B(n219), .Z(n230) );
  NOR2_X1 U249 ( .A1(n222), .A2(n221), .ZN(n220) );
  MUX2_X1 U250 ( .A(n350), .B(n220), .S(n292), .Z(n382) );
  NAND2_X1 U251 ( .A1(n222), .A2(n221), .ZN(n223) );
  MUX2_X1 U252 ( .A(n351), .B(n223), .S(n292), .Z(n384) );
  NAND2_X1 U253 ( .A1(n225), .A2(n224), .ZN(n226) );
  MUX2_X1 U254 ( .A(n354), .B(n226), .S(n292), .Z(n390) );
  NAND2_X1 U255 ( .A1(n228), .A2(n227), .ZN(n229) );
  MUX2_X1 U256 ( .A(n355), .B(n229), .S(n292), .Z(n392) );
  FA_X1 U257 ( .A(n232), .B(n231), .CI(n230), .CO(n221), .S(n260) );
  XNOR2_X1 U258 ( .A(n331), .B(\mult_x_1/n285 ), .ZN(n241) );
  OAI22_X1 U259 ( .A1(n250), .A2(n241), .B1(n233), .B2(n27), .ZN(n238) );
  AND2_X1 U260 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n237) );
  XNOR2_X1 U261 ( .A(n561), .B(\mult_x_1/n287 ), .ZN(n239) );
  OAI22_X1 U262 ( .A1(n245), .A2(n239), .B1(n247), .B2(n235), .ZN(n236) );
  FA_X1 U263 ( .A(n238), .B(n237), .CI(n236), .CO(n259), .S(n258) );
  XNOR2_X1 U264 ( .A(n332), .B(\mult_x_1/n288 ), .ZN(n240) );
  OAI22_X1 U265 ( .A1(n245), .A2(n240), .B1(n247), .B2(n239), .ZN(n243) );
  XNOR2_X1 U266 ( .A(n331), .B(\mult_x_1/n286 ), .ZN(n246) );
  OAI22_X1 U267 ( .A1(n250), .A2(n246), .B1(n241), .B2(n27), .ZN(n242) );
  NOR2_X1 U268 ( .A1(n258), .A2(n257), .ZN(n279) );
  HA_X1 U269 ( .A(n243), .B(n242), .CO(n257), .S(n255) );
  OR2_X1 U270 ( .A1(\mult_x_1/n288 ), .A2(n336), .ZN(n244) );
  OAI22_X1 U271 ( .A1(n17), .A2(n336), .B1(n244), .B2(n247), .ZN(n254) );
  OR2_X1 U272 ( .A1(n255), .A2(n254), .ZN(n275) );
  XNOR2_X1 U273 ( .A(n331), .B(\mult_x_1/n287 ), .ZN(n249) );
  OAI22_X1 U274 ( .A1(n250), .A2(n249), .B1(n246), .B2(n27), .ZN(n253) );
  INV_X1 U275 ( .A(n247), .ZN(n248) );
  AND2_X1 U276 ( .A1(\mult_x_1/n288 ), .A2(n248), .ZN(n252) );
  NOR2_X1 U277 ( .A1(n253), .A2(n252), .ZN(n268) );
  OAI22_X1 U278 ( .A1(n250), .A2(\mult_x_1/n288 ), .B1(n249), .B2(n27), .ZN(
        n265) );
  OR2_X1 U279 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n251) );
  NAND2_X1 U280 ( .A1(n251), .A2(n250), .ZN(n264) );
  NAND2_X1 U281 ( .A1(n265), .A2(n264), .ZN(n271) );
  NAND2_X1 U282 ( .A1(n253), .A2(n252), .ZN(n269) );
  OAI21_X1 U283 ( .B1(n268), .B2(n271), .A(n269), .ZN(n276) );
  NAND2_X1 U284 ( .A1(n255), .A2(n254), .ZN(n274) );
  INV_X1 U285 ( .A(n274), .ZN(n256) );
  AOI21_X1 U286 ( .B1(n275), .B2(n276), .A(n256), .ZN(n282) );
  NAND2_X1 U287 ( .A1(n258), .A2(n257), .ZN(n280) );
  OAI21_X1 U288 ( .B1(n279), .B2(n282), .A(n280), .ZN(n287) );
  NAND2_X1 U289 ( .A1(n260), .A2(n259), .ZN(n285) );
  INV_X1 U290 ( .A(n285), .ZN(n261) );
  AOI21_X1 U291 ( .B1(n286), .B2(n287), .A(n261), .ZN(n262) );
  MUX2_X1 U292 ( .A(n357), .B(n262), .S(n292), .Z(n396) );
  MUX2_X1 U293 ( .A(product[0]), .B(n523), .S(n292), .Z(n413) );
  MUX2_X1 U294 ( .A(n523), .B(n524), .S(n292), .Z(n415) );
  AND2_X1 U295 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n263) );
  MUX2_X1 U296 ( .A(n524), .B(n263), .S(n292), .Z(n417) );
  MUX2_X1 U297 ( .A(product[1]), .B(n526), .S(n292), .Z(n419) );
  MUX2_X1 U298 ( .A(n526), .B(n527), .S(n292), .Z(n421) );
  OR2_X1 U299 ( .A1(n265), .A2(n264), .ZN(n266) );
  AND2_X1 U300 ( .A1(n266), .A2(n271), .ZN(n267) );
  MUX2_X1 U301 ( .A(n527), .B(n267), .S(n292), .Z(n423) );
  MUX2_X1 U302 ( .A(product[2]), .B(n529), .S(n292), .Z(n425) );
  MUX2_X1 U303 ( .A(n529), .B(n530), .S(n292), .Z(n427) );
  INV_X1 U304 ( .A(n268), .ZN(n270) );
  NAND2_X1 U305 ( .A1(n270), .A2(n269), .ZN(n272) );
  XOR2_X1 U306 ( .A(n272), .B(n271), .Z(n273) );
  MUX2_X1 U307 ( .A(n530), .B(n273), .S(n292), .Z(n429) );
  MUX2_X1 U308 ( .A(product[3]), .B(n532), .S(n292), .Z(n431) );
  MUX2_X1 U309 ( .A(n532), .B(n533), .S(n292), .Z(n433) );
  NAND2_X1 U310 ( .A1(n275), .A2(n274), .ZN(n277) );
  XNOR2_X1 U311 ( .A(n277), .B(n276), .ZN(n278) );
  MUX2_X1 U312 ( .A(n533), .B(n278), .S(n292), .Z(n435) );
  MUX2_X1 U313 ( .A(product[4]), .B(n535), .S(n292), .Z(n437) );
  MUX2_X1 U314 ( .A(n535), .B(n536), .S(n292), .Z(n439) );
  INV_X1 U315 ( .A(n279), .ZN(n281) );
  NAND2_X1 U316 ( .A1(n281), .A2(n280), .ZN(n283) );
  XOR2_X1 U317 ( .A(n283), .B(n282), .Z(n284) );
  MUX2_X1 U318 ( .A(n536), .B(n284), .S(n292), .Z(n441) );
  MUX2_X1 U319 ( .A(product[5]), .B(n538), .S(n292), .Z(n443) );
  MUX2_X1 U320 ( .A(n538), .B(n539), .S(n292), .Z(n445) );
  NAND2_X1 U321 ( .A1(n286), .A2(n285), .ZN(n288) );
  MUX2_X1 U322 ( .A(product[6]), .B(n541), .S(n292), .Z(n449) );
  NAND2_X1 U323 ( .A1(n400), .A2(n351), .ZN(n289) );
  XOR2_X1 U324 ( .A(n289), .B(n357), .Z(n290) );
  MUX2_X1 U325 ( .A(n541), .B(n290), .S(n292), .Z(n451) );
  MUX2_X1 U326 ( .A(product[7]), .B(n543), .S(n292), .Z(n453) );
  OAI21_X1 U327 ( .B1(n350), .B2(n357), .A(n351), .ZN(n294) );
  NAND2_X1 U328 ( .A1(n340), .A2(n349), .ZN(n291) );
  XNOR2_X1 U329 ( .A(n294), .B(n291), .ZN(n293) );
  MUX2_X1 U330 ( .A(n543), .B(n293), .S(n292), .Z(n455) );
  MUX2_X1 U331 ( .A(product[8]), .B(n545), .S(n334), .Z(n457) );
  AOI21_X1 U332 ( .B1(n294), .B2(n340), .A(n401), .ZN(n297) );
  NAND2_X1 U333 ( .A1(n402), .A2(n348), .ZN(n295) );
  XOR2_X1 U334 ( .A(n297), .B(n295), .Z(n296) );
  MUX2_X1 U335 ( .A(n545), .B(n296), .S(n334), .Z(n459) );
  MUX2_X1 U336 ( .A(product[9]), .B(n547), .S(n334), .Z(n461) );
  OAI21_X1 U337 ( .B1(n297), .B2(n347), .A(n348), .ZN(n305) );
  INV_X1 U338 ( .A(n305), .ZN(n300) );
  NAND2_X1 U339 ( .A1(n403), .A2(n356), .ZN(n298) );
  XOR2_X1 U340 ( .A(n300), .B(n298), .Z(n299) );
  MUX2_X1 U341 ( .A(n547), .B(n299), .S(n334), .Z(n463) );
  MUX2_X1 U342 ( .A(product[10]), .B(n549), .S(n334), .Z(n465) );
  OAI21_X1 U343 ( .B1(n300), .B2(n346), .A(n356), .ZN(n302) );
  NAND2_X1 U344 ( .A1(n405), .A2(n353), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n303) );
  MUX2_X1 U346 ( .A(n549), .B(n303), .S(n334), .Z(n467) );
  MUX2_X1 U347 ( .A(product[11]), .B(n551), .S(n334), .Z(n469) );
  NOR2_X1 U348 ( .A1(n352), .A2(n346), .ZN(n306) );
  OAI21_X1 U349 ( .B1(n352), .B2(n356), .A(n353), .ZN(n304) );
  AOI21_X1 U350 ( .B1(n306), .B2(n305), .A(n304), .ZN(n328) );
  NAND2_X1 U351 ( .A1(n406), .A2(n345), .ZN(n307) );
  XOR2_X1 U352 ( .A(n328), .B(n307), .Z(n308) );
  MUX2_X1 U353 ( .A(n551), .B(n308), .S(n334), .Z(n471) );
  MUX2_X1 U354 ( .A(product[12]), .B(n553), .S(n334), .Z(n473) );
  OAI21_X1 U355 ( .B1(n328), .B2(n344), .A(n345), .ZN(n310) );
  NAND2_X1 U356 ( .A1(n339), .A2(n355), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  MUX2_X1 U358 ( .A(n553), .B(n311), .S(n334), .Z(n475) );
  MUX2_X1 U359 ( .A(product[13]), .B(n555), .S(n334), .Z(n477) );
  NAND2_X1 U360 ( .A1(n406), .A2(n339), .ZN(n313) );
  AOI21_X1 U361 ( .B1(n404), .B2(n339), .A(n407), .ZN(n312) );
  OAI21_X1 U362 ( .B1(n328), .B2(n313), .A(n312), .ZN(n315) );
  NAND2_X1 U363 ( .A1(n341), .A2(n354), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  MUX2_X1 U365 ( .A(n555), .B(n316), .S(n334), .Z(n479) );
  MUX2_X1 U366 ( .A(product[14]), .B(n557), .S(n334), .Z(n481) );
  NAND2_X1 U367 ( .A1(n339), .A2(n341), .ZN(n318) );
  NOR2_X1 U368 ( .A1(n344), .A2(n318), .ZN(n324) );
  INV_X1 U369 ( .A(n324), .ZN(n320) );
  AOI21_X1 U370 ( .B1(n407), .B2(n341), .A(n399), .ZN(n317) );
  OAI21_X1 U371 ( .B1(n318), .B2(n345), .A(n317), .ZN(n325) );
  INV_X1 U372 ( .A(n325), .ZN(n319) );
  OAI21_X1 U373 ( .B1(n328), .B2(n320), .A(n319), .ZN(n322) );
  NAND2_X1 U374 ( .A1(n338), .A2(n343), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  MUX2_X1 U376 ( .A(n557), .B(n323), .S(n334), .Z(n483) );
  MUX2_X1 U377 ( .A(product[15]), .B(n559), .S(n334), .Z(n485) );
  NAND2_X1 U378 ( .A1(n324), .A2(n338), .ZN(n327) );
  AOI21_X1 U379 ( .B1(n325), .B2(n338), .A(n398), .ZN(n326) );
  OAI21_X1 U380 ( .B1(n328), .B2(n327), .A(n326), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n329), .B(n342), .ZN(n330) );
  MUX2_X1 U382 ( .A(n559), .B(n330), .S(n334), .Z(n487) );
  MUX2_X1 U383 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n334), .Z(n489) );
  MUX2_X1 U384 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n334), .Z(n491) );
  MUX2_X1 U385 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n334), .Z(n493) );
  MUX2_X1 U386 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n334), .Z(n495) );
  MUX2_X1 U387 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n334), .Z(n497) );
  MUX2_X1 U388 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n334), .Z(n499) );
  MUX2_X1 U389 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n334), .Z(n501) );
  MUX2_X1 U390 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n334), .Z(n503) );
  MUX2_X1 U391 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n334), .Z(n505) );
  MUX2_X1 U392 ( .A(n331), .B(A_extended[1]), .S(n334), .Z(n507) );
  MUX2_X1 U393 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n334), .Z(n509) );
  MUX2_X1 U394 ( .A(n332), .B(A_extended[3]), .S(n334), .Z(n511) );
  MUX2_X1 U395 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n334), .Z(n513) );
  MUX2_X1 U396 ( .A(n333), .B(A_extended[5]), .S(n334), .Z(n515) );
  MUX2_X1 U397 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n334), .Z(n517) );
  MUX2_X1 U398 ( .A(n26), .B(A_extended[7]), .S(n334), .Z(n519) );
  OR2_X1 U399 ( .A1(n334), .A2(n563), .ZN(n521) );
endmodule


module conv_128_32_DW_mult_pipe_J1_25 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n352, n354, n356, n358, n360, n362, n364, n366,
         n368, n370, n372, n374, n376, n378, n380, n382, n384, n386, n388,
         n390, n392, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n407, n409, n411, n413, n415, n417, n419, n421,
         n423, n425, n427, n429, n431, n433, n435, n437, n439, n441, n443,
         n445, n447, n449, n451, n453, n455, n457, n459, n461, n463, n465,
         n467, n469, n471, n473, n475, n477, n479, n481, n483, n485, n487,
         n489, n491, n493, n495, n497, n499, n501, n503, n505, n507, n509,
         n511, n513, n515, n516, n518, n519, n521, n522, n524, n525, n527,
         n528, n530, n532, n534, n536, n538, n540, n542, n544, n546, n548,
         n550, n551, n552, n553;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n405), .SE(n513), .CK(clk), .Q(n552), 
        .QN(n28) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n405), .SE(n509), .CK(clk), .Q(
        \mult_x_1/a[6] ) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n405), .SE(n505), .CK(clk), .Q(
        \mult_x_1/a[4] ) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n405), .SE(n501), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n16) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n405), .SE(n499), .CK(clk), .Q(n551), 
        .QN(n30) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n405), .SE(n497), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n17) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n405), .SE(n495), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n20) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n405), .SE(n493), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n26) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n403), .SE(n491), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n27) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n404), .SE(n489), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n25) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n402), .SE(n487), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n24) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n405), .SE(n485), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n22) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n402), .SE(n483), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n23) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n402), .SE(n481), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n18) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n402), .SE(n479), .CK(clk), .Q(n550)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n402), .SE(n477), .CK(clk), .Q(
        product[15]) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n402), .SE(n475), .CK(clk), .Q(n548)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n402), .SE(n473), .CK(clk), .Q(
        product[14]) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n402), .SE(n471), .CK(clk), .Q(n546)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n404), .SE(n469), .CK(clk), .Q(
        product[13]) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n405), .SE(n467), .CK(clk), .Q(n544)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n403), .SE(n465), .CK(clk), .Q(
        product[12]) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n402), .SE(n463), .CK(clk), .Q(n542)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n402), .SE(n461), .CK(clk), .Q(
        product[11]) );
  SDFF_X1 clk_r_REG22_S3 ( .D(1'b0), .SI(n402), .SE(n459), .CK(clk), .Q(n540)
         );
  SDFF_X1 clk_r_REG23_S4 ( .D(1'b0), .SI(n402), .SE(n457), .CK(clk), .Q(
        product[10]) );
  SDFF_X1 clk_r_REG20_S3 ( .D(1'b0), .SI(n402), .SE(n455), .CK(clk), .Q(n538)
         );
  SDFF_X1 clk_r_REG21_S4 ( .D(1'b0), .SI(n402), .SE(n453), .CK(clk), .Q(
        product[9]) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n402), .SE(n451), .CK(clk), .Q(n536)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n404), .SE(n449), .CK(clk), .Q(
        product[8]) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n404), .SE(n447), .CK(clk), .Q(n534)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n404), .SE(n445), .CK(clk), .Q(
        product[7]) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n404), .SE(n443), .CK(clk), .Q(n532)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n404), .SE(n441), .CK(clk), .Q(
        product[6]) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n404), .SE(n439), .CK(clk), .Q(n530)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n404), .SE(n437), .CK(clk), .Q(
        product[5]) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n404), .SE(n435), .CK(clk), .Q(n528)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n404), .SE(n433), .CK(clk), .Q(n527)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n404), .SE(n431), .CK(clk), .Q(
        product[4]) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n404), .SE(n429), .CK(clk), .Q(n525)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n403), .SE(n427), .CK(clk), .Q(n524)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n403), .SE(n425), .CK(clk), .Q(
        product[3]) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n403), .SE(n423), .CK(clk), .Q(n522)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n403), .SE(n421), .CK(clk), .Q(n521)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n403), .SE(n419), .CK(clk), .Q(
        product[2]) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n403), .SE(n417), .CK(clk), .Q(n519)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n403), .SE(n415), .CK(clk), .Q(n518)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n403), .SE(n413), .CK(clk), .Q(
        product[1]) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n403), .SE(n411), .CK(clk), .Q(n516)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n403), .SE(n409), .CK(clk), .Q(n515)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n403), .SE(n407), .CK(clk), .Q(
        product[0]) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n553), .SE(n392), .CK(
        clk), .QN(n349) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2_IP  ( .D(1'b1), .SI(n553), .SE(n390), .CK(
        clk), .QN(n348) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2_IP  ( .D(1'b1), .SI(n553), .SE(n388), .CK(
        clk), .QN(n347) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n553), .SI(1'b1), .SE(n386), .CK(clk), 
        .Q(n346) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n553), .SE(n384), .CK(
        clk), .QN(n345) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n553), .SI(1'b1), .SE(n382), .CK(clk), 
        .Q(n344) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n553), .SI(1'b1), .SE(n380), .CK(clk), 
        .Q(n343), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n553), .SI(1'b1), .SE(n378), .CK(clk), 
        .Q(n342), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n553), .SE(n376), .CK(
        clk), .QN(n341) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n553), .SE(n374), .CK(
        clk), .Q(n400), .QN(n340) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n553), .SI(1'b1), .SE(n372), .CK(clk), 
        .Q(n339) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n553), .SI(1'b1), .SE(n370), .CK(clk), 
        .Q(n338) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n553), .SI(1'b1), .SE(n368), .CK(clk), 
        .Q(n337), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n553), .SI(1'b1), .SE(n366), .CK(clk), 
        .Q(n336), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n553), .SI(1'b1), .SE(n364), .CK(clk), 
        .Q(n335) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n553), .SI(1'b1), .SE(n362), .CK(clk), 
        .Q(n334), .QN(n399) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n553), .SI(1'b1), .SE(n360), .CK(clk), 
        .Q(n333), .QN(n394) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n553), .SE(n358), .CK(
        clk), .QN(n332) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n553), .SE(n356), .CK(
        clk), .QN(n331) );
  SDFF_X1 \mult_x_1/clk_r_REG17_S2  ( .D(n553), .SI(1'b1), .SE(n354), .CK(clk), 
        .Q(n330) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n553), .SI(1'b1), .SE(n352), .CK(clk), 
        .Q(n329) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n553), .SI(1'b1), .SE(n350), .CK(clk), 
        .Q(n328), .QN(n395) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n405), .SE(n507), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n327) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n405), .SE(n511), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n326) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n405), .SE(n503), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n19) );
  BUF_X1 U2 ( .A(en), .Z(n249) );
  INV_X1 U3 ( .A(rst_n), .ZN(n553) );
  INV_X1 U4 ( .A(n553), .ZN(n402) );
  CLKBUF_X2 U5 ( .A(n249), .Z(n14) );
  CLKBUF_X1 U6 ( .A(n402), .Z(n404) );
  CLKBUF_X1 U7 ( .A(n402), .Z(n405) );
  CLKBUF_X1 U8 ( .A(n402), .Z(n403) );
  BUF_X1 U9 ( .A(n551), .Z(n322) );
  BUF_X2 U10 ( .A(n249), .Z(n13) );
  BUF_X8 U11 ( .A(en), .Z(n325) );
  XNOR2_X1 U12 ( .A(n9), .B(n95), .ZN(n237) );
  XNOR2_X1 U13 ( .A(n97), .B(n96), .ZN(n9) );
  INV_X1 U14 ( .A(n36), .ZN(n212) );
  INV_X1 U15 ( .A(n39), .ZN(n160) );
  INV_X1 U16 ( .A(n196), .ZN(n148) );
  INV_X1 U17 ( .A(n19), .ZN(n15) );
  NAND2_X1 U18 ( .A1(n37), .A2(n38), .ZN(n159) );
  NAND2_X1 U19 ( .A1(n32), .A2(n33), .ZN(n150) );
  AND2_X1 U20 ( .A1(n552), .A2(\mult_x_1/n281 ), .ZN(n112) );
  INV_X1 U21 ( .A(n326), .ZN(n324) );
  XNOR2_X1 U22 ( .A(n133), .B(n5), .ZN(n109) );
  XNOR2_X1 U23 ( .A(n135), .B(n134), .ZN(n5) );
  OAI21_X1 U24 ( .B1(n8), .B2(n7), .A(n6), .ZN(n235) );
  NAND2_X1 U25 ( .A1(n97), .A2(n96), .ZN(n6) );
  NOR2_X1 U26 ( .A1(n97), .A2(n96), .ZN(n7) );
  INV_X1 U27 ( .A(n95), .ZN(n8) );
  OAI21_X1 U28 ( .B1(n202), .B2(n11), .A(n10), .ZN(n374) );
  NAND2_X1 U29 ( .A1(n60), .A2(n340), .ZN(n10) );
  NAND2_X1 U30 ( .A1(n12), .A2(n325), .ZN(n11) );
  INV_X1 U31 ( .A(n201), .ZN(n12) );
  NOR2_X1 U32 ( .A1(n102), .A2(n101), .ZN(n86) );
  NAND2_X1 U33 ( .A1(n130), .A2(n129), .ZN(n126) );
  OR2_X1 U34 ( .A1(n130), .A2(n129), .ZN(n125) );
  AND2_X1 U35 ( .A1(n202), .A2(n201), .ZN(n61) );
  OAI21_X1 U36 ( .B1(n109), .B2(n108), .A(n13), .ZN(n111) );
  NAND2_X1 U37 ( .A1(n111), .A2(n110), .ZN(n354) );
  XNOR2_X1 U38 ( .A(n16), .B(n30), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n61), .B2(n60), .A(n59), .ZN(n376) );
  NAND2_X1 U40 ( .A1(n60), .A2(n330), .ZN(n110) );
  NAND2_X1 U41 ( .A1(n60), .A2(n341), .ZN(n59) );
  AND2_X1 U42 ( .A1(n58), .A2(n57), .ZN(n21) );
  INV_X1 U43 ( .A(n249), .ZN(n60) );
  XOR2_X1 U44 ( .A(n58), .B(n57), .Z(n29) );
  NAND2_X1 U45 ( .A1(n102), .A2(n101), .ZN(n31) );
  XOR2_X1 U46 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n32) );
  XNOR2_X1 U47 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n33) );
  INV_X1 U48 ( .A(n327), .ZN(n323) );
  XNOR2_X1 U49 ( .A(n323), .B(\mult_x_1/n284 ), .ZN(n52) );
  INV_X1 U50 ( .A(n33), .ZN(n196) );
  XNOR2_X1 U51 ( .A(n323), .B(\mult_x_1/n283 ), .ZN(n40) );
  OAI22_X1 U52 ( .A1(n150), .A2(n52), .B1(n148), .B2(n40), .ZN(n43) );
  XNOR2_X1 U53 ( .A(n19), .B(\mult_x_1/a[2] ), .ZN(n34) );
  NAND2_X1 U54 ( .A1(n34), .A2(n35), .ZN(n210) );
  XNOR2_X1 U55 ( .A(n15), .B(\mult_x_1/n282 ), .ZN(n53) );
  INV_X1 U56 ( .A(n35), .ZN(n36) );
  XNOR2_X1 U57 ( .A(n15), .B(\mult_x_1/n281 ), .ZN(n92) );
  OAI22_X1 U58 ( .A1(n210), .A2(n53), .B1(n212), .B2(n92), .ZN(n42) );
  XNOR2_X1 U59 ( .A(n43), .B(n42), .ZN(n58) );
  XOR2_X1 U60 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n37) );
  XNOR2_X1 U61 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[6] ), .ZN(n38) );
  XNOR2_X1 U62 ( .A(n324), .B(\mult_x_1/n287 ), .ZN(n55) );
  INV_X1 U63 ( .A(n38), .ZN(n39) );
  XNOR2_X1 U64 ( .A(n324), .B(\mult_x_1/n286 ), .ZN(n47) );
  OAI22_X1 U65 ( .A1(n159), .A2(n55), .B1(n160), .B2(n47), .ZN(n64) );
  NAND2_X1 U66 ( .A1(n322), .A2(n17), .ZN(n214) );
  XNOR2_X1 U67 ( .A(n322), .B(\mult_x_1/n281 ), .ZN(n66) );
  XNOR2_X1 U68 ( .A(n112), .B(n322), .ZN(n44) );
  OAI22_X1 U69 ( .A1(n214), .A2(n66), .B1(n44), .B2(n17), .ZN(n63) );
  NAND2_X1 U70 ( .A1(n28), .A2(n324), .ZN(n162) );
  NOR2_X1 U71 ( .A1(n162), .A2(n18), .ZN(n62) );
  XNOR2_X1 U72 ( .A(n324), .B(\mult_x_1/n285 ), .ZN(n46) );
  XNOR2_X1 U73 ( .A(n324), .B(\mult_x_1/n284 ), .ZN(n91) );
  OAI22_X1 U74 ( .A1(n159), .A2(n46), .B1(n160), .B2(n91), .ZN(n84) );
  XNOR2_X1 U75 ( .A(n323), .B(\mult_x_1/n282 ), .ZN(n85) );
  OAI22_X1 U76 ( .A1(n150), .A2(n40), .B1(n148), .B2(n85), .ZN(n83) );
  XNOR2_X1 U77 ( .A(n112), .B(n15), .ZN(n93) );
  OAI22_X1 U78 ( .A1(n210), .A2(n92), .B1(n93), .B2(n212), .ZN(n41) );
  INV_X1 U79 ( .A(n41), .ZN(n82) );
  XNOR2_X1 U80 ( .A(n21), .B(n238), .ZN(n48) );
  OR2_X1 U81 ( .A1(n43), .A2(n42), .ZN(n97) );
  NOR2_X1 U82 ( .A1(n22), .A2(n162), .ZN(n96) );
  AOI21_X1 U83 ( .B1(n214), .B2(n17), .A(n44), .ZN(n45) );
  INV_X1 U84 ( .A(n45), .ZN(n51) );
  OAI22_X1 U85 ( .A1(n159), .A2(n47), .B1(n160), .B2(n46), .ZN(n50) );
  NOR2_X1 U86 ( .A1(n23), .A2(n162), .ZN(n49) );
  XNOR2_X1 U87 ( .A(n48), .B(n237), .ZN(n202) );
  FA_X1 U88 ( .A(n51), .B(n50), .CI(n49), .CO(n95), .S(n244) );
  XNOR2_X1 U89 ( .A(n323), .B(\mult_x_1/n285 ), .ZN(n65) );
  OAI22_X1 U90 ( .A1(n150), .A2(n65), .B1(n148), .B2(n52), .ZN(n70) );
  XNOR2_X1 U91 ( .A(n15), .B(\mult_x_1/n283 ), .ZN(n67) );
  OAI22_X1 U92 ( .A1(n210), .A2(n67), .B1(n212), .B2(n53), .ZN(n69) );
  OR2_X1 U93 ( .A1(\mult_x_1/n288 ), .A2(n326), .ZN(n54) );
  OAI22_X1 U94 ( .A1(n160), .A2(n54), .B1(n159), .B2(n326), .ZN(n75) );
  XNOR2_X1 U95 ( .A(n324), .B(\mult_x_1/n288 ), .ZN(n56) );
  OAI22_X1 U96 ( .A1(n159), .A2(n56), .B1(n160), .B2(n55), .ZN(n74) );
  FA_X1 U97 ( .A(n64), .B(n63), .CI(n62), .CO(n57), .S(n248) );
  XNOR2_X1 U98 ( .A(n323), .B(\mult_x_1/n286 ), .ZN(n147) );
  OAI22_X1 U99 ( .A1(n150), .A2(n147), .B1(n148), .B2(n65), .ZN(n78) );
  XNOR2_X1 U100 ( .A(n322), .B(\mult_x_1/n282 ), .ZN(n71) );
  OAI22_X1 U101 ( .A1(n214), .A2(n71), .B1(n66), .B2(n17), .ZN(n77) );
  XNOR2_X1 U102 ( .A(n15), .B(\mult_x_1/n284 ), .ZN(n73) );
  OAI22_X1 U103 ( .A1(n210), .A2(n73), .B1(n212), .B2(n67), .ZN(n76) );
  FA_X1 U104 ( .A(n70), .B(n69), .CI(n68), .CO(n243), .S(n246) );
  XNOR2_X1 U105 ( .A(n322), .B(\mult_x_1/n283 ), .ZN(n185) );
  OAI22_X1 U106 ( .A1(n214), .A2(n185), .B1(n71), .B2(n17), .ZN(n153) );
  INV_X1 U107 ( .A(n160), .ZN(n72) );
  AND2_X1 U108 ( .A1(\mult_x_1/n288 ), .A2(n72), .ZN(n152) );
  XNOR2_X1 U109 ( .A(n15), .B(\mult_x_1/n285 ), .ZN(n184) );
  OAI22_X1 U110 ( .A1(n210), .A2(n184), .B1(n212), .B2(n73), .ZN(n151) );
  HA_X1 U111 ( .A(n75), .B(n74), .CO(n68), .S(n143) );
  FA_X1 U112 ( .A(n78), .B(n77), .CI(n76), .CO(n247), .S(n142) );
  NAND2_X1 U113 ( .A1(n176), .A2(n175), .ZN(n79) );
  NAND2_X1 U114 ( .A1(n79), .A2(n325), .ZN(n81) );
  NAND2_X1 U115 ( .A1(n60), .A2(n335), .ZN(n80) );
  NAND2_X1 U116 ( .A1(n81), .A2(n80), .ZN(n364) );
  FA_X1 U117 ( .A(n84), .B(n83), .CI(n82), .CO(n104), .S(n238) );
  INV_X1 U118 ( .A(n104), .ZN(n87) );
  NOR2_X1 U119 ( .A1(n24), .A2(n162), .ZN(n102) );
  XNOR2_X1 U120 ( .A(n323), .B(\mult_x_1/n281 ), .ZN(n88) );
  OAI22_X1 U121 ( .A1(n150), .A2(n85), .B1(n148), .B2(n88), .ZN(n101) );
  OAI21_X1 U122 ( .B1(n87), .B2(n86), .A(n31), .ZN(n133) );
  NOR2_X1 U123 ( .A1(n25), .A2(n162), .ZN(n120) );
  XNOR2_X1 U124 ( .A(n324), .B(\mult_x_1/n283 ), .ZN(n90) );
  XNOR2_X1 U125 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n114) );
  OAI22_X1 U126 ( .A1(n159), .A2(n90), .B1(n160), .B2(n114), .ZN(n121) );
  XNOR2_X1 U127 ( .A(n120), .B(n121), .ZN(n89) );
  XNOR2_X1 U128 ( .A(n112), .B(\mult_x_1/n311 ), .ZN(n115) );
  OAI22_X1 U129 ( .A1(n150), .A2(n88), .B1(n115), .B2(n148), .ZN(n117) );
  INV_X1 U130 ( .A(n117), .ZN(n122) );
  XNOR2_X1 U131 ( .A(n89), .B(n122), .ZN(n135) );
  OAI22_X1 U132 ( .A1(n159), .A2(n91), .B1(n160), .B2(n90), .ZN(n100) );
  OAI22_X1 U133 ( .A1(n210), .A2(n92), .B1(n93), .B2(n212), .ZN(n99) );
  AOI21_X1 U134 ( .B1(n212), .B2(n210), .A(n93), .ZN(n94) );
  INV_X1 U135 ( .A(n94), .ZN(n98) );
  FA_X1 U136 ( .A(n100), .B(n99), .CI(n98), .CO(n134), .S(n234) );
  XOR2_X1 U137 ( .A(n102), .B(n101), .Z(n103) );
  XOR2_X1 U138 ( .A(n104), .B(n103), .Z(n233) );
  NAND2_X1 U139 ( .A1(n109), .A2(n108), .ZN(n105) );
  NAND2_X1 U140 ( .A1(n105), .A2(n325), .ZN(n107) );
  NAND2_X1 U141 ( .A1(n60), .A2(n343), .ZN(n106) );
  NAND2_X1 U142 ( .A1(n107), .A2(n106), .ZN(n380) );
  NOR2_X1 U165 ( .A1(n26), .A2(n162), .ZN(n157) );
  XNOR2_X1 U166 ( .A(n324), .B(\mult_x_1/n281 ), .ZN(n113) );
  XNOR2_X1 U167 ( .A(n112), .B(n324), .ZN(n158) );
  OAI22_X1 U168 ( .A1(n159), .A2(n113), .B1(n158), .B2(n160), .ZN(n166) );
  INV_X1 U169 ( .A(n166), .ZN(n156) );
  OAI22_X1 U170 ( .A1(n159), .A2(n114), .B1(n160), .B2(n113), .ZN(n119) );
  AOI21_X1 U171 ( .B1(n148), .B2(n150), .A(n115), .ZN(n116) );
  INV_X1 U172 ( .A(n116), .ZN(n118) );
  FA_X1 U173 ( .A(n119), .B(n118), .CI(n117), .CO(n155), .S(n131) );
  OAI21_X1 U174 ( .B1(n122), .B2(n121), .A(n120), .ZN(n124) );
  NAND2_X1 U175 ( .A1(n122), .A2(n121), .ZN(n123) );
  NAND2_X1 U176 ( .A1(n124), .A2(n123), .ZN(n130) );
  NOR2_X1 U177 ( .A1(n27), .A2(n162), .ZN(n129) );
  NAND2_X1 U178 ( .A1(n131), .A2(n125), .ZN(n127) );
  NAND2_X1 U179 ( .A1(n127), .A2(n126), .ZN(n172) );
  OR2_X1 U180 ( .A1(n173), .A2(n172), .ZN(n128) );
  MUX2_X1 U181 ( .A(n328), .B(n128), .S(n325), .Z(n350) );
  XNOR2_X1 U182 ( .A(n130), .B(n129), .ZN(n132) );
  XNOR2_X1 U183 ( .A(n132), .B(n131), .ZN(n204) );
  INV_X1 U184 ( .A(n204), .ZN(n140) );
  NAND2_X1 U185 ( .A1(n133), .A2(n135), .ZN(n138) );
  NAND2_X1 U186 ( .A1(n133), .A2(n134), .ZN(n137) );
  NAND2_X1 U187 ( .A1(n135), .A2(n134), .ZN(n136) );
  NAND3_X1 U188 ( .A1(n138), .A2(n137), .A3(n136), .ZN(n203) );
  INV_X1 U189 ( .A(n203), .ZN(n139) );
  NAND2_X1 U190 ( .A1(n140), .A2(n139), .ZN(n141) );
  MUX2_X1 U191 ( .A(n329), .B(n141), .S(n14), .Z(n352) );
  FA_X1 U192 ( .A(n144), .B(n143), .CI(n142), .CO(n175), .S(n179) );
  OR2_X1 U193 ( .A1(\mult_x_1/n288 ), .A2(n327), .ZN(n145) );
  OAI22_X1 U194 ( .A1(n150), .A2(n327), .B1(n145), .B2(n148), .ZN(n187) );
  XNOR2_X1 U195 ( .A(n323), .B(\mult_x_1/n288 ), .ZN(n146) );
  XNOR2_X1 U196 ( .A(n323), .B(\mult_x_1/n287 ), .ZN(n149) );
  OAI22_X1 U197 ( .A1(n150), .A2(n146), .B1(n148), .B2(n149), .ZN(n186) );
  OAI22_X1 U198 ( .A1(n150), .A2(n149), .B1(n148), .B2(n147), .ZN(n182) );
  FA_X1 U199 ( .A(n153), .B(n152), .CI(n151), .CO(n144), .S(n181) );
  OR2_X1 U200 ( .A1(n179), .A2(n178), .ZN(n154) );
  MUX2_X1 U201 ( .A(n331), .B(n154), .S(n325), .Z(n356) );
  FA_X1 U202 ( .A(n157), .B(n156), .CI(n155), .CO(n168), .S(n173) );
  AOI21_X1 U203 ( .B1(n160), .B2(n159), .A(n158), .ZN(n161) );
  INV_X1 U204 ( .A(n161), .ZN(n164) );
  NOR2_X1 U205 ( .A1(n20), .A2(n162), .ZN(n163) );
  XOR2_X1 U206 ( .A(n164), .B(n163), .Z(n165) );
  XOR2_X1 U207 ( .A(n166), .B(n165), .Z(n167) );
  OR2_X1 U208 ( .A1(n168), .A2(n167), .ZN(n170) );
  NAND2_X1 U209 ( .A1(n168), .A2(n167), .ZN(n169) );
  NAND2_X1 U210 ( .A1(n170), .A2(n169), .ZN(n171) );
  MUX2_X1 U211 ( .A(n332), .B(n171), .S(n14), .Z(n358) );
  NAND2_X1 U212 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2_X1 U213 ( .A(n333), .B(n174), .S(n325), .Z(n360) );
  NOR2_X1 U214 ( .A1(n176), .A2(n175), .ZN(n177) );
  MUX2_X1 U215 ( .A(n334), .B(n177), .S(n325), .Z(n362) );
  NAND2_X1 U216 ( .A1(n179), .A2(n178), .ZN(n180) );
  MUX2_X1 U217 ( .A(n336), .B(n180), .S(n13), .Z(n366) );
  FA_X1 U218 ( .A(n183), .B(n182), .CI(n181), .CO(n178), .S(n190) );
  XNOR2_X1 U219 ( .A(n15), .B(\mult_x_1/n286 ), .ZN(n197) );
  OAI22_X1 U220 ( .A1(n210), .A2(n197), .B1(n212), .B2(n184), .ZN(n194) );
  XNOR2_X1 U221 ( .A(n322), .B(\mult_x_1/n284 ), .ZN(n195) );
  OAI22_X1 U222 ( .A1(n214), .A2(n195), .B1(n185), .B2(n17), .ZN(n193) );
  HA_X1 U223 ( .A(n187), .B(n186), .CO(n183), .S(n192) );
  NOR2_X1 U224 ( .A1(n190), .A2(n189), .ZN(n188) );
  MUX2_X1 U225 ( .A(n337), .B(n188), .S(n325), .Z(n368) );
  NAND2_X1 U226 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2_X1 U227 ( .A(n338), .B(n191), .S(n325), .Z(n370) );
  FA_X1 U228 ( .A(n194), .B(n193), .CI(n192), .CO(n189), .S(n199) );
  XNOR2_X1 U229 ( .A(n322), .B(\mult_x_1/n285 ), .ZN(n208) );
  OAI22_X1 U230 ( .A1(n214), .A2(n208), .B1(n195), .B2(n17), .ZN(n223) );
  AND2_X1 U231 ( .A1(n196), .A2(\mult_x_1/n288 ), .ZN(n222) );
  XNOR2_X1 U232 ( .A(n15), .B(\mult_x_1/n287 ), .ZN(n206) );
  OAI22_X1 U233 ( .A1(n210), .A2(n206), .B1(n212), .B2(n197), .ZN(n221) );
  OR2_X1 U234 ( .A1(n199), .A2(n198), .ZN(n230) );
  NAND2_X1 U235 ( .A1(n199), .A2(n198), .ZN(n228) );
  NAND2_X1 U236 ( .A1(n230), .A2(n228), .ZN(n200) );
  MUX2_X1 U237 ( .A(n339), .B(n200), .S(n14), .Z(n372) );
  NAND2_X1 U238 ( .A1(n204), .A2(n203), .ZN(n205) );
  MUX2_X1 U239 ( .A(n342), .B(n205), .S(n325), .Z(n378) );
  XNOR2_X1 U240 ( .A(n15), .B(\mult_x_1/n288 ), .ZN(n207) );
  OAI22_X1 U241 ( .A1(n210), .A2(n207), .B1(n212), .B2(n206), .ZN(n225) );
  XNOR2_X1 U242 ( .A(n322), .B(\mult_x_1/n286 ), .ZN(n211) );
  OAI22_X1 U243 ( .A1(n214), .A2(n211), .B1(n208), .B2(n17), .ZN(n224) );
  OR2_X1 U244 ( .A1(\mult_x_1/n288 ), .A2(n19), .ZN(n209) );
  OAI22_X1 U245 ( .A1(n210), .A2(n19), .B1(n209), .B2(n212), .ZN(n218) );
  OR2_X1 U246 ( .A1(n219), .A2(n218), .ZN(n263) );
  XNOR2_X1 U247 ( .A(n322), .B(\mult_x_1/n287 ), .ZN(n213) );
  OAI22_X1 U248 ( .A1(n214), .A2(n213), .B1(n211), .B2(n17), .ZN(n217) );
  AND2_X1 U249 ( .A1(\mult_x_1/n288 ), .A2(n36), .ZN(n216) );
  NOR2_X1 U250 ( .A1(n217), .A2(n216), .ZN(n256) );
  OAI22_X1 U251 ( .A1(n214), .A2(\mult_x_1/n288 ), .B1(n213), .B2(n17), .ZN(
        n253) );
  OR2_X1 U252 ( .A1(\mult_x_1/n288 ), .A2(n30), .ZN(n215) );
  NAND2_X1 U253 ( .A1(n215), .A2(n214), .ZN(n252) );
  NAND2_X1 U254 ( .A1(n253), .A2(n252), .ZN(n259) );
  NAND2_X1 U255 ( .A1(n217), .A2(n216), .ZN(n257) );
  OAI21_X1 U256 ( .B1(n256), .B2(n259), .A(n257), .ZN(n264) );
  NAND2_X1 U257 ( .A1(n219), .A2(n218), .ZN(n262) );
  INV_X1 U258 ( .A(n262), .ZN(n220) );
  AOI21_X1 U259 ( .B1(n263), .B2(n264), .A(n220), .ZN(n270) );
  FA_X1 U260 ( .A(n223), .B(n222), .CI(n221), .CO(n198), .S(n227) );
  HA_X1 U261 ( .A(n225), .B(n224), .CO(n226), .S(n219) );
  NOR2_X1 U262 ( .A1(n227), .A2(n226), .ZN(n267) );
  NAND2_X1 U263 ( .A1(n227), .A2(n226), .ZN(n268) );
  OAI21_X1 U264 ( .B1(n270), .B2(n267), .A(n268), .ZN(n232) );
  INV_X1 U265 ( .A(n228), .ZN(n229) );
  AOI21_X1 U266 ( .B1(n230), .B2(n232), .A(n229), .ZN(n231) );
  MUX2_X1 U267 ( .A(n344), .B(n231), .S(n13), .Z(n382) );
  MUX2_X1 U268 ( .A(n345), .B(n232), .S(n325), .Z(n384) );
  FA_X1 U269 ( .A(n235), .B(n234), .CI(n233), .CO(n108), .S(n236) );
  MUX2_X1 U270 ( .A(n346), .B(n236), .S(n325), .Z(n386) );
  NAND2_X1 U271 ( .A1(n237), .A2(n21), .ZN(n241) );
  NAND2_X1 U272 ( .A1(n237), .A2(n238), .ZN(n240) );
  NAND2_X1 U273 ( .A1(n21), .A2(n238), .ZN(n239) );
  NAND3_X1 U274 ( .A1(n241), .A2(n240), .A3(n239), .ZN(n242) );
  MUX2_X1 U275 ( .A(n347), .B(n242), .S(n14), .Z(n388) );
  FA_X1 U276 ( .A(n244), .B(n243), .CI(n29), .CO(n201), .S(n245) );
  MUX2_X1 U277 ( .A(n348), .B(n245), .S(n325), .Z(n390) );
  FA_X1 U278 ( .A(n248), .B(n247), .CI(n246), .CO(n250), .S(n176) );
  MUX2_X1 U279 ( .A(n349), .B(n250), .S(n325), .Z(n392) );
  MUX2_X1 U280 ( .A(product[0]), .B(n515), .S(n325), .Z(n407) );
  MUX2_X1 U281 ( .A(n515), .B(n516), .S(n325), .Z(n409) );
  AND2_X1 U282 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n251) );
  MUX2_X1 U283 ( .A(n516), .B(n251), .S(n325), .Z(n411) );
  MUX2_X1 U284 ( .A(product[1]), .B(n518), .S(n13), .Z(n413) );
  MUX2_X1 U285 ( .A(n518), .B(n519), .S(n325), .Z(n415) );
  OR2_X1 U286 ( .A1(n253), .A2(n252), .ZN(n254) );
  AND2_X1 U287 ( .A1(n254), .A2(n259), .ZN(n255) );
  MUX2_X1 U288 ( .A(n519), .B(n255), .S(n14), .Z(n417) );
  MUX2_X1 U289 ( .A(product[2]), .B(n521), .S(n325), .Z(n419) );
  MUX2_X1 U290 ( .A(n521), .B(n522), .S(n13), .Z(n421) );
  INV_X1 U291 ( .A(n256), .ZN(n258) );
  NAND2_X1 U292 ( .A1(n258), .A2(n257), .ZN(n260) );
  XOR2_X1 U293 ( .A(n260), .B(n259), .Z(n261) );
  MUX2_X1 U294 ( .A(n522), .B(n261), .S(n325), .Z(n423) );
  MUX2_X1 U295 ( .A(product[3]), .B(n524), .S(n14), .Z(n425) );
  MUX2_X1 U296 ( .A(n524), .B(n525), .S(n325), .Z(n427) );
  NAND2_X1 U297 ( .A1(n263), .A2(n262), .ZN(n265) );
  XNOR2_X1 U298 ( .A(n265), .B(n264), .ZN(n266) );
  MUX2_X1 U299 ( .A(n525), .B(n266), .S(n13), .Z(n429) );
  MUX2_X1 U300 ( .A(product[4]), .B(n527), .S(n14), .Z(n431) );
  MUX2_X1 U301 ( .A(n527), .B(n528), .S(n13), .Z(n433) );
  INV_X1 U302 ( .A(n267), .ZN(n269) );
  NAND2_X1 U303 ( .A1(n269), .A2(n268), .ZN(n271) );
  XOR2_X1 U304 ( .A(n271), .B(n270), .Z(n272) );
  MUX2_X1 U305 ( .A(n528), .B(n272), .S(n14), .Z(n435) );
  MUX2_X1 U306 ( .A(product[5]), .B(n530), .S(n325), .Z(n437) );
  XNOR2_X1 U307 ( .A(n339), .B(n345), .ZN(n273) );
  MUX2_X1 U308 ( .A(n530), .B(n273), .S(n13), .Z(n439) );
  MUX2_X1 U309 ( .A(product[6]), .B(n532), .S(n325), .Z(n441) );
  NAND2_X1 U310 ( .A1(n396), .A2(n338), .ZN(n274) );
  XOR2_X1 U311 ( .A(n274), .B(n344), .Z(n275) );
  MUX2_X1 U312 ( .A(n532), .B(n275), .S(n14), .Z(n443) );
  MUX2_X1 U313 ( .A(product[7]), .B(n534), .S(n325), .Z(n445) );
  OAI21_X1 U314 ( .B1(n337), .B2(n344), .A(n338), .ZN(n278) );
  NAND2_X1 U315 ( .A1(n331), .A2(n336), .ZN(n276) );
  XNOR2_X1 U316 ( .A(n278), .B(n276), .ZN(n277) );
  MUX2_X1 U317 ( .A(n534), .B(n277), .S(n325), .Z(n447) );
  MUX2_X1 U318 ( .A(product[8]), .B(n536), .S(n13), .Z(n449) );
  AOI21_X1 U319 ( .B1(n278), .B2(n331), .A(n398), .ZN(n281) );
  NAND2_X1 U320 ( .A1(n399), .A2(n335), .ZN(n279) );
  XOR2_X1 U321 ( .A(n281), .B(n279), .Z(n280) );
  MUX2_X1 U322 ( .A(n536), .B(n280), .S(n325), .Z(n451) );
  MUX2_X1 U323 ( .A(product[9]), .B(n538), .S(n13), .Z(n453) );
  OAI21_X1 U324 ( .B1(n281), .B2(n334), .A(n335), .ZN(n292) );
  INV_X1 U325 ( .A(n292), .ZN(n285) );
  NOR2_X1 U326 ( .A1(n348), .A2(n349), .ZN(n289) );
  INV_X1 U327 ( .A(n289), .ZN(n282) );
  NAND2_X1 U328 ( .A1(n348), .A2(n349), .ZN(n290) );
  NAND2_X1 U329 ( .A1(n282), .A2(n290), .ZN(n283) );
  XOR2_X1 U330 ( .A(n285), .B(n283), .Z(n284) );
  MUX2_X1 U331 ( .A(n538), .B(n284), .S(n325), .Z(n455) );
  MUX2_X1 U332 ( .A(product[10]), .B(n540), .S(n325), .Z(n457) );
  OAI21_X1 U333 ( .B1(n285), .B2(n289), .A(n290), .ZN(n287) );
  NAND2_X1 U334 ( .A1(n400), .A2(n341), .ZN(n286) );
  XNOR2_X1 U335 ( .A(n287), .B(n286), .ZN(n288) );
  MUX2_X1 U336 ( .A(n540), .B(n288), .S(n13), .Z(n459) );
  MUX2_X1 U337 ( .A(product[11]), .B(n542), .S(n325), .Z(n461) );
  NOR2_X1 U338 ( .A1(n340), .A2(n289), .ZN(n293) );
  OAI21_X1 U339 ( .B1(n340), .B2(n290), .A(n341), .ZN(n291) );
  AOI21_X1 U340 ( .B1(n293), .B2(n292), .A(n291), .ZN(n319) );
  NOR2_X1 U341 ( .A1(n346), .A2(n347), .ZN(n305) );
  INV_X1 U342 ( .A(n305), .ZN(n315) );
  NAND2_X1 U343 ( .A1(n346), .A2(n347), .ZN(n307) );
  NAND2_X1 U344 ( .A1(n315), .A2(n307), .ZN(n294) );
  XOR2_X1 U345 ( .A(n319), .B(n294), .Z(n295) );
  MUX2_X1 U346 ( .A(n542), .B(n295), .S(n13), .Z(n463) );
  MUX2_X1 U347 ( .A(product[12]), .B(n544), .S(n325), .Z(n465) );
  OAI21_X1 U348 ( .B1(n319), .B2(n305), .A(n307), .ZN(n297) );
  NAND2_X1 U349 ( .A1(n330), .A2(n343), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  MUX2_X1 U351 ( .A(n544), .B(n298), .S(n14), .Z(n467) );
  MUX2_X1 U352 ( .A(product[13]), .B(n546), .S(n325), .Z(n469) );
  NAND2_X1 U353 ( .A1(n315), .A2(n330), .ZN(n301) );
  INV_X1 U354 ( .A(n307), .ZN(n299) );
  AOI21_X1 U355 ( .B1(n299), .B2(n330), .A(n401), .ZN(n300) );
  OAI21_X1 U356 ( .B1(n319), .B2(n301), .A(n300), .ZN(n303) );
  NAND2_X1 U357 ( .A1(n329), .A2(n342), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  MUX2_X1 U359 ( .A(n546), .B(n304), .S(n325), .Z(n471) );
  MUX2_X1 U360 ( .A(product[14]), .B(n548), .S(n14), .Z(n473) );
  NAND2_X1 U361 ( .A1(n330), .A2(n329), .ZN(n313) );
  OR2_X1 U362 ( .A1(n305), .A2(n313), .ZN(n309) );
  AOI21_X1 U363 ( .B1(n401), .B2(n329), .A(n397), .ZN(n306) );
  OAI21_X1 U364 ( .B1(n313), .B2(n307), .A(n306), .ZN(n316) );
  INV_X1 U365 ( .A(n316), .ZN(n308) );
  OAI21_X1 U366 ( .B1(n319), .B2(n309), .A(n308), .ZN(n311) );
  NAND2_X1 U367 ( .A1(n328), .A2(n333), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  MUX2_X1 U369 ( .A(n548), .B(n312), .S(n325), .Z(n475) );
  MUX2_X1 U370 ( .A(product[15]), .B(n550), .S(n325), .Z(n477) );
  NOR2_X1 U371 ( .A1(n313), .A2(n395), .ZN(n314) );
  NAND2_X1 U372 ( .A1(n315), .A2(n314), .ZN(n318) );
  AOI21_X1 U373 ( .B1(n316), .B2(n328), .A(n394), .ZN(n317) );
  OAI21_X1 U374 ( .B1(n319), .B2(n318), .A(n317), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n320), .B(n332), .ZN(n321) );
  MUX2_X1 U376 ( .A(n550), .B(n321), .S(n14), .Z(n479) );
  MUX2_X1 U377 ( .A(\mult_x_1/n288 ), .B(B_extended[0]), .S(n325), .Z(n481) );
  MUX2_X1 U378 ( .A(\mult_x_1/n287 ), .B(B_extended[1]), .S(n325), .Z(n483) );
  MUX2_X1 U379 ( .A(\mult_x_1/n286 ), .B(B_extended[2]), .S(n325), .Z(n485) );
  MUX2_X1 U380 ( .A(\mult_x_1/n285 ), .B(B_extended[3]), .S(n325), .Z(n487) );
  MUX2_X1 U381 ( .A(\mult_x_1/n284 ), .B(B_extended[4]), .S(n325), .Z(n489) );
  MUX2_X1 U382 ( .A(\mult_x_1/n283 ), .B(B_extended[5]), .S(n325), .Z(n491) );
  MUX2_X1 U383 ( .A(\mult_x_1/n282 ), .B(B_extended[6]), .S(n13), .Z(n493) );
  MUX2_X1 U384 ( .A(\mult_x_1/n281 ), .B(B_extended[7]), .S(n325), .Z(n495) );
  MUX2_X1 U385 ( .A(\mult_x_1/n180 ), .B(A_extended[0]), .S(n325), .Z(n497) );
  MUX2_X1 U386 ( .A(n322), .B(A_extended[1]), .S(n325), .Z(n499) );
  MUX2_X1 U387 ( .A(\mult_x_1/a[2] ), .B(A_extended[2]), .S(n325), .Z(n501) );
  MUX2_X1 U388 ( .A(n15), .B(A_extended[3]), .S(n14), .Z(n503) );
  MUX2_X1 U389 ( .A(\mult_x_1/a[4] ), .B(A_extended[4]), .S(n325), .Z(n505) );
  MUX2_X1 U390 ( .A(n323), .B(A_extended[5]), .S(n325), .Z(n507) );
  MUX2_X1 U391 ( .A(\mult_x_1/a[6] ), .B(A_extended[6]), .S(n13), .Z(n509) );
  MUX2_X1 U392 ( .A(n324), .B(A_extended[7]), .S(n325), .Z(n511) );
  OR2_X1 U393 ( .A1(n325), .A2(n552), .ZN(n513) );
endmodule


module conv_128_32_DW_mult_pipe_J1_26 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n394, n396, n398, n400, n402, n404, n406, n408, n410, n412,
         n414, n416, n418, n420, n422, n424, n426, n428, n430, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n508, n510, n512, n514,
         n516, n518, n520, n522, n524, n526, n528, n530, n532, n534, n536,
         n538, n540, n542, n544, n546, n548, n550, n552, n554, n556, n558,
         n560, n562, n564, n566, n568, n570, n572, n574, n576, n578, n580,
         n582, n584, n586, n588, n590, n592, n594, n596, n598, n600, n602,
         n604, n606, n608, n610, n612, n614, n616, n633, n634;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n616), .CK(clk), .Q(n633), 
        .QN(n452) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n612), .CK(clk), .QN(n454) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n608), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n456) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(rst_n), .SE(n606), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n457) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(rst_n), .SE(n604), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n458) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(rst_n), .SE(n600), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n460) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(rst_n), .SE(n598), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n461) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(rst_n), .SE(n596), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n462) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n594), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n463) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n592), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n464) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n451), .SE(n590), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n465) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n588), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n466) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n451), .SE(n586), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n467) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n451), .SE(n584), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n468) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n451), .SE(n582), .CK(clk), .QN(n469)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n451), .SE(n580), .CK(clk), .Q(
        product[15]), .QN(n470) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n451), .SE(n578), .CK(clk), .QN(n471)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n451), .SE(n576), .CK(clk), .Q(
        product[14]), .QN(n472) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n451), .SE(n574), .CK(clk), .QN(n473)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(rst_n), .SE(n572), .CK(clk), .Q(
        product[13]), .QN(n474) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(rst_n), .SE(n570), .CK(clk), .QN(n475) );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n568), .CK(clk), .Q(
        product[12]), .QN(n476) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n451), .SE(n566), .CK(clk), .QN(n477)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n451), .SE(n564), .CK(clk), .Q(
        product[11]), .QN(n478) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n451), .SE(n562), .CK(clk), .QN(n479)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n451), .SE(n560), .CK(clk), .Q(
        product[10]), .QN(n480) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n451), .SE(n558), .CK(clk), .QN(n481)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n451), .SE(n556), .CK(clk), .Q(
        product[9]), .QN(n482) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n451), .SE(n554), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n451), .SE(n552), .CK(clk), .Q(
        product[8]), .QN(n484) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n550), .CK(clk), .QN(n485) );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n548), .CK(clk), .Q(
        product[7]), .QN(n486) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n546), .CK(clk), .QN(n487) );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n544), .CK(clk), .Q(
        product[6]), .QN(n488) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n542), .CK(clk), .QN(n489) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n540), .CK(clk), .QN(n490) );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n538), .CK(clk), .Q(
        product[5]), .QN(n491) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n536), .CK(clk), .QN(n492) );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n534), .CK(clk), .QN(n493) );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n532), .CK(clk), .Q(
        product[4]), .QN(n494) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n530), .CK(clk), .QN(n495) );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n528), .CK(clk), .QN(n496) );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n526), .CK(clk), .Q(
        product[3]), .QN(n497) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n451), .SE(n524), .CK(clk), .QN(n498)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n522), .CK(clk), .QN(n499) );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n520), .CK(clk), .Q(
        product[2]), .QN(n500) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n518), .CK(clk), .QN(n501) );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n516), .CK(clk), .QN(n502) );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n514), .CK(clk), .Q(
        product[1]), .QN(n503) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n451), .SE(n512), .CK(clk), .QN(n504)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n510), .CK(clk), .QN(n505) );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n508), .CK(clk), .Q(
        product[0]), .QN(n506) );
  SDFF_X2 clk_r_REG0_S1 ( .D(1'b0), .SI(rst_n), .SE(n614), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n453) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(rst_n), .SE(n602), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n634), .SE(n426), .CK(
        clk), .Q(n434), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n634), .SI(1'b1), .SE(n430), .CK(clk), 
        .Q(n391), .QN(n432) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n634), .SI(1'b1), .SE(n428), .CK(clk), 
        .Q(n390), .QN(n433) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n634), .SI(1'b1), .SE(n424), .CK(clk), 
        .Q(n388), .QN(n435) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n634), .SE(n422), .CK(
        clk), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n634), .SE(n420), .CK(
        clk), .Q(n436), .QN(n386) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n634), .SI(1'b1), .SE(n418), .CK(clk), 
        .Q(n385), .QN(n437) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n634), .SI(1'b1), .SE(n416), .CK(clk), 
        .Q(n384), .QN(n438) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n634), .SI(1'b1), .SE(n414), .CK(clk), 
        .Q(n383), .QN(n439) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n634), .SI(1'b1), .SE(n412), .CK(clk), 
        .Q(n382), .QN(n440) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n634), .SI(1'b1), .SE(n410), .CK(clk), 
        .Q(n381), .QN(n441) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n634), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n380), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n634), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n379), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n634), .SI(1'b1), .SE(n404), .CK(clk), 
        .Q(n378), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n634), .SI(1'b1), .SE(n402), .CK(clk), 
        .Q(n377), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n634), .SE(n400), .CK(
        clk), .Q(n446), .QN(n376) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n634), .SE(n398), .CK(
        clk), .Q(n447), .QN(n375) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n634), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n374), .QN(n448) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n634), .SI(1'b1), .SE(n394), .CK(clk), 
        .Q(n373), .QN(n449) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n634), .SI(1'b1), .SE(n392), .CK(clk), 
        .Q(n372), .QN(n450) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n610), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n455) );
  BUF_X1 U2 ( .A(n344), .Z(n257) );
  INV_X1 U3 ( .A(rst_n), .ZN(n634) );
  BUF_X2 U4 ( .A(n344), .Z(n5) );
  CLKBUF_X2 U5 ( .A(n265), .Z(n326) );
  BUF_X1 U6 ( .A(n265), .Z(n273) );
  INV_X1 U7 ( .A(n634), .ZN(n451) );
  OAI21_X1 U8 ( .B1(n162), .B2(n161), .A(n287), .ZN(n101) );
  BUF_X1 U9 ( .A(n344), .Z(n287) );
  INV_X2 U10 ( .A(n273), .ZN(n371) );
  INV_X2 U11 ( .A(n265), .ZN(n344) );
  AOI22_X1 U12 ( .A1(n240), .A2(n181), .B1(n238), .B2(n237), .ZN(n229) );
  NAND2_X1 U13 ( .A1(n11), .A2(n10), .ZN(n233) );
  OAI21_X1 U14 ( .B1(n56), .B2(n55), .A(n54), .ZN(n11) );
  NAND2_X1 U15 ( .A1(n56), .A2(n55), .ZN(n10) );
  NAND2_X1 U16 ( .A1(n28), .A2(n29), .ZN(n18) );
  NAND2_X1 U17 ( .A1(n452), .A2(\mult_x_1/n310 ), .ZN(n176) );
  CLKBUF_X2 U18 ( .A(\mult_x_1/n313 ), .Z(n212) );
  AND2_X1 U19 ( .A1(\mult_x_1/n310 ), .A2(n633), .ZN(n6) );
  XNOR2_X1 U20 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n95) );
  NAND2_X1 U21 ( .A1(n7), .A2(n257), .ZN(n189) );
  NAND2_X1 U22 ( .A1(n242), .A2(n243), .ZN(n7) );
  NAND2_X1 U23 ( .A1(n8), .A2(n241), .ZN(n426) );
  NAND2_X1 U24 ( .A1(n16), .A2(n15), .ZN(n8) );
  XNOR2_X1 U25 ( .A(n9), .B(n171), .ZN(n230) );
  INV_X1 U26 ( .A(n172), .ZN(n9) );
  OAI21_X1 U27 ( .B1(n243), .B2(n242), .A(n5), .ZN(n244) );
  NOR2_X1 U28 ( .A1(n176), .A2(n467), .ZN(n173) );
  XNOR2_X1 U29 ( .A(n56), .B(n12), .ZN(n64) );
  XNOR2_X1 U30 ( .A(n55), .B(n54), .ZN(n12) );
  OR2_X1 U31 ( .A1(n13), .A2(n261), .ZN(n258) );
  NAND2_X1 U32 ( .A1(n14), .A2(n257), .ZN(n13) );
  XNOR2_X1 U33 ( .A(n237), .B(n238), .ZN(n239) );
  NOR2_X1 U34 ( .A1(n176), .A2(n466), .ZN(n238) );
  INV_X1 U35 ( .A(n260), .ZN(n14) );
  NOR2_X1 U36 ( .A1(n246), .A2(n326), .ZN(n15) );
  INV_X1 U37 ( .A(n247), .ZN(n16) );
  NAND2_X1 U38 ( .A1(n17), .A2(n249), .ZN(n404) );
  NAND2_X1 U39 ( .A1(n248), .A2(n344), .ZN(n17) );
  INV_X1 U40 ( .A(n63), .ZN(n59) );
  XNOR2_X1 U41 ( .A(n57), .B(n233), .ZN(n252) );
  NAND2_X1 U42 ( .A1(n66), .A2(n65), .ZN(n136) );
  NAND2_X1 U43 ( .A1(n64), .A2(n63), .ZN(n65) );
  NAND2_X1 U44 ( .A1(n62), .A2(n61), .ZN(n66) );
  NAND2_X1 U45 ( .A1(n60), .A2(n59), .ZN(n61) );
  XNOR2_X1 U46 ( .A(n62), .B(n37), .ZN(n141) );
  XNOR2_X1 U47 ( .A(n64), .B(n63), .ZN(n37) );
  NAND2_X1 U48 ( .A1(n256), .A2(n255), .ZN(n260) );
  NAND2_X1 U49 ( .A1(n254), .A2(n253), .ZN(n255) );
  OAI21_X1 U50 ( .B1(n254), .B2(n253), .A(n252), .ZN(n256) );
  NAND2_X1 U51 ( .A1(n29), .A2(n28), .ZN(n119) );
  INV_X1 U52 ( .A(n455), .ZN(n19) );
  INV_X1 U53 ( .A(n27), .ZN(n209) );
  XNOR2_X1 U54 ( .A(\mult_x_1/n310 ), .B(n454), .ZN(n28) );
  INV_X1 U55 ( .A(n64), .ZN(n60) );
  CLKBUF_X1 U56 ( .A(\mult_x_1/n311 ), .Z(n20) );
  INV_X2 U57 ( .A(n273), .ZN(n21) );
  INV_X2 U58 ( .A(n273), .ZN(n366) );
  AND2_X1 U59 ( .A1(n233), .A2(n232), .ZN(n22) );
  AND2_X1 U60 ( .A1(n141), .A2(n140), .ZN(n23) );
  XOR2_X1 U61 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n24) );
  XNOR2_X1 U62 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n312 ), .ZN(n25) );
  NAND2_X2 U63 ( .A1(n24), .A2(n25), .ZN(n109) );
  XNOR2_X1 U64 ( .A(n20), .B(\mult_x_1/n285 ), .ZN(n34) );
  BUF_X2 U65 ( .A(n25), .Z(n194) );
  XNOR2_X1 U66 ( .A(n20), .B(\mult_x_1/n284 ), .ZN(n52) );
  OAI22_X1 U67 ( .A1(n109), .A2(n34), .B1(n194), .B2(n52), .ZN(n51) );
  XNOR2_X1 U68 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n312 ), .ZN(n26) );
  XOR2_X1 U69 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .Z(n27) );
  OR2_X2 U70 ( .A1(n26), .A2(n27), .ZN(n207) );
  BUF_X2 U71 ( .A(\mult_x_1/n312 ), .Z(n205) );
  XNOR2_X1 U72 ( .A(n205), .B(\mult_x_1/n283 ), .ZN(n36) );
  XNOR2_X1 U73 ( .A(n205), .B(\mult_x_1/n282 ), .ZN(n53) );
  OAI22_X1 U74 ( .A1(n207), .A2(n36), .B1(n209), .B2(n53), .ZN(n50) );
  XNOR2_X1 U75 ( .A(n455), .B(n454), .ZN(n29) );
  INV_X1 U76 ( .A(n29), .ZN(n39) );
  INV_X2 U77 ( .A(n39), .ZN(n120) );
  OR2_X1 U78 ( .A1(\mult_x_1/n288 ), .A2(n453), .ZN(n30) );
  OAI22_X1 U79 ( .A1(n120), .A2(n30), .B1(n119), .B2(n453), .ZN(n42) );
  XNOR2_X1 U80 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n31) );
  XNOR2_X1 U81 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n32) );
  OAI22_X1 U82 ( .A1(n119), .A2(n31), .B1(n120), .B2(n32), .ZN(n41) );
  XNOR2_X1 U83 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n48) );
  OAI22_X1 U84 ( .A1(n119), .A2(n32), .B1(n120), .B2(n48), .ZN(n56) );
  NAND2_X1 U85 ( .A1(n212), .A2(n460), .ZN(n213) );
  XNOR2_X1 U86 ( .A(n212), .B(\mult_x_1/n281 ), .ZN(n35) );
  AND2_X1 U87 ( .A1(n633), .A2(\mult_x_1/n281 ), .ZN(n82) );
  XNOR2_X1 U88 ( .A(n82), .B(n212), .ZN(n46) );
  OAI22_X1 U89 ( .A1(n213), .A2(n35), .B1(n46), .B2(n460), .ZN(n55) );
  XOR2_X1 U90 ( .A(n6), .B(\mult_x_1/n310 ), .Z(n33) );
  AND2_X1 U91 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n54) );
  XNOR2_X1 U92 ( .A(n20), .B(\mult_x_1/n286 ), .ZN(n107) );
  OAI22_X1 U93 ( .A1(n109), .A2(n107), .B1(n194), .B2(n34), .ZN(n45) );
  XNOR2_X1 U94 ( .A(n212), .B(\mult_x_1/n282 ), .ZN(n38) );
  OAI22_X1 U95 ( .A1(n213), .A2(n38), .B1(n35), .B2(n460), .ZN(n44) );
  XNOR2_X1 U96 ( .A(n205), .B(\mult_x_1/n284 ), .ZN(n40) );
  OAI22_X1 U97 ( .A1(n207), .A2(n40), .B1(n209), .B2(n36), .ZN(n43) );
  XNOR2_X1 U98 ( .A(n212), .B(\mult_x_1/n283 ), .ZN(n152) );
  OAI22_X1 U99 ( .A1(n213), .A2(n152), .B1(n38), .B2(n460), .ZN(n112) );
  AND2_X1 U100 ( .A1(n39), .A2(\mult_x_1/n288 ), .ZN(n111) );
  XNOR2_X1 U101 ( .A(n205), .B(\mult_x_1/n285 ), .ZN(n151) );
  OAI22_X1 U102 ( .A1(n207), .A2(n151), .B1(n209), .B2(n40), .ZN(n110) );
  HA_X1 U103 ( .A(n42), .B(n41), .CO(n49), .S(n103) );
  FA_X1 U104 ( .A(n45), .B(n44), .CI(n43), .CO(n63), .S(n102) );
  INV_X1 U105 ( .A(en), .ZN(n265) );
  OAI22_X1 U106 ( .A1(n23), .A2(n326), .B1(n287), .B2(n440), .ZN(n412) );
  AOI21_X1 U107 ( .B1(n213), .B2(n460), .A(n46), .ZN(n47) );
  INV_X1 U108 ( .A(n47), .ZN(n175) );
  XNOR2_X1 U109 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n85) );
  OAI22_X1 U110 ( .A1(n18), .A2(n48), .B1(n120), .B2(n85), .ZN(n174) );
  FA_X1 U111 ( .A(n51), .B(n50), .CI(n49), .CO(n253), .S(n62) );
  XNOR2_X1 U112 ( .A(n254), .B(n253), .ZN(n58) );
  XNOR2_X1 U113 ( .A(n19), .B(\mult_x_1/n283 ), .ZN(n84) );
  OAI22_X1 U114 ( .A1(n109), .A2(n52), .B1(n194), .B2(n84), .ZN(n178) );
  XNOR2_X1 U115 ( .A(n205), .B(\mult_x_1/n281 ), .ZN(n83) );
  OAI22_X1 U116 ( .A1(n207), .A2(n53), .B1(n209), .B2(n83), .ZN(n177) );
  XNOR2_X1 U117 ( .A(n178), .B(n177), .ZN(n232) );
  INV_X1 U118 ( .A(n232), .ZN(n57) );
  XNOR2_X1 U119 ( .A(n58), .B(n252), .ZN(n137) );
  NOR2_X1 U120 ( .A1(n137), .A2(n136), .ZN(n67) );
  NAND2_X1 U121 ( .A1(n67), .A2(n257), .ZN(n69) );
  OR2_X1 U122 ( .A1(n344), .A2(n443), .ZN(n68) );
  NAND2_X1 U123 ( .A1(n69), .A2(n68), .ZN(n406) );
  NOR2_X1 U144 ( .A1(n462), .A2(n176), .ZN(n117) );
  XNOR2_X1 U145 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n70) );
  XNOR2_X1 U146 ( .A(n82), .B(\mult_x_1/n310 ), .ZN(n118) );
  OAI22_X1 U147 ( .A1(n18), .A2(n70), .B1(n118), .B2(n120), .ZN(n125) );
  INV_X1 U148 ( .A(n125), .ZN(n116) );
  XNOR2_X1 U149 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n73) );
  OAI22_X1 U150 ( .A1(n18), .A2(n73), .B1(n120), .B2(n70), .ZN(n76) );
  XNOR2_X1 U151 ( .A(n19), .B(\mult_x_1/n281 ), .ZN(n86) );
  XNOR2_X1 U152 ( .A(n82), .B(n19), .ZN(n71) );
  OAI22_X1 U153 ( .A1(n109), .A2(n86), .B1(n71), .B2(n194), .ZN(n75) );
  AOI21_X1 U154 ( .B1(n194), .B2(n109), .A(n71), .ZN(n72) );
  INV_X1 U155 ( .A(n72), .ZN(n74) );
  INV_X1 U156 ( .A(n75), .ZN(n93) );
  XNOR2_X1 U157 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n94) );
  OAI22_X1 U158 ( .A1(n18), .A2(n94), .B1(n120), .B2(n73), .ZN(n92) );
  NOR2_X1 U159 ( .A1(n464), .A2(n176), .ZN(n91) );
  NOR2_X1 U160 ( .A1(n463), .A2(n176), .ZN(n80) );
  FA_X1 U161 ( .A(n76), .B(n74), .CI(n75), .CO(n115), .S(n79) );
  OR2_X1 U162 ( .A1(n133), .A2(n132), .ZN(n77) );
  NAND2_X1 U163 ( .A1(n257), .A2(n77), .ZN(n78) );
  OAI21_X1 U164 ( .B1(n257), .B2(n450), .A(n78), .ZN(n392) );
  FA_X1 U165 ( .A(n81), .B(n80), .CI(n79), .CO(n132), .S(n162) );
  XNOR2_X1 U166 ( .A(n82), .B(n205), .ZN(n96) );
  OAI22_X1 U167 ( .A1(n207), .A2(n83), .B1(n96), .B2(n209), .ZN(n183) );
  INV_X1 U168 ( .A(n183), .ZN(n236) );
  XNOR2_X1 U169 ( .A(n20), .B(\mult_x_1/n282 ), .ZN(n87) );
  OAI22_X1 U170 ( .A1(n109), .A2(n84), .B1(n194), .B2(n87), .ZN(n235) );
  OAI22_X1 U171 ( .A1(n18), .A2(n85), .B1(n120), .B2(n95), .ZN(n234) );
  NOR2_X1 U172 ( .A1(n465), .A2(n176), .ZN(n170) );
  NAND2_X1 U173 ( .A1(n172), .A2(n170), .ZN(n90) );
  OAI22_X1 U174 ( .A1(n109), .A2(n87), .B1(n194), .B2(n86), .ZN(n169) );
  NAND2_X1 U175 ( .A1(n172), .A2(n169), .ZN(n89) );
  NAND2_X1 U176 ( .A1(n170), .A2(n169), .ZN(n88) );
  NAND3_X1 U177 ( .A1(n90), .A2(n89), .A3(n88), .ZN(n168) );
  FA_X1 U178 ( .A(n93), .B(n91), .CI(n92), .CO(n81), .S(n166) );
  NAND2_X1 U179 ( .A1(n168), .A2(n166), .ZN(n100) );
  OAI22_X1 U180 ( .A1(n18), .A2(n95), .B1(n120), .B2(n94), .ZN(n184) );
  AOI21_X1 U181 ( .B1(n209), .B2(n207), .A(n96), .ZN(n97) );
  INV_X1 U182 ( .A(n97), .ZN(n182) );
  NAND2_X1 U183 ( .A1(n168), .A2(n165), .ZN(n99) );
  NAND2_X1 U184 ( .A1(n166), .A2(n165), .ZN(n98) );
  NAND3_X1 U185 ( .A1(n100), .A2(n99), .A3(n98), .ZN(n161) );
  OAI21_X1 U186 ( .B1(n5), .B2(n449), .A(n101), .ZN(n394) );
  FA_X1 U187 ( .A(n104), .B(n103), .CI(n102), .CO(n140), .S(n145) );
  OR2_X1 U188 ( .A1(\mult_x_1/n288 ), .A2(n455), .ZN(n105) );
  OAI22_X1 U189 ( .A1(n109), .A2(n455), .B1(n105), .B2(n194), .ZN(n154) );
  XNOR2_X1 U190 ( .A(n20), .B(\mult_x_1/n288 ), .ZN(n106) );
  XNOR2_X1 U191 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n108) );
  OAI22_X1 U192 ( .A1(n109), .A2(n106), .B1(n194), .B2(n108), .ZN(n153) );
  OAI22_X1 U193 ( .A1(n109), .A2(n108), .B1(n194), .B2(n107), .ZN(n149) );
  FA_X1 U194 ( .A(n112), .B(n111), .CI(n110), .CO(n104), .S(n148) );
  OR2_X1 U195 ( .A1(n145), .A2(n144), .ZN(n113) );
  NAND2_X1 U196 ( .A1(n287), .A2(n113), .ZN(n114) );
  OAI21_X1 U197 ( .B1(n287), .B2(n447), .A(n114), .ZN(n398) );
  FA_X1 U198 ( .A(n117), .B(n116), .CI(n115), .CO(n127), .S(n133) );
  AOI21_X1 U199 ( .B1(n120), .B2(n18), .A(n118), .ZN(n121) );
  INV_X1 U200 ( .A(n121), .ZN(n123) );
  NOR2_X1 U201 ( .A1(n461), .A2(n176), .ZN(n122) );
  XOR2_X1 U202 ( .A(n123), .B(n122), .Z(n124) );
  XOR2_X1 U203 ( .A(n125), .B(n124), .Z(n126) );
  OR2_X1 U204 ( .A1(n127), .A2(n126), .ZN(n129) );
  NAND2_X1 U205 ( .A1(n127), .A2(n126), .ZN(n128) );
  NAND2_X1 U206 ( .A1(n129), .A2(n128), .ZN(n130) );
  NAND2_X1 U207 ( .A1(n5), .A2(n130), .ZN(n131) );
  OAI21_X1 U208 ( .B1(n287), .B2(n446), .A(n131), .ZN(n400) );
  NAND2_X1 U209 ( .A1(n133), .A2(n132), .ZN(n134) );
  NAND2_X1 U210 ( .A1(n344), .A2(n134), .ZN(n135) );
  OAI21_X1 U211 ( .B1(n257), .B2(n445), .A(n135), .ZN(n402) );
  NAND2_X1 U212 ( .A1(n137), .A2(n136), .ZN(n138) );
  NAND2_X1 U213 ( .A1(n344), .A2(n138), .ZN(n139) );
  OAI21_X1 U214 ( .B1(n5), .B2(n442), .A(n139), .ZN(n408) );
  NOR2_X1 U215 ( .A1(n141), .A2(n140), .ZN(n142) );
  NAND2_X1 U216 ( .A1(n344), .A2(n142), .ZN(n143) );
  OAI21_X1 U217 ( .B1(n287), .B2(n441), .A(n143), .ZN(n410) );
  NAND2_X1 U218 ( .A1(n145), .A2(n144), .ZN(n146) );
  NAND2_X1 U219 ( .A1(n5), .A2(n146), .ZN(n147) );
  OAI21_X1 U220 ( .B1(n287), .B2(n439), .A(n147), .ZN(n414) );
  FA_X1 U221 ( .A(n150), .B(n149), .CI(n148), .CO(n144), .S(n158) );
  XNOR2_X1 U222 ( .A(n205), .B(\mult_x_1/n286 ), .ZN(n196) );
  OAI22_X1 U223 ( .A1(n207), .A2(n196), .B1(n209), .B2(n151), .ZN(n192) );
  XNOR2_X1 U224 ( .A(n212), .B(\mult_x_1/n284 ), .ZN(n193) );
  OAI22_X1 U225 ( .A1(n213), .A2(n193), .B1(n152), .B2(n460), .ZN(n191) );
  HA_X1 U226 ( .A(n154), .B(n153), .CO(n150), .S(n190) );
  NOR2_X1 U227 ( .A1(n158), .A2(n157), .ZN(n155) );
  NAND2_X1 U228 ( .A1(n257), .A2(n155), .ZN(n156) );
  OAI21_X1 U229 ( .B1(n5), .B2(n438), .A(n156), .ZN(n416) );
  NAND2_X1 U230 ( .A1(n158), .A2(n157), .ZN(n159) );
  NAND2_X1 U231 ( .A1(n257), .A2(n159), .ZN(n160) );
  OAI21_X1 U232 ( .B1(n5), .B2(n437), .A(n160), .ZN(n418) );
  NAND2_X1 U233 ( .A1(n162), .A2(n161), .ZN(n163) );
  NAND2_X1 U234 ( .A1(n287), .A2(n163), .ZN(n164) );
  OAI21_X1 U235 ( .B1(n5), .B2(n435), .A(n164), .ZN(n424) );
  XNOR2_X1 U236 ( .A(n166), .B(n165), .ZN(n167) );
  XNOR2_X1 U237 ( .A(n168), .B(n167), .ZN(n243) );
  XOR2_X1 U238 ( .A(n170), .B(n169), .Z(n171) );
  FA_X1 U239 ( .A(n175), .B(n173), .CI(n174), .CO(n240), .S(n254) );
  INV_X1 U240 ( .A(n238), .ZN(n180) );
  OR2_X1 U241 ( .A1(n178), .A2(n177), .ZN(n237) );
  INV_X1 U242 ( .A(n237), .ZN(n179) );
  NAND2_X1 U243 ( .A1(n180), .A2(n179), .ZN(n181) );
  INV_X1 U244 ( .A(n229), .ZN(n185) );
  NAND2_X1 U245 ( .A1(n230), .A2(n185), .ZN(n188) );
  FA_X1 U246 ( .A(n182), .B(n183), .CI(n184), .CO(n165), .S(n227) );
  NAND2_X1 U247 ( .A1(n230), .A2(n227), .ZN(n187) );
  NAND2_X1 U248 ( .A1(n185), .A2(n227), .ZN(n186) );
  NAND3_X1 U249 ( .A1(n188), .A2(n187), .A3(n186), .ZN(n242) );
  OAI21_X1 U250 ( .B1(n257), .B2(n433), .A(n189), .ZN(n428) );
  FA_X1 U251 ( .A(n192), .B(n191), .CI(n190), .CO(n157), .S(n223) );
  XNOR2_X1 U252 ( .A(n212), .B(\mult_x_1/n285 ), .ZN(n202) );
  OAI22_X1 U253 ( .A1(n213), .A2(n202), .B1(n193), .B2(n460), .ZN(n199) );
  INV_X1 U254 ( .A(n194), .ZN(n195) );
  AND2_X1 U255 ( .A1(\mult_x_1/n288 ), .A2(n195), .ZN(n198) );
  XNOR2_X1 U256 ( .A(n205), .B(\mult_x_1/n287 ), .ZN(n200) );
  OAI22_X1 U257 ( .A1(n207), .A2(n200), .B1(n209), .B2(n196), .ZN(n197) );
  OR2_X1 U258 ( .A1(n223), .A2(n222), .ZN(n296) );
  FA_X1 U259 ( .A(n199), .B(n198), .CI(n197), .CO(n222), .S(n221) );
  XNOR2_X1 U260 ( .A(n205), .B(\mult_x_1/n288 ), .ZN(n201) );
  OAI22_X1 U261 ( .A1(n207), .A2(n201), .B1(n209), .B2(n200), .ZN(n204) );
  XNOR2_X1 U262 ( .A(n212), .B(\mult_x_1/n286 ), .ZN(n208) );
  OAI22_X1 U263 ( .A1(n213), .A2(n208), .B1(n202), .B2(n460), .ZN(n203) );
  NOR2_X1 U264 ( .A1(n221), .A2(n220), .ZN(n288) );
  HA_X1 U265 ( .A(n204), .B(n203), .CO(n220), .S(n218) );
  OR2_X1 U266 ( .A1(\mult_x_1/n288 ), .A2(n457), .ZN(n206) );
  OAI22_X1 U267 ( .A1(n207), .A2(n457), .B1(n206), .B2(n209), .ZN(n217) );
  OR2_X1 U268 ( .A1(n218), .A2(n217), .ZN(n282) );
  XNOR2_X1 U269 ( .A(n212), .B(\mult_x_1/n287 ), .ZN(n211) );
  OAI22_X1 U270 ( .A1(n213), .A2(n211), .B1(n208), .B2(n460), .ZN(n216) );
  INV_X1 U271 ( .A(n209), .ZN(n210) );
  AND2_X1 U272 ( .A1(\mult_x_1/n288 ), .A2(n210), .ZN(n215) );
  NOR2_X1 U273 ( .A1(n216), .A2(n215), .ZN(n274) );
  OAI22_X1 U274 ( .A1(n213), .A2(\mult_x_1/n288 ), .B1(n211), .B2(n460), .ZN(
        n269) );
  OR2_X1 U275 ( .A1(\mult_x_1/n288 ), .A2(n459), .ZN(n214) );
  NAND2_X1 U276 ( .A1(n214), .A2(n213), .ZN(n268) );
  NAND2_X1 U277 ( .A1(n269), .A2(n268), .ZN(n277) );
  NAND2_X1 U278 ( .A1(n216), .A2(n215), .ZN(n275) );
  OAI21_X1 U279 ( .B1(n274), .B2(n277), .A(n275), .ZN(n283) );
  NAND2_X1 U280 ( .A1(n218), .A2(n217), .ZN(n281) );
  INV_X1 U281 ( .A(n281), .ZN(n219) );
  AOI21_X1 U282 ( .B1(n282), .B2(n283), .A(n219), .ZN(n291) );
  NAND2_X1 U283 ( .A1(n221), .A2(n220), .ZN(n289) );
  OAI21_X1 U284 ( .B1(n288), .B2(n291), .A(n289), .ZN(n297) );
  NAND2_X1 U285 ( .A1(n223), .A2(n222), .ZN(n295) );
  INV_X1 U286 ( .A(n295), .ZN(n224) );
  AOI21_X1 U287 ( .B1(n296), .B2(n297), .A(n224), .ZN(n225) );
  NAND2_X1 U288 ( .A1(n5), .A2(n225), .ZN(n226) );
  OAI21_X1 U289 ( .B1(n5), .B2(n432), .A(n226), .ZN(n430) );
  OR2_X1 U290 ( .A1(n344), .A2(n434), .ZN(n241) );
  INV_X1 U291 ( .A(n227), .ZN(n228) );
  XNOR2_X1 U292 ( .A(n228), .B(n229), .ZN(n231) );
  XNOR2_X1 U293 ( .A(n231), .B(n230), .ZN(n247) );
  FA_X1 U294 ( .A(n236), .B(n235), .CI(n234), .CO(n172), .S(n251) );
  XNOR2_X1 U295 ( .A(n240), .B(n239), .ZN(n250) );
  OR2_X1 U296 ( .A1(n344), .A2(n448), .ZN(n245) );
  NAND2_X1 U297 ( .A1(n245), .A2(n244), .ZN(n396) );
  OR2_X1 U298 ( .A1(n344), .A2(n444), .ZN(n249) );
  NAND2_X1 U299 ( .A1(n247), .A2(n246), .ZN(n248) );
  OR2_X1 U300 ( .A1(n344), .A2(n436), .ZN(n259) );
  FA_X1 U301 ( .A(n22), .B(n251), .CI(n250), .CO(n246), .S(n261) );
  NAND2_X1 U302 ( .A1(n259), .A2(n258), .ZN(n420) );
  NAND2_X1 U303 ( .A1(n261), .A2(n260), .ZN(n262) );
  NAND2_X1 U304 ( .A1(n262), .A2(n366), .ZN(n264) );
  NAND2_X1 U305 ( .A1(n326), .A2(n387), .ZN(n263) );
  NAND2_X1 U306 ( .A1(n264), .A2(n263), .ZN(n422) );
  AOI22_X1 U307 ( .A1(n366), .A2(n505), .B1(n506), .B2(n326), .ZN(n508) );
  AOI22_X1 U308 ( .A1(n21), .A2(n504), .B1(n505), .B2(n326), .ZN(n510) );
  AND2_X1 U309 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n266) );
  NAND2_X1 U310 ( .A1(n5), .A2(n266), .ZN(n267) );
  OAI21_X1 U311 ( .B1(n371), .B2(n504), .A(n267), .ZN(n512) );
  AOI22_X1 U312 ( .A1(n5), .A2(n502), .B1(n503), .B2(n326), .ZN(n514) );
  AOI22_X1 U313 ( .A1(n371), .A2(n501), .B1(n502), .B2(n326), .ZN(n516) );
  OR2_X1 U314 ( .A1(n269), .A2(n268), .ZN(n270) );
  AND2_X1 U315 ( .A1(n270), .A2(n277), .ZN(n271) );
  NAND2_X1 U316 ( .A1(n366), .A2(n271), .ZN(n272) );
  OAI21_X1 U317 ( .B1(n371), .B2(n501), .A(n272), .ZN(n518) );
  AOI22_X1 U318 ( .A1(n366), .A2(n499), .B1(n500), .B2(n326), .ZN(n520) );
  AOI22_X1 U319 ( .A1(n21), .A2(n498), .B1(n499), .B2(n326), .ZN(n522) );
  INV_X1 U320 ( .A(n274), .ZN(n276) );
  NAND2_X1 U321 ( .A1(n276), .A2(n275), .ZN(n278) );
  XOR2_X1 U322 ( .A(n278), .B(n277), .Z(n279) );
  NAND2_X1 U323 ( .A1(n21), .A2(n279), .ZN(n280) );
  OAI21_X1 U324 ( .B1(n21), .B2(n498), .A(n280), .ZN(n524) );
  AOI22_X1 U325 ( .A1(n366), .A2(n496), .B1(n497), .B2(n326), .ZN(n526) );
  AOI22_X1 U326 ( .A1(n371), .A2(n495), .B1(n496), .B2(n326), .ZN(n528) );
  NAND2_X1 U327 ( .A1(n282), .A2(n281), .ZN(n284) );
  XNOR2_X1 U328 ( .A(n284), .B(n283), .ZN(n285) );
  NAND2_X1 U329 ( .A1(n21), .A2(n285), .ZN(n286) );
  OAI21_X1 U330 ( .B1(n21), .B2(n495), .A(n286), .ZN(n530) );
  AOI22_X1 U331 ( .A1(n5), .A2(n493), .B1(n494), .B2(n326), .ZN(n532) );
  AOI22_X1 U332 ( .A1(n5), .A2(n492), .B1(n493), .B2(n326), .ZN(n534) );
  INV_X1 U333 ( .A(n288), .ZN(n290) );
  NAND2_X1 U334 ( .A1(n290), .A2(n289), .ZN(n292) );
  XOR2_X1 U335 ( .A(n292), .B(n291), .Z(n293) );
  NAND2_X1 U336 ( .A1(n5), .A2(n293), .ZN(n294) );
  OAI21_X1 U337 ( .B1(n371), .B2(n492), .A(n294), .ZN(n536) );
  AOI22_X1 U338 ( .A1(n366), .A2(n490), .B1(n491), .B2(n326), .ZN(n538) );
  AOI22_X1 U339 ( .A1(n366), .A2(n489), .B1(n490), .B2(n326), .ZN(n540) );
  NAND2_X1 U340 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  NAND2_X1 U342 ( .A1(n371), .A2(n299), .ZN(n300) );
  OAI21_X1 U343 ( .B1(n371), .B2(n489), .A(n300), .ZN(n542) );
  AOI22_X1 U344 ( .A1(n366), .A2(n487), .B1(n488), .B2(n326), .ZN(n544) );
  NAND2_X1 U345 ( .A1(n438), .A2(n385), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(n391), .Z(n302) );
  NAND2_X1 U347 ( .A1(n371), .A2(n302), .ZN(n303) );
  OAI21_X1 U348 ( .B1(n5), .B2(n487), .A(n303), .ZN(n546) );
  AOI22_X1 U349 ( .A1(n21), .A2(n485), .B1(n486), .B2(n326), .ZN(n548) );
  OAI21_X1 U350 ( .B1(n384), .B2(n391), .A(n385), .ZN(n307) );
  NAND2_X1 U351 ( .A1(n375), .A2(n383), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n307), .B(n304), .ZN(n305) );
  NAND2_X1 U353 ( .A1(n287), .A2(n305), .ZN(n306) );
  OAI21_X1 U354 ( .B1(n21), .B2(n485), .A(n306), .ZN(n550) );
  AOI22_X1 U355 ( .A1(n21), .A2(n483), .B1(n484), .B2(n326), .ZN(n552) );
  AOI21_X1 U356 ( .B1(n307), .B2(n375), .A(n439), .ZN(n311) );
  NAND2_X1 U357 ( .A1(n441), .A2(n382), .ZN(n308) );
  XOR2_X1 U358 ( .A(n311), .B(n308), .Z(n309) );
  NAND2_X1 U359 ( .A1(n366), .A2(n309), .ZN(n310) );
  OAI21_X1 U360 ( .B1(n366), .B2(n483), .A(n310), .ZN(n554) );
  AOI22_X1 U361 ( .A1(n21), .A2(n481), .B1(n482), .B2(n326), .ZN(n556) );
  OAI21_X1 U362 ( .B1(n311), .B2(n381), .A(n382), .ZN(n321) );
  INV_X1 U363 ( .A(n321), .ZN(n315) );
  NAND2_X1 U364 ( .A1(n443), .A2(n380), .ZN(n312) );
  XOR2_X1 U365 ( .A(n315), .B(n312), .Z(n313) );
  NAND2_X1 U366 ( .A1(n366), .A2(n313), .ZN(n314) );
  OAI21_X1 U367 ( .B1(n371), .B2(n481), .A(n314), .ZN(n558) );
  AOI22_X1 U368 ( .A1(n371), .A2(n479), .B1(n480), .B2(n326), .ZN(n560) );
  OAI21_X1 U369 ( .B1(n315), .B2(n379), .A(n380), .ZN(n317) );
  NAND2_X1 U370 ( .A1(n436), .A2(n387), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  NAND2_X1 U372 ( .A1(n366), .A2(n318), .ZN(n319) );
  OAI21_X1 U373 ( .B1(n371), .B2(n479), .A(n319), .ZN(n562) );
  AOI22_X1 U374 ( .A1(n5), .A2(n477), .B1(n478), .B2(n326), .ZN(n564) );
  NOR2_X1 U375 ( .A1(n386), .A2(n379), .ZN(n322) );
  OAI21_X1 U376 ( .B1(n386), .B2(n380), .A(n387), .ZN(n320) );
  AOI21_X1 U377 ( .B1(n322), .B2(n321), .A(n320), .ZN(n350) );
  NAND2_X1 U378 ( .A1(n434), .A2(n378), .ZN(n323) );
  XOR2_X1 U379 ( .A(n350), .B(n323), .Z(n324) );
  NAND2_X1 U380 ( .A1(n21), .A2(n324), .ZN(n325) );
  OAI21_X1 U381 ( .B1(n366), .B2(n477), .A(n325), .ZN(n566) );
  AOI22_X1 U382 ( .A1(n21), .A2(n475), .B1(n476), .B2(n326), .ZN(n568) );
  OAI21_X1 U383 ( .B1(n350), .B2(n389), .A(n378), .ZN(n328) );
  NAND2_X1 U384 ( .A1(n374), .A2(n390), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  NAND2_X1 U386 ( .A1(n371), .A2(n329), .ZN(n330) );
  OAI21_X1 U387 ( .B1(n21), .B2(n475), .A(n330), .ZN(n570) );
  AOI22_X1 U388 ( .A1(n21), .A2(n473), .B1(n474), .B2(n326), .ZN(n572) );
  NAND2_X1 U389 ( .A1(n434), .A2(n374), .ZN(n332) );
  AOI21_X1 U390 ( .B1(n444), .B2(n374), .A(n433), .ZN(n331) );
  OAI21_X1 U391 ( .B1(n350), .B2(n332), .A(n331), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n373), .A2(n388), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  NAND2_X1 U394 ( .A1(n21), .A2(n335), .ZN(n336) );
  OAI21_X1 U395 ( .B1(n371), .B2(n473), .A(n336), .ZN(n574) );
  AOI22_X1 U396 ( .A1(n21), .A2(n471), .B1(n472), .B2(n326), .ZN(n576) );
  NAND2_X1 U397 ( .A1(n374), .A2(n373), .ZN(n345) );
  OR2_X1 U398 ( .A1(n389), .A2(n345), .ZN(n339) );
  AOI21_X1 U399 ( .B1(n433), .B2(n373), .A(n435), .ZN(n337) );
  OAI21_X1 U400 ( .B1(n345), .B2(n378), .A(n337), .ZN(n347) );
  INV_X1 U401 ( .A(n347), .ZN(n338) );
  OAI21_X1 U402 ( .B1(n350), .B2(n339), .A(n338), .ZN(n341) );
  NAND2_X1 U403 ( .A1(n372), .A2(n377), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n342) );
  NAND2_X1 U405 ( .A1(n5), .A2(n342), .ZN(n343) );
  OAI21_X1 U406 ( .B1(n371), .B2(n471), .A(n343), .ZN(n578) );
  AOI22_X1 U407 ( .A1(n371), .A2(n469), .B1(n470), .B2(n326), .ZN(n580) );
  NOR2_X1 U408 ( .A1(n345), .A2(n450), .ZN(n346) );
  NAND2_X1 U409 ( .A1(n434), .A2(n346), .ZN(n349) );
  AOI21_X1 U410 ( .B1(n347), .B2(n372), .A(n445), .ZN(n348) );
  OAI21_X1 U411 ( .B1(n350), .B2(n349), .A(n348), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n351), .B(n376), .ZN(n352) );
  NAND2_X1 U413 ( .A1(n366), .A2(n352), .ZN(n353) );
  OAI21_X1 U414 ( .B1(n366), .B2(n469), .A(n353), .ZN(n582) );
  NAND2_X1 U415 ( .A1(n366), .A2(B_extended[0]), .ZN(n354) );
  OAI21_X1 U416 ( .B1(n21), .B2(n468), .A(n354), .ZN(n584) );
  NAND2_X1 U417 ( .A1(n366), .A2(B_extended[1]), .ZN(n355) );
  OAI21_X1 U418 ( .B1(n21), .B2(n467), .A(n355), .ZN(n586) );
  NAND2_X1 U419 ( .A1(n21), .A2(B_extended[2]), .ZN(n356) );
  OAI21_X1 U420 ( .B1(n371), .B2(n466), .A(n356), .ZN(n588) );
  NAND2_X1 U421 ( .A1(n287), .A2(B_extended[3]), .ZN(n357) );
  OAI21_X1 U422 ( .B1(n366), .B2(n465), .A(n357), .ZN(n590) );
  NAND2_X1 U423 ( .A1(n371), .A2(B_extended[4]), .ZN(n358) );
  OAI21_X1 U424 ( .B1(n21), .B2(n464), .A(n358), .ZN(n592) );
  NAND2_X1 U425 ( .A1(n366), .A2(B_extended[5]), .ZN(n359) );
  OAI21_X1 U426 ( .B1(n366), .B2(n463), .A(n359), .ZN(n594) );
  NAND2_X1 U427 ( .A1(n21), .A2(B_extended[6]), .ZN(n360) );
  OAI21_X1 U428 ( .B1(n371), .B2(n462), .A(n360), .ZN(n596) );
  NAND2_X1 U429 ( .A1(n21), .A2(B_extended[7]), .ZN(n361) );
  OAI21_X1 U430 ( .B1(n366), .B2(n461), .A(n361), .ZN(n598) );
  NAND2_X1 U431 ( .A1(n5), .A2(A_extended[0]), .ZN(n362) );
  OAI21_X1 U432 ( .B1(n21), .B2(n460), .A(n362), .ZN(n600) );
  NAND2_X1 U433 ( .A1(n371), .A2(A_extended[1]), .ZN(n363) );
  OAI21_X1 U434 ( .B1(n366), .B2(n459), .A(n363), .ZN(n602) );
  NAND2_X1 U435 ( .A1(n366), .A2(A_extended[2]), .ZN(n364) );
  OAI21_X1 U436 ( .B1(n366), .B2(n458), .A(n364), .ZN(n604) );
  NAND2_X1 U437 ( .A1(n371), .A2(A_extended[3]), .ZN(n365) );
  OAI21_X1 U438 ( .B1(n21), .B2(n457), .A(n365), .ZN(n606) );
  NAND2_X1 U439 ( .A1(n21), .A2(A_extended[4]), .ZN(n367) );
  OAI21_X1 U440 ( .B1(n371), .B2(n456), .A(n367), .ZN(n608) );
  NAND2_X1 U441 ( .A1(n287), .A2(A_extended[5]), .ZN(n368) );
  OAI21_X1 U442 ( .B1(n287), .B2(n455), .A(n368), .ZN(n610) );
  NAND2_X1 U443 ( .A1(n371), .A2(A_extended[6]), .ZN(n369) );
  OAI21_X1 U444 ( .B1(n366), .B2(n454), .A(n369), .ZN(n612) );
  NAND2_X1 U445 ( .A1(n371), .A2(A_extended[7]), .ZN(n370) );
  OAI21_X1 U446 ( .B1(n371), .B2(n453), .A(n370), .ZN(n614) );
  NAND2_X1 U447 ( .A1(n452), .A2(n326), .ZN(n616) );
endmodule


module conv_128_32_DW_mult_pipe_J1_27 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[2] , \mult_x_1/n313 , \mult_x_1/n312 ,
         \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 , \mult_x_1/n286 ,
         \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 , \mult_x_1/n282 ,
         \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n408, n410, n412, n414, n416, n418, n420, n422, n424, n426,
         n428, n430, n432, n434, n436, n438, n440, n442, n444, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n521, n523, n525, n527, n529, n531,
         n533, n535, n537, n539, n541, n543, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n567, n569, n571, n573, n575,
         n577, n579, n581, n583, n585, n587, n589, n591, n593, n595, n597,
         n599, n601, n603, n605, n607, n609, n611, n613, n615, n617, n619,
         n621, n623, n625, n627, n629, n646, n647, n648;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n629), .CK(clk), .Q(n647), 
        .QN(n465) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n625), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n467) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(rst_n), .SE(n623), .CK(clk), .Q(n646), 
        .QN(n468) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(rst_n), .SE(n621), .CK(clk), .Q(n26), 
        .QN(n469) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n464), .SE(n617), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n471) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n464), .SE(n613), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n473) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n464), .SE(n609), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n475) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(rst_n), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n476) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(rst_n), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n477) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n464), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n478) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(rst_n), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n479) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n464), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n480) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n464), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n481) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n464), .SE(n595), .CK(clk), .QN(n482)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n464), .SE(n593), .CK(clk), .Q(
        product[15]), .QN(n483) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n464), .SE(n591), .CK(clk), .QN(n484)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n464), .SE(n589), .CK(clk), .Q(
        product[14]), .QN(n485) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n464), .SE(n587), .CK(clk), .QN(n486)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(rst_n), .SE(n585), .CK(clk), .Q(
        product[13]), .QN(n487) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n464), .SE(n583), .CK(clk), .QN(n488)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(rst_n), .SE(n581), .CK(clk), .Q(
        product[12]), .QN(n489) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n464), .SE(n579), .CK(clk), .QN(n490)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n464), .SE(n577), .CK(clk), .Q(
        product[11]), .QN(n491) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n464), .SE(n575), .CK(clk), .QN(n492)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n464), .SE(n573), .CK(clk), .Q(
        product[10]), .QN(n493) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n464), .SE(n571), .CK(clk), .QN(n494)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n464), .SE(n569), .CK(clk), .Q(
        product[9]), .QN(n495) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n464), .SE(n567), .CK(clk), .QN(n496)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n464), .SE(n565), .CK(clk), .Q(
        product[8]), .QN(n497) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(rst_n), .SE(n563), .CK(clk), .QN(n498) );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(rst_n), .SE(n561), .CK(clk), .Q(
        product[7]), .QN(n499) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(rst_n), .SE(n559), .CK(clk), .QN(n500) );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(rst_n), .SE(n557), .CK(clk), .Q(
        product[6]), .QN(n501) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(rst_n), .SE(n555), .CK(clk), .QN(n502) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(rst_n), .SE(n553), .CK(clk), .QN(n503) );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(rst_n), .SE(n551), .CK(clk), .Q(
        product[5]), .QN(n504) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(rst_n), .SE(n549), .CK(clk), .QN(n505) );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(rst_n), .SE(n547), .CK(clk), .QN(n506) );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(rst_n), .SE(n545), .CK(clk), .Q(
        product[4]), .QN(n507) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(rst_n), .SE(n543), .CK(clk), .QN(n508) );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(rst_n), .SE(n541), .CK(clk), .QN(n509) );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(rst_n), .SE(n539), .CK(clk), .Q(
        product[3]), .QN(n510) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(rst_n), .SE(n537), .CK(clk), .QN(n511) );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(rst_n), .SE(n535), .CK(clk), .QN(n512) );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(rst_n), .SE(n533), .CK(clk), .Q(
        product[2]), .QN(n513) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(rst_n), .SE(n531), .CK(clk), .QN(n514) );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(rst_n), .SE(n529), .CK(clk), .QN(n515) );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(rst_n), .SE(n527), .CK(clk), .Q(
        product[1]), .QN(n516) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(rst_n), .SE(n525), .CK(clk), .QN(n517) );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(rst_n), .SE(n523), .CK(clk), .QN(n518) );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(rst_n), .SE(n521), .CK(clk), .Q(
        product[0]), .QN(n519) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(rst_n), .SE(n615), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n472) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n648), .SI(1'b1), .SE(n444), .CK(clk), 
        .Q(n405), .QN(n446) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n648), .SI(1'b1), .SE(n442), .CK(clk), 
        .Q(n404), .QN(n447) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n648), .SI(1'b1), .SE(n440), .CK(clk), 
        .Q(n403), .QN(n448) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n648), .SE(n438), .CK(
        clk), .QN(n402) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n648), .SE(n436), .CK(
        clk), .Q(n449), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n648), .SI(1'b1), .SE(n434), .CK(clk), 
        .Q(n400), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n648), .SI(1'b1), .SE(n432), .CK(clk), 
        .Q(n399), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n648), .SI(1'b1), .SE(n430), .CK(clk), 
        .Q(n398), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n648), .SI(1'b1), .SE(n428), .CK(clk), 
        .Q(n397), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n648), .SI(1'b1), .SE(n426), .CK(clk), 
        .Q(n396), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n648), .SI(1'b1), .SE(n424), .CK(clk), 
        .Q(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n648), .SI(1'b1), .SE(n420), .CK(clk), 
        .Q(n393), .QN(n456) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n648), .SE(n418), .CK(
        clk), .Q(n457), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n648), .SI(1'b1), .SE(n416), .CK(clk), 
        .Q(n391), .QN(n458) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n648), .SE(n414), .CK(
        clk), .Q(n459), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n648), .SE(n412), .CK(
        clk), .Q(n460), .QN(n389) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n648), .SI(1'b1), .SE(n410), .CK(clk), 
        .Q(n388), .QN(n461) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n648), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n648), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n386), .QN(n463) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n464), .SE(n619), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n470) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n648), .SI(1'b1), .SE(n422), .CK(clk), 
        .Q(n394), .QN(n455) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n464), .SE(n627), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n466) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n464), .SE(n611), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n474) );
  INV_X1 U2 ( .A(en), .ZN(n290) );
  INV_X1 U3 ( .A(n648), .ZN(n464) );
  INV_X2 U4 ( .A(rst_n), .ZN(n648) );
  CLKBUF_X2 U5 ( .A(n646), .Z(n167) );
  BUF_X1 U6 ( .A(\mult_x_1/n313 ), .Z(n261) );
  XNOR2_X1 U7 ( .A(n8), .B(n82), .ZN(n117) );
  XNOR2_X1 U8 ( .A(n62), .B(n16), .ZN(n100) );
  XNOR2_X1 U9 ( .A(n12), .B(n11), .ZN(n115) );
  XNOR2_X1 U10 ( .A(n83), .B(n84), .ZN(n8) );
  XNOR2_X1 U11 ( .A(n64), .B(n63), .ZN(n16) );
  XNOR2_X1 U12 ( .A(n90), .B(n91), .ZN(n12) );
  OR2_X1 U13 ( .A1(n64), .A2(n63), .ZN(n15) );
  NAND2_X1 U14 ( .A1(n64), .A2(n63), .ZN(n13) );
  NAND2_X1 U15 ( .A1(n22), .A2(n43), .ZN(n171) );
  NAND2_X1 U16 ( .A1(n30), .A2(n31), .ZN(n181) );
  AND2_X1 U17 ( .A1(n647), .A2(\mult_x_1/n281 ), .ZN(n136) );
  NOR2_X1 U18 ( .A1(n465), .A2(n466), .ZN(n33) );
  NAND2_X1 U19 ( .A1(n5), .A2(n237), .ZN(n211) );
  NAND2_X1 U20 ( .A1(n210), .A2(n209), .ZN(n5) );
  NAND2_X1 U21 ( .A1(n7), .A2(n6), .ZN(n106) );
  NAND2_X1 U22 ( .A1(n83), .A2(n84), .ZN(n6) );
  OAI21_X1 U23 ( .B1(n83), .B2(n84), .A(n82), .ZN(n7) );
  NAND2_X1 U24 ( .A1(n10), .A2(n9), .ZN(n81) );
  NAND2_X1 U25 ( .A1(n91), .A2(n90), .ZN(n9) );
  OAI21_X1 U26 ( .B1(n90), .B2(n91), .A(n11), .ZN(n10) );
  NOR2_X1 U27 ( .A1(n49), .A2(n185), .ZN(n11) );
  NAND2_X1 U28 ( .A1(n14), .A2(n13), .ZN(n152) );
  NAND2_X1 U29 ( .A1(n62), .A2(n15), .ZN(n14) );
  XNOR2_X1 U30 ( .A(n470), .B(n469), .ZN(n22) );
  NAND2_X1 U31 ( .A1(n20), .A2(n17), .ZN(n408) );
  NAND2_X1 U32 ( .A1(n155), .A2(n237), .ZN(n17) );
  NAND2_X1 U33 ( .A1(n19), .A2(n18), .ZN(n144) );
  NAND2_X1 U34 ( .A1(n171), .A2(n244), .ZN(n18) );
  INV_X1 U35 ( .A(n139), .ZN(n19) );
  INV_X1 U36 ( .A(n78), .ZN(n54) );
  INV_X1 U37 ( .A(n79), .ZN(n55) );
  BUF_X1 U38 ( .A(\mult_x_1/n310 ), .Z(n27) );
  INV_X1 U39 ( .A(n239), .ZN(n223) );
  INV_X1 U40 ( .A(n240), .ZN(n224) );
  XNOR2_X1 U41 ( .A(n242), .B(n241), .ZN(n272) );
  XNOR2_X1 U42 ( .A(n240), .B(n239), .ZN(n241) );
  NAND2_X1 U43 ( .A1(n227), .A2(n226), .ZN(n230) );
  NAND2_X1 U44 ( .A1(n240), .A2(n239), .ZN(n226) );
  NAND2_X1 U45 ( .A1(n242), .A2(n225), .ZN(n227) );
  NAND2_X1 U46 ( .A1(n224), .A2(n223), .ZN(n225) );
  NAND2_X1 U47 ( .A1(n94), .A2(n93), .ZN(n109) );
  NAND2_X1 U48 ( .A1(n117), .A2(n92), .ZN(n94) );
  NAND2_X1 U49 ( .A1(n58), .A2(n57), .ZN(n102) );
  NAND2_X1 U50 ( .A1(n79), .A2(n78), .ZN(n57) );
  XNOR2_X1 U51 ( .A(n117), .B(n116), .ZN(n134) );
  NAND2_X1 U52 ( .A1(n128), .A2(n387), .ZN(n20) );
  OAI22_X1 U53 ( .A1(n134), .A2(n133), .B1(n279), .B2(n455), .ZN(n422) );
  NAND2_X1 U54 ( .A1(n132), .A2(n276), .ZN(n133) );
  INV_X1 U55 ( .A(n131), .ZN(n132) );
  INV_X1 U56 ( .A(n75), .ZN(n21) );
  XNOR2_X1 U57 ( .A(n468), .B(n26), .ZN(n43) );
  NAND2_X1 U58 ( .A1(n37), .A2(n36), .ZN(n23) );
  NAND2_X1 U59 ( .A1(n37), .A2(n36), .ZN(n24) );
  NAND2_X1 U60 ( .A1(n37), .A2(n36), .ZN(n257) );
  NAND2_X1 U61 ( .A1(n115), .A2(n114), .ZN(n93) );
  XNOR2_X1 U62 ( .A(n115), .B(n114), .ZN(n116) );
  OR2_X1 U63 ( .A1(n114), .A2(n115), .ZN(n92) );
  XNOR2_X1 U64 ( .A(n52), .B(n33), .ZN(n185) );
  OAI22_X1 U65 ( .A1(n171), .A2(n85), .B1(n244), .B2(n50), .ZN(n25) );
  XNOR2_X1 U66 ( .A(n26), .B(n470), .ZN(n42) );
  INV_X1 U67 ( .A(n38), .ZN(n259) );
  INV_X1 U68 ( .A(n38), .ZN(n37) );
  INV_X2 U69 ( .A(n290), .ZN(n380) );
  BUF_X2 U70 ( .A(en), .Z(n276) );
  INV_X2 U71 ( .A(n290), .ZN(n385) );
  INV_X2 U72 ( .A(n42), .ZN(n244) );
  XNOR2_X1 U73 ( .A(n136), .B(n167), .ZN(n139) );
  XNOR2_X1 U74 ( .A(n167), .B(\mult_x_1/n281 ), .ZN(n44) );
  INV_X1 U75 ( .A(n44), .ZN(n28) );
  NAND3_X1 U76 ( .A1(n244), .A2(n43), .A3(n28), .ZN(n29) );
  OAI21_X1 U77 ( .B1(n244), .B2(n139), .A(n29), .ZN(n145) );
  INV_X1 U78 ( .A(n145), .ZN(n142) );
  XOR2_X1 U79 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .Z(n30) );
  XNOR2_X1 U80 ( .A(\mult_x_1/a[6] ), .B(n646), .ZN(n31) );
  XNOR2_X1 U81 ( .A(n27), .B(\mult_x_1/n283 ), .ZN(n35) );
  INV_X1 U82 ( .A(n31), .ZN(n32) );
  INV_X2 U83 ( .A(n32), .ZN(n182) );
  XNOR2_X1 U84 ( .A(n27), .B(\mult_x_1/n282 ), .ZN(n138) );
  OAI22_X1 U85 ( .A1(n181), .A2(n35), .B1(n182), .B2(n138), .ZN(n141) );
  BUF_X2 U86 ( .A(n33), .Z(n184) );
  XNOR2_X1 U87 ( .A(n184), .B(\mult_x_1/n284 ), .ZN(n34) );
  INV_X1 U88 ( .A(n466), .ZN(n52) );
  NOR2_X1 U89 ( .A1(n34), .A2(n185), .ZN(n140) );
  XNOR2_X1 U90 ( .A(n27), .B(\mult_x_1/n284 ), .ZN(n46) );
  OAI22_X1 U91 ( .A1(n181), .A2(n46), .B1(n182), .B2(n35), .ZN(n61) );
  XOR2_X1 U92 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .Z(n38) );
  XNOR2_X1 U93 ( .A(\mult_x_1/n312 ), .B(n471), .ZN(n36) );
  XNOR2_X1 U94 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n51) );
  XNOR2_X1 U95 ( .A(n136), .B(\mult_x_1/n312 ), .ZN(n39) );
  OAI22_X1 U96 ( .A1(n257), .A2(n51), .B1(n39), .B2(n259), .ZN(n60) );
  AOI21_X1 U97 ( .B1(n259), .B2(n23), .A(n39), .ZN(n40) );
  INV_X1 U98 ( .A(n40), .ZN(n59) );
  XNOR2_X1 U99 ( .A(n184), .B(\mult_x_1/n285 ), .ZN(n41) );
  NOR2_X1 U100 ( .A1(n41), .A2(n185), .ZN(n64) );
  XNOR2_X1 U101 ( .A(n167), .B(\mult_x_1/n282 ), .ZN(n45) );
  OAI22_X1 U102 ( .A1(n171), .A2(n45), .B1(n244), .B2(n44), .ZN(n63) );
  XNOR2_X1 U103 ( .A(n167), .B(\mult_x_1/n283 ), .ZN(n50) );
  OAI22_X1 U104 ( .A1(n171), .A2(n50), .B1(n244), .B2(n45), .ZN(n77) );
  XNOR2_X1 U105 ( .A(n27), .B(\mult_x_1/n285 ), .ZN(n48) );
  OAI22_X1 U106 ( .A1(n181), .A2(n48), .B1(n182), .B2(n46), .ZN(n76) );
  INV_X1 U107 ( .A(n60), .ZN(n75) );
  NAND2_X1 U108 ( .A1(n261), .A2(n473), .ZN(n262) );
  XNOR2_X1 U109 ( .A(n136), .B(n261), .ZN(n73) );
  AOI21_X1 U110 ( .B1(n262), .B2(n473), .A(n73), .ZN(n47) );
  INV_X1 U111 ( .A(n47), .ZN(n91) );
  XNOR2_X1 U112 ( .A(n27), .B(\mult_x_1/n286 ), .ZN(n72) );
  OAI22_X1 U113 ( .A1(n181), .A2(n72), .B1(n182), .B2(n48), .ZN(n90) );
  XNOR2_X1 U114 ( .A(n184), .B(\mult_x_1/n287 ), .ZN(n49) );
  XNOR2_X1 U115 ( .A(n167), .B(\mult_x_1/n284 ), .ZN(n85) );
  OAI22_X1 U116 ( .A1(n171), .A2(n85), .B1(n244), .B2(n50), .ZN(n69) );
  XNOR2_X1 U117 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n86) );
  OAI22_X1 U118 ( .A1(n24), .A2(n86), .B1(n259), .B2(n51), .ZN(n68) );
  OR2_X1 U119 ( .A1(n25), .A2(n68), .ZN(n79) );
  XNOR2_X1 U120 ( .A(n184), .B(\mult_x_1/n286 ), .ZN(n53) );
  XNOR2_X1 U121 ( .A(n52), .B(n33), .ZN(n74) );
  NOR2_X1 U122 ( .A1(n53), .A2(n74), .ZN(n78) );
  NAND2_X1 U123 ( .A1(n55), .A2(n54), .ZN(n56) );
  NAND2_X1 U124 ( .A1(n81), .A2(n56), .ZN(n58) );
  FA_X1 U125 ( .A(n61), .B(n21), .CI(n59), .CO(n153), .S(n101) );
  NAND2_X1 U126 ( .A1(n157), .A2(n156), .ZN(n65) );
  BUF_X2 U127 ( .A(en), .Z(n279) );
  NAND2_X1 U128 ( .A1(n65), .A2(n237), .ZN(n67) );
  BUF_X2 U129 ( .A(en), .Z(n237) );
  NAND2_X1 U130 ( .A1(n97), .A2(n403), .ZN(n66) );
  NAND2_X1 U131 ( .A1(n67), .A2(n66), .ZN(n440) );
  XNOR2_X1 U132 ( .A(n69), .B(n68), .ZN(n84) );
  INV_X1 U133 ( .A(n184), .ZN(n70) );
  OR2_X1 U134 ( .A1(\mult_x_1/n288 ), .A2(n70), .ZN(n71) );
  NOR2_X1 U135 ( .A1(n71), .A2(n185), .ZN(n83) );
  XNOR2_X1 U136 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n88) );
  OAI22_X1 U137 ( .A1(n181), .A2(n88), .B1(n182), .B2(n72), .ZN(n120) );
  XNOR2_X1 U138 ( .A(n261), .B(\mult_x_1/n281 ), .ZN(n122) );
  OAI22_X1 U139 ( .A1(n262), .A2(n122), .B1(n73), .B2(n473), .ZN(n119) );
  NOR2_X1 U140 ( .A1(n74), .A2(n481), .ZN(n118) );
  FA_X1 U141 ( .A(n77), .B(n76), .CI(n75), .CO(n62), .S(n105) );
  XNOR2_X1 U142 ( .A(n79), .B(n78), .ZN(n80) );
  XNOR2_X1 U143 ( .A(n81), .B(n80), .ZN(n104) );
  INV_X1 U144 ( .A(n110), .ZN(n96) );
  XNOR2_X1 U145 ( .A(n167), .B(\mult_x_1/n285 ), .ZN(n121) );
  OAI22_X1 U146 ( .A1(n171), .A2(n121), .B1(n244), .B2(n85), .ZN(n126) );
  INV_X1 U147 ( .A(n470), .ZN(n255) );
  XNOR2_X1 U148 ( .A(n255), .B(\mult_x_1/n283 ), .ZN(n123) );
  OAI22_X1 U149 ( .A1(n24), .A2(n123), .B1(n259), .B2(n86), .ZN(n125) );
  OR2_X1 U150 ( .A1(\mult_x_1/n288 ), .A2(n466), .ZN(n87) );
  OAI22_X1 U151 ( .A1(n181), .A2(n466), .B1(n87), .B2(n182), .ZN(n162) );
  XNOR2_X1 U152 ( .A(n27), .B(\mult_x_1/n288 ), .ZN(n89) );
  OAI22_X1 U153 ( .A1(n181), .A2(n89), .B1(n182), .B2(n88), .ZN(n161) );
  NOR2_X1 U154 ( .A1(n109), .A2(n290), .ZN(n95) );
  NAND2_X1 U155 ( .A1(n96), .A2(n95), .ZN(n99) );
  INV_X1 U156 ( .A(n276), .ZN(n97) );
  NAND2_X1 U157 ( .A1(n97), .A2(n401), .ZN(n98) );
  NAND2_X1 U158 ( .A1(n99), .A2(n98), .ZN(n436) );
  FA_X1 U159 ( .A(n102), .B(n101), .CI(n100), .CO(n156), .S(n282) );
  INV_X1 U160 ( .A(n276), .ZN(n103) );
  NAND2_X1 U161 ( .A1(n103), .A2(n393), .ZN(n108) );
  FA_X1 U162 ( .A(n106), .B(n105), .CI(n104), .CO(n277), .S(n110) );
  NAND2_X1 U163 ( .A1(n278), .A2(n279), .ZN(n107) );
  OAI211_X1 U164 ( .C1(n282), .C2(n97), .A(n108), .B(n107), .ZN(n420) );
  NAND2_X1 U165 ( .A1(n110), .A2(n109), .ZN(n111) );
  NAND2_X1 U166 ( .A1(n111), .A2(n237), .ZN(n113) );
  NAND2_X1 U167 ( .A1(n128), .A2(n402), .ZN(n112) );
  NAND2_X1 U168 ( .A1(n113), .A2(n112), .ZN(n438) );
  FA_X1 U169 ( .A(n118), .B(n119), .CI(n120), .CO(n82), .S(n203) );
  XNOR2_X1 U170 ( .A(n167), .B(\mult_x_1/n286 ), .ZN(n169) );
  OAI22_X1 U171 ( .A1(n171), .A2(n169), .B1(n244), .B2(n121), .ZN(n165) );
  XNOR2_X1 U172 ( .A(n261), .B(\mult_x_1/n282 ), .ZN(n159) );
  OAI22_X1 U173 ( .A1(n262), .A2(n159), .B1(n122), .B2(n473), .ZN(n164) );
  XNOR2_X1 U174 ( .A(n255), .B(\mult_x_1/n284 ), .ZN(n160) );
  OAI22_X1 U175 ( .A1(n23), .A2(n160), .B1(n259), .B2(n123), .ZN(n163) );
  FA_X1 U176 ( .A(n126), .B(n125), .CI(n124), .CO(n114), .S(n201) );
  NAND2_X1 U177 ( .A1(n134), .A2(n131), .ZN(n127) );
  NAND2_X1 U178 ( .A1(n127), .A2(n237), .ZN(n130) );
  INV_X1 U179 ( .A(n276), .ZN(n128) );
  NAND2_X1 U180 ( .A1(n128), .A2(n395), .ZN(n129) );
  NAND2_X1 U181 ( .A1(n130), .A2(n129), .ZN(n424) );
  XNOR2_X1 U202 ( .A(n184), .B(\mult_x_1/n282 ), .ZN(n135) );
  NOR2_X1 U203 ( .A1(n135), .A2(n185), .ZN(n179) );
  XNOR2_X1 U204 ( .A(n27), .B(\mult_x_1/n281 ), .ZN(n137) );
  XNOR2_X1 U205 ( .A(n136), .B(n27), .ZN(n180) );
  OAI22_X1 U206 ( .A1(n181), .A2(n137), .B1(n180), .B2(n182), .ZN(n190) );
  INV_X1 U207 ( .A(n190), .ZN(n178) );
  OAI22_X1 U208 ( .A1(n181), .A2(n138), .B1(n182), .B2(n137), .ZN(n146) );
  FA_X1 U209 ( .A(n140), .B(n141), .CI(n142), .CO(n151), .S(n154) );
  XNOR2_X1 U210 ( .A(n184), .B(\mult_x_1/n283 ), .ZN(n143) );
  NOR2_X1 U211 ( .A1(n143), .A2(n185), .ZN(n150) );
  FA_X1 U212 ( .A(n146), .B(n144), .CI(n145), .CO(n177), .S(n149) );
  OR2_X1 U213 ( .A1(n198), .A2(n197), .ZN(n147) );
  NAND2_X1 U214 ( .A1(n237), .A2(n147), .ZN(n148) );
  OAI21_X1 U215 ( .B1(n237), .B2(n463), .A(n148), .ZN(n406) );
  FA_X1 U216 ( .A(n151), .B(n150), .CI(n149), .CO(n197), .S(n235) );
  FA_X1 U217 ( .A(n154), .B(n153), .CI(n152), .CO(n234), .S(n157) );
  OR2_X1 U218 ( .A1(n235), .A2(n234), .ZN(n155) );
  OAI21_X1 U219 ( .B1(n157), .B2(n156), .A(n237), .ZN(n158) );
  OAI21_X1 U220 ( .B1(n279), .B2(n461), .A(n158), .ZN(n410) );
  XNOR2_X1 U221 ( .A(n261), .B(\mult_x_1/n283 ), .ZN(n222) );
  OAI22_X1 U222 ( .A1(n262), .A2(n222), .B1(n159), .B2(n473), .ZN(n174) );
  AND2_X1 U223 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n173) );
  XNOR2_X1 U224 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n221) );
  OAI22_X1 U225 ( .A1(n24), .A2(n221), .B1(n259), .B2(n160), .ZN(n172) );
  HA_X1 U226 ( .A(n162), .B(n161), .CO(n124), .S(n205) );
  FA_X1 U227 ( .A(n165), .B(n164), .CI(n163), .CO(n202), .S(n204) );
  OR2_X1 U228 ( .A1(\mult_x_1/n288 ), .A2(n468), .ZN(n166) );
  OAI22_X1 U229 ( .A1(n171), .A2(n468), .B1(n166), .B2(n244), .ZN(n220) );
  XNOR2_X1 U230 ( .A(n167), .B(\mult_x_1/n288 ), .ZN(n168) );
  XNOR2_X1 U231 ( .A(n167), .B(\mult_x_1/n287 ), .ZN(n170) );
  OAI22_X1 U232 ( .A1(n171), .A2(n168), .B1(n244), .B2(n170), .ZN(n219) );
  OAI22_X1 U233 ( .A1(n171), .A2(n170), .B1(n244), .B2(n169), .ZN(n217) );
  FA_X1 U234 ( .A(n174), .B(n173), .CI(n172), .CO(n206), .S(n216) );
  OR2_X1 U235 ( .A1(n213), .A2(n212), .ZN(n175) );
  NAND2_X1 U236 ( .A1(n237), .A2(n175), .ZN(n176) );
  OAI21_X1 U237 ( .B1(n279), .B2(n460), .A(n176), .ZN(n412) );
  FA_X1 U238 ( .A(n179), .B(n178), .CI(n177), .CO(n192), .S(n198) );
  AOI21_X1 U239 ( .B1(n182), .B2(n181), .A(n180), .ZN(n183) );
  INV_X1 U240 ( .A(n183), .ZN(n188) );
  XNOR2_X1 U241 ( .A(n184), .B(\mult_x_1/n281 ), .ZN(n186) );
  NOR2_X1 U242 ( .A1(n186), .A2(n185), .ZN(n187) );
  XOR2_X1 U243 ( .A(n188), .B(n187), .Z(n189) );
  XOR2_X1 U244 ( .A(n190), .B(n189), .Z(n191) );
  OR2_X1 U245 ( .A1(n192), .A2(n191), .ZN(n194) );
  NAND2_X1 U246 ( .A1(n192), .A2(n191), .ZN(n193) );
  NAND2_X1 U247 ( .A1(n194), .A2(n193), .ZN(n195) );
  NAND2_X1 U248 ( .A1(n279), .A2(n195), .ZN(n196) );
  OAI21_X1 U249 ( .B1(n279), .B2(n459), .A(n196), .ZN(n414) );
  NAND2_X1 U250 ( .A1(n198), .A2(n197), .ZN(n199) );
  NAND2_X1 U251 ( .A1(n237), .A2(n199), .ZN(n200) );
  OAI21_X1 U252 ( .B1(n237), .B2(n458), .A(n200), .ZN(n416) );
  FA_X1 U253 ( .A(n203), .B(n202), .CI(n201), .CO(n131), .S(n210) );
  FA_X1 U254 ( .A(n206), .B(n205), .CI(n204), .CO(n209), .S(n213) );
  NOR2_X1 U255 ( .A1(n210), .A2(n209), .ZN(n207) );
  NAND2_X1 U256 ( .A1(n237), .A2(n207), .ZN(n208) );
  OAI21_X1 U257 ( .B1(n237), .B2(n454), .A(n208), .ZN(n426) );
  OAI21_X1 U258 ( .B1(n237), .B2(n453), .A(n211), .ZN(n428) );
  NAND2_X1 U259 ( .A1(n213), .A2(n212), .ZN(n214) );
  NAND2_X1 U260 ( .A1(n279), .A2(n214), .ZN(n215) );
  OAI21_X1 U261 ( .B1(n279), .B2(n452), .A(n215), .ZN(n430) );
  FA_X1 U262 ( .A(n218), .B(n217), .CI(n216), .CO(n212), .S(n231) );
  HA_X1 U263 ( .A(n220), .B(n219), .CO(n218), .S(n242) );
  XNOR2_X1 U264 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n246) );
  OAI22_X1 U265 ( .A1(n23), .A2(n246), .B1(n259), .B2(n221), .ZN(n240) );
  XNOR2_X1 U266 ( .A(n261), .B(\mult_x_1/n284 ), .ZN(n243) );
  OAI22_X1 U267 ( .A1(n262), .A2(n243), .B1(n222), .B2(n473), .ZN(n239) );
  NOR2_X1 U268 ( .A1(n231), .A2(n230), .ZN(n228) );
  NAND2_X1 U269 ( .A1(n279), .A2(n228), .ZN(n229) );
  OAI21_X1 U270 ( .B1(n237), .B2(n451), .A(n229), .ZN(n432) );
  NAND2_X1 U271 ( .A1(n231), .A2(n230), .ZN(n232) );
  NAND2_X1 U272 ( .A1(n237), .A2(n232), .ZN(n233) );
  OAI21_X1 U273 ( .B1(n237), .B2(n450), .A(n233), .ZN(n434) );
  NAND2_X1 U274 ( .A1(n235), .A2(n234), .ZN(n236) );
  NAND2_X1 U275 ( .A1(n279), .A2(n236), .ZN(n238) );
  OAI21_X1 U276 ( .B1(n279), .B2(n447), .A(n238), .ZN(n442) );
  XNOR2_X1 U277 ( .A(n261), .B(\mult_x_1/n285 ), .ZN(n252) );
  OAI22_X1 U278 ( .A1(n262), .A2(n252), .B1(n243), .B2(n473), .ZN(n249) );
  INV_X1 U279 ( .A(n244), .ZN(n245) );
  AND2_X1 U280 ( .A1(\mult_x_1/n288 ), .A2(n245), .ZN(n248) );
  XNOR2_X1 U281 ( .A(n255), .B(\mult_x_1/n287 ), .ZN(n250) );
  OAI22_X1 U282 ( .A1(n23), .A2(n250), .B1(n259), .B2(n246), .ZN(n247) );
  OR2_X1 U283 ( .A1(n272), .A2(n271), .ZN(n312) );
  FA_X1 U284 ( .A(n249), .B(n248), .CI(n247), .CO(n271), .S(n270) );
  XNOR2_X1 U285 ( .A(n255), .B(\mult_x_1/n288 ), .ZN(n251) );
  OAI22_X1 U286 ( .A1(n24), .A2(n251), .B1(n259), .B2(n250), .ZN(n254) );
  XNOR2_X1 U287 ( .A(n261), .B(\mult_x_1/n286 ), .ZN(n258) );
  OAI22_X1 U288 ( .A1(n262), .A2(n258), .B1(n252), .B2(n473), .ZN(n253) );
  NOR2_X1 U289 ( .A1(n270), .A2(n269), .ZN(n304) );
  HA_X1 U290 ( .A(n254), .B(n253), .CO(n269), .S(n267) );
  OR2_X1 U291 ( .A1(\mult_x_1/n288 ), .A2(n470), .ZN(n256) );
  OAI22_X1 U292 ( .A1(n24), .A2(n470), .B1(n256), .B2(n259), .ZN(n266) );
  OR2_X1 U293 ( .A1(n267), .A2(n266), .ZN(n299) );
  XNOR2_X1 U294 ( .A(n261), .B(\mult_x_1/n287 ), .ZN(n260) );
  OAI22_X1 U295 ( .A1(n262), .A2(n260), .B1(n258), .B2(n473), .ZN(n265) );
  AND2_X1 U296 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n264) );
  NOR2_X1 U297 ( .A1(n265), .A2(n264), .ZN(n291) );
  OAI22_X1 U298 ( .A1(n262), .A2(\mult_x_1/n288 ), .B1(n260), .B2(n473), .ZN(
        n286) );
  OR2_X1 U299 ( .A1(\mult_x_1/n288 ), .A2(n472), .ZN(n263) );
  NAND2_X1 U300 ( .A1(n263), .A2(n262), .ZN(n285) );
  NAND2_X1 U301 ( .A1(n286), .A2(n285), .ZN(n294) );
  NAND2_X1 U302 ( .A1(n265), .A2(n264), .ZN(n292) );
  OAI21_X1 U303 ( .B1(n291), .B2(n294), .A(n292), .ZN(n300) );
  NAND2_X1 U304 ( .A1(n267), .A2(n266), .ZN(n298) );
  INV_X1 U305 ( .A(n298), .ZN(n268) );
  AOI21_X1 U306 ( .B1(n299), .B2(n300), .A(n268), .ZN(n307) );
  NAND2_X1 U307 ( .A1(n270), .A2(n269), .ZN(n305) );
  OAI21_X1 U308 ( .B1(n304), .B2(n307), .A(n305), .ZN(n313) );
  NAND2_X1 U309 ( .A1(n272), .A2(n271), .ZN(n311) );
  INV_X1 U310 ( .A(n311), .ZN(n273) );
  AOI21_X1 U311 ( .B1(n312), .B2(n313), .A(n273), .ZN(n274) );
  NAND2_X1 U312 ( .A1(n237), .A2(n274), .ZN(n275) );
  OAI21_X1 U313 ( .B1(n279), .B2(n446), .A(n275), .ZN(n444) );
  INV_X1 U314 ( .A(n277), .ZN(n278) );
  NAND2_X1 U315 ( .A1(n278), .A2(n237), .ZN(n281) );
  OR2_X1 U316 ( .A1(n279), .A2(n457), .ZN(n280) );
  OAI21_X1 U317 ( .B1(n282), .B2(n281), .A(n280), .ZN(n418) );
  AOI22_X1 U318 ( .A1(n385), .A2(n518), .B1(n519), .B2(n128), .ZN(n521) );
  AOI22_X1 U319 ( .A1(n385), .A2(n517), .B1(n518), .B2(n97), .ZN(n523) );
  AND2_X1 U320 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n283) );
  NAND2_X1 U321 ( .A1(n237), .A2(n283), .ZN(n284) );
  OAI21_X1 U322 ( .B1(n385), .B2(n517), .A(n284), .ZN(n525) );
  AOI22_X1 U323 ( .A1(n380), .A2(n515), .B1(n516), .B2(n97), .ZN(n527) );
  AOI22_X1 U324 ( .A1(n380), .A2(n514), .B1(n515), .B2(n97), .ZN(n529) );
  OR2_X1 U325 ( .A1(n286), .A2(n285), .ZN(n287) );
  AND2_X1 U326 ( .A1(n287), .A2(n294), .ZN(n288) );
  NAND2_X1 U327 ( .A1(n279), .A2(n288), .ZN(n289) );
  OAI21_X1 U328 ( .B1(n385), .B2(n514), .A(n289), .ZN(n531) );
  AOI22_X1 U329 ( .A1(n385), .A2(n512), .B1(n513), .B2(n97), .ZN(n533) );
  AOI22_X1 U330 ( .A1(n385), .A2(n511), .B1(n512), .B2(n103), .ZN(n535) );
  INV_X1 U331 ( .A(n291), .ZN(n293) );
  NAND2_X1 U332 ( .A1(n293), .A2(n292), .ZN(n295) );
  XOR2_X1 U333 ( .A(n295), .B(n294), .Z(n296) );
  NAND2_X1 U334 ( .A1(n276), .A2(n296), .ZN(n297) );
  OAI21_X1 U335 ( .B1(n380), .B2(n511), .A(n297), .ZN(n537) );
  AOI22_X1 U336 ( .A1(n380), .A2(n509), .B1(n510), .B2(n128), .ZN(n539) );
  AOI22_X1 U337 ( .A1(n237), .A2(n508), .B1(n509), .B2(n128), .ZN(n541) );
  NAND2_X1 U338 ( .A1(n299), .A2(n298), .ZN(n301) );
  XNOR2_X1 U339 ( .A(n301), .B(n300), .ZN(n302) );
  NAND2_X1 U340 ( .A1(n279), .A2(n302), .ZN(n303) );
  OAI21_X1 U341 ( .B1(n380), .B2(n508), .A(n303), .ZN(n543) );
  AOI22_X1 U342 ( .A1(n385), .A2(n506), .B1(n507), .B2(n103), .ZN(n545) );
  AOI22_X1 U343 ( .A1(n380), .A2(n505), .B1(n506), .B2(n103), .ZN(n547) );
  INV_X1 U344 ( .A(n304), .ZN(n306) );
  NAND2_X1 U345 ( .A1(n306), .A2(n305), .ZN(n308) );
  XOR2_X1 U346 ( .A(n308), .B(n307), .Z(n309) );
  NAND2_X1 U347 ( .A1(n279), .A2(n309), .ZN(n310) );
  OAI21_X1 U348 ( .B1(n385), .B2(n505), .A(n310), .ZN(n549) );
  AOI22_X1 U349 ( .A1(n385), .A2(n503), .B1(n504), .B2(n128), .ZN(n551) );
  AOI22_X1 U350 ( .A1(n385), .A2(n502), .B1(n503), .B2(n97), .ZN(n553) );
  NAND2_X1 U351 ( .A1(n312), .A2(n311), .ZN(n314) );
  XNOR2_X1 U352 ( .A(n314), .B(n313), .ZN(n315) );
  NAND2_X1 U353 ( .A1(n315), .A2(n279), .ZN(n316) );
  OAI21_X1 U354 ( .B1(n380), .B2(n502), .A(n316), .ZN(n555) );
  AOI22_X1 U355 ( .A1(n385), .A2(n500), .B1(n501), .B2(n103), .ZN(n557) );
  NAND2_X1 U356 ( .A1(n451), .A2(n400), .ZN(n317) );
  XOR2_X1 U357 ( .A(n317), .B(n405), .Z(n318) );
  NAND2_X1 U358 ( .A1(n279), .A2(n318), .ZN(n319) );
  OAI21_X1 U359 ( .B1(n380), .B2(n500), .A(n319), .ZN(n559) );
  AOI22_X1 U360 ( .A1(n385), .A2(n498), .B1(n499), .B2(n128), .ZN(n561) );
  OAI21_X1 U361 ( .B1(n399), .B2(n405), .A(n400), .ZN(n323) );
  NAND2_X1 U362 ( .A1(n389), .A2(n398), .ZN(n320) );
  XNOR2_X1 U363 ( .A(n323), .B(n320), .ZN(n321) );
  NAND2_X1 U364 ( .A1(n279), .A2(n321), .ZN(n322) );
  OAI21_X1 U365 ( .B1(n385), .B2(n498), .A(n322), .ZN(n563) );
  AOI22_X1 U366 ( .A1(n385), .A2(n496), .B1(n497), .B2(n128), .ZN(n565) );
  AOI21_X1 U367 ( .B1(n323), .B2(n389), .A(n452), .ZN(n327) );
  NAND2_X1 U368 ( .A1(n454), .A2(n397), .ZN(n324) );
  XOR2_X1 U369 ( .A(n327), .B(n324), .Z(n325) );
  NAND2_X1 U370 ( .A1(n279), .A2(n325), .ZN(n326) );
  OAI21_X1 U371 ( .B1(n380), .B2(n496), .A(n326), .ZN(n567) );
  AOI22_X1 U372 ( .A1(n385), .A2(n494), .B1(n495), .B2(n103), .ZN(n569) );
  OAI21_X1 U373 ( .B1(n327), .B2(n396), .A(n397), .ZN(n337) );
  INV_X1 U374 ( .A(n337), .ZN(n331) );
  NAND2_X1 U375 ( .A1(n455), .A2(n395), .ZN(n328) );
  XOR2_X1 U376 ( .A(n331), .B(n328), .Z(n329) );
  NAND2_X1 U377 ( .A1(n237), .A2(n329), .ZN(n330) );
  OAI21_X1 U378 ( .B1(n385), .B2(n494), .A(n330), .ZN(n571) );
  AOI22_X1 U379 ( .A1(n385), .A2(n492), .B1(n493), .B2(n97), .ZN(n573) );
  OAI21_X1 U380 ( .B1(n331), .B2(n394), .A(n395), .ZN(n333) );
  NAND2_X1 U381 ( .A1(n449), .A2(n402), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  NAND2_X1 U383 ( .A1(n237), .A2(n334), .ZN(n335) );
  OAI21_X1 U384 ( .B1(n380), .B2(n492), .A(n335), .ZN(n575) );
  AOI22_X1 U385 ( .A1(n385), .A2(n490), .B1(n491), .B2(n97), .ZN(n577) );
  NOR2_X1 U386 ( .A1(n401), .A2(n394), .ZN(n338) );
  OAI21_X1 U387 ( .B1(n401), .B2(n395), .A(n402), .ZN(n336) );
  AOI21_X1 U388 ( .B1(n338), .B2(n337), .A(n336), .ZN(n364) );
  NAND2_X1 U389 ( .A1(n457), .A2(n393), .ZN(n339) );
  XOR2_X1 U390 ( .A(n364), .B(n339), .Z(n340) );
  NAND2_X1 U391 ( .A1(n279), .A2(n340), .ZN(n341) );
  OAI21_X1 U392 ( .B1(n380), .B2(n490), .A(n341), .ZN(n579) );
  AOI22_X1 U393 ( .A1(n385), .A2(n488), .B1(n489), .B2(n128), .ZN(n581) );
  OAI21_X1 U394 ( .B1(n364), .B2(n392), .A(n393), .ZN(n343) );
  NAND2_X1 U395 ( .A1(n388), .A2(n403), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  NAND2_X1 U397 ( .A1(n279), .A2(n344), .ZN(n345) );
  OAI21_X1 U398 ( .B1(n380), .B2(n488), .A(n345), .ZN(n583) );
  AOI22_X1 U399 ( .A1(n385), .A2(n486), .B1(n487), .B2(n128), .ZN(n585) );
  NAND2_X1 U400 ( .A1(n457), .A2(n388), .ZN(n347) );
  AOI21_X1 U401 ( .B1(n456), .B2(n388), .A(n448), .ZN(n346) );
  OAI21_X1 U402 ( .B1(n364), .B2(n347), .A(n346), .ZN(n349) );
  NAND2_X1 U403 ( .A1(n387), .A2(n404), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  NAND2_X1 U405 ( .A1(n276), .A2(n350), .ZN(n351) );
  OAI21_X1 U406 ( .B1(n380), .B2(n486), .A(n351), .ZN(n587) );
  AOI22_X1 U407 ( .A1(n380), .A2(n484), .B1(n485), .B2(n103), .ZN(n589) );
  NAND2_X1 U408 ( .A1(n388), .A2(n387), .ZN(n353) );
  NOR2_X1 U409 ( .A1(n392), .A2(n353), .ZN(n360) );
  INV_X1 U410 ( .A(n360), .ZN(n355) );
  AOI21_X1 U411 ( .B1(n448), .B2(n387), .A(n447), .ZN(n352) );
  OAI21_X1 U412 ( .B1(n353), .B2(n393), .A(n352), .ZN(n361) );
  INV_X1 U413 ( .A(n361), .ZN(n354) );
  OAI21_X1 U414 ( .B1(n364), .B2(n355), .A(n354), .ZN(n357) );
  NAND2_X1 U415 ( .A1(n386), .A2(n391), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  NAND2_X1 U417 ( .A1(n237), .A2(n358), .ZN(n359) );
  OAI21_X1 U418 ( .B1(n380), .B2(n484), .A(n359), .ZN(n591) );
  AOI22_X1 U419 ( .A1(n380), .A2(n482), .B1(n483), .B2(n103), .ZN(n593) );
  NAND2_X1 U420 ( .A1(n360), .A2(n386), .ZN(n363) );
  AOI21_X1 U421 ( .B1(n361), .B2(n386), .A(n458), .ZN(n362) );
  OAI21_X1 U422 ( .B1(n364), .B2(n363), .A(n362), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n365), .B(n390), .ZN(n366) );
  NAND2_X1 U424 ( .A1(n279), .A2(n366), .ZN(n367) );
  OAI21_X1 U425 ( .B1(n380), .B2(n482), .A(n367), .ZN(n595) );
  NAND2_X1 U426 ( .A1(n276), .A2(B_extended[0]), .ZN(n368) );
  OAI21_X1 U427 ( .B1(n380), .B2(n481), .A(n368), .ZN(n597) );
  NAND2_X1 U428 ( .A1(n237), .A2(B_extended[1]), .ZN(n369) );
  OAI21_X1 U429 ( .B1(n380), .B2(n480), .A(n369), .ZN(n599) );
  NAND2_X1 U430 ( .A1(n276), .A2(B_extended[2]), .ZN(n370) );
  OAI21_X1 U431 ( .B1(n380), .B2(n479), .A(n370), .ZN(n601) );
  NAND2_X1 U432 ( .A1(n276), .A2(B_extended[3]), .ZN(n371) );
  OAI21_X1 U433 ( .B1(n380), .B2(n478), .A(n371), .ZN(n603) );
  NAND2_X1 U434 ( .A1(n279), .A2(B_extended[4]), .ZN(n372) );
  OAI21_X1 U435 ( .B1(n380), .B2(n477), .A(n372), .ZN(n605) );
  NAND2_X1 U436 ( .A1(n276), .A2(B_extended[5]), .ZN(n373) );
  OAI21_X1 U437 ( .B1(n380), .B2(n476), .A(n373), .ZN(n607) );
  NAND2_X1 U438 ( .A1(n279), .A2(B_extended[6]), .ZN(n374) );
  OAI21_X1 U439 ( .B1(n380), .B2(n475), .A(n374), .ZN(n609) );
  NAND2_X1 U440 ( .A1(n237), .A2(B_extended[7]), .ZN(n375) );
  OAI21_X1 U441 ( .B1(n385), .B2(n474), .A(n375), .ZN(n611) );
  NAND2_X1 U442 ( .A1(n279), .A2(A_extended[0]), .ZN(n376) );
  OAI21_X1 U443 ( .B1(n385), .B2(n473), .A(n376), .ZN(n613) );
  NAND2_X1 U444 ( .A1(n279), .A2(A_extended[1]), .ZN(n377) );
  OAI21_X1 U445 ( .B1(n385), .B2(n472), .A(n377), .ZN(n615) );
  NAND2_X1 U446 ( .A1(n276), .A2(A_extended[2]), .ZN(n378) );
  OAI21_X1 U447 ( .B1(n380), .B2(n471), .A(n378), .ZN(n617) );
  NAND2_X1 U448 ( .A1(n279), .A2(A_extended[3]), .ZN(n379) );
  OAI21_X1 U449 ( .B1(n380), .B2(n470), .A(n379), .ZN(n619) );
  NAND2_X1 U450 ( .A1(n237), .A2(A_extended[4]), .ZN(n381) );
  OAI21_X1 U451 ( .B1(n385), .B2(n469), .A(n381), .ZN(n621) );
  NAND2_X1 U452 ( .A1(n279), .A2(A_extended[5]), .ZN(n382) );
  OAI21_X1 U453 ( .B1(n385), .B2(n468), .A(n382), .ZN(n623) );
  NAND2_X1 U454 ( .A1(n279), .A2(A_extended[6]), .ZN(n383) );
  OAI21_X1 U455 ( .B1(n385), .B2(n467), .A(n383), .ZN(n625) );
  NAND2_X1 U456 ( .A1(n279), .A2(A_extended[7]), .ZN(n384) );
  OAI21_X1 U457 ( .B1(n385), .B2(n466), .A(n384), .ZN(n627) );
  NAND2_X1 U458 ( .A1(n465), .A2(n97), .ZN(n629) );
endmodule


module conv_128_32_DW_mult_pipe_J1_28 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n402, n404,
         n406, n408, n410, n412, n414, n416, n418, n420, n422, n424, n426,
         n428, n430, n432, n434, n436, n438, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n515, n517, n519, n521, n523, n525, n527, n529, n531,
         n533, n535, n537, n539, n541, n543, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n567, n569, n571, n573, n575,
         n577, n579, n581, n583, n585, n587, n589, n591, n593, n595, n597,
         n599, n601, n603, n605, n607, n609, n611, n613, n615, n617, n619,
         n621, n623, n640, n641;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n458), .SE(n623), .CK(clk), .Q(n640), 
        .QN(n459) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n458), .SE(n619), .CK(clk), .QN(n461)
         );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n458), .SE(n611), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n465) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n458), .SE(n609), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n466) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n458), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n467) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n458), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n468) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n458), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n469) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n458), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n470) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n458), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n471) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n472) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n458), .SE(n595), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n473) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n593), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n474) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n591), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n475) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n589), .CK(clk), .QN(n476)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n587), .CK(clk), .Q(
        product[15]), .QN(n477) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(rst_n), .SE(n585), .CK(clk), .QN(n478)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(rst_n), .SE(n583), .CK(clk), .Q(
        product[14]), .QN(n479) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(rst_n), .SE(n581), .CK(clk), .QN(n480)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n458), .SE(n579), .CK(clk), .Q(
        product[13]), .QN(n481) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n458), .SE(n577), .CK(clk), .QN(n482)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n458), .SE(n575), .CK(clk), .Q(
        product[12]), .QN(n483) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(rst_n), .SE(n573), .CK(clk), .QN(n484) );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(rst_n), .SE(n571), .CK(clk), .Q(
        product[11]), .QN(n485) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(rst_n), .SE(n569), .CK(clk), .QN(n486) );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(rst_n), .SE(n567), .CK(clk), .Q(
        product[10]), .QN(n487) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(rst_n), .SE(n565), .CK(clk), .QN(n488) );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(rst_n), .SE(n563), .CK(clk), .Q(
        product[9]), .QN(n489) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(rst_n), .SE(n561), .CK(clk), .QN(n490) );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(rst_n), .SE(n559), .CK(clk), .Q(
        product[8]), .QN(n491) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n458), .SE(n557), .CK(clk), .QN(n492)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n458), .SE(n555), .CK(clk), .Q(
        product[7]), .QN(n493) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n458), .SE(n553), .CK(clk), .QN(n494)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n458), .SE(n551), .CK(clk), .Q(
        product[6]), .QN(n495) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n458), .SE(n549), .CK(clk), .QN(n496)
         );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n458), .SE(n547), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n458), .SE(n545), .CK(clk), .Q(
        product[5]), .QN(n498) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n458), .SE(n543), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n458), .SE(n541), .CK(clk), .QN(n500)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n458), .SE(n539), .CK(clk), .Q(
        product[4]), .QN(n501) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n458), .SE(n537), .CK(clk), .QN(n502)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n458), .SE(n535), .CK(clk), .QN(n503)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n458), .SE(n533), .CK(clk), .Q(
        product[3]), .QN(n504) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n458), .SE(n531), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n458), .SE(n529), .CK(clk), .QN(n506)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n458), .SE(n527), .CK(clk), .Q(
        product[2]), .QN(n507) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n458), .SE(n525), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n458), .SE(n523), .CK(clk), .QN(n509)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n458), .SE(n521), .CK(clk), .Q(
        product[1]), .QN(n510) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n458), .SE(n519), .CK(clk), .QN(n511)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n458), .SE(n517), .CK(clk), .QN(n512)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n458), .SE(n515), .CK(clk), .Q(
        product[0]), .QN(n513) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n641), .SI(1'b1), .SE(n438), .CK(clk), 
        .Q(n399), .QN(n440) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2_IP  ( .D(1'b1), .SI(n641), .SE(n436), .CK(
        clk), .Q(n441), .QN(n398) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n641), .SI(1'b1), .SE(n434), .CK(clk), 
        .Q(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n641), .SI(1'b1), .SE(n432), .CK(clk), 
        .Q(n396), .QN(n442) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n641), .SI(1'b1), .SE(n430), .CK(clk), 
        .Q(n395), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n641), .SI(1'b1), .SE(n428), .CK(clk), 
        .Q(n394), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n641), .SI(1'b1), .SE(n426), .CK(clk), 
        .Q(n393), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n641), .SE(n424), .CK(
        clk), .QN(n392) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n641), .SE(n422), .CK(
        clk), .Q(n446), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n641), .SI(1'b1), .SE(n420), .CK(clk), 
        .Q(n390), .QN(n447) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n641), .SI(1'b1), .SE(n418), .CK(clk), 
        .Q(n389), .QN(n448) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n641), .SI(1'b1), .SE(n416), .CK(clk), 
        .Q(n388), .QN(n449) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n641), .SI(1'b1), .SE(n414), .CK(clk), 
        .Q(n387), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n641), .SI(1'b1), .SE(n412), .CK(clk), 
        .Q(n386), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n641), .SI(1'b1), .SE(n410), .CK(clk), 
        .Q(n385) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n641), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n383), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n641), .SE(n404), .CK(
        clk), .Q(n455), .QN(n382) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n641), .SE(n402), .CK(
        clk), .Q(n456), .QN(n381) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n641), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n380), .QN(n457) );
  SDFF_X2 clk_r_REG50_S1 ( .D(1'b0), .SI(n458), .SE(n613), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n464) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n458), .SE(n621), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n460) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n458), .SE(n617), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n462) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n641), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n384), .QN(n453) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n458), .SE(n615), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n463) );
  BUF_X1 U2 ( .A(en), .Z(n351) );
  INV_X1 U3 ( .A(rst_n), .ZN(n641) );
  BUF_X2 U4 ( .A(n25), .Z(n19) );
  BUF_X1 U5 ( .A(n273), .Z(n332) );
  BUF_X1 U6 ( .A(en), .Z(n270) );
  CLKBUF_X1 U7 ( .A(en), .Z(n266) );
  BUF_X1 U8 ( .A(\mult_x_1/n313 ), .Z(n251) );
  INV_X1 U9 ( .A(n273), .ZN(n379) );
  INV_X1 U10 ( .A(n273), .ZN(n372) );
  INV_X1 U11 ( .A(n273), .ZN(n374) );
  INV_X1 U12 ( .A(n273), .ZN(n377) );
  XNOR2_X1 U13 ( .A(n11), .B(n104), .ZN(n120) );
  XNOR2_X1 U14 ( .A(n14), .B(n137), .ZN(n217) );
  XNOR2_X1 U15 ( .A(n105), .B(n103), .ZN(n11) );
  CLKBUF_X2 U16 ( .A(rst_n), .Z(n458) );
  XNOR2_X1 U17 ( .A(n136), .B(n135), .ZN(n14) );
  NAND2_X1 U18 ( .A1(n71), .A2(n70), .ZN(n22) );
  NAND2_X1 U19 ( .A1(n105), .A2(n103), .ZN(n9) );
  INV_X1 U20 ( .A(n26), .ZN(n16) );
  BUF_X2 U21 ( .A(n39), .Z(n5) );
  NAND2_X1 U22 ( .A1(n6), .A2(n74), .ZN(n219) );
  NAND2_X1 U23 ( .A1(n69), .A2(n22), .ZN(n6) );
  NAND2_X1 U24 ( .A1(n7), .A2(n266), .ZN(n224) );
  NAND2_X1 U25 ( .A1(n223), .A2(n222), .ZN(n7) );
  NAND2_X1 U26 ( .A1(n8), .A2(n269), .ZN(n194) );
  NAND2_X1 U27 ( .A1(n193), .A2(n192), .ZN(n8) );
  AND2_X2 U28 ( .A1(n640), .A2(\mult_x_1/n281 ), .ZN(n130) );
  NAND2_X1 U29 ( .A1(n10), .A2(n9), .ZN(n43) );
  OAI21_X1 U30 ( .B1(n103), .B2(n105), .A(n104), .ZN(n10) );
  NAND2_X1 U31 ( .A1(n13), .A2(n12), .ZN(n216) );
  NAND2_X1 U32 ( .A1(n137), .A2(n136), .ZN(n12) );
  OAI21_X1 U33 ( .B1(n137), .B2(n136), .A(n135), .ZN(n13) );
  OAI21_X1 U34 ( .B1(n86), .B2(n87), .A(n85), .ZN(n53) );
  INV_X1 U35 ( .A(n120), .ZN(n117) );
  INV_X1 U36 ( .A(n26), .ZN(n166) );
  INV_X1 U37 ( .A(n31), .ZN(n33) );
  XNOR2_X1 U38 ( .A(n205), .B(n204), .ZN(n232) );
  XNOR2_X1 U39 ( .A(n233), .B(n232), .ZN(n262) );
  XNOR2_X1 U40 ( .A(n231), .B(n230), .ZN(n233) );
  INV_X1 U41 ( .A(n229), .ZN(n230) );
  XNOR2_X1 U42 ( .A(n88), .B(n87), .ZN(n184) );
  OAI21_X1 U43 ( .B1(n207), .B2(n232), .A(n206), .ZN(n210) );
  NOR2_X1 U44 ( .A1(n231), .A2(n229), .ZN(n207) );
  NAND2_X1 U45 ( .A1(n231), .A2(n229), .ZN(n206) );
  NAND2_X1 U46 ( .A1(n122), .A2(n121), .ZN(n267) );
  NAND2_X1 U47 ( .A1(n21), .A2(n118), .ZN(n122) );
  NAND2_X1 U48 ( .A1(n117), .A2(n116), .ZN(n118) );
  NAND2_X1 U49 ( .A1(n124), .A2(n123), .ZN(n59) );
  XNOR2_X1 U50 ( .A(n21), .B(n106), .ZN(n112) );
  OR2_X1 U51 ( .A1(n270), .A2(n450), .ZN(n15) );
  NAND2_X1 U52 ( .A1(n15), .A2(n194), .ZN(n414) );
  XNOR2_X1 U53 ( .A(n73), .B(n72), .ZN(n34) );
  INV_X1 U54 ( .A(n73), .ZN(n71) );
  NAND2_X1 U55 ( .A1(n73), .A2(n72), .ZN(n74) );
  XNOR2_X1 U56 ( .A(n462), .B(n461), .ZN(n17) );
  INV_X1 U57 ( .A(n460), .ZN(n18) );
  XNOR2_X1 U58 ( .A(\mult_x_1/a[4] ), .B(n462), .ZN(n24) );
  NAND2_X1 U59 ( .A1(n459), .A2(\mult_x_1/n310 ), .ZN(n50) );
  XNOR2_X1 U60 ( .A(n464), .B(n463), .ZN(n25) );
  INV_X1 U61 ( .A(n270), .ZN(n20) );
  BUF_X1 U62 ( .A(en), .Z(n269) );
  INV_X1 U63 ( .A(en), .ZN(n273) );
  XOR2_X1 U64 ( .A(n99), .B(n98), .Z(n21) );
  INV_X1 U65 ( .A(n23), .ZN(n124) );
  NAND2_X1 U66 ( .A1(n98), .A2(n99), .ZN(n23) );
  NAND2_X2 U67 ( .A1(n25), .A2(n24), .ZN(n155) );
  XNOR2_X1 U68 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n29) );
  XNOR2_X1 U69 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n281 ), .ZN(n78) );
  OAI22_X1 U70 ( .A1(n155), .A2(n29), .B1(n19), .B2(n78), .ZN(n73) );
  NOR2_X1 U71 ( .A1(n472), .A2(n50), .ZN(n72) );
  XNOR2_X1 U72 ( .A(n462), .B(n461), .ZN(n28) );
  INV_X1 U73 ( .A(n28), .ZN(n26) );
  XNOR2_X1 U74 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n35) );
  XNOR2_X1 U75 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n42) );
  XNOR2_X1 U76 ( .A(n461), .B(\mult_x_1/n310 ), .ZN(n27) );
  NAND2_X2 U77 ( .A1(n27), .A2(n17), .ZN(n165) );
  OAI22_X1 U78 ( .A1(n166), .A2(n35), .B1(n42), .B2(n165), .ZN(n56) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n38) );
  OAI22_X1 U80 ( .A1(n155), .A2(n38), .B1(n19), .B2(n29), .ZN(n55) );
  NOR2_X1 U81 ( .A1(\mult_x_1/a[2] ), .A2(\mult_x_1/n313 ), .ZN(n31) );
  NAND2_X1 U82 ( .A1(\mult_x_1/a[2] ), .A2(\mult_x_1/n313 ), .ZN(n32) );
  NAND2_X1 U83 ( .A1(n32), .A2(n464), .ZN(n30) );
  OAI21_X1 U84 ( .B1(n31), .B2(n246), .A(n30), .ZN(n39) );
  XNOR2_X1 U85 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n40) );
  XNOR2_X1 U86 ( .A(n130), .B(\mult_x_1/n312 ), .ZN(n36) );
  NAND2_X2 U87 ( .A1(n33), .A2(n32), .ZN(n248) );
  OAI22_X1 U88 ( .A1(n39), .A2(n40), .B1(n36), .B2(n248), .ZN(n76) );
  INV_X1 U89 ( .A(n76), .ZN(n54) );
  XNOR2_X1 U90 ( .A(n69), .B(n34), .ZN(n82) );
  XNOR2_X1 U91 ( .A(n18), .B(\mult_x_1/n283 ), .ZN(n79) );
  OAI22_X1 U92 ( .A1(n165), .A2(n35), .B1(n16), .B2(n79), .ZN(n77) );
  AOI21_X1 U93 ( .B1(n248), .B2(n5), .A(n36), .ZN(n37) );
  INV_X1 U94 ( .A(n37), .ZN(n75) );
  XNOR2_X1 U95 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n284 ), .ZN(n90) );
  OAI22_X1 U96 ( .A1(n155), .A2(n90), .B1(n19), .B2(n38), .ZN(n47) );
  XNOR2_X1 U97 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n92) );
  OAI22_X1 U98 ( .A1(n5), .A2(n92), .B1(n248), .B2(n40), .ZN(n46) );
  OR2_X1 U99 ( .A1(n47), .A2(n46), .ZN(n45) );
  NOR2_X1 U100 ( .A1(n473), .A2(n50), .ZN(n44) );
  NAND2_X1 U101 ( .A1(n467), .A2(\mult_x_1/n313 ), .ZN(n252) );
  XNOR2_X1 U102 ( .A(n130), .B(n251), .ZN(n49) );
  AOI21_X1 U103 ( .B1(n252), .B2(n467), .A(n49), .ZN(n41) );
  INV_X1 U104 ( .A(n41), .ZN(n105) );
  XNOR2_X1 U105 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n48) );
  OAI22_X1 U106 ( .A1(n165), .A2(n48), .B1(n166), .B2(n42), .ZN(n104) );
  NOR2_X1 U107 ( .A1(n474), .A2(n50), .ZN(n103) );
  FA_X1 U108 ( .A(n45), .B(n44), .CI(n43), .CO(n80), .S(n125) );
  XNOR2_X1 U109 ( .A(n47), .B(n46), .ZN(n99) );
  XNOR2_X1 U110 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n95) );
  OAI22_X1 U111 ( .A1(n16), .A2(n48), .B1(n95), .B2(n165), .ZN(n86) );
  XNOR2_X1 U112 ( .A(n251), .B(\mult_x_1/n281 ), .ZN(n89) );
  OAI22_X1 U113 ( .A1(n252), .A2(n89), .B1(n49), .B2(n467), .ZN(n87) );
  INV_X1 U114 ( .A(n50), .ZN(n51) );
  AND2_X1 U115 ( .A1(\mult_x_1/n288 ), .A2(n51), .ZN(n85) );
  NAND2_X1 U116 ( .A1(n87), .A2(n86), .ZN(n52) );
  NAND2_X1 U117 ( .A1(n53), .A2(n52), .ZN(n98) );
  FA_X1 U118 ( .A(n56), .B(n55), .CI(n54), .CO(n69), .S(n123) );
  INV_X1 U119 ( .A(n123), .ZN(n57) );
  NAND2_X1 U120 ( .A1(n23), .A2(n57), .ZN(n58) );
  NAND2_X1 U121 ( .A1(n125), .A2(n58), .ZN(n60) );
  NAND2_X1 U122 ( .A1(n60), .A2(n59), .ZN(n64) );
  NAND2_X1 U123 ( .A1(n65), .A2(n64), .ZN(n61) );
  NAND2_X1 U124 ( .A1(n61), .A2(n269), .ZN(n63) );
  NAND2_X1 U125 ( .A1(n20), .A2(n396), .ZN(n62) );
  NAND2_X1 U126 ( .A1(n63), .A2(n62), .ZN(n432) );
  NOR2_X1 U127 ( .A1(n65), .A2(n64), .ZN(n66) );
  NAND2_X1 U128 ( .A1(n66), .A2(n269), .ZN(n68) );
  OR2_X1 U129 ( .A1(n266), .A2(n441), .ZN(n67) );
  NAND2_X1 U130 ( .A1(n68), .A2(n67), .ZN(n436) );
  INV_X1 U131 ( .A(n72), .ZN(n70) );
  FA_X1 U132 ( .A(n77), .B(n76), .CI(n75), .CO(n218), .S(n81) );
  XNOR2_X1 U133 ( .A(n130), .B(\mult_x_1/n311 ), .ZN(n133) );
  OAI22_X1 U134 ( .A1(n155), .A2(n78), .B1(n133), .B2(n19), .ZN(n139) );
  INV_X1 U135 ( .A(n139), .ZN(n137) );
  XNOR2_X1 U136 ( .A(n18), .B(\mult_x_1/n282 ), .ZN(n132) );
  OAI22_X1 U137 ( .A1(n165), .A2(n79), .B1(n16), .B2(n132), .ZN(n136) );
  NOR2_X1 U138 ( .A1(n471), .A2(n50), .ZN(n135) );
  FA_X1 U139 ( .A(n82), .B(n81), .CI(n80), .CO(n222), .S(n65) );
  OAI21_X1 U140 ( .B1(n223), .B2(n222), .A(n269), .ZN(n84) );
  NAND2_X1 U141 ( .A1(n20), .A2(n397), .ZN(n83) );
  NAND2_X1 U142 ( .A1(n84), .A2(n83), .ZN(n434) );
  XNOR2_X1 U143 ( .A(n86), .B(n85), .ZN(n88) );
  XNOR2_X1 U144 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n286 ), .ZN(n153) );
  XNOR2_X1 U145 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n285 ), .ZN(n91) );
  OAI22_X1 U146 ( .A1(n155), .A2(n153), .B1(n19), .B2(n91), .ZN(n149) );
  XNOR2_X1 U147 ( .A(n251), .B(\mult_x_1/n282 ), .ZN(n143) );
  OAI22_X1 U148 ( .A1(n252), .A2(n143), .B1(n89), .B2(n467), .ZN(n148) );
  XNOR2_X1 U149 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n144) );
  XNOR2_X1 U150 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n93) );
  OAI22_X1 U151 ( .A1(n5), .A2(n144), .B1(n248), .B2(n93), .ZN(n147) );
  OAI22_X1 U152 ( .A1(n155), .A2(n91), .B1(n19), .B2(n90), .ZN(n102) );
  OAI22_X1 U153 ( .A1(n5), .A2(n93), .B1(n248), .B2(n92), .ZN(n101) );
  OR2_X1 U154 ( .A1(\mult_x_1/n288 ), .A2(n460), .ZN(n94) );
  OAI22_X1 U155 ( .A1(n165), .A2(n460), .B1(n94), .B2(n166), .ZN(n146) );
  XNOR2_X1 U156 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n96) );
  OAI22_X1 U157 ( .A1(n165), .A2(n96), .B1(n166), .B2(n95), .ZN(n145) );
  INV_X1 U158 ( .A(n111), .ZN(n97) );
  AND2_X1 U159 ( .A1(n269), .A2(n97), .ZN(n108) );
  FA_X1 U160 ( .A(n102), .B(n101), .CI(n100), .CO(n119), .S(n182) );
  XNOR2_X1 U161 ( .A(n119), .B(n120), .ZN(n106) );
  INV_X1 U162 ( .A(n112), .ZN(n107) );
  NAND2_X1 U163 ( .A1(n108), .A2(n107), .ZN(n110) );
  OR2_X1 U164 ( .A1(n270), .A2(n453), .ZN(n109) );
  NAND2_X1 U165 ( .A1(n110), .A2(n109), .ZN(n408) );
  NAND2_X1 U166 ( .A1(n112), .A2(n111), .ZN(n113) );
  NAND2_X1 U167 ( .A1(n113), .A2(n269), .ZN(n115) );
  NAND2_X1 U168 ( .A1(n20), .A2(n385), .ZN(n114) );
  NAND2_X1 U169 ( .A1(n115), .A2(n114), .ZN(n410) );
  INV_X1 U170 ( .A(n119), .ZN(n116) );
  NAND2_X1 U171 ( .A1(n120), .A2(n119), .ZN(n121) );
  XNOR2_X1 U172 ( .A(n124), .B(n123), .ZN(n126) );
  XNOR2_X1 U173 ( .A(n126), .B(n125), .ZN(n271) );
  NAND2_X1 U174 ( .A1(n267), .A2(n271), .ZN(n127) );
  NAND2_X1 U175 ( .A1(n127), .A2(n266), .ZN(n129) );
  NAND2_X1 U176 ( .A1(n20), .A2(n392), .ZN(n128) );
  NAND2_X1 U177 ( .A1(n129), .A2(n128), .ZN(n424) );
  NOR2_X1 U198 ( .A1(n469), .A2(n50), .ZN(n163) );
  XNOR2_X1 U199 ( .A(n18), .B(\mult_x_1/n281 ), .ZN(n131) );
  XNOR2_X1 U200 ( .A(n130), .B(n18), .ZN(n164) );
  OAI22_X1 U201 ( .A1(n165), .A2(n131), .B1(n164), .B2(n16), .ZN(n171) );
  INV_X1 U202 ( .A(n171), .ZN(n162) );
  OAI22_X1 U203 ( .A1(n165), .A2(n132), .B1(n16), .B2(n131), .ZN(n140) );
  AOI21_X1 U204 ( .B1(n19), .B2(n155), .A(n133), .ZN(n134) );
  INV_X1 U205 ( .A(n134), .ZN(n138) );
  NOR2_X1 U206 ( .A1(n470), .A2(n50), .ZN(n215) );
  FA_X1 U207 ( .A(n140), .B(n139), .CI(n138), .CO(n161), .S(n214) );
  OR2_X1 U208 ( .A1(n179), .A2(n178), .ZN(n141) );
  NAND2_X1 U209 ( .A1(n351), .A2(n141), .ZN(n142) );
  OAI21_X1 U210 ( .B1(n270), .B2(n457), .A(n142), .ZN(n400) );
  XNOR2_X1 U211 ( .A(n251), .B(\mult_x_1/n283 ), .ZN(n203) );
  OAI22_X1 U212 ( .A1(n252), .A2(n203), .B1(n143), .B2(n467), .ZN(n158) );
  AND2_X1 U213 ( .A1(\mult_x_1/n288 ), .A2(n26), .ZN(n157) );
  XNOR2_X1 U214 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n202) );
  OAI22_X1 U215 ( .A1(n5), .A2(n202), .B1(n248), .B2(n144), .ZN(n156) );
  HA_X1 U216 ( .A(n146), .B(n145), .CO(n100), .S(n186) );
  FA_X1 U217 ( .A(n149), .B(n148), .CI(n147), .CO(n183), .S(n185) );
  INV_X1 U218 ( .A(\mult_x_1/n311 ), .ZN(n151) );
  OR2_X1 U219 ( .A1(\mult_x_1/n288 ), .A2(n151), .ZN(n150) );
  OAI22_X1 U220 ( .A1(n155), .A2(n151), .B1(n150), .B2(n19), .ZN(n205) );
  XNOR2_X1 U221 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n288 ), .ZN(n152) );
  XNOR2_X1 U222 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n154) );
  OAI22_X1 U223 ( .A1(n155), .A2(n152), .B1(n19), .B2(n154), .ZN(n204) );
  AND2_X1 U224 ( .A1(n205), .A2(n204), .ZN(n201) );
  OAI22_X1 U225 ( .A1(n155), .A2(n154), .B1(n19), .B2(n153), .ZN(n200) );
  FA_X1 U226 ( .A(n158), .B(n157), .CI(n156), .CO(n187), .S(n199) );
  OR2_X1 U227 ( .A1(n196), .A2(n195), .ZN(n159) );
  NAND2_X1 U228 ( .A1(n351), .A2(n159), .ZN(n160) );
  OAI21_X1 U229 ( .B1(n270), .B2(n456), .A(n160), .ZN(n402) );
  FA_X1 U230 ( .A(n163), .B(n162), .CI(n161), .CO(n173), .S(n179) );
  AOI21_X1 U231 ( .B1(n16), .B2(n165), .A(n164), .ZN(n167) );
  INV_X1 U232 ( .A(n167), .ZN(n169) );
  NOR2_X1 U233 ( .A1(n468), .A2(n50), .ZN(n168) );
  XOR2_X1 U234 ( .A(n169), .B(n168), .Z(n170) );
  XOR2_X1 U235 ( .A(n171), .B(n170), .Z(n172) );
  OR2_X1 U236 ( .A1(n173), .A2(n172), .ZN(n175) );
  NAND2_X1 U237 ( .A1(n173), .A2(n172), .ZN(n174) );
  NAND2_X1 U238 ( .A1(n175), .A2(n174), .ZN(n176) );
  NAND2_X1 U239 ( .A1(n351), .A2(n176), .ZN(n177) );
  OAI21_X1 U240 ( .B1(n270), .B2(n455), .A(n177), .ZN(n404) );
  NAND2_X1 U241 ( .A1(n179), .A2(n178), .ZN(n180) );
  NAND2_X1 U242 ( .A1(n269), .A2(n180), .ZN(n181) );
  OAI21_X1 U243 ( .B1(n270), .B2(n454), .A(n181), .ZN(n406) );
  FA_X1 U244 ( .A(n184), .B(n183), .CI(n182), .CO(n111), .S(n193) );
  INV_X1 U245 ( .A(n193), .ZN(n190) );
  FA_X1 U246 ( .A(n187), .B(n186), .CI(n185), .CO(n192), .S(n196) );
  INV_X1 U247 ( .A(n192), .ZN(n188) );
  AND2_X1 U248 ( .A1(n269), .A2(n188), .ZN(n189) );
  NAND2_X1 U249 ( .A1(n190), .A2(n189), .ZN(n191) );
  OAI21_X1 U250 ( .B1(n270), .B2(n451), .A(n191), .ZN(n412) );
  NAND2_X1 U251 ( .A1(n196), .A2(n195), .ZN(n197) );
  NAND2_X1 U252 ( .A1(n269), .A2(n197), .ZN(n198) );
  OAI21_X1 U253 ( .B1(n270), .B2(n449), .A(n198), .ZN(n416) );
  FA_X1 U254 ( .A(n201), .B(n200), .CI(n199), .CO(n195), .S(n211) );
  XNOR2_X1 U255 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n236) );
  OAI22_X1 U256 ( .A1(n5), .A2(n236), .B1(n248), .B2(n202), .ZN(n231) );
  XNOR2_X1 U257 ( .A(n251), .B(\mult_x_1/n284 ), .ZN(n234) );
  OAI22_X1 U258 ( .A1(n252), .A2(n234), .B1(n203), .B2(n467), .ZN(n229) );
  NOR2_X1 U259 ( .A1(n211), .A2(n210), .ZN(n208) );
  NAND2_X1 U260 ( .A1(n266), .A2(n208), .ZN(n209) );
  OAI21_X1 U261 ( .B1(n270), .B2(n448), .A(n209), .ZN(n418) );
  NAND2_X1 U262 ( .A1(n211), .A2(n210), .ZN(n212) );
  NAND2_X1 U263 ( .A1(n269), .A2(n212), .ZN(n213) );
  OAI21_X1 U264 ( .B1(n270), .B2(n447), .A(n213), .ZN(n420) );
  FA_X1 U265 ( .A(n216), .B(n215), .CI(n214), .CO(n178), .S(n226) );
  FA_X1 U266 ( .A(n219), .B(n218), .CI(n217), .CO(n225), .S(n223) );
  NAND2_X1 U267 ( .A1(n226), .A2(n225), .ZN(n220) );
  NAND2_X1 U268 ( .A1(n266), .A2(n220), .ZN(n221) );
  OAI21_X1 U269 ( .B1(n266), .B2(n445), .A(n221), .ZN(n426) );
  OAI21_X1 U270 ( .B1(n266), .B2(n444), .A(n224), .ZN(n428) );
  OR2_X1 U271 ( .A1(n226), .A2(n225), .ZN(n227) );
  NAND2_X1 U272 ( .A1(n269), .A2(n227), .ZN(n228) );
  OAI21_X1 U273 ( .B1(n266), .B2(n443), .A(n228), .ZN(n430) );
  XNOR2_X1 U274 ( .A(n251), .B(\mult_x_1/n285 ), .ZN(n242) );
  OAI22_X1 U275 ( .A1(n252), .A2(n242), .B1(n234), .B2(n467), .ZN(n239) );
  INV_X1 U276 ( .A(n19), .ZN(n235) );
  AND2_X1 U277 ( .A1(\mult_x_1/n288 ), .A2(n235), .ZN(n238) );
  XNOR2_X1 U278 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n240) );
  OAI22_X1 U279 ( .A1(n5), .A2(n240), .B1(n248), .B2(n236), .ZN(n237) );
  OR2_X1 U280 ( .A1(n262), .A2(n261), .ZN(n302) );
  FA_X1 U281 ( .A(n239), .B(n238), .CI(n237), .CO(n261), .S(n260) );
  XNOR2_X1 U282 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n241) );
  OAI22_X1 U283 ( .A1(n5), .A2(n241), .B1(n248), .B2(n240), .ZN(n244) );
  XNOR2_X1 U284 ( .A(n251), .B(\mult_x_1/n286 ), .ZN(n247) );
  OAI22_X1 U285 ( .A1(n252), .A2(n247), .B1(n242), .B2(n467), .ZN(n243) );
  NOR2_X1 U286 ( .A1(n260), .A2(n259), .ZN(n294) );
  HA_X1 U287 ( .A(n244), .B(n243), .CO(n259), .S(n257) );
  INV_X1 U288 ( .A(\mult_x_1/n312 ), .ZN(n246) );
  OR2_X1 U289 ( .A1(\mult_x_1/n288 ), .A2(n246), .ZN(n245) );
  OAI22_X1 U290 ( .A1(n5), .A2(n246), .B1(n245), .B2(n248), .ZN(n256) );
  OR2_X1 U291 ( .A1(n257), .A2(n256), .ZN(n289) );
  XNOR2_X1 U292 ( .A(n251), .B(\mult_x_1/n287 ), .ZN(n250) );
  OAI22_X1 U293 ( .A1(n252), .A2(n250), .B1(n247), .B2(n467), .ZN(n255) );
  INV_X1 U294 ( .A(n248), .ZN(n249) );
  AND2_X1 U295 ( .A1(\mult_x_1/n288 ), .A2(n249), .ZN(n254) );
  NOR2_X1 U296 ( .A1(n255), .A2(n254), .ZN(n281) );
  OAI22_X1 U297 ( .A1(n252), .A2(\mult_x_1/n288 ), .B1(n250), .B2(n467), .ZN(
        n277) );
  OR2_X1 U298 ( .A1(\mult_x_1/n288 ), .A2(n466), .ZN(n253) );
  NAND2_X1 U299 ( .A1(n253), .A2(n252), .ZN(n276) );
  NAND2_X1 U300 ( .A1(n277), .A2(n276), .ZN(n284) );
  NAND2_X1 U301 ( .A1(n255), .A2(n254), .ZN(n282) );
  OAI21_X1 U302 ( .B1(n281), .B2(n284), .A(n282), .ZN(n290) );
  NAND2_X1 U303 ( .A1(n257), .A2(n256), .ZN(n288) );
  INV_X1 U304 ( .A(n288), .ZN(n258) );
  AOI21_X1 U305 ( .B1(n289), .B2(n290), .A(n258), .ZN(n297) );
  NAND2_X1 U306 ( .A1(n260), .A2(n259), .ZN(n295) );
  OAI21_X1 U307 ( .B1(n294), .B2(n297), .A(n295), .ZN(n303) );
  NAND2_X1 U308 ( .A1(n262), .A2(n261), .ZN(n301) );
  INV_X1 U309 ( .A(n301), .ZN(n263) );
  AOI21_X1 U310 ( .B1(n302), .B2(n303), .A(n263), .ZN(n264) );
  NAND2_X1 U311 ( .A1(n351), .A2(n264), .ZN(n265) );
  OAI21_X1 U312 ( .B1(n266), .B2(n440), .A(n265), .ZN(n438) );
  INV_X1 U313 ( .A(n267), .ZN(n268) );
  NAND2_X1 U314 ( .A1(n269), .A2(n268), .ZN(n272) );
  OAI22_X1 U315 ( .A1(n272), .A2(n271), .B1(n270), .B2(n446), .ZN(n422) );
  AOI22_X1 U316 ( .A1(n351), .A2(n512), .B1(n513), .B2(n332), .ZN(n515) );
  AOI22_X1 U317 ( .A1(n351), .A2(n511), .B1(n512), .B2(n332), .ZN(n517) );
  AND2_X1 U318 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n274) );
  NAND2_X1 U319 ( .A1(n379), .A2(n274), .ZN(n275) );
  OAI21_X1 U320 ( .B1(n379), .B2(n511), .A(n275), .ZN(n519) );
  AOI22_X1 U321 ( .A1(n351), .A2(n509), .B1(n510), .B2(n332), .ZN(n521) );
  AOI22_X1 U322 ( .A1(n351), .A2(n508), .B1(n509), .B2(n332), .ZN(n523) );
  OR2_X1 U323 ( .A1(n277), .A2(n276), .ZN(n278) );
  AND2_X1 U324 ( .A1(n278), .A2(n284), .ZN(n279) );
  NAND2_X1 U325 ( .A1(n377), .A2(n279), .ZN(n280) );
  OAI21_X1 U326 ( .B1(n377), .B2(n508), .A(n280), .ZN(n525) );
  AOI22_X1 U327 ( .A1(n351), .A2(n506), .B1(n507), .B2(n332), .ZN(n527) );
  AOI22_X1 U328 ( .A1(n351), .A2(n505), .B1(n506), .B2(n332), .ZN(n529) );
  INV_X1 U329 ( .A(n281), .ZN(n283) );
  NAND2_X1 U330 ( .A1(n283), .A2(n282), .ZN(n285) );
  XOR2_X1 U331 ( .A(n285), .B(n284), .Z(n286) );
  NAND2_X1 U332 ( .A1(n374), .A2(n286), .ZN(n287) );
  OAI21_X1 U333 ( .B1(n377), .B2(n505), .A(n287), .ZN(n531) );
  AOI22_X1 U334 ( .A1(n351), .A2(n503), .B1(n504), .B2(n332), .ZN(n533) );
  AOI22_X1 U335 ( .A1(n351), .A2(n502), .B1(n503), .B2(n332), .ZN(n535) );
  NAND2_X1 U336 ( .A1(n289), .A2(n288), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n292) );
  NAND2_X1 U338 ( .A1(n374), .A2(n292), .ZN(n293) );
  OAI21_X1 U339 ( .B1(n372), .B2(n502), .A(n293), .ZN(n537) );
  AOI22_X1 U340 ( .A1(n351), .A2(n500), .B1(n501), .B2(n332), .ZN(n539) );
  AOI22_X1 U341 ( .A1(n351), .A2(n499), .B1(n500), .B2(n332), .ZN(n541) );
  INV_X1 U342 ( .A(n294), .ZN(n296) );
  NAND2_X1 U343 ( .A1(n296), .A2(n295), .ZN(n298) );
  XOR2_X1 U344 ( .A(n298), .B(n297), .Z(n299) );
  NAND2_X1 U345 ( .A1(n374), .A2(n299), .ZN(n300) );
  OAI21_X1 U346 ( .B1(n377), .B2(n499), .A(n300), .ZN(n543) );
  AOI22_X1 U347 ( .A1(n351), .A2(n497), .B1(n498), .B2(n332), .ZN(n545) );
  AOI22_X1 U348 ( .A1(n379), .A2(n496), .B1(n497), .B2(n332), .ZN(n547) );
  NAND2_X1 U349 ( .A1(n302), .A2(n301), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  NAND2_X1 U351 ( .A1(n305), .A2(n374), .ZN(n306) );
  OAI21_X1 U352 ( .B1(n377), .B2(n496), .A(n306), .ZN(n549) );
  AOI22_X1 U353 ( .A1(n379), .A2(n494), .B1(n495), .B2(n332), .ZN(n551) );
  NAND2_X1 U354 ( .A1(n448), .A2(n390), .ZN(n307) );
  XOR2_X1 U355 ( .A(n307), .B(n399), .Z(n308) );
  NAND2_X1 U356 ( .A1(n374), .A2(n308), .ZN(n309) );
  OAI21_X1 U357 ( .B1(n372), .B2(n494), .A(n309), .ZN(n553) );
  AOI22_X1 U358 ( .A1(n379), .A2(n492), .B1(n493), .B2(n332), .ZN(n555) );
  OAI21_X1 U359 ( .B1(n389), .B2(n399), .A(n390), .ZN(n313) );
  NAND2_X1 U360 ( .A1(n381), .A2(n388), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n313), .B(n310), .ZN(n311) );
  NAND2_X1 U362 ( .A1(n374), .A2(n311), .ZN(n312) );
  OAI21_X1 U363 ( .B1(n377), .B2(n492), .A(n312), .ZN(n557) );
  AOI22_X1 U364 ( .A1(n379), .A2(n490), .B1(n491), .B2(n332), .ZN(n559) );
  AOI21_X1 U365 ( .B1(n313), .B2(n381), .A(n449), .ZN(n317) );
  NAND2_X1 U366 ( .A1(n451), .A2(n387), .ZN(n314) );
  XOR2_X1 U367 ( .A(n317), .B(n314), .Z(n315) );
  NAND2_X1 U368 ( .A1(n377), .A2(n315), .ZN(n316) );
  OAI21_X1 U369 ( .B1(n377), .B2(n490), .A(n316), .ZN(n561) );
  AOI22_X1 U370 ( .A1(n379), .A2(n488), .B1(n489), .B2(n20), .ZN(n563) );
  OAI21_X1 U371 ( .B1(n317), .B2(n386), .A(n387), .ZN(n327) );
  INV_X1 U372 ( .A(n327), .ZN(n321) );
  NAND2_X1 U373 ( .A1(n453), .A2(n385), .ZN(n318) );
  XOR2_X1 U374 ( .A(n321), .B(n318), .Z(n319) );
  NAND2_X1 U375 ( .A1(n377), .A2(n319), .ZN(n320) );
  OAI21_X1 U376 ( .B1(n377), .B2(n488), .A(n320), .ZN(n565) );
  AOI22_X1 U377 ( .A1(n379), .A2(n486), .B1(n487), .B2(n20), .ZN(n567) );
  OAI21_X1 U378 ( .B1(n321), .B2(n384), .A(n385), .ZN(n323) );
  NAND2_X1 U379 ( .A1(n446), .A2(n392), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  NAND2_X1 U381 ( .A1(n377), .A2(n324), .ZN(n325) );
  OAI21_X1 U382 ( .B1(n372), .B2(n486), .A(n325), .ZN(n569) );
  AOI22_X1 U383 ( .A1(n379), .A2(n484), .B1(n485), .B2(n20), .ZN(n571) );
  NOR2_X1 U384 ( .A1(n391), .A2(n384), .ZN(n328) );
  OAI21_X1 U385 ( .B1(n391), .B2(n385), .A(n392), .ZN(n326) );
  AOI21_X1 U386 ( .B1(n328), .B2(n327), .A(n326), .ZN(n356) );
  NAND2_X1 U387 ( .A1(n441), .A2(n396), .ZN(n329) );
  XOR2_X1 U388 ( .A(n356), .B(n329), .Z(n330) );
  NAND2_X1 U389 ( .A1(n377), .A2(n330), .ZN(n331) );
  OAI21_X1 U390 ( .B1(n372), .B2(n484), .A(n331), .ZN(n573) );
  AOI22_X1 U391 ( .A1(n351), .A2(n482), .B1(n483), .B2(n332), .ZN(n575) );
  OAI21_X1 U392 ( .B1(n356), .B2(n398), .A(n396), .ZN(n334) );
  NAND2_X1 U393 ( .A1(n397), .A2(n394), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  NAND2_X1 U395 ( .A1(n377), .A2(n335), .ZN(n336) );
  OAI21_X1 U396 ( .B1(n372), .B2(n482), .A(n336), .ZN(n577) );
  AOI22_X1 U397 ( .A1(n379), .A2(n480), .B1(n481), .B2(n332), .ZN(n579) );
  NAND2_X1 U398 ( .A1(n441), .A2(n397), .ZN(n338) );
  AOI21_X1 U399 ( .B1(n442), .B2(n397), .A(n444), .ZN(n337) );
  OAI21_X1 U400 ( .B1(n356), .B2(n338), .A(n337), .ZN(n340) );
  NAND2_X1 U401 ( .A1(n395), .A2(n393), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  NAND2_X1 U403 ( .A1(n377), .A2(n341), .ZN(n342) );
  OAI21_X1 U404 ( .B1(n372), .B2(n480), .A(n342), .ZN(n581) );
  AOI22_X1 U405 ( .A1(n351), .A2(n478), .B1(n479), .B2(n332), .ZN(n583) );
  NAND2_X1 U406 ( .A1(n397), .A2(n395), .ZN(n344) );
  NOR2_X1 U407 ( .A1(n398), .A2(n344), .ZN(n352) );
  INV_X1 U408 ( .A(n352), .ZN(n346) );
  AOI21_X1 U409 ( .B1(n444), .B2(n395), .A(n445), .ZN(n343) );
  OAI21_X1 U410 ( .B1(n344), .B2(n396), .A(n343), .ZN(n353) );
  INV_X1 U411 ( .A(n353), .ZN(n345) );
  OAI21_X1 U412 ( .B1(n356), .B2(n346), .A(n345), .ZN(n348) );
  NAND2_X1 U413 ( .A1(n380), .A2(n383), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n349) );
  NAND2_X1 U415 ( .A1(n377), .A2(n349), .ZN(n350) );
  OAI21_X1 U416 ( .B1(n372), .B2(n478), .A(n350), .ZN(n585) );
  AOI22_X1 U417 ( .A1(n351), .A2(n476), .B1(n477), .B2(n332), .ZN(n587) );
  NAND2_X1 U418 ( .A1(n352), .A2(n380), .ZN(n355) );
  AOI21_X1 U419 ( .B1(n353), .B2(n380), .A(n454), .ZN(n354) );
  OAI21_X1 U420 ( .B1(n356), .B2(n355), .A(n354), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n357), .B(n382), .ZN(n358) );
  NAND2_X1 U422 ( .A1(n377), .A2(n358), .ZN(n359) );
  OAI21_X1 U423 ( .B1(n372), .B2(n476), .A(n359), .ZN(n589) );
  NAND2_X1 U424 ( .A1(n374), .A2(B_extended[0]), .ZN(n360) );
  OAI21_X1 U425 ( .B1(n372), .B2(n475), .A(n360), .ZN(n591) );
  NAND2_X1 U426 ( .A1(n377), .A2(B_extended[1]), .ZN(n361) );
  OAI21_X1 U427 ( .B1(n372), .B2(n474), .A(n361), .ZN(n593) );
  NAND2_X1 U428 ( .A1(n374), .A2(B_extended[2]), .ZN(n362) );
  OAI21_X1 U429 ( .B1(n372), .B2(n473), .A(n362), .ZN(n595) );
  NAND2_X1 U430 ( .A1(n374), .A2(B_extended[3]), .ZN(n363) );
  OAI21_X1 U431 ( .B1(n372), .B2(n472), .A(n363), .ZN(n597) );
  NAND2_X1 U432 ( .A1(n374), .A2(B_extended[4]), .ZN(n364) );
  OAI21_X1 U433 ( .B1(n372), .B2(n471), .A(n364), .ZN(n599) );
  NAND2_X1 U434 ( .A1(n374), .A2(B_extended[5]), .ZN(n365) );
  OAI21_X1 U435 ( .B1(n372), .B2(n470), .A(n365), .ZN(n601) );
  NAND2_X1 U436 ( .A1(n374), .A2(B_extended[6]), .ZN(n366) );
  OAI21_X1 U437 ( .B1(n372), .B2(n469), .A(n366), .ZN(n603) );
  NAND2_X1 U438 ( .A1(n374), .A2(B_extended[7]), .ZN(n367) );
  OAI21_X1 U439 ( .B1(n379), .B2(n468), .A(n367), .ZN(n605) );
  NAND2_X1 U440 ( .A1(n374), .A2(A_extended[0]), .ZN(n368) );
  OAI21_X1 U441 ( .B1(n379), .B2(n467), .A(n368), .ZN(n607) );
  NAND2_X1 U442 ( .A1(n374), .A2(A_extended[1]), .ZN(n369) );
  OAI21_X1 U443 ( .B1(n379), .B2(n466), .A(n369), .ZN(n609) );
  NAND2_X1 U444 ( .A1(n374), .A2(A_extended[2]), .ZN(n370) );
  OAI21_X1 U445 ( .B1(n372), .B2(n465), .A(n370), .ZN(n611) );
  NAND2_X1 U446 ( .A1(n374), .A2(A_extended[3]), .ZN(n371) );
  OAI21_X1 U447 ( .B1(n372), .B2(n464), .A(n371), .ZN(n613) );
  NAND2_X1 U448 ( .A1(n372), .A2(A_extended[4]), .ZN(n373) );
  OAI21_X1 U449 ( .B1(n379), .B2(n463), .A(n373), .ZN(n615) );
  NAND2_X1 U450 ( .A1(n374), .A2(A_extended[5]), .ZN(n375) );
  OAI21_X1 U451 ( .B1(n379), .B2(n151), .A(n375), .ZN(n617) );
  NAND2_X1 U452 ( .A1(n379), .A2(A_extended[6]), .ZN(n376) );
  OAI21_X1 U453 ( .B1(n379), .B2(n461), .A(n376), .ZN(n619) );
  NAND2_X1 U454 ( .A1(n377), .A2(A_extended[7]), .ZN(n378) );
  OAI21_X1 U455 ( .B1(n379), .B2(n460), .A(n378), .ZN(n621) );
  NAND2_X1 U456 ( .A1(n459), .A2(n20), .ZN(n623) );
endmodule


module conv_128_32_DW_mult_pipe_J1_29 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n415, n417, n419, n421, n423, n425, n427, n429, n431,
         n433, n435, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n530, n532,
         n534, n536, n538, n540, n542, n544, n546, n548, n550, n552, n554,
         n556, n558, n560, n562, n564, n566, n568, n570, n572, n574, n576,
         n578, n580, n582, n584, n586, n588, n590, n592, n594, n596, n598,
         n600, n602, n604, n606, n608, n610, n612, n614, n616, n618, n620,
         n622, n624, n626, n628, n630, n632, n634, n636, n638, n655, n656;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n473), .SE(n630), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n478) );
  SDFF_X1 clk_r_REG54_S1 ( .D(1'b0), .SI(n473), .SE(n626), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n480) );
  SDFF_X1 clk_r_REG58_S1 ( .D(1'b0), .SI(n473), .SE(n624), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n481) );
  SDFF_X1 clk_r_REG62_S1 ( .D(1'b0), .SI(n473), .SE(n622), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n482) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n473), .SE(n618), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n484) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n473), .SE(n616), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n485) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n473), .SE(n614), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n486) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(rst_n), .SE(n612), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n487) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n473), .SE(n610), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n488) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(rst_n), .SE(n608), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n489) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(rst_n), .SE(n606), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n490) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(rst_n), .SE(n604), .CK(clk), .QN(n491) );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(rst_n), .SE(n602), .CK(clk), .Q(
        product[15]), .QN(n492) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(rst_n), .SE(n600), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(rst_n), .SE(n598), .CK(clk), .Q(
        product[14]), .QN(n494) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(rst_n), .SE(n596), .CK(clk), .QN(n495) );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n473), .SE(n594), .CK(clk), .Q(
        product[13]), .QN(n496) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n473), .SE(n592), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n473), .SE(n590), .CK(clk), .Q(
        product[12]), .QN(n498) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(rst_n), .SE(n588), .CK(clk), .QN(n499) );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(rst_n), .SE(n586), .CK(clk), .Q(
        product[11]), .QN(n500) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(rst_n), .SE(n584), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(rst_n), .SE(n582), .CK(clk), .Q(
        product[10]), .QN(n502) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(rst_n), .SE(n580), .CK(clk), .QN(n503)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(rst_n), .SE(n578), .CK(clk), .Q(
        product[9]), .QN(n504) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(rst_n), .SE(n576), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(rst_n), .SE(n574), .CK(clk), .Q(
        product[8]), .QN(n506) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n473), .SE(n572), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n473), .SE(n570), .CK(clk), .Q(
        product[7]), .QN(n508) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n473), .SE(n568), .CK(clk), .QN(n509)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n473), .SE(n566), .CK(clk), .Q(
        product[6]), .QN(n510) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n473), .SE(n562), .CK(clk), .QN(n512)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n473), .SE(n560), .CK(clk), .Q(
        product[5]), .QN(n513) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n473), .SE(n558), .CK(clk), .QN(n514)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n473), .SE(n556), .CK(clk), .QN(n515)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n473), .SE(n554), .CK(clk), .Q(
        product[4]), .QN(n516) );
  SDFF_X1 clk_r_REG51_S2 ( .D(1'b0), .SI(n473), .SE(n552), .CK(clk), .QN(n517)
         );
  SDFF_X1 clk_r_REG52_S3 ( .D(1'b0), .SI(n473), .SE(n550), .CK(clk), .QN(n518)
         );
  SDFF_X1 clk_r_REG53_S4 ( .D(1'b0), .SI(n473), .SE(n548), .CK(clk), .Q(
        product[3]), .QN(n519) );
  SDFF_X1 clk_r_REG55_S2 ( .D(1'b0), .SI(n473), .SE(n546), .CK(clk), .QN(n520)
         );
  SDFF_X1 clk_r_REG56_S3 ( .D(1'b0), .SI(n473), .SE(n544), .CK(clk), .QN(n521)
         );
  SDFF_X1 clk_r_REG57_S4 ( .D(1'b0), .SI(n473), .SE(n542), .CK(clk), .Q(
        product[2]), .QN(n522) );
  SDFF_X1 clk_r_REG59_S2 ( .D(1'b0), .SI(n473), .SE(n540), .CK(clk), .QN(n523)
         );
  SDFF_X1 clk_r_REG60_S3 ( .D(1'b0), .SI(n473), .SE(n538), .CK(clk), .QN(n524)
         );
  SDFF_X1 clk_r_REG61_S4 ( .D(1'b0), .SI(n473), .SE(n536), .CK(clk), .Q(
        product[1]), .QN(n525) );
  SDFF_X1 clk_r_REG63_S2 ( .D(1'b0), .SI(n473), .SE(n534), .CK(clk), .QN(n526)
         );
  SDFF_X1 clk_r_REG64_S3 ( .D(1'b0), .SI(n473), .SE(n532), .CK(clk), .QN(n527)
         );
  SDFF_X1 clk_r_REG65_S4 ( .D(1'b0), .SI(n473), .SE(n530), .CK(clk), .Q(
        product[0]), .QN(n528) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n656), .SE(n429), .CK(
        clk), .Q(n464), .QN(n401) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n656), .SI(1'b1), .SE(n451), .CK(clk), 
        .Q(n412), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n656), .SI(1'b1), .SE(n449), .CK(clk), 
        .Q(n411), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n656), .SE(n447), .CK(
        clk), .Q(n455), .QN(n410) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n656), .SE(n445), .CK(
        clk), .Q(n456), .QN(n409) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n656), .SI(1'b1), .SE(n443), .CK(clk), 
        .Q(n408), .QN(n457) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n656), .SI(1'b1), .SE(n441), .CK(clk), 
        .Q(n407), .QN(n458) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n656), .SI(1'b1), .SE(n439), .CK(clk), 
        .Q(n406), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n656), .SI(1'b1), .SE(n437), .CK(clk), 
        .Q(n405), .QN(n460) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n656), .SI(1'b1), .SE(n435), .CK(clk), 
        .Q(n404), .QN(n461) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n656), .SI(1'b1), .SE(n433), .CK(clk), 
        .Q(n403), .QN(n462) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n656), .SI(1'b1), .SE(n427), .CK(clk), 
        .Q(n400), .QN(n465) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n656), .SI(1'b1), .SE(n425), .CK(clk), 
        .Q(n399), .QN(n466) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n656), .SI(1'b1), .SE(n423), .CK(clk), 
        .Q(n398), .QN(n467) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2_IP  ( .D(1'b1), .SI(n656), .SE(n421), .CK(
        clk), .Q(n468), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n656), .SE(n419), .CK(
        clk), .Q(n469), .QN(n396) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n656), .SI(1'b1), .SE(n417), .CK(clk), 
        .Q(n395), .QN(n470) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n656), .SI(1'b1), .SE(n415), .CK(clk), 
        .Q(n394), .QN(n471) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n656), .SI(1'b1), .SE(n413), .CK(clk), 
        .Q(n393), .QN(n472) );
  SDFF_X1 clk_r_REG50_S1 ( .D(1'b0), .SI(n473), .SE(n628), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n479) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n473), .SE(n632), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n477) );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n473), .SE(n636), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n475) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(rst_n), .SE(n634), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n476) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(rst_n), .SE(n638), .CK(clk), .Q(n655), 
        .QN(n474) );
  SDFF_X1 clk_r_REG66_S1 ( .D(1'b0), .SI(n473), .SE(n620), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n483) );
  SDFF_X1 clk_r_REG42_S2 ( .D(1'b0), .SI(n473), .SE(n564), .CK(clk), .QN(n511)
         );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2  ( .D(n656), .SI(1'b1), .SE(n431), .CK(clk), 
        .Q(n402), .QN(n463) );
  INV_X1 U2 ( .A(rst_n), .ZN(n656) );
  OR2_X1 U3 ( .A1(n384), .A2(n461), .ZN(n6) );
  CLKBUF_X1 U4 ( .A(n362), .Z(n244) );
  BUF_X2 U5 ( .A(n362), .Z(n7) );
  INV_X1 U6 ( .A(n48), .ZN(n249) );
  OR2_X1 U7 ( .A1(n387), .A2(n465), .ZN(n25) );
  OAI21_X1 U8 ( .B1(n229), .B2(n228), .A(n387), .ZN(n170) );
  NAND2_X1 U9 ( .A1(n10), .A2(n9), .ZN(n224) );
  NAND2_X1 U10 ( .A1(n152), .A2(n151), .ZN(n29) );
  NAND2_X1 U11 ( .A1(n220), .A2(n11), .ZN(n10) );
  NAND2_X1 U12 ( .A1(n13), .A2(n12), .ZN(n11) );
  NAND2_X1 U13 ( .A1(n28), .A2(n27), .ZN(n148) );
  XNOR2_X1 U14 ( .A(n220), .B(n14), .ZN(n229) );
  XNOR2_X1 U15 ( .A(n245), .B(n23), .ZN(n277) );
  NAND2_X1 U16 ( .A1(n222), .A2(n221), .ZN(n9) );
  INV_X1 U17 ( .A(n222), .ZN(n13) );
  XNOR2_X1 U18 ( .A(n222), .B(n221), .ZN(n14) );
  OAI21_X1 U19 ( .B1(n144), .B2(n145), .A(n143), .ZN(n28) );
  NAND2_X1 U20 ( .A1(n145), .A2(n144), .ZN(n27) );
  INV_X1 U21 ( .A(n221), .ZN(n12) );
  CLKBUF_X2 U22 ( .A(rst_n), .Z(n473) );
  XNOR2_X1 U23 ( .A(n247), .B(n246), .ZN(n23) );
  OAI22_X1 U24 ( .A1(n166), .A2(n164), .B1(n249), .B2(n156), .ZN(n211) );
  INV_X1 U25 ( .A(n43), .ZN(n176) );
  CLKBUF_X1 U26 ( .A(\mult_x_1/n310 ), .Z(n41) );
  BUF_X1 U27 ( .A(\mult_x_1/n311 ), .Z(n44) );
  XNOR2_X1 U28 ( .A(n92), .B(n8), .ZN(n88) );
  XNOR2_X1 U29 ( .A(n94), .B(n93), .ZN(n8) );
  INV_X1 U30 ( .A(n15), .ZN(n439) );
  AOI21_X1 U31 ( .B1(n230), .B2(n387), .A(n16), .ZN(n15) );
  NOR2_X1 U32 ( .A1(n382), .A2(n459), .ZN(n16) );
  NAND2_X1 U33 ( .A1(n17), .A2(n6), .ZN(n435) );
  NAND2_X1 U34 ( .A1(n223), .A2(n387), .ZN(n17) );
  NAND2_X1 U35 ( .A1(n19), .A2(n18), .ZN(n240) );
  NAND2_X1 U36 ( .A1(n247), .A2(n246), .ZN(n18) );
  NAND2_X1 U37 ( .A1(n245), .A2(n20), .ZN(n19) );
  NAND2_X1 U38 ( .A1(n22), .A2(n21), .ZN(n20) );
  INV_X1 U39 ( .A(n246), .ZN(n21) );
  INV_X1 U40 ( .A(n247), .ZN(n22) );
  NAND2_X1 U41 ( .A1(n24), .A2(n382), .ZN(n318) );
  XNOR2_X1 U42 ( .A(n317), .B(n316), .ZN(n24) );
  OAI21_X1 U43 ( .B1(n151), .B2(n152), .A(n31), .ZN(n30) );
  NAND2_X1 U44 ( .A1(n30), .A2(n29), .ZN(n199) );
  NAND2_X1 U45 ( .A1(n26), .A2(n25), .ZN(n427) );
  NAND2_X1 U46 ( .A1(n201), .A2(n7), .ZN(n26) );
  BUF_X2 U47 ( .A(n98), .Z(n257) );
  INV_X2 U48 ( .A(n286), .ZN(n382) );
  XNOR2_X1 U49 ( .A(n33), .B(n31), .ZN(n111) );
  XNOR2_X1 U50 ( .A(n32), .B(n143), .ZN(n31) );
  XNOR2_X1 U51 ( .A(n144), .B(n145), .ZN(n32) );
  XNOR2_X1 U52 ( .A(n152), .B(n151), .ZN(n33) );
  OR2_X2 U53 ( .A1(n54), .A2(n53), .ZN(n175) );
  OR2_X2 U54 ( .A1(n47), .A2(n48), .ZN(n166) );
  AND2_X1 U55 ( .A1(n655), .A2(\mult_x_1/n281 ), .ZN(n34) );
  XNOR2_X1 U56 ( .A(\mult_x_1/n312 ), .B(n34), .ZN(n37) );
  OR2_X1 U57 ( .A1(\mult_x_1/n288 ), .A2(n479), .ZN(n262) );
  CLKBUF_X1 U58 ( .A(n179), .Z(n42) );
  NAND2_X1 U59 ( .A1(n203), .A2(n202), .ZN(n69) );
  OAI21_X1 U60 ( .B1(n200), .B2(n199), .A(n7), .ZN(n153) );
  OR2_X1 U61 ( .A1(n277), .A2(n276), .ZN(n35) );
  INV_X1 U62 ( .A(n286), .ZN(n362) );
  AND2_X1 U63 ( .A1(n655), .A2(\mult_x_1/n281 ), .ZN(n36) );
  XOR2_X1 U64 ( .A(\mult_x_1/n312 ), .B(n483), .Z(n77) );
  XNOR2_X1 U65 ( .A(n178), .B(n63), .ZN(n38) );
  INV_X1 U66 ( .A(n51), .ZN(n39) );
  NOR2_X2 U67 ( .A1(n474), .A2(n475), .ZN(n178) );
  XNOR2_X2 U68 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n40) );
  BUF_X2 U69 ( .A(\mult_x_1/n313 ), .Z(n266) );
  INV_X1 U70 ( .A(n55), .ZN(n179) );
  XNOR2_X1 U71 ( .A(n477), .B(\mult_x_1/a[6] ), .ZN(n43) );
  CLKBUF_X1 U72 ( .A(\mult_x_1/n310 ), .Z(n45) );
  XNOR2_X1 U73 ( .A(n205), .B(n204), .ZN(n282) );
  INV_X1 U74 ( .A(n286), .ZN(n391) );
  INV_X1 U75 ( .A(n286), .ZN(n384) );
  INV_X1 U76 ( .A(n286), .ZN(n389) );
  OR2_X1 U77 ( .A1(n94), .A2(n93), .ZN(n46) );
  INV_X1 U78 ( .A(en), .ZN(n286) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/a[4] ), .ZN(n47) );
  XNOR2_X1 U80 ( .A(\mult_x_1/n312 ), .B(n478), .ZN(n48) );
  XNOR2_X1 U81 ( .A(n44), .B(\mult_x_1/n284 ), .ZN(n60) );
  XNOR2_X1 U82 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n283 ), .ZN(n76) );
  OAI22_X1 U83 ( .A1(n60), .A2(n166), .B1(n249), .B2(n76), .ZN(n82) );
  XOR2_X1 U84 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[2] ), .Z(n49) );
  XNOR2_X1 U85 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .ZN(n50) );
  NAND2_X1 U86 ( .A1(n49), .A2(n50), .ZN(n98) );
  INV_X1 U87 ( .A(n479), .ZN(n261) );
  XNOR2_X1 U88 ( .A(n261), .B(\mult_x_1/n282 ), .ZN(n61) );
  OAI22_X1 U89 ( .A1(n98), .A2(n61), .B1(n40), .B2(n77), .ZN(n81) );
  XNOR2_X1 U90 ( .A(n82), .B(n81), .ZN(n74) );
  INV_X1 U91 ( .A(n178), .ZN(n51) );
  OR2_X1 U92 ( .A1(\mult_x_1/n288 ), .A2(n51), .ZN(n52) );
  INV_X1 U93 ( .A(\mult_x_1/n310 ), .ZN(n63) );
  XNOR2_X1 U94 ( .A(n178), .B(n63), .ZN(n55) );
  NOR2_X1 U95 ( .A1(n52), .A2(n42), .ZN(n73) );
  XNOR2_X1 U96 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n53) );
  XNOR2_X1 U97 ( .A(n477), .B(\mult_x_1/a[6] ), .ZN(n54) );
  XNOR2_X1 U98 ( .A(n41), .B(\mult_x_1/n287 ), .ZN(n64) );
  XNOR2_X1 U99 ( .A(n41), .B(\mult_x_1/n286 ), .ZN(n58) );
  OAI22_X1 U100 ( .A1(n175), .A2(n64), .B1(n176), .B2(n58), .ZN(n208) );
  NAND2_X1 U101 ( .A1(n266), .A2(n482), .ZN(n267) );
  XNOR2_X1 U102 ( .A(n266), .B(\mult_x_1/n281 ), .ZN(n157) );
  XNOR2_X1 U103 ( .A(n36), .B(n266), .ZN(n56) );
  OAI22_X1 U104 ( .A1(n267), .A2(n157), .B1(n56), .B2(n482), .ZN(n207) );
  AND2_X1 U105 ( .A1(\mult_x_1/n288 ), .A2(n38), .ZN(n206) );
  AOI21_X1 U106 ( .B1(n267), .B2(n482), .A(n56), .ZN(n57) );
  INV_X1 U107 ( .A(n57), .ZN(n80) );
  XNOR2_X1 U108 ( .A(n41), .B(\mult_x_1/n285 ), .ZN(n75) );
  OAI22_X1 U109 ( .A1(n175), .A2(n58), .B1(n176), .B2(n75), .ZN(n79) );
  XNOR2_X1 U110 ( .A(n178), .B(\mult_x_1/n287 ), .ZN(n59) );
  NOR2_X1 U111 ( .A1(n59), .A2(n179), .ZN(n78) );
  INV_X1 U112 ( .A(n203), .ZN(n67) );
  XNOR2_X1 U113 ( .A(n44), .B(\mult_x_1/n285 ), .ZN(n156) );
  OAI22_X1 U114 ( .A1(n166), .A2(n156), .B1(n249), .B2(n60), .ZN(n214) );
  XNOR2_X1 U115 ( .A(n261), .B(\mult_x_1/n283 ), .ZN(n159) );
  OAI22_X1 U116 ( .A1(n257), .A2(n159), .B1(n40), .B2(n61), .ZN(n213) );
  OR2_X1 U117 ( .A1(\mult_x_1/n288 ), .A2(n63), .ZN(n62) );
  OAI22_X1 U118 ( .A1(n175), .A2(n63), .B1(n62), .B2(n176), .ZN(n155) );
  XNOR2_X1 U119 ( .A(n45), .B(\mult_x_1/n288 ), .ZN(n65) );
  OAI22_X1 U120 ( .A1(n175), .A2(n65), .B1(n176), .B2(n64), .ZN(n154) );
  INV_X1 U121 ( .A(n202), .ZN(n66) );
  NAND2_X1 U122 ( .A1(n67), .A2(n66), .ZN(n68) );
  NAND2_X1 U123 ( .A1(n205), .A2(n68), .ZN(n70) );
  NAND2_X1 U124 ( .A1(n70), .A2(n69), .ZN(n115) );
  INV_X1 U125 ( .A(n115), .ZN(n71) );
  AND2_X1 U126 ( .A1(n7), .A2(n71), .ZN(n85) );
  FA_X1 U127 ( .A(n74), .B(n73), .CI(n72), .CO(n90), .S(n205) );
  XNOR2_X1 U128 ( .A(n41), .B(\mult_x_1/n284 ), .ZN(n97) );
  OAI22_X1 U129 ( .A1(n175), .A2(n75), .B1(n176), .B2(n97), .ZN(n105) );
  XNOR2_X1 U130 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n282 ), .ZN(n102) );
  OAI22_X1 U131 ( .A1(n166), .A2(n76), .B1(n249), .B2(n102), .ZN(n104) );
  XNOR2_X1 U132 ( .A(n36), .B(n261), .ZN(n99) );
  OAI22_X1 U133 ( .A1(n98), .A2(n77), .B1(n37), .B2(n40), .ZN(n141) );
  INV_X1 U134 ( .A(n141), .ZN(n103) );
  FA_X1 U135 ( .A(n80), .B(n79), .CI(n78), .CO(n92), .S(n203) );
  OR2_X1 U136 ( .A1(n82), .A2(n81), .ZN(n94) );
  XNOR2_X1 U137 ( .A(n178), .B(\mult_x_1/n286 ), .ZN(n83) );
  NOR2_X1 U138 ( .A1(n83), .A2(n179), .ZN(n93) );
  INV_X1 U139 ( .A(n116), .ZN(n84) );
  NAND2_X1 U140 ( .A1(n85), .A2(n84), .ZN(n87) );
  OR2_X1 U141 ( .A1(n387), .A2(n456), .ZN(n86) );
  NAND2_X1 U142 ( .A1(n87), .A2(n86), .ZN(n445) );
  FA_X1 U143 ( .A(n90), .B(n89), .CI(n88), .CO(n110), .S(n116) );
  INV_X1 U144 ( .A(n110), .ZN(n91) );
  AND2_X1 U145 ( .A1(n91), .A2(n7), .ZN(n107) );
  NAND2_X1 U146 ( .A1(n92), .A2(n46), .ZN(n96) );
  NAND2_X1 U147 ( .A1(n94), .A2(n93), .ZN(n95) );
  NAND2_X1 U148 ( .A1(n96), .A2(n95), .ZN(n152) );
  XNOR2_X1 U149 ( .A(n45), .B(\mult_x_1/n283 ), .ZN(n126) );
  OAI22_X1 U150 ( .A1(n175), .A2(n97), .B1(n176), .B2(n126), .ZN(n142) );
  AOI21_X1 U151 ( .B1(n40), .B2(n257), .A(n99), .ZN(n100) );
  INV_X1 U152 ( .A(n100), .ZN(n140) );
  XNOR2_X1 U153 ( .A(n39), .B(\mult_x_1/n285 ), .ZN(n101) );
  NOR2_X1 U154 ( .A1(n101), .A2(n179), .ZN(n145) );
  XNOR2_X1 U155 ( .A(n44), .B(\mult_x_1/n281 ), .ZN(n122) );
  OAI22_X1 U156 ( .A1(n166), .A2(n102), .B1(n249), .B2(n122), .ZN(n144) );
  FA_X1 U157 ( .A(n104), .B(n105), .CI(n103), .CO(n143), .S(n89) );
  INV_X1 U158 ( .A(n111), .ZN(n106) );
  NAND2_X1 U159 ( .A1(n107), .A2(n106), .ZN(n109) );
  OR2_X1 U160 ( .A1(n362), .A2(n464), .ZN(n108) );
  NAND2_X1 U161 ( .A1(n109), .A2(n108), .ZN(n429) );
  NAND2_X1 U162 ( .A1(n111), .A2(n110), .ZN(n112) );
  NAND2_X1 U163 ( .A1(n112), .A2(n382), .ZN(n114) );
  OR2_X1 U164 ( .A1(n7), .A2(n463), .ZN(n113) );
  NAND2_X1 U165 ( .A1(n114), .A2(n113), .ZN(n431) );
  NAND2_X1 U166 ( .A1(n116), .A2(n115), .ZN(n117) );
  NAND2_X1 U167 ( .A1(n117), .A2(n391), .ZN(n119) );
  OR2_X1 U168 ( .A1(n7), .A2(n455), .ZN(n118) );
  NAND2_X1 U169 ( .A1(n119), .A2(n118), .ZN(n447) );
  XNOR2_X1 U190 ( .A(n39), .B(\mult_x_1/n282 ), .ZN(n120) );
  NOR2_X1 U191 ( .A1(n120), .A2(n42), .ZN(n173) );
  XNOR2_X1 U192 ( .A(n45), .B(\mult_x_1/n281 ), .ZN(n121) );
  XNOR2_X1 U193 ( .A(n36), .B(n45), .ZN(n174) );
  OAI22_X1 U194 ( .A1(n175), .A2(n121), .B1(n174), .B2(n176), .ZN(n184) );
  INV_X1 U195 ( .A(n184), .ZN(n172) );
  XNOR2_X1 U196 ( .A(n45), .B(\mult_x_1/n282 ), .ZN(n125) );
  OAI22_X1 U197 ( .A1(n175), .A2(n125), .B1(n176), .B2(n121), .ZN(n131) );
  XNOR2_X1 U198 ( .A(\mult_x_1/n311 ), .B(n36), .ZN(n123) );
  OAI22_X1 U199 ( .A1(n122), .A2(n166), .B1(n123), .B2(n249), .ZN(n130) );
  AOI21_X1 U200 ( .B1(n166), .B2(n249), .A(n123), .ZN(n124) );
  INV_X1 U201 ( .A(n124), .ZN(n129) );
  INV_X1 U202 ( .A(n130), .ZN(n139) );
  OAI22_X1 U203 ( .A1(n175), .A2(n126), .B1(n176), .B2(n125), .ZN(n138) );
  XNOR2_X1 U204 ( .A(n178), .B(\mult_x_1/n284 ), .ZN(n127) );
  NOR2_X1 U205 ( .A1(n127), .A2(n179), .ZN(n137) );
  XNOR2_X1 U206 ( .A(n39), .B(\mult_x_1/n283 ), .ZN(n128) );
  NOR2_X1 U207 ( .A1(n128), .A2(n42), .ZN(n135) );
  FA_X1 U208 ( .A(n131), .B(n129), .CI(n130), .CO(n171), .S(n134) );
  OR2_X1 U209 ( .A1(n192), .A2(n191), .ZN(n132) );
  NAND2_X1 U210 ( .A1(n387), .A2(n132), .ZN(n133) );
  OAI21_X1 U211 ( .B1(n362), .B2(n472), .A(n133), .ZN(n413) );
  FA_X1 U212 ( .A(n136), .B(n135), .CI(n134), .CO(n191), .S(n196) );
  FA_X1 U213 ( .A(n139), .B(n138), .CI(n137), .CO(n136), .S(n150) );
  FA_X1 U214 ( .A(n142), .B(n141), .CI(n140), .CO(n149), .S(n151) );
  OR2_X1 U215 ( .A1(n196), .A2(n195), .ZN(n146) );
  NAND2_X1 U216 ( .A1(n387), .A2(n146), .ZN(n147) );
  OAI21_X1 U217 ( .B1(n244), .B2(n471), .A(n147), .ZN(n415) );
  FA_X1 U218 ( .A(n150), .B(n149), .CI(n148), .CO(n195), .S(n200) );
  OAI21_X1 U219 ( .B1(n384), .B2(n470), .A(n153), .ZN(n417) );
  XNOR2_X1 U220 ( .A(n266), .B(\mult_x_1/n283 ), .ZN(n235) );
  XNOR2_X1 U221 ( .A(n266), .B(\mult_x_1/n282 ), .ZN(n158) );
  OAI22_X1 U222 ( .A1(n267), .A2(n235), .B1(n158), .B2(n482), .ZN(n169) );
  AND2_X1 U223 ( .A1(\mult_x_1/n288 ), .A2(n54), .ZN(n168) );
  XNOR2_X1 U224 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n234) );
  XNOR2_X1 U225 ( .A(n261), .B(\mult_x_1/n284 ), .ZN(n160) );
  OAI22_X1 U226 ( .A1(n257), .A2(n234), .B1(n40), .B2(n160), .ZN(n167) );
  HA_X1 U227 ( .A(n155), .B(n154), .CO(n212), .S(n221) );
  XNOR2_X1 U228 ( .A(n44), .B(\mult_x_1/n286 ), .ZN(n164) );
  OAI22_X1 U229 ( .A1(n267), .A2(n158), .B1(n157), .B2(n482), .ZN(n210) );
  OAI22_X1 U230 ( .A1(n257), .A2(n160), .B1(n50), .B2(n159), .ZN(n209) );
  INV_X1 U231 ( .A(\mult_x_1/n311 ), .ZN(n162) );
  OR2_X1 U232 ( .A1(\mult_x_1/n288 ), .A2(n162), .ZN(n161) );
  OAI22_X1 U233 ( .A1(n166), .A2(n162), .B1(n161), .B2(n249), .ZN(n237) );
  XNOR2_X1 U234 ( .A(n44), .B(\mult_x_1/n288 ), .ZN(n163) );
  XNOR2_X1 U235 ( .A(\mult_x_1/n311 ), .B(\mult_x_1/n287 ), .ZN(n165) );
  OAI22_X1 U236 ( .A1(n163), .A2(n166), .B1(n249), .B2(n165), .ZN(n236) );
  OAI22_X1 U237 ( .A1(n166), .A2(n165), .B1(n249), .B2(n164), .ZN(n232) );
  FA_X1 U238 ( .A(n169), .B(n168), .CI(n167), .CO(n222), .S(n231) );
  OAI21_X1 U239 ( .B1(n389), .B2(n469), .A(n170), .ZN(n419) );
  FA_X1 U240 ( .A(n173), .B(n172), .CI(n171), .CO(n186), .S(n192) );
  AOI21_X1 U241 ( .B1(n176), .B2(n175), .A(n174), .ZN(n177) );
  INV_X1 U242 ( .A(n177), .ZN(n182) );
  XNOR2_X1 U243 ( .A(n39), .B(\mult_x_1/n281 ), .ZN(n180) );
  NOR2_X1 U244 ( .A1(n180), .A2(n42), .ZN(n181) );
  XOR2_X1 U245 ( .A(n182), .B(n181), .Z(n183) );
  XOR2_X1 U246 ( .A(n184), .B(n183), .Z(n185) );
  OR2_X1 U247 ( .A1(n186), .A2(n185), .ZN(n188) );
  NAND2_X1 U248 ( .A1(n186), .A2(n185), .ZN(n187) );
  NAND2_X1 U249 ( .A1(n188), .A2(n187), .ZN(n189) );
  NAND2_X1 U250 ( .A1(n7), .A2(n189), .ZN(n190) );
  OAI21_X1 U251 ( .B1(n7), .B2(n468), .A(n190), .ZN(n421) );
  NAND2_X1 U252 ( .A1(n192), .A2(n191), .ZN(n193) );
  NAND2_X1 U253 ( .A1(n244), .A2(n193), .ZN(n194) );
  OAI21_X1 U254 ( .B1(n7), .B2(n467), .A(n194), .ZN(n423) );
  NAND2_X1 U255 ( .A1(n196), .A2(n195), .ZN(n197) );
  NAND2_X1 U256 ( .A1(n387), .A2(n197), .ZN(n198) );
  OAI21_X1 U257 ( .B1(n384), .B2(n466), .A(n198), .ZN(n425) );
  NAND2_X1 U258 ( .A1(n200), .A2(n199), .ZN(n201) );
  XNOR2_X1 U259 ( .A(n203), .B(n202), .ZN(n204) );
  FA_X1 U260 ( .A(n208), .B(n206), .CI(n207), .CO(n72), .S(n219) );
  FA_X1 U261 ( .A(n209), .B(n210), .CI(n211), .CO(n218), .S(n220) );
  FA_X1 U262 ( .A(n212), .B(n213), .CI(n214), .CO(n202), .S(n217) );
  NAND2_X1 U263 ( .A1(n282), .A2(n281), .ZN(n215) );
  NAND2_X1 U264 ( .A1(n382), .A2(n215), .ZN(n216) );
  OAI21_X1 U265 ( .B1(n389), .B2(n462), .A(n216), .ZN(n433) );
  FA_X1 U266 ( .A(n219), .B(n218), .CI(n217), .CO(n281), .S(n225) );
  NOR2_X1 U267 ( .A1(n225), .A2(n224), .ZN(n223) );
  NAND2_X1 U268 ( .A1(n225), .A2(n224), .ZN(n226) );
  NAND2_X1 U269 ( .A1(n244), .A2(n226), .ZN(n227) );
  OAI21_X1 U270 ( .B1(n382), .B2(n460), .A(n227), .ZN(n437) );
  NAND2_X1 U271 ( .A1(n229), .A2(n228), .ZN(n230) );
  FA_X1 U272 ( .A(n233), .B(n232), .CI(n231), .CO(n228), .S(n241) );
  XNOR2_X1 U273 ( .A(n261), .B(\mult_x_1/n286 ), .ZN(n251) );
  OAI22_X1 U274 ( .A1(n257), .A2(n251), .B1(n40), .B2(n234), .ZN(n247) );
  XNOR2_X1 U275 ( .A(n266), .B(\mult_x_1/n284 ), .ZN(n248) );
  OAI22_X1 U276 ( .A1(n267), .A2(n248), .B1(n235), .B2(n482), .ZN(n246) );
  HA_X1 U277 ( .A(n236), .B(n237), .CO(n233), .S(n245) );
  NOR2_X1 U278 ( .A1(n241), .A2(n240), .ZN(n238) );
  NAND2_X1 U279 ( .A1(n244), .A2(n238), .ZN(n239) );
  OAI21_X1 U280 ( .B1(n244), .B2(n458), .A(n239), .ZN(n441) );
  NAND2_X1 U281 ( .A1(n241), .A2(n240), .ZN(n242) );
  NAND2_X1 U282 ( .A1(n244), .A2(n242), .ZN(n243) );
  OAI21_X1 U283 ( .B1(n382), .B2(n457), .A(n243), .ZN(n443) );
  XNOR2_X1 U284 ( .A(n266), .B(\mult_x_1/n285 ), .ZN(n258) );
  OAI22_X1 U285 ( .A1(n267), .A2(n258), .B1(n248), .B2(n482), .ZN(n254) );
  INV_X1 U286 ( .A(n249), .ZN(n250) );
  AND2_X1 U287 ( .A1(\mult_x_1/n288 ), .A2(n250), .ZN(n253) );
  XNOR2_X1 U288 ( .A(n261), .B(\mult_x_1/n287 ), .ZN(n255) );
  OAI22_X1 U289 ( .A1(n257), .A2(n255), .B1(n40), .B2(n251), .ZN(n252) );
  OR2_X1 U290 ( .A1(n277), .A2(n276), .ZN(n315) );
  FA_X1 U291 ( .A(n254), .B(n253), .CI(n252), .CO(n276), .S(n275) );
  XNOR2_X1 U292 ( .A(n261), .B(\mult_x_1/n288 ), .ZN(n256) );
  OAI22_X1 U293 ( .A1(n257), .A2(n256), .B1(n40), .B2(n255), .ZN(n260) );
  XNOR2_X1 U294 ( .A(n266), .B(\mult_x_1/n286 ), .ZN(n263) );
  OAI22_X1 U295 ( .A1(n267), .A2(n263), .B1(n258), .B2(n482), .ZN(n259) );
  NOR2_X1 U296 ( .A1(n275), .A2(n274), .ZN(n307) );
  HA_X1 U297 ( .A(n260), .B(n259), .CO(n274), .S(n272) );
  OAI22_X1 U298 ( .A1(n257), .A2(n479), .B1(n262), .B2(n40), .ZN(n271) );
  OR2_X1 U299 ( .A1(n272), .A2(n271), .ZN(n302) );
  XNOR2_X1 U300 ( .A(n266), .B(\mult_x_1/n287 ), .ZN(n265) );
  OAI22_X1 U301 ( .A1(n267), .A2(n265), .B1(n263), .B2(n482), .ZN(n270) );
  INV_X1 U302 ( .A(n50), .ZN(n264) );
  AND2_X1 U303 ( .A1(\mult_x_1/n288 ), .A2(n264), .ZN(n269) );
  NOR2_X1 U304 ( .A1(n270), .A2(n269), .ZN(n294) );
  OAI22_X1 U305 ( .A1(n267), .A2(\mult_x_1/n288 ), .B1(n265), .B2(n482), .ZN(
        n290) );
  OR2_X1 U306 ( .A1(\mult_x_1/n288 ), .A2(n481), .ZN(n268) );
  NAND2_X1 U307 ( .A1(n268), .A2(n267), .ZN(n289) );
  NAND2_X1 U308 ( .A1(n290), .A2(n289), .ZN(n297) );
  NAND2_X1 U309 ( .A1(n270), .A2(n269), .ZN(n295) );
  OAI21_X1 U310 ( .B1(n294), .B2(n297), .A(n295), .ZN(n303) );
  NAND2_X1 U311 ( .A1(n272), .A2(n271), .ZN(n301) );
  INV_X1 U312 ( .A(n301), .ZN(n273) );
  AOI21_X1 U313 ( .B1(n302), .B2(n303), .A(n273), .ZN(n310) );
  NAND2_X1 U314 ( .A1(n275), .A2(n274), .ZN(n308) );
  OAI21_X1 U315 ( .B1(n307), .B2(n310), .A(n308), .ZN(n316) );
  NAND2_X1 U316 ( .A1(n277), .A2(n276), .ZN(n314) );
  INV_X1 U317 ( .A(n314), .ZN(n278) );
  AOI21_X1 U318 ( .B1(n315), .B2(n316), .A(n278), .ZN(n279) );
  NAND2_X1 U319 ( .A1(n391), .A2(n279), .ZN(n280) );
  OAI21_X1 U320 ( .B1(n7), .B2(n453), .A(n280), .ZN(n451) );
  OR2_X1 U321 ( .A1(n387), .A2(n454), .ZN(n285) );
  NOR2_X1 U322 ( .A1(n282), .A2(n281), .ZN(n283) );
  NAND2_X1 U323 ( .A1(n389), .A2(n283), .ZN(n284) );
  NAND2_X1 U324 ( .A1(n285), .A2(n284), .ZN(n449) );
  BUF_X2 U325 ( .A(n286), .Z(n392) );
  AOI22_X1 U326 ( .A1(n362), .A2(n527), .B1(n528), .B2(n392), .ZN(n530) );
  AOI22_X1 U327 ( .A1(n362), .A2(n526), .B1(n527), .B2(n392), .ZN(n532) );
  INV_X1 U328 ( .A(n286), .ZN(n387) );
  AND2_X1 U329 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n287) );
  NAND2_X1 U330 ( .A1(n387), .A2(n287), .ZN(n288) );
  OAI21_X1 U331 ( .B1(n391), .B2(n526), .A(n288), .ZN(n534) );
  AOI22_X1 U332 ( .A1(n387), .A2(n524), .B1(n525), .B2(n392), .ZN(n536) );
  AOI22_X1 U333 ( .A1(n391), .A2(n523), .B1(n524), .B2(n392), .ZN(n538) );
  OR2_X1 U334 ( .A1(n290), .A2(n289), .ZN(n291) );
  AND2_X1 U335 ( .A1(n291), .A2(n297), .ZN(n292) );
  NAND2_X1 U336 ( .A1(n387), .A2(n292), .ZN(n293) );
  OAI21_X1 U337 ( .B1(n389), .B2(n523), .A(n293), .ZN(n540) );
  AOI22_X1 U338 ( .A1(n387), .A2(n521), .B1(n522), .B2(n392), .ZN(n542) );
  AOI22_X1 U339 ( .A1(n387), .A2(n520), .B1(n521), .B2(n392), .ZN(n544) );
  INV_X1 U340 ( .A(n294), .ZN(n296) );
  NAND2_X1 U341 ( .A1(n296), .A2(n295), .ZN(n298) );
  XOR2_X1 U342 ( .A(n298), .B(n297), .Z(n299) );
  NAND2_X1 U343 ( .A1(n382), .A2(n299), .ZN(n300) );
  OAI21_X1 U344 ( .B1(n389), .B2(n520), .A(n300), .ZN(n546) );
  AOI22_X1 U345 ( .A1(n391), .A2(n518), .B1(n519), .B2(n392), .ZN(n548) );
  AOI22_X1 U346 ( .A1(n387), .A2(n517), .B1(n518), .B2(n392), .ZN(n550) );
  NAND2_X1 U347 ( .A1(n302), .A2(n301), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  NAND2_X1 U349 ( .A1(n382), .A2(n305), .ZN(n306) );
  OAI21_X1 U350 ( .B1(n384), .B2(n517), .A(n306), .ZN(n552) );
  AOI22_X1 U351 ( .A1(n244), .A2(n515), .B1(n516), .B2(n392), .ZN(n554) );
  AOI22_X1 U352 ( .A1(n384), .A2(n514), .B1(n515), .B2(n392), .ZN(n556) );
  INV_X1 U353 ( .A(n307), .ZN(n309) );
  NAND2_X1 U354 ( .A1(n309), .A2(n308), .ZN(n311) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n312) );
  NAND2_X1 U356 ( .A1(n382), .A2(n312), .ZN(n313) );
  OAI21_X1 U357 ( .B1(n389), .B2(n514), .A(n313), .ZN(n558) );
  AOI22_X1 U358 ( .A1(n391), .A2(n512), .B1(n513), .B2(n392), .ZN(n560) );
  AOI22_X1 U359 ( .A1(n391), .A2(n511), .B1(n512), .B2(n392), .ZN(n562) );
  NAND2_X1 U360 ( .A1(n35), .A2(n314), .ZN(n317) );
  OAI21_X1 U361 ( .B1(n389), .B2(n511), .A(n318), .ZN(n564) );
  AOI22_X1 U362 ( .A1(n391), .A2(n509), .B1(n510), .B2(n392), .ZN(n566) );
  NAND2_X1 U363 ( .A1(n458), .A2(n408), .ZN(n319) );
  XOR2_X1 U364 ( .A(n319), .B(n412), .Z(n320) );
  NAND2_X1 U365 ( .A1(n382), .A2(n320), .ZN(n321) );
  OAI21_X1 U366 ( .B1(n384), .B2(n509), .A(n321), .ZN(n568) );
  AOI22_X1 U367 ( .A1(n391), .A2(n507), .B1(n508), .B2(n392), .ZN(n570) );
  OAI21_X1 U368 ( .B1(n407), .B2(n412), .A(n408), .ZN(n325) );
  NAND2_X1 U369 ( .A1(n396), .A2(n406), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n325), .B(n322), .ZN(n323) );
  NAND2_X1 U371 ( .A1(n382), .A2(n323), .ZN(n324) );
  OAI21_X1 U372 ( .B1(n389), .B2(n507), .A(n324), .ZN(n572) );
  AOI22_X1 U373 ( .A1(n391), .A2(n505), .B1(n506), .B2(n392), .ZN(n574) );
  AOI21_X1 U374 ( .B1(n325), .B2(n396), .A(n459), .ZN(n329) );
  NAND2_X1 U375 ( .A1(n461), .A2(n405), .ZN(n326) );
  XOR2_X1 U376 ( .A(n329), .B(n326), .Z(n327) );
  NAND2_X1 U377 ( .A1(n389), .A2(n327), .ZN(n328) );
  OAI21_X1 U378 ( .B1(n389), .B2(n505), .A(n328), .ZN(n576) );
  AOI22_X1 U379 ( .A1(n391), .A2(n503), .B1(n504), .B2(n392), .ZN(n578) );
  OAI21_X1 U380 ( .B1(n329), .B2(n404), .A(n405), .ZN(n339) );
  INV_X1 U381 ( .A(n339), .ZN(n333) );
  NAND2_X1 U382 ( .A1(n454), .A2(n403), .ZN(n330) );
  XOR2_X1 U383 ( .A(n333), .B(n330), .Z(n331) );
  NAND2_X1 U384 ( .A1(n389), .A2(n331), .ZN(n332) );
  OAI21_X1 U385 ( .B1(n389), .B2(n503), .A(n332), .ZN(n580) );
  AOI22_X1 U386 ( .A1(n391), .A2(n501), .B1(n502), .B2(n392), .ZN(n582) );
  OAI21_X1 U387 ( .B1(n333), .B2(n411), .A(n403), .ZN(n335) );
  NAND2_X1 U388 ( .A1(n456), .A2(n410), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n336) );
  NAND2_X1 U390 ( .A1(n389), .A2(n336), .ZN(n337) );
  OAI21_X1 U391 ( .B1(n384), .B2(n501), .A(n337), .ZN(n584) );
  AOI22_X1 U392 ( .A1(n391), .A2(n499), .B1(n500), .B2(n392), .ZN(n586) );
  NOR2_X1 U393 ( .A1(n409), .A2(n411), .ZN(n340) );
  OAI21_X1 U394 ( .B1(n409), .B2(n403), .A(n410), .ZN(n338) );
  AOI21_X1 U395 ( .B1(n340), .B2(n339), .A(n338), .ZN(n367) );
  NAND2_X1 U396 ( .A1(n464), .A2(n402), .ZN(n341) );
  XOR2_X1 U397 ( .A(n367), .B(n341), .Z(n342) );
  NAND2_X1 U398 ( .A1(n389), .A2(n342), .ZN(n343) );
  OAI21_X1 U399 ( .B1(n384), .B2(n499), .A(n343), .ZN(n588) );
  AOI22_X1 U400 ( .A1(n387), .A2(n497), .B1(n498), .B2(n392), .ZN(n590) );
  OAI21_X1 U401 ( .B1(n367), .B2(n401), .A(n402), .ZN(n345) );
  NAND2_X1 U402 ( .A1(n395), .A2(n400), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U404 ( .A1(n389), .A2(n346), .ZN(n347) );
  OAI21_X1 U405 ( .B1(n384), .B2(n497), .A(n347), .ZN(n592) );
  AOI22_X1 U406 ( .A1(n391), .A2(n495), .B1(n496), .B2(n392), .ZN(n594) );
  NAND2_X1 U407 ( .A1(n464), .A2(n395), .ZN(n349) );
  AOI21_X1 U408 ( .B1(n463), .B2(n395), .A(n465), .ZN(n348) );
  OAI21_X1 U409 ( .B1(n367), .B2(n349), .A(n348), .ZN(n351) );
  NAND2_X1 U410 ( .A1(n394), .A2(n399), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  NAND2_X1 U412 ( .A1(n389), .A2(n352), .ZN(n353) );
  OAI21_X1 U413 ( .B1(n384), .B2(n495), .A(n353), .ZN(n596) );
  AOI22_X1 U414 ( .A1(n7), .A2(n493), .B1(n494), .B2(n392), .ZN(n598) );
  NAND2_X1 U415 ( .A1(n395), .A2(n394), .ZN(n355) );
  NOR2_X1 U416 ( .A1(n401), .A2(n355), .ZN(n363) );
  INV_X1 U417 ( .A(n363), .ZN(n357) );
  AOI21_X1 U418 ( .B1(n465), .B2(n394), .A(n466), .ZN(n354) );
  OAI21_X1 U419 ( .B1(n355), .B2(n402), .A(n354), .ZN(n364) );
  INV_X1 U420 ( .A(n364), .ZN(n356) );
  OAI21_X1 U421 ( .B1(n367), .B2(n357), .A(n356), .ZN(n359) );
  NAND2_X1 U422 ( .A1(n393), .A2(n398), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  NAND2_X1 U424 ( .A1(n389), .A2(n360), .ZN(n361) );
  OAI21_X1 U425 ( .B1(n384), .B2(n493), .A(n361), .ZN(n600) );
  AOI22_X1 U426 ( .A1(n7), .A2(n491), .B1(n492), .B2(n392), .ZN(n602) );
  NAND2_X1 U427 ( .A1(n363), .A2(n393), .ZN(n366) );
  AOI21_X1 U428 ( .B1(n364), .B2(n393), .A(n467), .ZN(n365) );
  OAI21_X1 U429 ( .B1(n367), .B2(n366), .A(n365), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n368), .B(n397), .ZN(n369) );
  NAND2_X1 U431 ( .A1(n389), .A2(n369), .ZN(n370) );
  OAI21_X1 U432 ( .B1(n384), .B2(n491), .A(n370), .ZN(n604) );
  NAND2_X1 U433 ( .A1(n382), .A2(B_extended[0]), .ZN(n371) );
  OAI21_X1 U434 ( .B1(n384), .B2(n490), .A(n371), .ZN(n606) );
  NAND2_X1 U435 ( .A1(n389), .A2(B_extended[1]), .ZN(n372) );
  OAI21_X1 U436 ( .B1(n384), .B2(n489), .A(n372), .ZN(n608) );
  NAND2_X1 U437 ( .A1(n382), .A2(B_extended[2]), .ZN(n373) );
  OAI21_X1 U438 ( .B1(n384), .B2(n488), .A(n373), .ZN(n610) );
  NAND2_X1 U439 ( .A1(n382), .A2(B_extended[3]), .ZN(n374) );
  OAI21_X1 U440 ( .B1(n384), .B2(n487), .A(n374), .ZN(n612) );
  NAND2_X1 U441 ( .A1(n382), .A2(B_extended[4]), .ZN(n375) );
  OAI21_X1 U442 ( .B1(n384), .B2(n486), .A(n375), .ZN(n614) );
  NAND2_X1 U443 ( .A1(n382), .A2(B_extended[5]), .ZN(n376) );
  OAI21_X1 U444 ( .B1(n384), .B2(n485), .A(n376), .ZN(n616) );
  NAND2_X1 U445 ( .A1(n382), .A2(B_extended[6]), .ZN(n377) );
  OAI21_X1 U446 ( .B1(n384), .B2(n484), .A(n377), .ZN(n618) );
  NAND2_X1 U447 ( .A1(n382), .A2(B_extended[7]), .ZN(n378) );
  OAI21_X1 U448 ( .B1(n391), .B2(n483), .A(n378), .ZN(n620) );
  NAND2_X1 U449 ( .A1(n382), .A2(A_extended[0]), .ZN(n379) );
  OAI21_X1 U450 ( .B1(n391), .B2(n482), .A(n379), .ZN(n622) );
  NAND2_X1 U451 ( .A1(n382), .A2(A_extended[1]), .ZN(n380) );
  OAI21_X1 U452 ( .B1(n391), .B2(n481), .A(n380), .ZN(n624) );
  NAND2_X1 U453 ( .A1(n382), .A2(A_extended[2]), .ZN(n381) );
  OAI21_X1 U454 ( .B1(n384), .B2(n480), .A(n381), .ZN(n626) );
  NAND2_X1 U455 ( .A1(n382), .A2(A_extended[3]), .ZN(n383) );
  OAI21_X1 U456 ( .B1(n384), .B2(n479), .A(n383), .ZN(n628) );
  NAND2_X1 U457 ( .A1(n387), .A2(A_extended[4]), .ZN(n385) );
  OAI21_X1 U458 ( .B1(n391), .B2(n478), .A(n385), .ZN(n630) );
  NAND2_X1 U459 ( .A1(n387), .A2(A_extended[5]), .ZN(n386) );
  OAI21_X1 U460 ( .B1(n391), .B2(n477), .A(n386), .ZN(n632) );
  NAND2_X1 U461 ( .A1(n387), .A2(A_extended[6]), .ZN(n388) );
  OAI21_X1 U462 ( .B1(n391), .B2(n476), .A(n388), .ZN(n634) );
  NAND2_X1 U463 ( .A1(n389), .A2(A_extended[7]), .ZN(n390) );
  OAI21_X1 U464 ( .B1(n391), .B2(n475), .A(n390), .ZN(n636) );
  NAND2_X1 U465 ( .A1(n474), .A2(n392), .ZN(n638) );
endmodule


module conv_128_32_DW_mult_pipe_J1_30 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/a[2] , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 ,
         \mult_x_1/n287 , \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 ,
         \mult_x_1/n283 , \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 ,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n400,
         n402, n404, n406, n408, n410, n412, n414, n416, n418, n420, n422,
         n424, n426, n428, n430, n432, n434, n436, n438, n440, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n523, n525, n527, n529, n531, n533, n535, n537, n539, n541,
         n543, n545, n547, n549, n551, n553, n555, n557, n559, n561, n563,
         n565, n567, n569, n571, n573, n575, n577, n579, n581, n583, n585,
         n587, n589, n591, n593, n595, n597, n599, n601, n603, n605, n607,
         n609, n611, n613, n615, n617, n619, n621, n623, n625, n627, n629,
         n646, n647;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n467), .SE(n629), .CK(clk), .Q(n646), 
        .QN(n468) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n467), .SE(n625), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n470) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n467), .SE(n621), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n472) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n467), .SE(n617), .CK(clk), .Q(
        \mult_x_1/a[2] ), .QN(n474) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n467), .SE(n613), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n476) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n467), .SE(n611), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n477) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n467), .SE(n609), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n478) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n465), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n479) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n466), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n480) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n464), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n481) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n467), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n482) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n464), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n483) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n464), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n484) );
  SDFF_X1 clk_r_REG10_S3 ( .D(1'b0), .SI(n464), .SE(n595), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG11_S4 ( .D(1'b0), .SI(n464), .SE(n593), .CK(clk), .Q(
        product[15]), .QN(n486) );
  SDFF_X1 clk_r_REG12_S3 ( .D(1'b0), .SI(n464), .SE(n591), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG13_S4 ( .D(1'b0), .SI(n464), .SE(n589), .CK(clk), .Q(
        product[14]), .QN(n488) );
  SDFF_X1 clk_r_REG14_S3 ( .D(1'b0), .SI(n464), .SE(n587), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG15_S4 ( .D(1'b0), .SI(n466), .SE(n585), .CK(clk), .Q(
        product[13]), .QN(n490) );
  SDFF_X1 clk_r_REG16_S3 ( .D(1'b0), .SI(n467), .SE(n583), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG17_S4 ( .D(1'b0), .SI(n465), .SE(n581), .CK(clk), .Q(
        product[12]), .QN(n492) );
  SDFF_X1 clk_r_REG8_S3 ( .D(1'b0), .SI(n464), .SE(n579), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG9_S4 ( .D(1'b0), .SI(n464), .SE(n577), .CK(clk), .Q(
        product[11]), .QN(n494) );
  SDFF_X1 clk_r_REG4_S3 ( .D(1'b0), .SI(n464), .SE(n575), .CK(clk), .QN(n495)
         );
  SDFF_X1 clk_r_REG5_S4 ( .D(1'b0), .SI(n464), .SE(n573), .CK(clk), .Q(
        product[10]), .QN(n496) );
  SDFF_X1 clk_r_REG6_S3 ( .D(1'b0), .SI(n464), .SE(n571), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG7_S4 ( .D(1'b0), .SI(n464), .SE(n569), .CK(clk), .Q(
        product[9]), .QN(n498) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n464), .SE(n567), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n466), .SE(n565), .CK(clk), .Q(
        product[8]), .QN(n500) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n466), .SE(n563), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n466), .SE(n561), .CK(clk), .Q(
        product[7]), .QN(n502) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n466), .SE(n559), .CK(clk), .QN(n503)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n466), .SE(n557), .CK(clk), .Q(
        product[6]), .QN(n504) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n466), .SE(n555), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n466), .SE(n553), .CK(clk), .Q(
        product[5]), .QN(n506) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n466), .SE(n551), .CK(clk), .QN(n507)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n466), .SE(n549), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n466), .SE(n547), .CK(clk), .Q(
        product[4]), .QN(n509) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n466), .SE(n545), .CK(clk), .QN(n510)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n465), .SE(n543), .CK(clk), .QN(n511)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n465), .SE(n541), .CK(clk), .Q(
        product[3]), .QN(n512) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n465), .SE(n539), .CK(clk), .QN(n513)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n465), .SE(n537), .CK(clk), .QN(n514)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n465), .SE(n535), .CK(clk), .Q(
        product[2]), .QN(n515) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n465), .SE(n533), .CK(clk), .QN(n516)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n465), .SE(n531), .CK(clk), .QN(n517)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n465), .SE(n529), .CK(clk), .Q(
        product[1]), .QN(n518) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n465), .SE(n527), .CK(clk), .QN(n519)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n465), .SE(n525), .CK(clk), .QN(n520)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n465), .SE(n523), .CK(clk), .Q(
        product[0]), .QN(n521) );
  SDFF_X2 clk_r_REG0_S1 ( .D(1'b0), .SI(n467), .SE(n627), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n469) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n467), .SE(n615), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n475) );
  SDFF_X1 \mult_x_1/clk_r_REG19_S2  ( .D(n647), .SI(1'b1), .SE(n412), .CK(clk), 
        .Q(n383), .QN(n456) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n647), .SE(n440), .CK(
        clk), .Q(n442), .QN(n397) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2  ( .D(n647), .SI(1'b1), .SE(n438), .CK(clk), 
        .Q(n396), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n647), .SE(n436), .CK(
        clk), .Q(n444), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n647), .SI(1'b1), .SE(n434), .CK(clk), 
        .Q(n394), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG20_S2  ( .D(n647), .SI(1'b1), .SE(n432), .CK(clk), 
        .Q(n393), .QN(n446) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n647), .SI(1'b1), .SE(n430), .CK(clk), 
        .Q(n392), .QN(n447) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2_IP  ( .D(1'b1), .SI(n647), .SE(n428), .CK(
        clk), .Q(n448), .QN(n391) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n647), .SE(n426), .CK(
        clk), .Q(n449), .QN(n390) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n647), .SI(1'b1), .SE(n424), .CK(clk), 
        .Q(n389), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n647), .SI(1'b1), .SE(n422), .CK(clk), 
        .Q(n388), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n647), .SI(1'b1), .SE(n420), .CK(clk), 
        .Q(n387), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n647), .SI(1'b1), .SE(n418), .CK(clk), 
        .Q(n386), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2  ( .D(n647), .SI(1'b1), .SE(n416), .CK(clk), 
        .Q(n385), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG18_S2  ( .D(n647), .SI(1'b1), .SE(n414), .CK(clk), 
        .Q(n384), .QN(n455) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n647), .SI(1'b1), .SE(n410), .CK(clk), 
        .Q(n382), .QN(n457) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n647), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n381), .QN(n458) );
  SDFF_X1 \mult_x_1/clk_r_REG29_S2  ( .D(n647), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n380), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2_IP  ( .D(1'b1), .SI(n647), .SE(n404), .CK(
        clk), .Q(n460), .QN(n379) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n647), .SI(1'b1), .SE(n402), .CK(clk), 
        .Q(n378), .QN(n461) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n647), .SE(n400), .CK(
        clk), .Q(n462), .QN(n377) );
  SDFF_X1 \mult_x_1/clk_r_REG30_S2  ( .D(n647), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n376), .QN(n463) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n467), .SE(n619), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n473) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n467), .SE(n623), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n471) );
  INV_X1 U2 ( .A(rst_n), .ZN(n647) );
  INV_X1 U3 ( .A(n647), .ZN(n464) );
  CLKBUF_X1 U4 ( .A(n464), .Z(n467) );
  CLKBUF_X1 U5 ( .A(n464), .Z(n465) );
  CLKBUF_X1 U6 ( .A(n464), .Z(n466) );
  INV_X1 U7 ( .A(n33), .ZN(n239) );
  OR2_X1 U8 ( .A1(n263), .A2(n461), .ZN(n13) );
  NAND2_X1 U9 ( .A1(n15), .A2(n14), .ZN(n187) );
  OAI21_X1 U10 ( .B1(n162), .B2(n163), .A(n16), .ZN(n15) );
  NAND2_X1 U11 ( .A1(n163), .A2(n162), .ZN(n14) );
  XNOR2_X1 U12 ( .A(n51), .B(n12), .ZN(n259) );
  XNOR2_X1 U13 ( .A(n53), .B(n52), .ZN(n12) );
  NAND2_X1 U14 ( .A1(n25), .A2(n24), .ZN(n156) );
  INV_X1 U15 ( .A(n28), .ZN(n174) );
  BUF_X1 U16 ( .A(\mult_x_1/n311 ), .Z(n152) );
  CLKBUF_X2 U17 ( .A(\mult_x_1/n313 ), .Z(n241) );
  OAI22_X1 U18 ( .A1(n302), .A2(n5), .B1(n374), .B2(n469), .ZN(n627) );
  INV_X1 U19 ( .A(A_extended[7]), .ZN(n5) );
  NAND2_X1 U20 ( .A1(n20), .A2(n6), .ZN(n438) );
  NAND2_X1 U21 ( .A1(n262), .A2(n269), .ZN(n6) );
  NAND2_X1 U22 ( .A1(n8), .A2(n7), .ZN(n164) );
  NAND2_X1 U23 ( .A1(n53), .A2(n52), .ZN(n7) );
  NAND2_X1 U24 ( .A1(n51), .A2(n9), .ZN(n8) );
  NAND2_X1 U25 ( .A1(n11), .A2(n10), .ZN(n9) );
  INV_X1 U26 ( .A(n52), .ZN(n10) );
  INV_X1 U27 ( .A(n53), .ZN(n11) );
  NAND2_X1 U28 ( .A1(n168), .A2(n13), .ZN(n402) );
  XNOR2_X1 U29 ( .A(n17), .B(n16), .ZN(n192) );
  XNOR2_X1 U30 ( .A(n144), .B(n145), .ZN(n16) );
  XNOR2_X1 U31 ( .A(n163), .B(n162), .ZN(n17) );
  INV_X1 U32 ( .A(n118), .ZN(n115) );
  AND2_X1 U33 ( .A1(\mult_x_1/n310 ), .A2(n646), .ZN(n29) );
  NAND2_X1 U34 ( .A1(n92), .A2(n91), .ZN(n93) );
  NAND2_X1 U35 ( .A1(n47), .A2(n46), .ZN(n261) );
  INV_X1 U36 ( .A(n110), .ZN(n44) );
  INV_X1 U37 ( .A(n141), .ZN(n145) );
  NAND2_X1 U38 ( .A1(n120), .A2(n119), .ZN(n128) );
  XNOR2_X1 U39 ( .A(n66), .B(n89), .ZN(n99) );
  XNOR2_X1 U40 ( .A(n92), .B(n91), .ZN(n66) );
  OAI21_X1 U41 ( .B1(n264), .B2(n447), .A(n54), .ZN(n430) );
  NAND2_X1 U42 ( .A1(n32), .A2(n31), .ZN(n18) );
  NAND2_X1 U43 ( .A1(n32), .A2(n31), .ZN(n19) );
  NAND2_X1 U44 ( .A1(n32), .A2(n31), .ZN(n237) );
  OR2_X1 U45 ( .A1(n264), .A2(n443), .ZN(n20) );
  BUF_X2 U46 ( .A(n375), .Z(n337) );
  INV_X2 U47 ( .A(n337), .ZN(n370) );
  INV_X2 U48 ( .A(n337), .ZN(n374) );
  INV_X1 U49 ( .A(n473), .ZN(n235) );
  XOR2_X1 U50 ( .A(n106), .B(n105), .Z(n21) );
  AND2_X1 U51 ( .A1(n105), .A2(n106), .ZN(n22) );
  XNOR2_X1 U52 ( .A(\mult_x_1/n311 ), .B(n470), .ZN(n28) );
  INV_X1 U53 ( .A(en), .ZN(n375) );
  INV_X2 U54 ( .A(n375), .ZN(n348) );
  BUF_X2 U55 ( .A(n348), .Z(n264) );
  XNOR2_X1 U56 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/a[4] ), .ZN(n24) );
  INV_X1 U57 ( .A(n24), .ZN(n23) );
  INV_X2 U58 ( .A(n23), .ZN(n220) );
  AND2_X1 U59 ( .A1(n646), .A2(\mult_x_1/n281 ), .ZN(n132) );
  XNOR2_X1 U60 ( .A(n132), .B(n152), .ZN(n133) );
  XNOR2_X1 U61 ( .A(n152), .B(\mult_x_1/n281 ), .ZN(n36) );
  XOR2_X1 U62 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n25) );
  OAI22_X1 U63 ( .A1(n220), .A2(n133), .B1(n36), .B2(n156), .ZN(n26) );
  INV_X1 U64 ( .A(n26), .ZN(n141) );
  XNOR2_X1 U65 ( .A(\mult_x_1/a[6] ), .B(\mult_x_1/n310 ), .ZN(n27) );
  OR2_X2 U66 ( .A1(n27), .A2(n28), .ZN(n173) );
  XNOR2_X1 U67 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n30) );
  XNOR2_X1 U68 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n136) );
  OAI22_X1 U69 ( .A1(n173), .A2(n30), .B1(n174), .B2(n136), .ZN(n140) );
  XNOR2_X1 U70 ( .A(n29), .B(n469), .ZN(n57) );
  INV_X1 U71 ( .A(n57), .ZN(n176) );
  NOR2_X1 U72 ( .A1(n480), .A2(n176), .ZN(n139) );
  XNOR2_X1 U73 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n37) );
  OAI22_X1 U74 ( .A1(n173), .A2(n37), .B1(n174), .B2(n30), .ZN(n50) );
  XOR2_X1 U75 ( .A(\mult_x_1/a[2] ), .B(\mult_x_1/n313 ), .Z(n33) );
  INV_X1 U76 ( .A(n33), .ZN(n32) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n312 ), .B(n474), .ZN(n31) );
  XNOR2_X1 U78 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n42) );
  XNOR2_X1 U79 ( .A(n132), .B(\mult_x_1/n312 ), .ZN(n34) );
  OAI22_X1 U80 ( .A1(n237), .A2(n42), .B1(n34), .B2(n239), .ZN(n49) );
  AOI21_X1 U81 ( .B1(n239), .B2(n18), .A(n34), .ZN(n35) );
  INV_X1 U82 ( .A(n35), .ZN(n48) );
  NOR2_X1 U83 ( .A1(n481), .A2(n176), .ZN(n53) );
  XNOR2_X1 U84 ( .A(n152), .B(\mult_x_1/n282 ), .ZN(n38) );
  OAI22_X1 U85 ( .A1(n156), .A2(n38), .B1(n220), .B2(n36), .ZN(n52) );
  XNOR2_X1 U86 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n40) );
  OAI22_X1 U87 ( .A1(n173), .A2(n40), .B1(n174), .B2(n37), .ZN(n109) );
  XNOR2_X1 U88 ( .A(n152), .B(\mult_x_1/n283 ), .ZN(n41) );
  OAI22_X1 U89 ( .A1(n156), .A2(n41), .B1(n220), .B2(n38), .ZN(n108) );
  INV_X1 U90 ( .A(n49), .ZN(n107) );
  NAND2_X1 U91 ( .A1(n241), .A2(n476), .ZN(n242) );
  XNOR2_X1 U92 ( .A(n132), .B(n241), .ZN(n56) );
  AOI21_X1 U93 ( .B1(n242), .B2(n476), .A(n56), .ZN(n39) );
  INV_X1 U94 ( .A(n39), .ZN(n97) );
  XNOR2_X1 U95 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n55) );
  OAI22_X1 U96 ( .A1(n173), .A2(n55), .B1(n174), .B2(n40), .ZN(n96) );
  NOR2_X1 U97 ( .A1(n483), .A2(n176), .ZN(n95) );
  XNOR2_X1 U98 ( .A(n152), .B(\mult_x_1/n284 ), .ZN(n59) );
  OAI22_X1 U99 ( .A1(n156), .A2(n59), .B1(n220), .B2(n41), .ZN(n83) );
  XNOR2_X1 U100 ( .A(n235), .B(\mult_x_1/n282 ), .ZN(n61) );
  OAI22_X1 U101 ( .A1(n18), .A2(n61), .B1(n239), .B2(n42), .ZN(n82) );
  OR2_X1 U102 ( .A1(n83), .A2(n82), .ZN(n110) );
  NOR2_X1 U103 ( .A1(n482), .A2(n176), .ZN(n111) );
  INV_X1 U104 ( .A(n111), .ZN(n43) );
  NAND2_X1 U105 ( .A1(n44), .A2(n43), .ZN(n45) );
  NAND2_X1 U106 ( .A1(n113), .A2(n45), .ZN(n47) );
  NAND2_X1 U107 ( .A1(n110), .A2(n111), .ZN(n46) );
  FA_X1 U108 ( .A(n50), .B(n49), .CI(n48), .CO(n165), .S(n260) );
  BUF_X2 U109 ( .A(n348), .Z(n255) );
  OAI21_X1 U110 ( .B1(n78), .B2(n77), .A(n255), .ZN(n54) );
  XNOR2_X1 U111 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n63) );
  OAI22_X1 U112 ( .A1(n173), .A2(n63), .B1(n174), .B2(n55), .ZN(n86) );
  XNOR2_X1 U113 ( .A(n241), .B(\mult_x_1/n281 ), .ZN(n58) );
  OAI22_X1 U114 ( .A1(n242), .A2(n58), .B1(n56), .B2(n476), .ZN(n85) );
  AND2_X1 U115 ( .A1(\mult_x_1/n288 ), .A2(n57), .ZN(n84) );
  XNOR2_X1 U116 ( .A(n152), .B(\mult_x_1/n286 ), .ZN(n154) );
  XNOR2_X1 U117 ( .A(n152), .B(\mult_x_1/n285 ), .ZN(n60) );
  OAI22_X1 U118 ( .A1(n156), .A2(n154), .B1(n220), .B2(n60), .ZN(n73) );
  XNOR2_X1 U119 ( .A(n241), .B(\mult_x_1/n282 ), .ZN(n67) );
  OAI22_X1 U120 ( .A1(n242), .A2(n67), .B1(n58), .B2(n476), .ZN(n72) );
  XNOR2_X1 U121 ( .A(n235), .B(\mult_x_1/n284 ), .ZN(n68) );
  XNOR2_X1 U122 ( .A(n235), .B(\mult_x_1/n283 ), .ZN(n62) );
  OAI22_X1 U123 ( .A1(n18), .A2(n68), .B1(n239), .B2(n62), .ZN(n71) );
  OAI22_X1 U124 ( .A1(n156), .A2(n60), .B1(n220), .B2(n59), .ZN(n92) );
  OAI22_X1 U125 ( .A1(n237), .A2(n62), .B1(n239), .B2(n61), .ZN(n91) );
  XNOR2_X1 U126 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n64) );
  OAI22_X1 U127 ( .A1(n173), .A2(n64), .B1(n174), .B2(n63), .ZN(n70) );
  OR2_X1 U128 ( .A1(\mult_x_1/n288 ), .A2(n469), .ZN(n65) );
  OAI22_X1 U129 ( .A1(n173), .A2(n469), .B1(n65), .B2(n174), .ZN(n69) );
  AND2_X1 U130 ( .A1(n70), .A2(n69), .ZN(n89) );
  XNOR2_X1 U131 ( .A(n241), .B(\mult_x_1/n283 ), .ZN(n207) );
  OAI22_X1 U132 ( .A1(n242), .A2(n207), .B1(n67), .B2(n476), .ZN(n159) );
  AND2_X1 U133 ( .A1(\mult_x_1/n288 ), .A2(n28), .ZN(n158) );
  XNOR2_X1 U134 ( .A(n235), .B(\mult_x_1/n285 ), .ZN(n206) );
  OAI22_X1 U135 ( .A1(n19), .A2(n206), .B1(n239), .B2(n68), .ZN(n157) );
  XOR2_X1 U136 ( .A(n70), .B(n69), .Z(n149) );
  FA_X1 U137 ( .A(n73), .B(n72), .CI(n71), .CO(n100), .S(n148) );
  NAND2_X1 U138 ( .A1(n196), .A2(n195), .ZN(n74) );
  NAND2_X1 U139 ( .A1(n269), .A2(n74), .ZN(n76) );
  BUF_X2 U140 ( .A(n348), .Z(n263) );
  OR2_X1 U141 ( .A1(n255), .A2(n454), .ZN(n75) );
  NAND2_X1 U142 ( .A1(n76), .A2(n75), .ZN(n416) );
  NAND2_X1 U143 ( .A1(n78), .A2(n77), .ZN(n79) );
  NAND2_X1 U144 ( .A1(n79), .A2(n263), .ZN(n81) );
  BUF_X2 U145 ( .A(n348), .Z(n269) );
  OR2_X1 U146 ( .A1(n255), .A2(n457), .ZN(n80) );
  NAND2_X1 U147 ( .A1(n81), .A2(n80), .ZN(n410) );
  XNOR2_X1 U148 ( .A(n83), .B(n82), .ZN(n106) );
  FA_X1 U149 ( .A(n86), .B(n85), .CI(n84), .CO(n105), .S(n101) );
  INV_X1 U150 ( .A(n92), .ZN(n88) );
  INV_X1 U151 ( .A(n91), .ZN(n87) );
  NAND2_X1 U152 ( .A1(n88), .A2(n87), .ZN(n90) );
  NAND2_X1 U153 ( .A1(n90), .A2(n89), .ZN(n94) );
  NAND2_X1 U154 ( .A1(n94), .A2(n93), .ZN(n118) );
  FA_X1 U155 ( .A(n97), .B(n96), .CI(n95), .CO(n113), .S(n117) );
  XNOR2_X1 U156 ( .A(n118), .B(n117), .ZN(n98) );
  XNOR2_X1 U157 ( .A(n21), .B(n98), .ZN(n127) );
  FA_X1 U158 ( .A(n101), .B(n100), .CI(n99), .CO(n124), .S(n196) );
  NAND2_X1 U159 ( .A1(n127), .A2(n124), .ZN(n102) );
  NAND2_X1 U160 ( .A1(n102), .A2(n264), .ZN(n104) );
  OR2_X1 U161 ( .A1(n255), .A2(n446), .ZN(n103) );
  NAND2_X1 U162 ( .A1(n104), .A2(n103), .ZN(n432) );
  FA_X1 U163 ( .A(n108), .B(n109), .CI(n107), .CO(n51), .S(n266) );
  XNOR2_X1 U164 ( .A(n111), .B(n110), .ZN(n112) );
  XNOR2_X1 U165 ( .A(n113), .B(n112), .ZN(n265) );
  INV_X1 U166 ( .A(n117), .ZN(n114) );
  NAND2_X1 U167 ( .A1(n115), .A2(n114), .ZN(n116) );
  NAND2_X1 U168 ( .A1(n21), .A2(n116), .ZN(n120) );
  NAND2_X1 U169 ( .A1(n118), .A2(n117), .ZN(n119) );
  NAND2_X1 U170 ( .A1(n131), .A2(n128), .ZN(n121) );
  NAND2_X1 U171 ( .A1(n121), .A2(n264), .ZN(n123) );
  OR2_X1 U172 ( .A1(n255), .A2(n448), .ZN(n122) );
  NAND2_X1 U173 ( .A1(n123), .A2(n122), .ZN(n428) );
  INV_X1 U174 ( .A(n124), .ZN(n125) );
  NAND2_X1 U175 ( .A1(n255), .A2(n125), .ZN(n126) );
  OAI22_X1 U176 ( .A1(n127), .A2(n126), .B1(n263), .B2(n456), .ZN(n412) );
  INV_X1 U177 ( .A(n128), .ZN(n129) );
  NAND2_X1 U178 ( .A1(n255), .A2(n129), .ZN(n130) );
  OAI22_X1 U179 ( .A1(n131), .A2(n130), .B1(n264), .B2(n449), .ZN(n426) );
  NOR2_X1 U202 ( .A1(n478), .A2(n176), .ZN(n171) );
  XNOR2_X1 U203 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n135) );
  XNOR2_X1 U204 ( .A(n132), .B(\mult_x_1/n310 ), .ZN(n172) );
  OAI22_X1 U205 ( .A1(n173), .A2(n135), .B1(n172), .B2(n174), .ZN(n180) );
  INV_X1 U206 ( .A(n180), .ZN(n170) );
  AOI21_X1 U207 ( .B1(n220), .B2(n156), .A(n133), .ZN(n134) );
  INV_X1 U208 ( .A(n134), .ZN(n143) );
  OAI22_X1 U209 ( .A1(n173), .A2(n136), .B1(n174), .B2(n135), .ZN(n142) );
  NOR2_X1 U210 ( .A1(n143), .A2(n142), .ZN(n138) );
  NAND2_X1 U211 ( .A1(n143), .A2(n142), .ZN(n137) );
  OAI21_X1 U212 ( .B1(n138), .B2(n141), .A(n137), .ZN(n169) );
  FA_X1 U213 ( .A(n141), .B(n140), .CI(n139), .CO(n163), .S(n166) );
  NOR2_X1 U214 ( .A1(n479), .A2(n176), .ZN(n162) );
  XNOR2_X1 U215 ( .A(n143), .B(n142), .ZN(n144) );
  OR2_X1 U216 ( .A1(n188), .A2(n187), .ZN(n146) );
  NAND2_X1 U217 ( .A1(n255), .A2(n146), .ZN(n147) );
  OAI21_X1 U218 ( .B1(n263), .B2(n463), .A(n147), .ZN(n398) );
  FA_X1 U219 ( .A(n150), .B(n149), .CI(n148), .CO(n195), .S(n200) );
  OR2_X1 U220 ( .A1(\mult_x_1/n288 ), .A2(n471), .ZN(n151) );
  OAI22_X1 U221 ( .A1(n156), .A2(n471), .B1(n151), .B2(n220), .ZN(n209) );
  XNOR2_X1 U222 ( .A(n152), .B(\mult_x_1/n288 ), .ZN(n153) );
  XNOR2_X1 U223 ( .A(n152), .B(\mult_x_1/n287 ), .ZN(n155) );
  OAI22_X1 U224 ( .A1(n156), .A2(n153), .B1(n220), .B2(n155), .ZN(n208) );
  OAI22_X1 U225 ( .A1(n156), .A2(n155), .B1(n220), .B2(n154), .ZN(n204) );
  FA_X1 U226 ( .A(n159), .B(n158), .CI(n157), .CO(n150), .S(n203) );
  OR2_X1 U227 ( .A1(n200), .A2(n199), .ZN(n160) );
  NAND2_X1 U228 ( .A1(n269), .A2(n160), .ZN(n161) );
  OAI21_X1 U229 ( .B1(n263), .B2(n462), .A(n161), .ZN(n400) );
  FA_X1 U230 ( .A(n166), .B(n165), .CI(n164), .CO(n191), .S(n78) );
  OR2_X1 U231 ( .A1(n192), .A2(n191), .ZN(n167) );
  NAND2_X1 U232 ( .A1(n263), .A2(n167), .ZN(n168) );
  FA_X1 U233 ( .A(n171), .B(n170), .CI(n169), .CO(n182), .S(n188) );
  AOI21_X1 U234 ( .B1(n174), .B2(n173), .A(n172), .ZN(n175) );
  INV_X1 U235 ( .A(n175), .ZN(n178) );
  NOR2_X1 U236 ( .A1(n477), .A2(n176), .ZN(n177) );
  XOR2_X1 U237 ( .A(n178), .B(n177), .Z(n179) );
  XOR2_X1 U238 ( .A(n180), .B(n179), .Z(n181) );
  OR2_X1 U239 ( .A1(n182), .A2(n181), .ZN(n184) );
  NAND2_X1 U240 ( .A1(n182), .A2(n181), .ZN(n183) );
  NAND2_X1 U241 ( .A1(n184), .A2(n183), .ZN(n185) );
  NAND2_X1 U242 ( .A1(n264), .A2(n185), .ZN(n186) );
  OAI21_X1 U243 ( .B1(n269), .B2(n460), .A(n186), .ZN(n404) );
  NAND2_X1 U244 ( .A1(n188), .A2(n187), .ZN(n189) );
  NAND2_X1 U245 ( .A1(n264), .A2(n189), .ZN(n190) );
  OAI21_X1 U246 ( .B1(n269), .B2(n459), .A(n190), .ZN(n406) );
  NAND2_X1 U247 ( .A1(n192), .A2(n191), .ZN(n193) );
  NAND2_X1 U248 ( .A1(n264), .A2(n193), .ZN(n194) );
  OAI21_X1 U249 ( .B1(n269), .B2(n458), .A(n194), .ZN(n408) );
  NOR2_X1 U250 ( .A1(n196), .A2(n195), .ZN(n197) );
  NAND2_X1 U251 ( .A1(n264), .A2(n197), .ZN(n198) );
  OAI21_X1 U252 ( .B1(n264), .B2(n455), .A(n198), .ZN(n414) );
  NAND2_X1 U253 ( .A1(n200), .A2(n199), .ZN(n201) );
  NAND2_X1 U254 ( .A1(n264), .A2(n201), .ZN(n202) );
  OAI21_X1 U255 ( .B1(n263), .B2(n453), .A(n202), .ZN(n418) );
  FA_X1 U256 ( .A(n205), .B(n204), .CI(n203), .CO(n199), .S(n213) );
  XNOR2_X1 U257 ( .A(n235), .B(\mult_x_1/n286 ), .ZN(n222) );
  OAI22_X1 U258 ( .A1(n19), .A2(n222), .B1(n239), .B2(n206), .ZN(n218) );
  XNOR2_X1 U259 ( .A(n241), .B(\mult_x_1/n284 ), .ZN(n219) );
  OAI22_X1 U260 ( .A1(n242), .A2(n219), .B1(n207), .B2(n476), .ZN(n217) );
  HA_X1 U261 ( .A(n209), .B(n208), .CO(n205), .S(n216) );
  NOR2_X1 U262 ( .A1(n213), .A2(n212), .ZN(n210) );
  NAND2_X1 U263 ( .A1(n263), .A2(n210), .ZN(n211) );
  OAI21_X1 U264 ( .B1(n263), .B2(n452), .A(n211), .ZN(n420) );
  NAND2_X1 U265 ( .A1(n213), .A2(n212), .ZN(n214) );
  NAND2_X1 U266 ( .A1(n269), .A2(n214), .ZN(n215) );
  OAI21_X1 U267 ( .B1(n263), .B2(n451), .A(n215), .ZN(n422) );
  FA_X1 U268 ( .A(n218), .B(n217), .CI(n216), .CO(n212), .S(n224) );
  XNOR2_X1 U269 ( .A(n241), .B(\mult_x_1/n285 ), .ZN(n232) );
  OAI22_X1 U270 ( .A1(n242), .A2(n232), .B1(n219), .B2(n476), .ZN(n229) );
  INV_X1 U271 ( .A(n220), .ZN(n221) );
  AND2_X1 U272 ( .A1(\mult_x_1/n288 ), .A2(n221), .ZN(n228) );
  XNOR2_X1 U273 ( .A(n235), .B(\mult_x_1/n287 ), .ZN(n230) );
  OAI22_X1 U274 ( .A1(n19), .A2(n230), .B1(n239), .B2(n222), .ZN(n227) );
  OR2_X1 U275 ( .A1(n224), .A2(n223), .ZN(n253) );
  NAND2_X1 U276 ( .A1(n224), .A2(n223), .ZN(n251) );
  NAND2_X1 U277 ( .A1(n253), .A2(n251), .ZN(n225) );
  NAND2_X1 U278 ( .A1(n255), .A2(n225), .ZN(n226) );
  OAI21_X1 U279 ( .B1(n269), .B2(n450), .A(n226), .ZN(n424) );
  FA_X1 U280 ( .A(n229), .B(n228), .CI(n227), .CO(n223), .S(n250) );
  XNOR2_X1 U281 ( .A(n235), .B(\mult_x_1/n288 ), .ZN(n231) );
  OAI22_X1 U282 ( .A1(n19), .A2(n231), .B1(n239), .B2(n230), .ZN(n234) );
  XNOR2_X1 U283 ( .A(n241), .B(\mult_x_1/n286 ), .ZN(n238) );
  OAI22_X1 U284 ( .A1(n242), .A2(n238), .B1(n232), .B2(n476), .ZN(n233) );
  NOR2_X1 U285 ( .A1(n250), .A2(n249), .ZN(n290) );
  HA_X1 U286 ( .A(n234), .B(n233), .CO(n249), .S(n247) );
  OR2_X1 U287 ( .A1(\mult_x_1/n288 ), .A2(n473), .ZN(n236) );
  OAI22_X1 U288 ( .A1(n18), .A2(n473), .B1(n236), .B2(n239), .ZN(n246) );
  OR2_X1 U289 ( .A1(n247), .A2(n246), .ZN(n285) );
  XNOR2_X1 U290 ( .A(n241), .B(\mult_x_1/n287 ), .ZN(n240) );
  OAI22_X1 U291 ( .A1(n242), .A2(n240), .B1(n238), .B2(n476), .ZN(n245) );
  AND2_X1 U292 ( .A1(\mult_x_1/n288 ), .A2(n33), .ZN(n244) );
  NOR2_X1 U293 ( .A1(n245), .A2(n244), .ZN(n277) );
  OAI22_X1 U294 ( .A1(n242), .A2(\mult_x_1/n288 ), .B1(n240), .B2(n476), .ZN(
        n273) );
  OR2_X1 U295 ( .A1(\mult_x_1/n288 ), .A2(n475), .ZN(n243) );
  NAND2_X1 U296 ( .A1(n243), .A2(n242), .ZN(n272) );
  NAND2_X1 U297 ( .A1(n273), .A2(n272), .ZN(n280) );
  NAND2_X1 U298 ( .A1(n245), .A2(n244), .ZN(n278) );
  OAI21_X1 U299 ( .B1(n277), .B2(n280), .A(n278), .ZN(n286) );
  NAND2_X1 U300 ( .A1(n247), .A2(n246), .ZN(n284) );
  INV_X1 U301 ( .A(n284), .ZN(n248) );
  AOI21_X1 U302 ( .B1(n285), .B2(n286), .A(n248), .ZN(n293) );
  NAND2_X1 U303 ( .A1(n250), .A2(n249), .ZN(n291) );
  OAI21_X1 U304 ( .B1(n290), .B2(n293), .A(n291), .ZN(n257) );
  INV_X1 U305 ( .A(n251), .ZN(n252) );
  AOI21_X1 U306 ( .B1(n253), .B2(n257), .A(n252), .ZN(n254) );
  NAND2_X1 U307 ( .A1(n263), .A2(n254), .ZN(n256) );
  OAI21_X1 U308 ( .B1(n269), .B2(n445), .A(n256), .ZN(n434) );
  NAND2_X1 U309 ( .A1(n269), .A2(n257), .ZN(n258) );
  OAI21_X1 U310 ( .B1(n269), .B2(n444), .A(n258), .ZN(n436) );
  FA_X1 U311 ( .A(n261), .B(n260), .CI(n259), .CO(n77), .S(n262) );
  FA_X1 U312 ( .A(n22), .B(n266), .CI(n265), .CO(n267), .S(n131) );
  NAND2_X1 U313 ( .A1(n255), .A2(n267), .ZN(n268) );
  OAI21_X1 U314 ( .B1(n264), .B2(n442), .A(n268), .ZN(n440) );
  INV_X1 U315 ( .A(en), .ZN(n302) );
  AOI22_X1 U316 ( .A1(n348), .A2(n520), .B1(n521), .B2(n302), .ZN(n523) );
  AOI22_X1 U317 ( .A1(n348), .A2(n519), .B1(n520), .B2(n302), .ZN(n525) );
  AND2_X1 U318 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n270) );
  NAND2_X1 U319 ( .A1(n373), .A2(n270), .ZN(n271) );
  OAI21_X1 U320 ( .B1(n374), .B2(n519), .A(n271), .ZN(n527) );
  AOI22_X1 U321 ( .A1(n348), .A2(n517), .B1(n518), .B2(n302), .ZN(n529) );
  AOI22_X1 U322 ( .A1(n348), .A2(n516), .B1(n517), .B2(n302), .ZN(n531) );
  INV_X2 U323 ( .A(n337), .ZN(n373) );
  OR2_X1 U324 ( .A1(n273), .A2(n272), .ZN(n274) );
  AND2_X1 U325 ( .A1(n274), .A2(n280), .ZN(n275) );
  NAND2_X1 U326 ( .A1(n373), .A2(n275), .ZN(n276) );
  OAI21_X1 U327 ( .B1(n370), .B2(n516), .A(n276), .ZN(n533) );
  AOI22_X1 U328 ( .A1(n348), .A2(n514), .B1(n515), .B2(n302), .ZN(n535) );
  AOI22_X1 U329 ( .A1(n348), .A2(n513), .B1(n514), .B2(n302), .ZN(n537) );
  INV_X1 U330 ( .A(n277), .ZN(n279) );
  NAND2_X1 U331 ( .A1(n279), .A2(n278), .ZN(n281) );
  XOR2_X1 U332 ( .A(n281), .B(n280), .Z(n282) );
  NAND2_X1 U333 ( .A1(n370), .A2(n282), .ZN(n283) );
  OAI21_X1 U334 ( .B1(n374), .B2(n513), .A(n283), .ZN(n539) );
  AOI22_X1 U335 ( .A1(n348), .A2(n511), .B1(n512), .B2(n302), .ZN(n541) );
  AOI22_X1 U336 ( .A1(n348), .A2(n510), .B1(n511), .B2(n302), .ZN(n543) );
  NAND2_X1 U337 ( .A1(n285), .A2(n284), .ZN(n287) );
  XNOR2_X1 U338 ( .A(n287), .B(n286), .ZN(n288) );
  NAND2_X1 U339 ( .A1(n373), .A2(n288), .ZN(n289) );
  OAI21_X1 U340 ( .B1(n370), .B2(n510), .A(n289), .ZN(n545) );
  AOI22_X1 U341 ( .A1(n348), .A2(n508), .B1(n509), .B2(n302), .ZN(n547) );
  AOI22_X1 U342 ( .A1(n348), .A2(n507), .B1(n508), .B2(n302), .ZN(n549) );
  INV_X1 U343 ( .A(n290), .ZN(n292) );
  NAND2_X1 U344 ( .A1(n292), .A2(n291), .ZN(n294) );
  XOR2_X1 U345 ( .A(n294), .B(n293), .Z(n295) );
  NAND2_X1 U346 ( .A1(n374), .A2(n295), .ZN(n296) );
  OAI21_X1 U347 ( .B1(n374), .B2(n507), .A(n296), .ZN(n551) );
  AOI22_X1 U348 ( .A1(n348), .A2(n505), .B1(n506), .B2(n302), .ZN(n553) );
  XNOR2_X1 U349 ( .A(n389), .B(n395), .ZN(n297) );
  NAND2_X1 U350 ( .A1(n269), .A2(n297), .ZN(n298) );
  OAI21_X1 U351 ( .B1(n374), .B2(n505), .A(n298), .ZN(n555) );
  AOI22_X1 U352 ( .A1(n374), .A2(n503), .B1(n504), .B2(n302), .ZN(n557) );
  NAND2_X1 U353 ( .A1(n452), .A2(n388), .ZN(n299) );
  XOR2_X1 U354 ( .A(n299), .B(n394), .Z(n300) );
  NAND2_X1 U355 ( .A1(n370), .A2(n300), .ZN(n301) );
  OAI21_X1 U356 ( .B1(n370), .B2(n503), .A(n301), .ZN(n559) );
  AOI22_X1 U357 ( .A1(n374), .A2(n501), .B1(n502), .B2(n302), .ZN(n561) );
  OAI21_X1 U358 ( .B1(n387), .B2(n394), .A(n388), .ZN(n306) );
  NAND2_X1 U359 ( .A1(n377), .A2(n386), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n306), .B(n303), .ZN(n304) );
  NAND2_X1 U361 ( .A1(n263), .A2(n304), .ZN(n305) );
  OAI21_X1 U362 ( .B1(n374), .B2(n501), .A(n305), .ZN(n563) );
  AOI22_X1 U363 ( .A1(n374), .A2(n499), .B1(n500), .B2(n337), .ZN(n565) );
  AOI21_X1 U364 ( .B1(n306), .B2(n377), .A(n453), .ZN(n310) );
  NAND2_X1 U365 ( .A1(n455), .A2(n385), .ZN(n307) );
  XOR2_X1 U366 ( .A(n310), .B(n307), .Z(n308) );
  NAND2_X1 U367 ( .A1(n373), .A2(n308), .ZN(n309) );
  OAI21_X1 U368 ( .B1(n374), .B2(n499), .A(n309), .ZN(n567) );
  AOI22_X1 U369 ( .A1(n374), .A2(n497), .B1(n498), .B2(n337), .ZN(n569) );
  OAI21_X1 U370 ( .B1(n310), .B2(n384), .A(n385), .ZN(n320) );
  INV_X1 U371 ( .A(n320), .ZN(n314) );
  NAND2_X1 U372 ( .A1(n456), .A2(n393), .ZN(n311) );
  XOR2_X1 U373 ( .A(n314), .B(n311), .Z(n312) );
  NAND2_X1 U374 ( .A1(n373), .A2(n312), .ZN(n313) );
  OAI21_X1 U375 ( .B1(n370), .B2(n497), .A(n313), .ZN(n571) );
  AOI22_X1 U376 ( .A1(n374), .A2(n495), .B1(n496), .B2(n337), .ZN(n573) );
  OAI21_X1 U377 ( .B1(n314), .B2(n383), .A(n393), .ZN(n316) );
  NAND2_X1 U378 ( .A1(n449), .A2(n391), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n316), .B(n315), .ZN(n317) );
  NAND2_X1 U380 ( .A1(n373), .A2(n317), .ZN(n318) );
  OAI21_X1 U381 ( .B1(n370), .B2(n495), .A(n318), .ZN(n575) );
  AOI22_X1 U382 ( .A1(n374), .A2(n493), .B1(n494), .B2(n337), .ZN(n577) );
  NOR2_X1 U383 ( .A1(n390), .A2(n383), .ZN(n321) );
  OAI21_X1 U384 ( .B1(n390), .B2(n393), .A(n391), .ZN(n319) );
  AOI21_X1 U385 ( .B1(n321), .B2(n320), .A(n319), .ZN(n353) );
  NOR2_X1 U386 ( .A1(n396), .A2(n397), .ZN(n338) );
  INV_X1 U387 ( .A(n338), .ZN(n329) );
  NAND2_X1 U388 ( .A1(n396), .A2(n397), .ZN(n340) );
  NAND2_X1 U389 ( .A1(n329), .A2(n340), .ZN(n322) );
  XOR2_X1 U390 ( .A(n353), .B(n322), .Z(n323) );
  NAND2_X1 U391 ( .A1(n373), .A2(n323), .ZN(n324) );
  OAI21_X1 U392 ( .B1(n370), .B2(n493), .A(n324), .ZN(n579) );
  AOI22_X1 U393 ( .A1(n348), .A2(n491), .B1(n492), .B2(n337), .ZN(n581) );
  OAI21_X1 U394 ( .B1(n353), .B2(n338), .A(n340), .ZN(n326) );
  NAND2_X1 U395 ( .A1(n392), .A2(n382), .ZN(n325) );
  XNOR2_X1 U396 ( .A(n326), .B(n325), .ZN(n327) );
  NAND2_X1 U397 ( .A1(n373), .A2(n327), .ZN(n328) );
  OAI21_X1 U398 ( .B1(n370), .B2(n491), .A(n328), .ZN(n583) );
  AOI22_X1 U399 ( .A1(n374), .A2(n489), .B1(n490), .B2(n337), .ZN(n585) );
  NAND2_X1 U400 ( .A1(n329), .A2(n392), .ZN(n332) );
  INV_X1 U401 ( .A(n340), .ZN(n330) );
  AOI21_X1 U402 ( .B1(n330), .B2(n392), .A(n457), .ZN(n331) );
  OAI21_X1 U403 ( .B1(n353), .B2(n332), .A(n331), .ZN(n334) );
  NAND2_X1 U404 ( .A1(n378), .A2(n381), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n334), .B(n333), .ZN(n335) );
  NAND2_X1 U406 ( .A1(n373), .A2(n335), .ZN(n336) );
  OAI21_X1 U407 ( .B1(n370), .B2(n489), .A(n336), .ZN(n587) );
  AOI22_X1 U408 ( .A1(n348), .A2(n487), .B1(n488), .B2(n337), .ZN(n589) );
  NAND2_X1 U409 ( .A1(n392), .A2(n378), .ZN(n341) );
  NOR2_X1 U410 ( .A1(n338), .A2(n341), .ZN(n349) );
  INV_X1 U411 ( .A(n349), .ZN(n343) );
  AOI21_X1 U412 ( .B1(n457), .B2(n378), .A(n458), .ZN(n339) );
  OAI21_X1 U413 ( .B1(n341), .B2(n340), .A(n339), .ZN(n350) );
  INV_X1 U414 ( .A(n350), .ZN(n342) );
  OAI21_X1 U415 ( .B1(n353), .B2(n343), .A(n342), .ZN(n345) );
  NAND2_X1 U416 ( .A1(n376), .A2(n380), .ZN(n344) );
  XNOR2_X1 U417 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U418 ( .A1(n373), .A2(n346), .ZN(n347) );
  OAI21_X1 U419 ( .B1(n370), .B2(n487), .A(n347), .ZN(n591) );
  AOI22_X1 U420 ( .A1(n348), .A2(n485), .B1(n486), .B2(n375), .ZN(n593) );
  NAND2_X1 U421 ( .A1(n349), .A2(n376), .ZN(n352) );
  AOI21_X1 U422 ( .B1(n350), .B2(n376), .A(n459), .ZN(n351) );
  OAI21_X1 U423 ( .B1(n353), .B2(n352), .A(n351), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n354), .B(n379), .ZN(n355) );
  NAND2_X1 U425 ( .A1(n373), .A2(n355), .ZN(n356) );
  OAI21_X1 U426 ( .B1(n370), .B2(n485), .A(n356), .ZN(n595) );
  NAND2_X1 U427 ( .A1(n373), .A2(B_extended[0]), .ZN(n357) );
  OAI21_X1 U428 ( .B1(n370), .B2(n484), .A(n357), .ZN(n597) );
  NAND2_X1 U429 ( .A1(n373), .A2(B_extended[1]), .ZN(n358) );
  OAI21_X1 U430 ( .B1(n370), .B2(n483), .A(n358), .ZN(n599) );
  NAND2_X1 U431 ( .A1(n373), .A2(B_extended[2]), .ZN(n359) );
  OAI21_X1 U432 ( .B1(n370), .B2(n482), .A(n359), .ZN(n601) );
  NAND2_X1 U433 ( .A1(n370), .A2(B_extended[3]), .ZN(n360) );
  OAI21_X1 U434 ( .B1(n370), .B2(n481), .A(n360), .ZN(n603) );
  NAND2_X1 U435 ( .A1(n373), .A2(B_extended[4]), .ZN(n361) );
  OAI21_X1 U436 ( .B1(n370), .B2(n480), .A(n361), .ZN(n605) );
  NAND2_X1 U437 ( .A1(n263), .A2(B_extended[5]), .ZN(n362) );
  OAI21_X1 U438 ( .B1(n370), .B2(n479), .A(n362), .ZN(n607) );
  NAND2_X1 U439 ( .A1(n373), .A2(B_extended[6]), .ZN(n363) );
  OAI21_X1 U440 ( .B1(n374), .B2(n478), .A(n363), .ZN(n609) );
  NAND2_X1 U441 ( .A1(n373), .A2(B_extended[7]), .ZN(n364) );
  OAI21_X1 U442 ( .B1(n370), .B2(n477), .A(n364), .ZN(n611) );
  NAND2_X1 U443 ( .A1(n255), .A2(A_extended[0]), .ZN(n365) );
  OAI21_X1 U444 ( .B1(n374), .B2(n476), .A(n365), .ZN(n613) );
  NAND2_X1 U445 ( .A1(n264), .A2(A_extended[1]), .ZN(n366) );
  OAI21_X1 U446 ( .B1(n374), .B2(n475), .A(n366), .ZN(n615) );
  NAND2_X1 U447 ( .A1(n269), .A2(A_extended[2]), .ZN(n367) );
  OAI21_X1 U448 ( .B1(n374), .B2(n474), .A(n367), .ZN(n617) );
  NAND2_X1 U449 ( .A1(n373), .A2(A_extended[3]), .ZN(n368) );
  OAI21_X1 U450 ( .B1(n374), .B2(n473), .A(n368), .ZN(n619) );
  NAND2_X1 U451 ( .A1(n370), .A2(A_extended[4]), .ZN(n369) );
  OAI21_X1 U452 ( .B1(n370), .B2(n472), .A(n369), .ZN(n621) );
  NAND2_X1 U453 ( .A1(n373), .A2(A_extended[5]), .ZN(n371) );
  OAI21_X1 U454 ( .B1(n374), .B2(n471), .A(n371), .ZN(n623) );
  NAND2_X1 U455 ( .A1(n373), .A2(A_extended[6]), .ZN(n372) );
  OAI21_X1 U456 ( .B1(n374), .B2(n470), .A(n372), .ZN(n625) );
  NAND2_X1 U457 ( .A1(n468), .A2(n302), .ZN(n629) );
endmodule


module conv_128_32_DW_mult_pipe_J1_31 ( clk, rst_n, en, tc, a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  input clk, rst_n, en, tc;
  wire   \mult_x_1/a[6] , \mult_x_1/a[4] , \mult_x_1/n313 , \mult_x_1/n312 ,
         \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n288 , \mult_x_1/n287 ,
         \mult_x_1/n286 , \mult_x_1/n285 , \mult_x_1/n284 , \mult_x_1/n283 ,
         \mult_x_1/n282 , \mult_x_1/n281 , \mult_x_1/n180 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n398, n400, n402, n404, n406, n408,
         n410, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n521, n523, n525, n527, n529,
         n531, n533, n535, n537, n539, n541, n543, n545, n547, n549, n551,
         n553, n555, n557, n559, n561, n563, n565, n567, n569, n571, n573,
         n575, n577, n579, n581, n583, n585, n587, n589, n591, n593, n595,
         n597, n599, n601, n603, n605, n607, n609, n611, n613, n615, n617,
         n619, n621, n623, n625, n627, n644, n645;
  wire   [8:0] A_extended;
  wire   [8:0] B_extended;
  assign A_extended[7] = a[7];
  assign A_extended[6] = a[6];
  assign A_extended[5] = a[5];
  assign A_extended[4] = a[4];
  assign A_extended[3] = a[3];
  assign A_extended[2] = a[2];
  assign A_extended[1] = a[1];
  assign A_extended[0] = a[0];
  assign B_extended[7] = b[7];
  assign B_extended[6] = b[6];
  assign B_extended[5] = b[5];
  assign B_extended[4] = b[4];
  assign B_extended[3] = b[3];
  assign B_extended[2] = b[2];
  assign B_extended[1] = b[1];
  assign B_extended[0] = b[0];

  SDFF_X1 clk_r_REG75_S1 ( .D(1'b0), .SI(n465), .SE(n627), .CK(clk), .Q(n644), 
        .QN(n466) );
  SDFF_X1 clk_r_REG36_S1 ( .D(1'b0), .SI(n465), .SE(n623), .CK(clk), .Q(
        \mult_x_1/a[6] ), .QN(n468) );
  SDFF_X1 clk_r_REG63_S1 ( .D(1'b0), .SI(n465), .SE(n611), .CK(clk), .Q(
        \mult_x_1/n180 ), .QN(n474) );
  SDFF_X1 clk_r_REG67_S1 ( .D(1'b0), .SI(n465), .SE(n609), .CK(clk), .Q(
        \mult_x_1/n281 ), .QN(n475) );
  SDFF_X1 clk_r_REG68_S1 ( .D(1'b0), .SI(n465), .SE(n607), .CK(clk), .Q(
        \mult_x_1/n282 ), .QN(n476) );
  SDFF_X1 clk_r_REG69_S1 ( .D(1'b0), .SI(n463), .SE(n605), .CK(clk), .Q(
        \mult_x_1/n283 ), .QN(n477) );
  SDFF_X1 clk_r_REG70_S1 ( .D(1'b0), .SI(n464), .SE(n603), .CK(clk), .Q(
        \mult_x_1/n284 ), .QN(n478) );
  SDFF_X1 clk_r_REG71_S1 ( .D(1'b0), .SI(n462), .SE(n601), .CK(clk), .Q(
        \mult_x_1/n285 ), .QN(n479) );
  SDFF_X1 clk_r_REG72_S1 ( .D(1'b0), .SI(n465), .SE(n599), .CK(clk), .Q(
        \mult_x_1/n286 ), .QN(n480) );
  SDFF_X1 clk_r_REG73_S1 ( .D(1'b0), .SI(n462), .SE(n597), .CK(clk), .Q(
        \mult_x_1/n287 ), .QN(n481) );
  SDFF_X1 clk_r_REG74_S1 ( .D(1'b0), .SI(n462), .SE(n595), .CK(clk), .Q(
        \mult_x_1/n288 ), .QN(n482) );
  SDFF_X1 clk_r_REG2_S3 ( .D(1'b0), .SI(n462), .SE(n593), .CK(clk), .QN(n483)
         );
  SDFF_X1 clk_r_REG3_S4 ( .D(1'b0), .SI(n462), .SE(n591), .CK(clk), .Q(
        product[15]), .QN(n484) );
  SDFF_X1 clk_r_REG5_S3 ( .D(1'b0), .SI(n462), .SE(n589), .CK(clk), .QN(n485)
         );
  SDFF_X1 clk_r_REG6_S4 ( .D(1'b0), .SI(n462), .SE(n587), .CK(clk), .Q(
        product[14]), .QN(n486) );
  SDFF_X1 clk_r_REG9_S3 ( .D(1'b0), .SI(n462), .SE(n585), .CK(clk), .QN(n487)
         );
  SDFF_X1 clk_r_REG10_S4 ( .D(1'b0), .SI(n464), .SE(n583), .CK(clk), .Q(
        product[13]), .QN(n488) );
  SDFF_X1 clk_r_REG15_S3 ( .D(1'b0), .SI(n465), .SE(n581), .CK(clk), .QN(n489)
         );
  SDFF_X1 clk_r_REG16_S4 ( .D(1'b0), .SI(n463), .SE(n579), .CK(clk), .Q(
        product[12]), .QN(n490) );
  SDFF_X1 clk_r_REG17_S3 ( .D(1'b0), .SI(n462), .SE(n577), .CK(clk), .QN(n491)
         );
  SDFF_X1 clk_r_REG18_S4 ( .D(1'b0), .SI(n462), .SE(n575), .CK(clk), .Q(
        product[11]), .QN(n492) );
  SDFF_X1 clk_r_REG19_S3 ( .D(1'b0), .SI(n462), .SE(n573), .CK(clk), .QN(n493)
         );
  SDFF_X1 clk_r_REG20_S4 ( .D(1'b0), .SI(n462), .SE(n571), .CK(clk), .Q(
        product[10]), .QN(n494) );
  SDFF_X1 clk_r_REG13_S3 ( .D(1'b0), .SI(n462), .SE(n569), .CK(clk), .QN(n495)
         );
  SDFF_X1 clk_r_REG14_S4 ( .D(1'b0), .SI(n462), .SE(n567), .CK(clk), .Q(
        product[9]), .QN(n496) );
  SDFF_X1 clk_r_REG29_S3 ( .D(1'b0), .SI(n462), .SE(n565), .CK(clk), .QN(n497)
         );
  SDFF_X1 clk_r_REG30_S4 ( .D(1'b0), .SI(n464), .SE(n563), .CK(clk), .Q(
        product[8]), .QN(n498) );
  SDFF_X1 clk_r_REG33_S3 ( .D(1'b0), .SI(n464), .SE(n561), .CK(clk), .QN(n499)
         );
  SDFF_X1 clk_r_REG34_S4 ( .D(1'b0), .SI(n464), .SE(n559), .CK(clk), .Q(
        product[7]), .QN(n500) );
  SDFF_X1 clk_r_REG38_S3 ( .D(1'b0), .SI(n464), .SE(n557), .CK(clk), .QN(n501)
         );
  SDFF_X1 clk_r_REG39_S4 ( .D(1'b0), .SI(n464), .SE(n555), .CK(clk), .Q(
        product[6]), .QN(n502) );
  SDFF_X1 clk_r_REG43_S3 ( .D(1'b0), .SI(n464), .SE(n553), .CK(clk), .QN(n503)
         );
  SDFF_X1 clk_r_REG44_S4 ( .D(1'b0), .SI(n464), .SE(n551), .CK(clk), .Q(
        product[5]), .QN(n504) );
  SDFF_X1 clk_r_REG47_S2 ( .D(1'b0), .SI(n464), .SE(n549), .CK(clk), .QN(n505)
         );
  SDFF_X1 clk_r_REG48_S3 ( .D(1'b0), .SI(n464), .SE(n547), .CK(clk), .QN(n506)
         );
  SDFF_X1 clk_r_REG49_S4 ( .D(1'b0), .SI(n464), .SE(n545), .CK(clk), .Q(
        product[4]), .QN(n507) );
  SDFF_X1 clk_r_REG52_S2 ( .D(1'b0), .SI(n464), .SE(n543), .CK(clk), .QN(n508)
         );
  SDFF_X1 clk_r_REG53_S3 ( .D(1'b0), .SI(n463), .SE(n541), .CK(clk), .QN(n509)
         );
  SDFF_X1 clk_r_REG54_S4 ( .D(1'b0), .SI(n463), .SE(n539), .CK(clk), .Q(
        product[3]), .QN(n510) );
  SDFF_X1 clk_r_REG56_S2 ( .D(1'b0), .SI(n463), .SE(n537), .CK(clk), .QN(n511)
         );
  SDFF_X1 clk_r_REG57_S3 ( .D(1'b0), .SI(n463), .SE(n535), .CK(clk), .QN(n512)
         );
  SDFF_X1 clk_r_REG58_S4 ( .D(1'b0), .SI(n463), .SE(n533), .CK(clk), .Q(
        product[2]), .QN(n513) );
  SDFF_X1 clk_r_REG60_S2 ( .D(1'b0), .SI(n463), .SE(n531), .CK(clk), .QN(n514)
         );
  SDFF_X1 clk_r_REG61_S3 ( .D(1'b0), .SI(n463), .SE(n529), .CK(clk), .QN(n515)
         );
  SDFF_X1 clk_r_REG62_S4 ( .D(1'b0), .SI(n463), .SE(n527), .CK(clk), .Q(
        product[1]), .QN(n516) );
  SDFF_X1 clk_r_REG64_S2 ( .D(1'b0), .SI(n463), .SE(n525), .CK(clk), .QN(n517)
         );
  SDFF_X1 clk_r_REG65_S3 ( .D(1'b0), .SI(n463), .SE(n523), .CK(clk), .QN(n518)
         );
  SDFF_X1 clk_r_REG66_S4 ( .D(1'b0), .SI(n463), .SE(n521), .CK(clk), .Q(
        product[0]), .QN(n519) );
  SDFF_X1 \mult_x_1/clk_r_REG24_S2_IP  ( .D(1'b1), .SI(n645), .SE(n438), .CK(
        clk), .Q(n440), .QN(n395) );
  SDFF_X1 \mult_x_1/clk_r_REG25_S2  ( .D(n645), .SI(1'b1), .SE(n436), .CK(clk), 
        .Q(n394), .QN(n441) );
  SDFF_X1 \mult_x_1/clk_r_REG50_S2_IP  ( .D(1'b1), .SI(n645), .SE(n434), .CK(
        clk), .Q(n442), .QN(n393) );
  SDFF_X1 \mult_x_1/clk_r_REG45_S2  ( .D(n645), .SI(1'b1), .SE(n432), .CK(clk), 
        .Q(n392), .QN(n443) );
  SDFF_X1 \mult_x_1/clk_r_REG21_S2  ( .D(n645), .SI(1'b1), .SE(n430), .CK(clk), 
        .Q(n391), .QN(n444) );
  SDFF_X1 \mult_x_1/clk_r_REG27_S2  ( .D(n645), .SI(1'b1), .SE(n428), .CK(clk), 
        .Q(n390), .QN(n445) );
  SDFF_X1 \mult_x_1/clk_r_REG11_S2  ( .D(n645), .SI(1'b1), .SE(n426), .CK(clk), 
        .Q(n389), .QN(n446) );
  SDFF_X1 \mult_x_1/clk_r_REG22_S2_IP  ( .D(1'b1), .SI(n645), .SE(n424), .CK(
        clk), .Q(n447), .QN(n388) );
  SDFF_X1 \mult_x_1/clk_r_REG23_S2_IP  ( .D(1'b1), .SI(n645), .SE(n422), .CK(
        clk), .Q(n448), .QN(n387) );
  SDFF_X1 \mult_x_1/clk_r_REG42_S2  ( .D(n645), .SI(1'b1), .SE(n420), .CK(clk), 
        .Q(n386), .QN(n449) );
  SDFF_X1 \mult_x_1/clk_r_REG37_S2  ( .D(n645), .SI(1'b1), .SE(n418), .CK(clk), 
        .Q(n385), .QN(n450) );
  SDFF_X1 \mult_x_1/clk_r_REG40_S2  ( .D(n645), .SI(1'b1), .SE(n416), .CK(clk), 
        .Q(n384), .QN(n451) );
  SDFF_X1 \mult_x_1/clk_r_REG32_S2  ( .D(n645), .SI(1'b1), .SE(n414), .CK(clk), 
        .Q(n383), .QN(n452) );
  SDFF_X1 \mult_x_1/clk_r_REG28_S2  ( .D(n645), .SI(1'b1), .SE(n412), .CK(clk), 
        .Q(n382), .QN(n453) );
  SDFF_X1 \mult_x_1/clk_r_REG31_S2  ( .D(n645), .SI(1'b1), .SE(n410), .CK(clk), 
        .Q(n381), .QN(n454) );
  SDFF_X1 \mult_x_1/clk_r_REG12_S2  ( .D(n645), .SI(1'b1), .SE(n408), .CK(clk), 
        .Q(n380), .QN(n455) );
  SDFF_X1 \mult_x_1/clk_r_REG4_S2  ( .D(n645), .SI(1'b1), .SE(n406), .CK(clk), 
        .Q(n379), .QN(n456) );
  SDFF_X1 \mult_x_1/clk_r_REG1_S2_IP  ( .D(1'b1), .SI(n645), .SE(n404), .CK(
        clk), .Q(n457), .QN(n378) );
  SDFF_X1 \mult_x_1/clk_r_REG35_S2_IP  ( .D(1'b1), .SI(n645), .SE(n402), .CK(
        clk), .Q(n458), .QN(n377) );
  SDFF_X1 \mult_x_1/clk_r_REG26_S2  ( .D(n645), .SI(1'b1), .SE(n400), .CK(clk), 
        .Q(n376), .QN(n459) );
  SDFF_X1 \mult_x_1/clk_r_REG8_S2  ( .D(n645), .SI(1'b1), .SE(n398), .CK(clk), 
        .Q(n375) );
  SDFF_X1 \mult_x_1/clk_r_REG7_S2  ( .D(n645), .SI(1'b1), .SE(n396), .CK(clk), 
        .Q(n374), .QN(n461) );
  SDFF_X1 clk_r_REG51_S1 ( .D(1'b0), .SI(n465), .SE(n617), .CK(clk), .Q(
        \mult_x_1/n312 ), .QN(n471) );
  SDFF_X1 clk_r_REG41_S1 ( .D(1'b0), .SI(n465), .SE(n621), .CK(clk), .Q(
        \mult_x_1/n311 ), .QN(n469) );
  SDFF_X1 clk_r_REG46_S1 ( .D(1'b0), .SI(n465), .SE(n619), .CK(clk), .Q(
        \mult_x_1/a[4] ), .QN(n470) );
  SDFF_X1 clk_r_REG55_S1 ( .D(1'b0), .SI(n465), .SE(n615), .CK(clk), .QN(n472)
         );
  SDFF_X1 clk_r_REG0_S1 ( .D(1'b0), .SI(n465), .SE(n625), .CK(clk), .Q(
        \mult_x_1/n310 ), .QN(n467) );
  SDFF_X1 clk_r_REG59_S1 ( .D(1'b0), .SI(n465), .SE(n613), .CK(clk), .Q(
        \mult_x_1/n313 ), .QN(n473) );
  BUF_X1 U2 ( .A(n268), .Z(n373) );
  INV_X1 U3 ( .A(n268), .ZN(n371) );
  INV_X1 U4 ( .A(rst_n), .ZN(n645) );
  INV_X1 U5 ( .A(n645), .ZN(n462) );
  AND2_X1 U6 ( .A1(n248), .A2(n249), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(n462), .Z(n465) );
  CLKBUF_X1 U8 ( .A(n462), .Z(n463) );
  CLKBUF_X1 U9 ( .A(n462), .Z(n464) );
  NAND2_X1 U10 ( .A1(n8), .A2(n7), .ZN(n206) );
  OAI21_X1 U11 ( .B1(n140), .B2(n139), .A(n9), .ZN(n8) );
  NAND2_X1 U12 ( .A1(n140), .A2(n139), .ZN(n7) );
  OAI22_X1 U13 ( .A1(n47), .A2(n45), .B1(n33), .B2(n25), .ZN(n57) );
  INV_X1 U14 ( .A(n32), .ZN(n220) );
  NAND2_X1 U15 ( .A1(n31), .A2(n25), .ZN(n24) );
  XNOR2_X1 U16 ( .A(n6), .B(n9), .ZN(n249) );
  XNOR2_X1 U17 ( .A(n140), .B(n139), .ZN(n6) );
  INV_X1 U18 ( .A(\mult_x_1/n311 ), .ZN(n16) );
  NAND2_X1 U19 ( .A1(n46), .A2(n31), .ZN(n47) );
  XNOR2_X1 U20 ( .A(n472), .B(\mult_x_1/n312 ), .ZN(n31) );
  OAI21_X1 U21 ( .B1(n5), .B2(n21), .A(n63), .ZN(n428) );
  NAND2_X1 U22 ( .A1(n42), .A2(n41), .ZN(n9) );
  NAND2_X1 U23 ( .A1(n37), .A2(n36), .ZN(n40) );
  INV_X1 U24 ( .A(n59), .ZN(n36) );
  INV_X1 U25 ( .A(n60), .ZN(n37) );
  OAI21_X1 U26 ( .B1(n23), .B2(n90), .A(n92), .ZN(n55) );
  NAND2_X1 U27 ( .A1(n23), .A2(n90), .ZN(n54) );
  XNOR2_X1 U28 ( .A(\mult_x_1/a[6] ), .B(n469), .ZN(n49) );
  NAND2_X1 U29 ( .A1(n60), .A2(n59), .ZN(n41) );
  NAND2_X1 U30 ( .A1(n55), .A2(n54), .ZN(n240) );
  XNOR2_X1 U31 ( .A(n60), .B(n59), .ZN(n61) );
  BUF_X2 U32 ( .A(n366), .Z(n262) );
  XNOR2_X1 U33 ( .A(\mult_x_1/a[4] ), .B(n471), .ZN(n10) );
  XOR2_X1 U34 ( .A(n258), .B(n257), .Z(n11) );
  XOR2_X1 U35 ( .A(n256), .B(n11), .Z(n86) );
  NAND2_X1 U36 ( .A1(n256), .A2(n258), .ZN(n12) );
  NAND2_X1 U37 ( .A1(n256), .A2(n257), .ZN(n13) );
  NAND2_X1 U38 ( .A1(n258), .A2(n257), .ZN(n14) );
  NAND3_X1 U39 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n264) );
  NAND2_X1 U40 ( .A1(n29), .A2(n50), .ZN(n15) );
  NAND2_X1 U41 ( .A1(n29), .A2(n50), .ZN(n161) );
  INV_X2 U42 ( .A(n16), .ZN(n17) );
  INV_X1 U43 ( .A(n49), .ZN(n162) );
  OR2_X1 U44 ( .A1(n262), .A2(n443), .ZN(n18) );
  NAND2_X1 U45 ( .A1(n18), .A2(n235), .ZN(n432) );
  XNOR2_X1 U46 ( .A(\mult_x_1/a[6] ), .B(n467), .ZN(n50) );
  NAND2_X1 U47 ( .A1(n466), .A2(\mult_x_1/n310 ), .ZN(n164) );
  XNOR2_X1 U48 ( .A(n62), .B(n61), .ZN(n238) );
  INV_X1 U49 ( .A(n10), .ZN(n19) );
  INV_X1 U50 ( .A(n10), .ZN(n20) );
  NAND2_X1 U51 ( .A1(n21), .A2(n375), .ZN(n22) );
  NAND2_X1 U52 ( .A1(n22), .A2(n142), .ZN(n398) );
  INV_X1 U53 ( .A(n366), .ZN(n21) );
  OR2_X1 U54 ( .A1(n101), .A2(n100), .ZN(n23) );
  OR2_X1 U55 ( .A1(n101), .A2(n100), .ZN(n91) );
  XNOR2_X1 U56 ( .A(n472), .B(n473), .ZN(n25) );
  OAI22_X1 U57 ( .A1(n147), .A2(n39), .B1(n20), .B2(n35), .ZN(n60) );
  XNOR2_X1 U58 ( .A(n472), .B(n473), .ZN(n46) );
  INV_X4 U59 ( .A(n268), .ZN(n369) );
  INV_X4 U60 ( .A(n268), .ZN(n345) );
  AND2_X1 U61 ( .A1(n28), .A2(n19), .ZN(n26) );
  INV_X2 U62 ( .A(en), .ZN(n268) );
  INV_X1 U63 ( .A(n268), .ZN(n366) );
  AND2_X1 U64 ( .A1(n103), .A2(n102), .ZN(n27) );
  XOR2_X1 U65 ( .A(\mult_x_1/a[4] ), .B(\mult_x_1/n311 ), .Z(n28) );
  INV_X1 U66 ( .A(n26), .ZN(n44) );
  XNOR2_X1 U67 ( .A(n17), .B(\mult_x_1/n281 ), .ZN(n35) );
  AND2_X1 U68 ( .A1(n644), .A2(\mult_x_1/n281 ), .ZN(n123) );
  XNOR2_X1 U69 ( .A(n123), .B(n17), .ZN(n126) );
  OAI22_X1 U70 ( .A1(n44), .A2(n35), .B1(n126), .B2(n20), .ZN(n132) );
  INV_X1 U71 ( .A(n132), .ZN(n130) );
  INV_X1 U72 ( .A(n49), .ZN(n29) );
  XNOR2_X1 U73 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n283 ), .ZN(n30) );
  XNOR2_X1 U74 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n282 ), .ZN(n125) );
  OAI22_X1 U75 ( .A1(n15), .A2(n30), .B1(n162), .B2(n125), .ZN(n129) );
  NOR2_X1 U76 ( .A1(n478), .A2(n164), .ZN(n128) );
  XNOR2_X1 U77 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n284 ), .ZN(n38) );
  OAI22_X1 U78 ( .A1(n15), .A2(n38), .B1(n162), .B2(n30), .ZN(n58) );
  XNOR2_X1 U79 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n281 ), .ZN(n45) );
  XNOR2_X1 U80 ( .A(n123), .B(\mult_x_1/n312 ), .ZN(n33) );
  INV_X1 U81 ( .A(n46), .ZN(n32) );
  AOI21_X1 U82 ( .B1(n220), .B2(n24), .A(n33), .ZN(n34) );
  INV_X1 U83 ( .A(n34), .ZN(n56) );
  INV_X1 U84 ( .A(n26), .ZN(n147) );
  XNOR2_X1 U85 ( .A(n17), .B(\mult_x_1/n282 ), .ZN(n39) );
  NOR2_X1 U86 ( .A1(n479), .A2(n164), .ZN(n59) );
  XNOR2_X1 U87 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n285 ), .ZN(n53) );
  OAI22_X1 U88 ( .A1(n15), .A2(n53), .B1(n162), .B2(n38), .ZN(n96) );
  INV_X1 U89 ( .A(n26), .ZN(n151) );
  XNOR2_X1 U90 ( .A(n17), .B(\mult_x_1/n283 ), .ZN(n43) );
  OAI22_X1 U91 ( .A1(n151), .A2(n43), .B1(n20), .B2(n39), .ZN(n95) );
  INV_X1 U92 ( .A(n57), .ZN(n94) );
  NAND2_X1 U93 ( .A1(n40), .A2(n62), .ZN(n42) );
  XNOR2_X1 U94 ( .A(n17), .B(\mult_x_1/n284 ), .ZN(n68) );
  OAI22_X1 U95 ( .A1(n44), .A2(n68), .B1(n20), .B2(n43), .ZN(n101) );
  XNOR2_X1 U96 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n282 ), .ZN(n70) );
  OAI22_X1 U97 ( .A1(n47), .A2(n70), .B1(n25), .B2(n45), .ZN(n100) );
  NOR2_X1 U98 ( .A1(n480), .A2(n164), .ZN(n90) );
  NAND2_X1 U99 ( .A1(\mult_x_1/n313 ), .A2(n474), .ZN(n222) );
  XNOR2_X1 U100 ( .A(n123), .B(\mult_x_1/n313 ), .ZN(n65) );
  AOI21_X1 U101 ( .B1(n222), .B2(n474), .A(n65), .ZN(n48) );
  INV_X1 U102 ( .A(n48), .ZN(n110) );
  XNOR2_X1 U103 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n286 ), .ZN(n64) );
  NOR2_X1 U104 ( .A1(n49), .A2(n64), .ZN(n51) );
  NAND2_X1 U105 ( .A1(n51), .A2(n50), .ZN(n52) );
  OAI21_X1 U106 ( .B1(n162), .B2(n53), .A(n52), .ZN(n109) );
  NOR2_X1 U107 ( .A1(n481), .A2(n164), .ZN(n108) );
  FA_X1 U108 ( .A(n58), .B(n57), .CI(n56), .CO(n139), .S(n239) );
  OR2_X1 U109 ( .A1(n262), .A2(n445), .ZN(n63) );
  XNOR2_X1 U110 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n287 ), .ZN(n72) );
  OAI22_X1 U111 ( .A1(n161), .A2(n72), .B1(n162), .B2(n64), .ZN(n99) );
  XNOR2_X1 U112 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n281 ), .ZN(n67) );
  OAI22_X1 U113 ( .A1(n222), .A2(n67), .B1(n65), .B2(n474), .ZN(n98) );
  INV_X1 U114 ( .A(n164), .ZN(n66) );
  AND2_X1 U115 ( .A1(\mult_x_1/n288 ), .A2(n66), .ZN(n97) );
  XNOR2_X1 U116 ( .A(n17), .B(\mult_x_1/n286 ), .ZN(n149) );
  XNOR2_X1 U117 ( .A(n17), .B(\mult_x_1/n285 ), .ZN(n69) );
  OAI22_X1 U118 ( .A1(n151), .A2(n149), .B1(n20), .B2(n69), .ZN(n81) );
  XNOR2_X1 U119 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n282 ), .ZN(n75) );
  OAI22_X1 U120 ( .A1(n222), .A2(n75), .B1(n67), .B2(n474), .ZN(n80) );
  XNOR2_X1 U121 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n284 ), .ZN(n76) );
  XNOR2_X1 U122 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n283 ), .ZN(n71) );
  OAI22_X1 U123 ( .A1(n24), .A2(n76), .B1(n220), .B2(n71), .ZN(n79) );
  OAI22_X1 U124 ( .A1(n147), .A2(n69), .B1(n20), .B2(n68), .ZN(n107) );
  OAI22_X1 U125 ( .A1(n24), .A2(n71), .B1(n220), .B2(n70), .ZN(n106) );
  XNOR2_X1 U126 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n288 ), .ZN(n73) );
  OAI22_X1 U127 ( .A1(n15), .A2(n73), .B1(n162), .B2(n72), .ZN(n78) );
  OR2_X1 U128 ( .A1(\mult_x_1/n288 ), .A2(n467), .ZN(n74) );
  OAI22_X1 U129 ( .A1(n161), .A2(n467), .B1(n74), .B2(n162), .ZN(n77) );
  XNOR2_X1 U130 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n283 ), .ZN(n187) );
  OAI22_X1 U131 ( .A1(n222), .A2(n187), .B1(n75), .B2(n474), .ZN(n154) );
  AND2_X1 U132 ( .A1(\mult_x_1/n288 ), .A2(n49), .ZN(n153) );
  XNOR2_X1 U133 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n285 ), .ZN(n186) );
  OAI22_X1 U134 ( .A1(n24), .A2(n186), .B1(n220), .B2(n76), .ZN(n152) );
  HA_X1 U135 ( .A(n78), .B(n77), .CO(n105), .S(n144) );
  FA_X1 U136 ( .A(n81), .B(n80), .CI(n79), .CO(n257), .S(n143) );
  NAND2_X1 U137 ( .A1(n86), .A2(n85), .ZN(n82) );
  NAND2_X1 U138 ( .A1(n82), .A2(n369), .ZN(n84) );
  OR2_X1 U139 ( .A1(n262), .A2(n453), .ZN(n83) );
  NAND2_X1 U140 ( .A1(n84), .A2(n83), .ZN(n412) );
  NOR2_X1 U141 ( .A1(n86), .A2(n85), .ZN(n87) );
  NAND2_X1 U142 ( .A1(n87), .A2(n345), .ZN(n89) );
  OR2_X1 U143 ( .A1(n262), .A2(n454), .ZN(n88) );
  NAND2_X1 U144 ( .A1(n89), .A2(n88), .ZN(n410) );
  XNOR2_X1 U145 ( .A(n91), .B(n90), .ZN(n93) );
  XNOR2_X1 U146 ( .A(n93), .B(n92), .ZN(n244) );
  FA_X1 U147 ( .A(n96), .B(n95), .CI(n94), .CO(n62), .S(n243) );
  FA_X1 U148 ( .A(n99), .B(n98), .CI(n97), .CO(n103), .S(n258) );
  XNOR2_X1 U149 ( .A(n101), .B(n100), .ZN(n102) );
  INV_X1 U150 ( .A(n102), .ZN(n104) );
  XNOR2_X1 U151 ( .A(n104), .B(n103), .ZN(n254) );
  FA_X1 U152 ( .A(n107), .B(n106), .CI(n105), .CO(n253), .S(n256) );
  NAND2_X1 U153 ( .A1(n254), .A2(n253), .ZN(n113) );
  FA_X1 U154 ( .A(n110), .B(n109), .CI(n108), .CO(n92), .S(n252) );
  NAND2_X1 U155 ( .A1(n254), .A2(n252), .ZN(n112) );
  NAND2_X1 U156 ( .A1(n253), .A2(n252), .ZN(n111) );
  NAND3_X1 U157 ( .A1(n113), .A2(n112), .A3(n111), .ZN(n118) );
  NAND2_X1 U158 ( .A1(n117), .A2(n118), .ZN(n114) );
  NAND2_X1 U159 ( .A1(n114), .A2(n262), .ZN(n116) );
  OR2_X1 U160 ( .A1(n262), .A2(n447), .ZN(n115) );
  NAND2_X1 U161 ( .A1(n116), .A2(n115), .ZN(n424) );
  INV_X1 U162 ( .A(n117), .ZN(n120) );
  INV_X1 U163 ( .A(n118), .ZN(n119) );
  NAND3_X1 U164 ( .A1(n120), .A2(n262), .A3(n119), .ZN(n122) );
  OR2_X1 U165 ( .A1(n262), .A2(n448), .ZN(n121) );
  NAND2_X1 U166 ( .A1(n122), .A2(n121), .ZN(n422) );
  BUF_X2 U189 ( .A(n366), .Z(n247) );
  NOR2_X1 U190 ( .A1(n476), .A2(n164), .ZN(n159) );
  XNOR2_X1 U191 ( .A(\mult_x_1/n310 ), .B(\mult_x_1/n281 ), .ZN(n124) );
  XNOR2_X1 U192 ( .A(n123), .B(\mult_x_1/n310 ), .ZN(n160) );
  OAI22_X1 U193 ( .A1(n15), .A2(n124), .B1(n160), .B2(n162), .ZN(n168) );
  INV_X1 U194 ( .A(n168), .ZN(n158) );
  OAI22_X1 U195 ( .A1(n15), .A2(n125), .B1(n162), .B2(n124), .ZN(n133) );
  AOI21_X1 U196 ( .B1(n20), .B2(n147), .A(n126), .ZN(n127) );
  INV_X1 U197 ( .A(n127), .ZN(n131) );
  FA_X1 U198 ( .A(n128), .B(n129), .CI(n130), .CO(n138), .S(n140) );
  NOR2_X1 U199 ( .A1(n477), .A2(n164), .ZN(n137) );
  FA_X1 U200 ( .A(n133), .B(n132), .CI(n131), .CO(n157), .S(n136) );
  OR2_X1 U201 ( .A1(n176), .A2(n175), .ZN(n134) );
  NAND2_X1 U202 ( .A1(n247), .A2(n134), .ZN(n135) );
  OAI21_X1 U203 ( .B1(n345), .B2(n461), .A(n135), .ZN(n396) );
  FA_X1 U204 ( .A(n138), .B(n137), .CI(n136), .CO(n175), .S(n207) );
  OR2_X1 U205 ( .A1(n207), .A2(n206), .ZN(n141) );
  NAND2_X1 U206 ( .A1(n247), .A2(n141), .ZN(n142) );
  FA_X1 U207 ( .A(n145), .B(n144), .CI(n143), .CO(n85), .S(n180) );
  OR2_X1 U208 ( .A1(\mult_x_1/n288 ), .A2(n16), .ZN(n146) );
  OAI22_X1 U209 ( .A1(n147), .A2(n16), .B1(n146), .B2(n20), .ZN(n189) );
  XNOR2_X1 U210 ( .A(n17), .B(\mult_x_1/n288 ), .ZN(n148) );
  XNOR2_X1 U211 ( .A(n17), .B(\mult_x_1/n287 ), .ZN(n150) );
  OAI22_X1 U212 ( .A1(n151), .A2(n148), .B1(n20), .B2(n150), .ZN(n188) );
  OAI22_X1 U213 ( .A1(n151), .A2(n150), .B1(n20), .B2(n149), .ZN(n184) );
  FA_X1 U214 ( .A(n154), .B(n153), .CI(n152), .CO(n145), .S(n183) );
  OR2_X1 U215 ( .A1(n180), .A2(n179), .ZN(n155) );
  NAND2_X1 U216 ( .A1(n247), .A2(n155), .ZN(n156) );
  OAI21_X1 U217 ( .B1(n369), .B2(n458), .A(n156), .ZN(n402) );
  FA_X1 U218 ( .A(n159), .B(n158), .CI(n157), .CO(n170), .S(n176) );
  AOI21_X1 U219 ( .B1(n162), .B2(n15), .A(n160), .ZN(n163) );
  INV_X1 U220 ( .A(n163), .ZN(n166) );
  NOR2_X1 U221 ( .A1(n475), .A2(n164), .ZN(n165) );
  XOR2_X1 U222 ( .A(n166), .B(n165), .Z(n167) );
  XOR2_X1 U223 ( .A(n168), .B(n167), .Z(n169) );
  OR2_X1 U224 ( .A1(n170), .A2(n169), .ZN(n172) );
  NAND2_X1 U225 ( .A1(n170), .A2(n169), .ZN(n171) );
  NAND2_X1 U226 ( .A1(n172), .A2(n171), .ZN(n173) );
  NAND2_X1 U227 ( .A1(n247), .A2(n173), .ZN(n174) );
  OAI21_X1 U228 ( .B1(n369), .B2(n457), .A(n174), .ZN(n404) );
  NAND2_X1 U229 ( .A1(n176), .A2(n175), .ZN(n177) );
  NAND2_X1 U230 ( .A1(n247), .A2(n177), .ZN(n178) );
  OAI21_X1 U231 ( .B1(n345), .B2(n456), .A(n178), .ZN(n406) );
  NAND2_X1 U232 ( .A1(n180), .A2(n179), .ZN(n181) );
  NAND2_X1 U233 ( .A1(n247), .A2(n181), .ZN(n182) );
  OAI21_X1 U234 ( .B1(n371), .B2(n452), .A(n182), .ZN(n414) );
  FA_X1 U235 ( .A(n185), .B(n184), .CI(n183), .CO(n179), .S(n193) );
  XNOR2_X1 U236 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n286 ), .ZN(n201) );
  OAI22_X1 U237 ( .A1(n24), .A2(n201), .B1(n220), .B2(n186), .ZN(n198) );
  XNOR2_X1 U238 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n284 ), .ZN(n199) );
  OAI22_X1 U239 ( .A1(n222), .A2(n199), .B1(n187), .B2(n474), .ZN(n197) );
  HA_X1 U240 ( .A(n189), .B(n188), .CO(n185), .S(n196) );
  NOR2_X1 U241 ( .A1(n193), .A2(n192), .ZN(n190) );
  NAND2_X1 U242 ( .A1(n247), .A2(n190), .ZN(n191) );
  OAI21_X1 U243 ( .B1(n369), .B2(n451), .A(n191), .ZN(n416) );
  NAND2_X1 U244 ( .A1(n193), .A2(n192), .ZN(n194) );
  NAND2_X1 U245 ( .A1(n247), .A2(n194), .ZN(n195) );
  OAI21_X1 U246 ( .B1(n345), .B2(n450), .A(n195), .ZN(n418) );
  FA_X1 U247 ( .A(n198), .B(n197), .CI(n196), .CO(n192), .S(n203) );
  XNOR2_X1 U248 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n285 ), .ZN(n215) );
  OAI22_X1 U249 ( .A1(n222), .A2(n215), .B1(n199), .B2(n474), .ZN(n212) );
  INV_X1 U250 ( .A(n20), .ZN(n200) );
  AND2_X1 U251 ( .A1(\mult_x_1/n288 ), .A2(n200), .ZN(n211) );
  XNOR2_X1 U252 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n287 ), .ZN(n213) );
  OAI22_X1 U253 ( .A1(n24), .A2(n213), .B1(n220), .B2(n201), .ZN(n210) );
  OR2_X1 U254 ( .A1(n203), .A2(n202), .ZN(n233) );
  NAND2_X1 U255 ( .A1(n203), .A2(n202), .ZN(n231) );
  NAND2_X1 U256 ( .A1(n233), .A2(n231), .ZN(n204) );
  NAND2_X1 U257 ( .A1(n371), .A2(n204), .ZN(n205) );
  OAI21_X1 U258 ( .B1(n262), .B2(n449), .A(n205), .ZN(n420) );
  NAND2_X1 U259 ( .A1(n207), .A2(n206), .ZN(n208) );
  NAND2_X1 U260 ( .A1(n247), .A2(n208), .ZN(n209) );
  OAI21_X1 U261 ( .B1(n262), .B2(n446), .A(n209), .ZN(n426) );
  FA_X1 U262 ( .A(n212), .B(n211), .CI(n210), .CO(n202), .S(n230) );
  XNOR2_X1 U263 ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n288 ), .ZN(n214) );
  OAI22_X1 U264 ( .A1(n24), .A2(n214), .B1(n220), .B2(n213), .ZN(n217) );
  XNOR2_X1 U265 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n286 ), .ZN(n219) );
  OAI22_X1 U266 ( .A1(n222), .A2(n219), .B1(n215), .B2(n474), .ZN(n216) );
  NOR2_X1 U267 ( .A1(n230), .A2(n229), .ZN(n289) );
  HA_X1 U268 ( .A(n217), .B(n216), .CO(n229), .S(n227) );
  OR2_X1 U269 ( .A1(\mult_x_1/n288 ), .A2(n471), .ZN(n218) );
  OAI22_X1 U270 ( .A1(n24), .A2(n471), .B1(n218), .B2(n220), .ZN(n226) );
  OR2_X1 U271 ( .A1(n227), .A2(n226), .ZN(n284) );
  XNOR2_X1 U272 ( .A(\mult_x_1/n313 ), .B(\mult_x_1/n287 ), .ZN(n221) );
  OAI22_X1 U273 ( .A1(n222), .A2(n221), .B1(n219), .B2(n474), .ZN(n225) );
  AND2_X1 U274 ( .A1(\mult_x_1/n288 ), .A2(n32), .ZN(n224) );
  NOR2_X1 U275 ( .A1(n225), .A2(n224), .ZN(n276) );
  OAI22_X1 U276 ( .A1(n222), .A2(\mult_x_1/n288 ), .B1(n221), .B2(n474), .ZN(
        n272) );
  OR2_X1 U277 ( .A1(\mult_x_1/n288 ), .A2(n473), .ZN(n223) );
  NAND2_X1 U278 ( .A1(n223), .A2(n222), .ZN(n271) );
  NAND2_X1 U279 ( .A1(n272), .A2(n271), .ZN(n279) );
  NAND2_X1 U280 ( .A1(n225), .A2(n224), .ZN(n277) );
  OAI21_X1 U281 ( .B1(n276), .B2(n279), .A(n277), .ZN(n285) );
  NAND2_X1 U282 ( .A1(n227), .A2(n226), .ZN(n283) );
  INV_X1 U283 ( .A(n283), .ZN(n228) );
  AOI21_X1 U284 ( .B1(n284), .B2(n285), .A(n228), .ZN(n292) );
  NAND2_X1 U285 ( .A1(n230), .A2(n229), .ZN(n290) );
  OAI21_X1 U286 ( .B1(n289), .B2(n292), .A(n290), .ZN(n236) );
  INV_X1 U287 ( .A(n231), .ZN(n232) );
  AOI21_X1 U288 ( .B1(n233), .B2(n236), .A(n232), .ZN(n234) );
  NAND2_X1 U289 ( .A1(n234), .A2(n369), .ZN(n235) );
  NAND2_X1 U290 ( .A1(n247), .A2(n236), .ZN(n237) );
  OAI21_X1 U291 ( .B1(n262), .B2(n442), .A(n237), .ZN(n434) );
  FA_X1 U292 ( .A(n240), .B(n239), .CI(n238), .CO(n248), .S(n241) );
  NAND2_X1 U293 ( .A1(n247), .A2(n241), .ZN(n242) );
  OAI21_X1 U294 ( .B1(n262), .B2(n441), .A(n242), .ZN(n436) );
  FA_X1 U295 ( .A(n27), .B(n243), .CI(n244), .CO(n245), .S(n117) );
  NAND2_X1 U296 ( .A1(n247), .A2(n245), .ZN(n246) );
  OAI21_X1 U297 ( .B1(n262), .B2(n440), .A(n246), .ZN(n438) );
  OR2_X1 U298 ( .A1(n371), .A2(n459), .ZN(n251) );
  OAI21_X1 U299 ( .B1(n248), .B2(n249), .A(n247), .ZN(n250) );
  NAND2_X1 U300 ( .A1(n251), .A2(n250), .ZN(n400) );
  OR2_X1 U301 ( .A1(en), .A2(n455), .ZN(n261) );
  XNOR2_X1 U302 ( .A(n253), .B(n252), .ZN(n255) );
  XNOR2_X1 U303 ( .A(n255), .B(n254), .ZN(n263) );
  NOR2_X1 U304 ( .A1(n263), .A2(n264), .ZN(n259) );
  NAND2_X1 U305 ( .A1(n371), .A2(n259), .ZN(n260) );
  NAND2_X1 U306 ( .A1(n261), .A2(n260), .ZN(n408) );
  OR2_X1 U307 ( .A1(n262), .A2(n444), .ZN(n267) );
  NAND2_X1 U308 ( .A1(n264), .A2(n263), .ZN(n265) );
  NAND2_X1 U309 ( .A1(n371), .A2(n265), .ZN(n266) );
  NAND2_X1 U310 ( .A1(n267), .A2(n266), .ZN(n430) );
  AOI22_X1 U311 ( .A1(n369), .A2(n518), .B1(n519), .B2(n373), .ZN(n521) );
  AOI22_X1 U312 ( .A1(n369), .A2(n517), .B1(n518), .B2(n373), .ZN(n523) );
  AND2_X1 U313 ( .A1(\mult_x_1/n288 ), .A2(\mult_x_1/n180 ), .ZN(n269) );
  NAND2_X1 U314 ( .A1(n369), .A2(n269), .ZN(n270) );
  OAI21_X1 U315 ( .B1(n369), .B2(n517), .A(n270), .ZN(n525) );
  AOI22_X1 U316 ( .A1(n369), .A2(n515), .B1(n516), .B2(n268), .ZN(n527) );
  AOI22_X1 U317 ( .A1(n345), .A2(n514), .B1(n515), .B2(n373), .ZN(n529) );
  OR2_X1 U318 ( .A1(n272), .A2(n271), .ZN(n273) );
  AND2_X1 U319 ( .A1(n273), .A2(n279), .ZN(n274) );
  NAND2_X1 U320 ( .A1(n371), .A2(n274), .ZN(n275) );
  OAI21_X1 U321 ( .B1(n369), .B2(n514), .A(n275), .ZN(n531) );
  AOI22_X1 U322 ( .A1(n369), .A2(n512), .B1(n513), .B2(n373), .ZN(n533) );
  AOI22_X1 U323 ( .A1(n371), .A2(n511), .B1(n512), .B2(n373), .ZN(n535) );
  INV_X1 U324 ( .A(n276), .ZN(n278) );
  NAND2_X1 U325 ( .A1(n278), .A2(n277), .ZN(n280) );
  XOR2_X1 U326 ( .A(n280), .B(n279), .Z(n281) );
  NAND2_X1 U327 ( .A1(n345), .A2(n281), .ZN(n282) );
  OAI21_X1 U328 ( .B1(n371), .B2(n511), .A(n282), .ZN(n537) );
  AOI22_X1 U329 ( .A1(n345), .A2(n509), .B1(n510), .B2(n373), .ZN(n539) );
  AOI22_X1 U330 ( .A1(n369), .A2(n508), .B1(n509), .B2(n373), .ZN(n541) );
  NAND2_X1 U331 ( .A1(n284), .A2(n283), .ZN(n286) );
  XNOR2_X1 U332 ( .A(n286), .B(n285), .ZN(n287) );
  NAND2_X1 U333 ( .A1(n345), .A2(n287), .ZN(n288) );
  OAI21_X1 U334 ( .B1(n369), .B2(n508), .A(n288), .ZN(n543) );
  AOI22_X1 U335 ( .A1(n345), .A2(n506), .B1(n507), .B2(n373), .ZN(n545) );
  AOI22_X1 U336 ( .A1(n345), .A2(n505), .B1(n506), .B2(n373), .ZN(n547) );
  INV_X1 U337 ( .A(n289), .ZN(n291) );
  NAND2_X1 U338 ( .A1(n291), .A2(n290), .ZN(n293) );
  XOR2_X1 U339 ( .A(n293), .B(n292), .Z(n294) );
  NAND2_X1 U340 ( .A1(n371), .A2(n294), .ZN(n295) );
  OAI21_X1 U341 ( .B1(n345), .B2(n505), .A(n295), .ZN(n549) );
  AOI22_X1 U342 ( .A1(n369), .A2(n503), .B1(n504), .B2(n373), .ZN(n551) );
  XNOR2_X1 U343 ( .A(n386), .B(n393), .ZN(n296) );
  NAND2_X1 U344 ( .A1(n369), .A2(n296), .ZN(n297) );
  OAI21_X1 U345 ( .B1(n369), .B2(n503), .A(n297), .ZN(n553) );
  AOI22_X1 U346 ( .A1(n371), .A2(n501), .B1(n502), .B2(n373), .ZN(n555) );
  NAND2_X1 U347 ( .A1(n451), .A2(n385), .ZN(n298) );
  XOR2_X1 U348 ( .A(n298), .B(n392), .Z(n299) );
  NAND2_X1 U349 ( .A1(n369), .A2(n299), .ZN(n300) );
  OAI21_X1 U350 ( .B1(n371), .B2(n501), .A(n300), .ZN(n557) );
  AOI22_X1 U351 ( .A1(n345), .A2(n499), .B1(n500), .B2(n373), .ZN(n559) );
  OAI21_X1 U352 ( .B1(n384), .B2(n392), .A(n385), .ZN(n304) );
  NAND2_X1 U353 ( .A1(n377), .A2(n383), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n304), .B(n301), .ZN(n302) );
  NAND2_X1 U355 ( .A1(n345), .A2(n302), .ZN(n303) );
  OAI21_X1 U356 ( .B1(n369), .B2(n499), .A(n303), .ZN(n561) );
  AOI22_X1 U357 ( .A1(n345), .A2(n497), .B1(n498), .B2(n268), .ZN(n563) );
  AOI21_X1 U358 ( .B1(n304), .B2(n377), .A(n452), .ZN(n308) );
  NAND2_X1 U359 ( .A1(n454), .A2(n382), .ZN(n305) );
  XOR2_X1 U360 ( .A(n308), .B(n305), .Z(n306) );
  NAND2_X1 U361 ( .A1(n345), .A2(n306), .ZN(n307) );
  OAI21_X1 U362 ( .B1(n345), .B2(n497), .A(n307), .ZN(n565) );
  AOI22_X1 U363 ( .A1(n369), .A2(n495), .B1(n496), .B2(n268), .ZN(n567) );
  OAI21_X1 U364 ( .B1(n308), .B2(n381), .A(n382), .ZN(n318) );
  INV_X1 U365 ( .A(n318), .ZN(n312) );
  NAND2_X1 U366 ( .A1(n455), .A2(n391), .ZN(n309) );
  XOR2_X1 U367 ( .A(n312), .B(n309), .Z(n310) );
  NAND2_X1 U368 ( .A1(n345), .A2(n310), .ZN(n311) );
  OAI21_X1 U369 ( .B1(n345), .B2(n495), .A(n311), .ZN(n569) );
  AOI22_X1 U370 ( .A1(n345), .A2(n493), .B1(n494), .B2(n268), .ZN(n571) );
  OAI21_X1 U371 ( .B1(n312), .B2(n380), .A(n391), .ZN(n314) );
  NAND2_X1 U372 ( .A1(n448), .A2(n388), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  NAND2_X1 U374 ( .A1(n369), .A2(n315), .ZN(n316) );
  OAI21_X1 U375 ( .B1(n369), .B2(n493), .A(n316), .ZN(n573) );
  AOI22_X1 U376 ( .A1(n369), .A2(n491), .B1(n492), .B2(n268), .ZN(n575) );
  NOR2_X1 U377 ( .A1(n387), .A2(n380), .ZN(n319) );
  OAI21_X1 U378 ( .B1(n387), .B2(n391), .A(n388), .ZN(n317) );
  AOI21_X1 U379 ( .B1(n319), .B2(n318), .A(n317), .ZN(n350) );
  NOR2_X1 U380 ( .A1(n394), .A2(n395), .ZN(n335) );
  INV_X1 U381 ( .A(n335), .ZN(n327) );
  NAND2_X1 U382 ( .A1(n394), .A2(n395), .ZN(n337) );
  NAND2_X1 U383 ( .A1(n327), .A2(n337), .ZN(n320) );
  XOR2_X1 U384 ( .A(n350), .B(n320), .Z(n321) );
  NAND2_X1 U385 ( .A1(n369), .A2(n321), .ZN(n322) );
  OAI21_X1 U386 ( .B1(n369), .B2(n491), .A(n322), .ZN(n577) );
  AOI22_X1 U387 ( .A1(n345), .A2(n489), .B1(n490), .B2(n268), .ZN(n579) );
  OAI21_X1 U388 ( .B1(n350), .B2(n335), .A(n337), .ZN(n324) );
  NAND2_X1 U389 ( .A1(n376), .A2(n390), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n325) );
  NAND2_X1 U391 ( .A1(n369), .A2(n325), .ZN(n326) );
  OAI21_X1 U392 ( .B1(n366), .B2(n489), .A(n326), .ZN(n581) );
  AOI22_X1 U393 ( .A1(n369), .A2(n487), .B1(n488), .B2(n373), .ZN(n583) );
  NAND2_X1 U394 ( .A1(n327), .A2(n376), .ZN(n330) );
  INV_X1 U395 ( .A(n337), .ZN(n328) );
  AOI21_X1 U396 ( .B1(n328), .B2(n376), .A(n445), .ZN(n329) );
  OAI21_X1 U397 ( .B1(n350), .B2(n330), .A(n329), .ZN(n332) );
  NAND2_X1 U398 ( .A1(n375), .A2(n389), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n333) );
  NAND2_X1 U400 ( .A1(n371), .A2(n333), .ZN(n334) );
  OAI21_X1 U401 ( .B1(n345), .B2(n487), .A(n334), .ZN(n585) );
  AOI22_X1 U402 ( .A1(n371), .A2(n485), .B1(n486), .B2(n373), .ZN(n587) );
  NAND2_X1 U403 ( .A1(n376), .A2(n375), .ZN(n338) );
  NOR2_X1 U404 ( .A1(n335), .A2(n338), .ZN(n346) );
  INV_X1 U405 ( .A(n346), .ZN(n340) );
  AOI21_X1 U406 ( .B1(n445), .B2(n375), .A(n446), .ZN(n336) );
  OAI21_X1 U407 ( .B1(n338), .B2(n337), .A(n336), .ZN(n347) );
  INV_X1 U408 ( .A(n347), .ZN(n339) );
  OAI21_X1 U409 ( .B1(n350), .B2(n340), .A(n339), .ZN(n342) );
  NAND2_X1 U410 ( .A1(n374), .A2(n379), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n342), .B(n341), .ZN(n343) );
  NAND2_X1 U412 ( .A1(n345), .A2(n343), .ZN(n344) );
  OAI21_X1 U413 ( .B1(n369), .B2(n485), .A(n344), .ZN(n589) );
  AOI22_X1 U414 ( .A1(n345), .A2(n483), .B1(n484), .B2(n373), .ZN(n591) );
  NAND2_X1 U415 ( .A1(n346), .A2(n374), .ZN(n349) );
  AOI21_X1 U416 ( .B1(n347), .B2(n374), .A(n456), .ZN(n348) );
  OAI21_X1 U417 ( .B1(n350), .B2(n349), .A(n348), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n351), .B(n378), .ZN(n352) );
  NAND2_X1 U419 ( .A1(n369), .A2(n352), .ZN(n353) );
  OAI21_X1 U420 ( .B1(n371), .B2(n483), .A(n353), .ZN(n593) );
  NAND2_X1 U421 ( .A1(n371), .A2(B_extended[0]), .ZN(n354) );
  OAI21_X1 U422 ( .B1(n345), .B2(n482), .A(n354), .ZN(n595) );
  NAND2_X1 U423 ( .A1(n371), .A2(B_extended[1]), .ZN(n355) );
  OAI21_X1 U424 ( .B1(n345), .B2(n481), .A(n355), .ZN(n597) );
  NAND2_X1 U425 ( .A1(n371), .A2(B_extended[2]), .ZN(n356) );
  OAI21_X1 U426 ( .B1(n369), .B2(n480), .A(n356), .ZN(n599) );
  NAND2_X1 U427 ( .A1(n345), .A2(B_extended[3]), .ZN(n357) );
  OAI21_X1 U428 ( .B1(n366), .B2(n479), .A(n357), .ZN(n601) );
  NAND2_X1 U429 ( .A1(n369), .A2(B_extended[4]), .ZN(n358) );
  OAI21_X1 U430 ( .B1(n345), .B2(n478), .A(n358), .ZN(n603) );
  NAND2_X1 U431 ( .A1(n345), .A2(B_extended[5]), .ZN(n359) );
  OAI21_X1 U432 ( .B1(n345), .B2(n477), .A(n359), .ZN(n605) );
  NAND2_X1 U433 ( .A1(n369), .A2(B_extended[6]), .ZN(n360) );
  OAI21_X1 U434 ( .B1(n371), .B2(n476), .A(n360), .ZN(n607) );
  NAND2_X1 U435 ( .A1(n345), .A2(B_extended[7]), .ZN(n361) );
  OAI21_X1 U436 ( .B1(n369), .B2(n475), .A(n361), .ZN(n609) );
  NAND2_X1 U437 ( .A1(n371), .A2(A_extended[0]), .ZN(n362) );
  OAI21_X1 U438 ( .B1(n345), .B2(n474), .A(n362), .ZN(n611) );
  NAND2_X1 U439 ( .A1(n345), .A2(A_extended[1]), .ZN(n363) );
  OAI21_X1 U440 ( .B1(n369), .B2(n473), .A(n363), .ZN(n613) );
  NAND2_X1 U441 ( .A1(n369), .A2(A_extended[2]), .ZN(n364) );
  OAI21_X1 U442 ( .B1(n345), .B2(n472), .A(n364), .ZN(n615) );
  NAND2_X1 U443 ( .A1(n369), .A2(A_extended[3]), .ZN(n365) );
  OAI21_X1 U444 ( .B1(n369), .B2(n471), .A(n365), .ZN(n617) );
  NAND2_X1 U445 ( .A1(n369), .A2(A_extended[4]), .ZN(n367) );
  OAI21_X1 U446 ( .B1(n369), .B2(n470), .A(n367), .ZN(n619) );
  NAND2_X1 U447 ( .A1(n345), .A2(A_extended[5]), .ZN(n368) );
  OAI21_X1 U448 ( .B1(n371), .B2(n469), .A(n368), .ZN(n621) );
  NAND2_X1 U449 ( .A1(n345), .A2(A_extended[6]), .ZN(n370) );
  OAI21_X1 U450 ( .B1(n345), .B2(n468), .A(n370), .ZN(n623) );
  NAND2_X1 U451 ( .A1(n345), .A2(A_extended[7]), .ZN(n372) );
  OAI21_X1 U452 ( .B1(n345), .B2(n467), .A(n372), .ZN(n625) );
  NAND2_X1 U453 ( .A1(n466), .A2(n373), .ZN(n627) );
endmodule


module conv_128_32 ( clk, reset, s_valid_x, s_valid_f, m_ready_y, s_data_in_x, 
        s_data_in_f, s_ready_f, s_ready_x, m_valid_y, m_data_out_y );
  input [7:0] s_data_in_x;
  input [7:0] s_data_in_f;
  output [20:0] m_data_out_y;
  input clk, reset, s_valid_x, s_valid_f, m_ready_y;
  output s_ready_f, s_ready_x, m_valid_y;
  wire   conv_done, xmem_full, \xmem_data[31][7] , \xmem_data[31][6] ,
         \xmem_data[31][5] , \xmem_data[31][4] , \xmem_data[31][3] ,
         \xmem_data[31][2] , \xmem_data[31][1] , \xmem_data[31][0] ,
         \xmem_data[30][7] , \xmem_data[30][6] , \xmem_data[30][5] ,
         \xmem_data[30][4] , \xmem_data[30][3] , \xmem_data[30][2] ,
         \xmem_data[30][1] , \xmem_data[30][0] , \xmem_data[29][7] ,
         \xmem_data[29][6] , \xmem_data[29][5] , \xmem_data[29][4] ,
         \xmem_data[29][3] , \xmem_data[29][2] , \xmem_data[29][1] ,
         \xmem_data[29][0] , \xmem_data[28][7] , \xmem_data[28][6] ,
         \xmem_data[28][5] , \xmem_data[28][4] , \xmem_data[28][3] ,
         \xmem_data[28][2] , \xmem_data[28][1] , \xmem_data[28][0] ,
         \xmem_data[27][7] , \xmem_data[27][6] , \xmem_data[27][5] ,
         \xmem_data[27][4] , \xmem_data[27][3] , \xmem_data[27][2] ,
         \xmem_data[27][1] , \xmem_data[27][0] , \xmem_data[26][7] ,
         \xmem_data[26][6] , \xmem_data[26][5] , \xmem_data[26][4] ,
         \xmem_data[26][3] , \xmem_data[26][2] , \xmem_data[26][1] ,
         \xmem_data[26][0] , \xmem_data[25][7] , \xmem_data[25][6] ,
         \xmem_data[25][5] , \xmem_data[25][4] , \xmem_data[25][3] ,
         \xmem_data[25][2] , \xmem_data[25][1] , \xmem_data[25][0] ,
         \xmem_data[24][7] , \xmem_data[24][6] , \xmem_data[24][5] ,
         \xmem_data[24][4] , \xmem_data[24][3] , \xmem_data[24][2] ,
         \xmem_data[24][1] , \xmem_data[24][0] , \xmem_data[23][7] ,
         \xmem_data[23][6] , \xmem_data[23][5] , \xmem_data[23][4] ,
         \xmem_data[23][3] , \xmem_data[23][2] , \xmem_data[23][1] ,
         \xmem_data[23][0] , \xmem_data[22][7] , \xmem_data[22][6] ,
         \xmem_data[22][5] , \xmem_data[22][4] , \xmem_data[22][3] ,
         \xmem_data[22][2] , \xmem_data[22][1] , \xmem_data[22][0] ,
         \xmem_data[21][7] , \xmem_data[21][6] , \xmem_data[21][5] ,
         \xmem_data[21][4] , \xmem_data[21][3] , \xmem_data[21][2] ,
         \xmem_data[21][1] , \xmem_data[21][0] , \xmem_data[20][7] ,
         \xmem_data[20][6] , \xmem_data[20][5] , \xmem_data[20][4] ,
         \xmem_data[20][3] , \xmem_data[20][2] , \xmem_data[20][1] ,
         \xmem_data[20][0] , \xmem_data[19][7] , \xmem_data[19][6] ,
         \xmem_data[19][5] , \xmem_data[19][4] , \xmem_data[19][3] ,
         \xmem_data[19][2] , \xmem_data[19][1] , \xmem_data[19][0] ,
         \xmem_data[18][7] , \xmem_data[18][6] , \xmem_data[18][5] ,
         \xmem_data[18][4] , \xmem_data[18][3] , \xmem_data[18][2] ,
         \xmem_data[18][1] , \xmem_data[18][0] , \xmem_data[17][7] ,
         \xmem_data[17][6] , \xmem_data[17][5] , \xmem_data[17][4] ,
         \xmem_data[17][3] , \xmem_data[17][2] , \xmem_data[17][1] ,
         \xmem_data[17][0] , \xmem_data[16][7] , \xmem_data[16][6] ,
         \xmem_data[16][5] , \xmem_data[16][4] , \xmem_data[16][3] ,
         \xmem_data[16][2] , \xmem_data[16][1] , \xmem_data[16][0] ,
         \xmem_data[15][7] , \xmem_data[15][6] , \xmem_data[15][5] ,
         \xmem_data[15][4] , \xmem_data[15][3] , \xmem_data[15][2] ,
         \xmem_data[15][1] , \xmem_data[15][0] , \xmem_data[14][7] ,
         \xmem_data[14][6] , \xmem_data[14][5] , \xmem_data[14][4] ,
         \xmem_data[14][3] , \xmem_data[14][2] , \xmem_data[14][1] ,
         \xmem_data[14][0] , \xmem_data[13][7] , \xmem_data[13][6] ,
         \xmem_data[13][5] , \xmem_data[13][4] , \xmem_data[13][3] ,
         \xmem_data[13][2] , \xmem_data[13][1] , \xmem_data[13][0] ,
         \xmem_data[12][7] , \xmem_data[12][6] , \xmem_data[12][5] ,
         \xmem_data[12][4] , \xmem_data[12][3] , \xmem_data[12][2] ,
         \xmem_data[12][1] , \xmem_data[12][0] , \xmem_data[11][7] ,
         \xmem_data[11][6] , \xmem_data[11][5] , \xmem_data[11][4] ,
         \xmem_data[11][3] , \xmem_data[11][2] , \xmem_data[11][1] ,
         \xmem_data[11][0] , \xmem_data[10][7] , \xmem_data[10][6] ,
         \xmem_data[10][5] , \xmem_data[10][4] , \xmem_data[10][3] ,
         \xmem_data[10][2] , \xmem_data[10][1] , \xmem_data[10][0] ,
         \xmem_data[9][7] , \xmem_data[9][6] , \xmem_data[9][5] ,
         \xmem_data[9][4] , \xmem_data[9][3] , \xmem_data[9][2] ,
         \xmem_data[9][1] , \xmem_data[9][0] , \xmem_data[8][7] ,
         \xmem_data[8][6] , \xmem_data[8][5] , \xmem_data[8][4] ,
         \xmem_data[8][3] , \xmem_data[8][2] , \xmem_data[8][1] ,
         \xmem_data[8][0] , \xmem_data[7][7] , \xmem_data[7][6] ,
         \xmem_data[7][5] , \xmem_data[7][4] , \xmem_data[7][3] ,
         \xmem_data[7][2] , \xmem_data[7][1] , \xmem_data[7][0] ,
         \xmem_data[6][7] , \xmem_data[6][6] , \xmem_data[6][5] ,
         \xmem_data[6][4] , \xmem_data[6][3] , \xmem_data[6][2] ,
         \xmem_data[6][1] , \xmem_data[6][0] , \xmem_data[5][7] ,
         \xmem_data[5][6] , \xmem_data[5][5] , \xmem_data[5][4] ,
         \xmem_data[5][3] , \xmem_data[5][2] , \xmem_data[5][1] ,
         \xmem_data[5][0] , \xmem_data[4][7] , \xmem_data[4][6] ,
         \xmem_data[4][5] , \xmem_data[4][4] , \xmem_data[4][3] ,
         \xmem_data[4][2] , \xmem_data[4][1] , \xmem_data[4][0] ,
         \xmem_data[3][7] , \xmem_data[3][6] , \xmem_data[3][5] ,
         \xmem_data[3][4] , \xmem_data[3][3] , \xmem_data[3][2] ,
         \xmem_data[3][1] , \xmem_data[3][0] , \xmem_data[2][7] ,
         \xmem_data[2][6] , \xmem_data[2][5] , \xmem_data[2][4] ,
         \xmem_data[2][3] , \xmem_data[2][2] , \xmem_data[2][1] ,
         \xmem_data[2][0] , \xmem_data[1][7] , \xmem_data[1][6] ,
         \xmem_data[1][5] , \xmem_data[1][4] , \xmem_data[1][3] ,
         \xmem_data[1][2] , \xmem_data[1][1] , \xmem_data[1][0] ,
         \xmem_data[0][7] , \xmem_data[0][6] , \xmem_data[0][5] ,
         \xmem_data[0][4] , \xmem_data[0][3] , \xmem_data[0][2] ,
         \xmem_data[0][1] , \xmem_data[0][0] , \fmem_data[31][7] ,
         \fmem_data[31][6] , \fmem_data[31][5] , \fmem_data[31][4] ,
         \fmem_data[31][3] , \fmem_data[31][2] , \fmem_data[31][1] ,
         \fmem_data[31][0] , \fmem_data[30][7] , \fmem_data[30][6] ,
         \fmem_data[30][5] , \fmem_data[30][4] , \fmem_data[30][3] ,
         \fmem_data[30][2] , \fmem_data[30][1] , \fmem_data[30][0] ,
         \fmem_data[29][7] , \fmem_data[29][6] , \fmem_data[29][5] ,
         \fmem_data[29][4] , \fmem_data[29][3] , \fmem_data[29][2] ,
         \fmem_data[29][1] , \fmem_data[29][0] , \fmem_data[28][7] ,
         \fmem_data[28][6] , \fmem_data[28][5] , \fmem_data[28][4] ,
         \fmem_data[28][3] , \fmem_data[28][2] , \fmem_data[28][1] ,
         \fmem_data[28][0] , \fmem_data[27][7] , \fmem_data[27][6] ,
         \fmem_data[27][5] , \fmem_data[27][4] , \fmem_data[27][3] ,
         \fmem_data[27][2] , \fmem_data[27][1] , \fmem_data[27][0] ,
         \fmem_data[26][7] , \fmem_data[26][6] , \fmem_data[26][5] ,
         \fmem_data[26][4] , \fmem_data[26][3] , \fmem_data[26][2] ,
         \fmem_data[26][1] , \fmem_data[26][0] , \fmem_data[25][7] ,
         \fmem_data[25][6] , \fmem_data[25][5] , \fmem_data[25][4] ,
         \fmem_data[25][3] , \fmem_data[25][2] , \fmem_data[25][1] ,
         \fmem_data[25][0] , \fmem_data[24][7] , \fmem_data[24][6] ,
         \fmem_data[24][5] , \fmem_data[24][4] , \fmem_data[24][3] ,
         \fmem_data[24][2] , \fmem_data[24][1] , \fmem_data[24][0] ,
         \fmem_data[23][7] , \fmem_data[23][6] , \fmem_data[23][5] ,
         \fmem_data[23][4] , \fmem_data[23][3] , \fmem_data[23][2] ,
         \fmem_data[23][1] , \fmem_data[23][0] , \fmem_data[22][7] ,
         \fmem_data[22][6] , \fmem_data[22][5] , \fmem_data[22][4] ,
         \fmem_data[22][3] , \fmem_data[22][2] , \fmem_data[22][1] ,
         \fmem_data[22][0] , \fmem_data[21][7] , \fmem_data[21][6] ,
         \fmem_data[21][5] , \fmem_data[21][4] , \fmem_data[21][3] ,
         \fmem_data[21][2] , \fmem_data[21][1] , \fmem_data[21][0] ,
         \fmem_data[20][7] , \fmem_data[20][6] , \fmem_data[20][5] ,
         \fmem_data[20][4] , \fmem_data[20][3] , \fmem_data[20][2] ,
         \fmem_data[20][1] , \fmem_data[20][0] , \fmem_data[19][7] ,
         \fmem_data[19][6] , \fmem_data[19][5] , \fmem_data[19][4] ,
         \fmem_data[19][3] , \fmem_data[19][2] , \fmem_data[19][1] ,
         \fmem_data[19][0] , \fmem_data[18][7] , \fmem_data[18][6] ,
         \fmem_data[18][5] , \fmem_data[18][4] , \fmem_data[18][3] ,
         \fmem_data[18][2] , \fmem_data[18][1] , \fmem_data[18][0] ,
         \fmem_data[17][7] , \fmem_data[17][6] , \fmem_data[17][5] ,
         \fmem_data[17][4] , \fmem_data[17][3] , \fmem_data[17][2] ,
         \fmem_data[17][1] , \fmem_data[17][0] , \fmem_data[16][7] ,
         \fmem_data[16][6] , \fmem_data[16][5] , \fmem_data[16][4] ,
         \fmem_data[16][3] , \fmem_data[16][2] , \fmem_data[16][1] ,
         \fmem_data[16][0] , \fmem_data[15][7] , \fmem_data[15][6] ,
         \fmem_data[15][5] , \fmem_data[15][4] , \fmem_data[15][3] ,
         \fmem_data[15][2] , \fmem_data[15][1] , \fmem_data[15][0] ,
         \fmem_data[14][7] , \fmem_data[14][6] , \fmem_data[14][5] ,
         \fmem_data[14][4] , \fmem_data[14][3] , \fmem_data[14][2] ,
         \fmem_data[14][1] , \fmem_data[14][0] , \fmem_data[13][7] ,
         \fmem_data[13][6] , \fmem_data[13][5] , \fmem_data[13][4] ,
         \fmem_data[13][3] , \fmem_data[13][2] , \fmem_data[13][1] ,
         \fmem_data[13][0] , \fmem_data[12][7] , \fmem_data[12][6] ,
         \fmem_data[12][5] , \fmem_data[12][4] , \fmem_data[12][3] ,
         \fmem_data[12][2] , \fmem_data[12][1] , \fmem_data[12][0] ,
         \fmem_data[11][7] , \fmem_data[11][6] , \fmem_data[11][5] ,
         \fmem_data[11][4] , \fmem_data[11][3] , \fmem_data[11][2] ,
         \fmem_data[11][1] , \fmem_data[11][0] , \fmem_data[10][7] ,
         \fmem_data[10][6] , \fmem_data[10][5] , \fmem_data[10][4] ,
         \fmem_data[10][3] , \fmem_data[10][2] , \fmem_data[10][1] ,
         \fmem_data[10][0] , \fmem_data[9][7] , \fmem_data[9][6] ,
         \fmem_data[9][5] , \fmem_data[9][4] , \fmem_data[9][3] ,
         \fmem_data[9][2] , \fmem_data[9][1] , \fmem_data[9][0] ,
         \fmem_data[8][7] , \fmem_data[8][6] , \fmem_data[8][5] ,
         \fmem_data[8][4] , \fmem_data[8][3] , \fmem_data[8][2] ,
         \fmem_data[8][1] , \fmem_data[8][0] , \fmem_data[7][7] ,
         \fmem_data[7][6] , \fmem_data[7][5] , \fmem_data[7][4] ,
         \fmem_data[7][3] , \fmem_data[7][2] , \fmem_data[7][1] ,
         \fmem_data[7][0] , \fmem_data[6][7] , \fmem_data[6][6] ,
         \fmem_data[6][5] , \fmem_data[6][4] , \fmem_data[6][3] ,
         \fmem_data[6][2] , \fmem_data[6][1] , \fmem_data[6][0] ,
         \fmem_data[5][7] , \fmem_data[5][6] , \fmem_data[5][5] ,
         \fmem_data[5][4] , \fmem_data[5][3] , \fmem_data[5][2] ,
         \fmem_data[5][1] , \fmem_data[5][0] , \fmem_data[4][7] ,
         \fmem_data[4][6] , \fmem_data[4][5] , \fmem_data[4][4] ,
         \fmem_data[4][3] , \fmem_data[4][2] , \fmem_data[4][1] ,
         \fmem_data[4][0] , \fmem_data[3][7] , \fmem_data[3][6] ,
         \fmem_data[3][5] , \fmem_data[3][4] , \fmem_data[3][3] ,
         \fmem_data[3][2] , \fmem_data[3][1] , \fmem_data[3][0] ,
         \fmem_data[2][7] , \fmem_data[2][6] , \fmem_data[2][5] ,
         \fmem_data[2][4] , \fmem_data[2][3] , \fmem_data[2][2] ,
         \fmem_data[2][1] , \fmem_data[2][0] , \fmem_data[1][7] ,
         \fmem_data[1][6] , \fmem_data[1][5] , \fmem_data[1][4] ,
         \fmem_data[1][3] , \fmem_data[1][2] , \fmem_data[1][1] ,
         \fmem_data[1][0] , \fmem_data[0][7] , \fmem_data[0][6] ,
         \fmem_data[0][5] , \fmem_data[0][4] , \fmem_data[0][3] ,
         \fmem_data[0][2] , \fmem_data[0][1] , \fmem_data[0][0] ,
         \x_mult_f_int[31][15] , \x_mult_f_int[31][14] ,
         \x_mult_f_int[31][13] , \x_mult_f_int[31][12] ,
         \x_mult_f_int[31][11] , \x_mult_f_int[31][10] , \x_mult_f_int[31][9] ,
         \x_mult_f_int[31][8] , \x_mult_f_int[31][7] , \x_mult_f_int[31][6] ,
         \x_mult_f_int[31][5] , \x_mult_f_int[31][4] , \x_mult_f_int[31][3] ,
         \x_mult_f_int[31][2] , \x_mult_f_int[31][1] , \x_mult_f_int[31][0] ,
         \x_mult_f_int[30][15] , \x_mult_f_int[30][14] ,
         \x_mult_f_int[30][13] , \x_mult_f_int[30][12] ,
         \x_mult_f_int[30][11] , \x_mult_f_int[30][10] , \x_mult_f_int[30][9] ,
         \x_mult_f_int[30][8] , \x_mult_f_int[30][7] , \x_mult_f_int[30][6] ,
         \x_mult_f_int[30][5] , \x_mult_f_int[30][4] , \x_mult_f_int[30][3] ,
         \x_mult_f_int[30][2] , \x_mult_f_int[30][1] , \x_mult_f_int[30][0] ,
         \x_mult_f_int[29][15] , \x_mult_f_int[29][14] ,
         \x_mult_f_int[29][13] , \x_mult_f_int[29][12] ,
         \x_mult_f_int[29][11] , \x_mult_f_int[29][10] , \x_mult_f_int[29][9] ,
         \x_mult_f_int[29][8] , \x_mult_f_int[29][7] , \x_mult_f_int[29][6] ,
         \x_mult_f_int[29][5] , \x_mult_f_int[29][4] , \x_mult_f_int[29][3] ,
         \x_mult_f_int[29][2] , \x_mult_f_int[29][1] , \x_mult_f_int[29][0] ,
         \x_mult_f_int[28][15] , \x_mult_f_int[28][14] ,
         \x_mult_f_int[28][13] , \x_mult_f_int[28][12] ,
         \x_mult_f_int[28][11] , \x_mult_f_int[28][10] , \x_mult_f_int[28][9] ,
         \x_mult_f_int[28][8] , \x_mult_f_int[28][7] , \x_mult_f_int[28][6] ,
         \x_mult_f_int[28][5] , \x_mult_f_int[28][4] , \x_mult_f_int[28][3] ,
         \x_mult_f_int[28][2] , \x_mult_f_int[28][1] , \x_mult_f_int[28][0] ,
         \x_mult_f_int[27][15] , \x_mult_f_int[27][14] ,
         \x_mult_f_int[27][13] , \x_mult_f_int[27][12] ,
         \x_mult_f_int[27][11] , \x_mult_f_int[27][10] , \x_mult_f_int[27][9] ,
         \x_mult_f_int[27][8] , \x_mult_f_int[27][7] , \x_mult_f_int[27][6] ,
         \x_mult_f_int[27][5] , \x_mult_f_int[27][4] , \x_mult_f_int[27][3] ,
         \x_mult_f_int[27][2] , \x_mult_f_int[27][1] , \x_mult_f_int[27][0] ,
         \x_mult_f_int[26][15] , \x_mult_f_int[26][14] ,
         \x_mult_f_int[26][13] , \x_mult_f_int[26][12] ,
         \x_mult_f_int[26][11] , \x_mult_f_int[26][10] , \x_mult_f_int[26][9] ,
         \x_mult_f_int[26][8] , \x_mult_f_int[26][7] , \x_mult_f_int[26][6] ,
         \x_mult_f_int[26][5] , \x_mult_f_int[26][4] , \x_mult_f_int[26][3] ,
         \x_mult_f_int[26][2] , \x_mult_f_int[26][1] , \x_mult_f_int[26][0] ,
         \x_mult_f_int[25][15] , \x_mult_f_int[25][14] ,
         \x_mult_f_int[25][13] , \x_mult_f_int[25][12] ,
         \x_mult_f_int[25][11] , \x_mult_f_int[25][10] , \x_mult_f_int[25][9] ,
         \x_mult_f_int[25][8] , \x_mult_f_int[25][7] , \x_mult_f_int[25][6] ,
         \x_mult_f_int[25][5] , \x_mult_f_int[25][4] , \x_mult_f_int[25][3] ,
         \x_mult_f_int[25][2] , \x_mult_f_int[25][1] , \x_mult_f_int[25][0] ,
         \x_mult_f_int[24][15] , \x_mult_f_int[24][14] ,
         \x_mult_f_int[24][13] , \x_mult_f_int[24][12] ,
         \x_mult_f_int[24][11] , \x_mult_f_int[24][10] , \x_mult_f_int[24][9] ,
         \x_mult_f_int[24][8] , \x_mult_f_int[24][7] , \x_mult_f_int[24][6] ,
         \x_mult_f_int[24][5] , \x_mult_f_int[24][4] , \x_mult_f_int[24][3] ,
         \x_mult_f_int[24][2] , \x_mult_f_int[24][1] , \x_mult_f_int[24][0] ,
         \x_mult_f_int[23][15] , \x_mult_f_int[23][14] ,
         \x_mult_f_int[23][13] , \x_mult_f_int[23][12] ,
         \x_mult_f_int[23][11] , \x_mult_f_int[23][10] , \x_mult_f_int[23][9] ,
         \x_mult_f_int[23][8] , \x_mult_f_int[23][7] , \x_mult_f_int[23][6] ,
         \x_mult_f_int[23][5] , \x_mult_f_int[23][4] , \x_mult_f_int[23][3] ,
         \x_mult_f_int[23][2] , \x_mult_f_int[23][1] , \x_mult_f_int[23][0] ,
         \x_mult_f_int[22][15] , \x_mult_f_int[22][14] ,
         \x_mult_f_int[22][13] , \x_mult_f_int[22][12] ,
         \x_mult_f_int[22][11] , \x_mult_f_int[22][10] , \x_mult_f_int[22][9] ,
         \x_mult_f_int[22][8] , \x_mult_f_int[22][7] , \x_mult_f_int[22][6] ,
         \x_mult_f_int[22][5] , \x_mult_f_int[22][4] , \x_mult_f_int[22][3] ,
         \x_mult_f_int[22][2] , \x_mult_f_int[22][1] , \x_mult_f_int[22][0] ,
         \x_mult_f_int[21][15] , \x_mult_f_int[21][14] ,
         \x_mult_f_int[21][13] , \x_mult_f_int[21][12] ,
         \x_mult_f_int[21][11] , \x_mult_f_int[21][10] , \x_mult_f_int[21][9] ,
         \x_mult_f_int[21][8] , \x_mult_f_int[21][7] , \x_mult_f_int[21][6] ,
         \x_mult_f_int[21][5] , \x_mult_f_int[21][4] , \x_mult_f_int[21][3] ,
         \x_mult_f_int[21][2] , \x_mult_f_int[21][1] , \x_mult_f_int[21][0] ,
         \x_mult_f_int[20][15] , \x_mult_f_int[20][14] ,
         \x_mult_f_int[20][13] , \x_mult_f_int[20][12] ,
         \x_mult_f_int[20][11] , \x_mult_f_int[20][10] , \x_mult_f_int[20][9] ,
         \x_mult_f_int[20][8] , \x_mult_f_int[20][7] , \x_mult_f_int[20][6] ,
         \x_mult_f_int[20][5] , \x_mult_f_int[20][4] , \x_mult_f_int[20][3] ,
         \x_mult_f_int[20][2] , \x_mult_f_int[20][1] , \x_mult_f_int[20][0] ,
         \x_mult_f_int[19][15] , \x_mult_f_int[19][14] ,
         \x_mult_f_int[19][13] , \x_mult_f_int[19][12] ,
         \x_mult_f_int[19][11] , \x_mult_f_int[19][10] , \x_mult_f_int[19][9] ,
         \x_mult_f_int[19][8] , \x_mult_f_int[19][7] , \x_mult_f_int[19][6] ,
         \x_mult_f_int[19][5] , \x_mult_f_int[19][4] , \x_mult_f_int[19][3] ,
         \x_mult_f_int[19][2] , \x_mult_f_int[19][1] , \x_mult_f_int[19][0] ,
         \x_mult_f_int[18][15] , \x_mult_f_int[18][14] ,
         \x_mult_f_int[18][13] , \x_mult_f_int[18][12] ,
         \x_mult_f_int[18][11] , \x_mult_f_int[18][10] , \x_mult_f_int[18][9] ,
         \x_mult_f_int[18][8] , \x_mult_f_int[18][7] , \x_mult_f_int[18][6] ,
         \x_mult_f_int[18][5] , \x_mult_f_int[18][4] , \x_mult_f_int[18][3] ,
         \x_mult_f_int[18][2] , \x_mult_f_int[18][1] , \x_mult_f_int[18][0] ,
         \x_mult_f_int[17][15] , \x_mult_f_int[17][14] ,
         \x_mult_f_int[17][13] , \x_mult_f_int[17][12] ,
         \x_mult_f_int[17][11] , \x_mult_f_int[17][10] , \x_mult_f_int[17][9] ,
         \x_mult_f_int[17][8] , \x_mult_f_int[17][7] , \x_mult_f_int[17][6] ,
         \x_mult_f_int[17][5] , \x_mult_f_int[17][4] , \x_mult_f_int[17][3] ,
         \x_mult_f_int[17][2] , \x_mult_f_int[17][1] , \x_mult_f_int[17][0] ,
         \x_mult_f_int[16][15] , \x_mult_f_int[16][14] ,
         \x_mult_f_int[16][13] , \x_mult_f_int[16][12] ,
         \x_mult_f_int[16][11] , \x_mult_f_int[16][10] , \x_mult_f_int[16][9] ,
         \x_mult_f_int[16][8] , \x_mult_f_int[16][7] , \x_mult_f_int[16][6] ,
         \x_mult_f_int[16][5] , \x_mult_f_int[16][4] , \x_mult_f_int[16][3] ,
         \x_mult_f_int[16][2] , \x_mult_f_int[16][1] , \x_mult_f_int[16][0] ,
         \x_mult_f_int[15][15] , \x_mult_f_int[15][14] ,
         \x_mult_f_int[15][13] , \x_mult_f_int[15][12] ,
         \x_mult_f_int[15][11] , \x_mult_f_int[15][10] , \x_mult_f_int[15][9] ,
         \x_mult_f_int[15][8] , \x_mult_f_int[15][7] , \x_mult_f_int[15][6] ,
         \x_mult_f_int[15][5] , \x_mult_f_int[15][4] , \x_mult_f_int[15][3] ,
         \x_mult_f_int[15][2] , \x_mult_f_int[15][1] , \x_mult_f_int[15][0] ,
         \x_mult_f_int[14][15] , \x_mult_f_int[14][14] ,
         \x_mult_f_int[14][13] , \x_mult_f_int[14][12] ,
         \x_mult_f_int[14][11] , \x_mult_f_int[14][10] , \x_mult_f_int[14][9] ,
         \x_mult_f_int[14][8] , \x_mult_f_int[14][7] , \x_mult_f_int[14][6] ,
         \x_mult_f_int[14][5] , \x_mult_f_int[14][4] , \x_mult_f_int[14][3] ,
         \x_mult_f_int[14][2] , \x_mult_f_int[14][1] , \x_mult_f_int[14][0] ,
         \x_mult_f_int[13][15] , \x_mult_f_int[13][14] ,
         \x_mult_f_int[13][13] , \x_mult_f_int[13][12] ,
         \x_mult_f_int[13][11] , \x_mult_f_int[13][10] , \x_mult_f_int[13][9] ,
         \x_mult_f_int[13][8] , \x_mult_f_int[13][7] , \x_mult_f_int[13][6] ,
         \x_mult_f_int[13][5] , \x_mult_f_int[13][4] , \x_mult_f_int[13][3] ,
         \x_mult_f_int[13][2] , \x_mult_f_int[13][1] , \x_mult_f_int[13][0] ,
         \x_mult_f_int[12][15] , \x_mult_f_int[12][14] ,
         \x_mult_f_int[12][13] , \x_mult_f_int[12][12] ,
         \x_mult_f_int[12][11] , \x_mult_f_int[12][10] , \x_mult_f_int[12][9] ,
         \x_mult_f_int[12][8] , \x_mult_f_int[12][7] , \x_mult_f_int[12][6] ,
         \x_mult_f_int[12][5] , \x_mult_f_int[12][4] , \x_mult_f_int[12][3] ,
         \x_mult_f_int[12][2] , \x_mult_f_int[12][1] , \x_mult_f_int[12][0] ,
         \x_mult_f_int[11][15] , \x_mult_f_int[11][14] ,
         \x_mult_f_int[11][13] , \x_mult_f_int[11][12] ,
         \x_mult_f_int[11][11] , \x_mult_f_int[11][10] , \x_mult_f_int[11][9] ,
         \x_mult_f_int[11][8] , \x_mult_f_int[11][7] , \x_mult_f_int[11][6] ,
         \x_mult_f_int[11][5] , \x_mult_f_int[11][4] , \x_mult_f_int[11][3] ,
         \x_mult_f_int[11][2] , \x_mult_f_int[11][1] , \x_mult_f_int[11][0] ,
         \x_mult_f_int[10][15] , \x_mult_f_int[10][14] ,
         \x_mult_f_int[10][13] , \x_mult_f_int[10][12] ,
         \x_mult_f_int[10][11] , \x_mult_f_int[10][10] , \x_mult_f_int[10][9] ,
         \x_mult_f_int[10][8] , \x_mult_f_int[10][7] , \x_mult_f_int[10][6] ,
         \x_mult_f_int[10][5] , \x_mult_f_int[10][4] , \x_mult_f_int[10][3] ,
         \x_mult_f_int[10][2] , \x_mult_f_int[10][1] , \x_mult_f_int[10][0] ,
         \x_mult_f_int[9][15] , \x_mult_f_int[9][14] , \x_mult_f_int[9][13] ,
         \x_mult_f_int[9][12] , \x_mult_f_int[9][11] , \x_mult_f_int[9][10] ,
         \x_mult_f_int[9][9] , \x_mult_f_int[9][8] , \x_mult_f_int[9][7] ,
         \x_mult_f_int[9][6] , \x_mult_f_int[9][5] , \x_mult_f_int[9][4] ,
         \x_mult_f_int[9][3] , \x_mult_f_int[9][2] , \x_mult_f_int[9][1] ,
         \x_mult_f_int[9][0] , \x_mult_f_int[8][15] , \x_mult_f_int[8][14] ,
         \x_mult_f_int[8][13] , \x_mult_f_int[8][12] , \x_mult_f_int[8][11] ,
         \x_mult_f_int[8][10] , \x_mult_f_int[8][9] , \x_mult_f_int[8][8] ,
         \x_mult_f_int[8][7] , \x_mult_f_int[8][6] , \x_mult_f_int[8][5] ,
         \x_mult_f_int[8][4] , \x_mult_f_int[8][3] , \x_mult_f_int[8][2] ,
         \x_mult_f_int[8][1] , \x_mult_f_int[8][0] , \x_mult_f_int[7][15] ,
         \x_mult_f_int[7][14] , \x_mult_f_int[7][13] , \x_mult_f_int[7][12] ,
         \x_mult_f_int[7][11] , \x_mult_f_int[7][10] , \x_mult_f_int[7][9] ,
         \x_mult_f_int[7][8] , \x_mult_f_int[7][7] , \x_mult_f_int[7][6] ,
         \x_mult_f_int[7][5] , \x_mult_f_int[7][4] , \x_mult_f_int[7][3] ,
         \x_mult_f_int[7][2] , \x_mult_f_int[7][1] , \x_mult_f_int[7][0] ,
         \x_mult_f_int[6][15] , \x_mult_f_int[6][14] , \x_mult_f_int[6][13] ,
         \x_mult_f_int[6][12] , \x_mult_f_int[6][11] , \x_mult_f_int[6][10] ,
         \x_mult_f_int[6][9] , \x_mult_f_int[6][8] , \x_mult_f_int[6][7] ,
         \x_mult_f_int[6][6] , \x_mult_f_int[6][5] , \x_mult_f_int[6][4] ,
         \x_mult_f_int[6][3] , \x_mult_f_int[6][2] , \x_mult_f_int[6][1] ,
         \x_mult_f_int[6][0] , \x_mult_f_int[5][15] , \x_mult_f_int[5][14] ,
         \x_mult_f_int[5][13] , \x_mult_f_int[5][12] , \x_mult_f_int[5][11] ,
         \x_mult_f_int[5][10] , \x_mult_f_int[5][9] , \x_mult_f_int[5][8] ,
         \x_mult_f_int[5][7] , \x_mult_f_int[5][6] , \x_mult_f_int[5][5] ,
         \x_mult_f_int[5][4] , \x_mult_f_int[5][3] , \x_mult_f_int[5][2] ,
         \x_mult_f_int[5][1] , \x_mult_f_int[5][0] , \x_mult_f_int[4][15] ,
         \x_mult_f_int[4][14] , \x_mult_f_int[4][13] , \x_mult_f_int[4][12] ,
         \x_mult_f_int[4][11] , \x_mult_f_int[4][10] , \x_mult_f_int[4][9] ,
         \x_mult_f_int[4][8] , \x_mult_f_int[4][7] , \x_mult_f_int[4][6] ,
         \x_mult_f_int[4][5] , \x_mult_f_int[4][4] , \x_mult_f_int[4][3] ,
         \x_mult_f_int[4][2] , \x_mult_f_int[4][1] , \x_mult_f_int[4][0] ,
         \x_mult_f_int[3][15] , \x_mult_f_int[3][14] , \x_mult_f_int[3][13] ,
         \x_mult_f_int[3][12] , \x_mult_f_int[3][11] , \x_mult_f_int[3][10] ,
         \x_mult_f_int[3][9] , \x_mult_f_int[3][8] , \x_mult_f_int[3][7] ,
         \x_mult_f_int[3][6] , \x_mult_f_int[3][5] , \x_mult_f_int[3][4] ,
         \x_mult_f_int[3][3] , \x_mult_f_int[3][2] , \x_mult_f_int[3][1] ,
         \x_mult_f_int[3][0] , \x_mult_f_int[2][15] , \x_mult_f_int[2][14] ,
         \x_mult_f_int[2][13] , \x_mult_f_int[2][12] , \x_mult_f_int[2][11] ,
         \x_mult_f_int[2][10] , \x_mult_f_int[2][9] , \x_mult_f_int[2][8] ,
         \x_mult_f_int[2][7] , \x_mult_f_int[2][6] , \x_mult_f_int[2][5] ,
         \x_mult_f_int[2][4] , \x_mult_f_int[2][3] , \x_mult_f_int[2][2] ,
         \x_mult_f_int[2][1] , \x_mult_f_int[2][0] , \x_mult_f_int[1][15] ,
         \x_mult_f_int[1][14] , \x_mult_f_int[1][13] , \x_mult_f_int[1][12] ,
         \x_mult_f_int[1][11] , \x_mult_f_int[1][10] , \x_mult_f_int[1][9] ,
         \x_mult_f_int[1][8] , \x_mult_f_int[1][7] , \x_mult_f_int[1][6] ,
         \x_mult_f_int[1][5] , \x_mult_f_int[1][4] , \x_mult_f_int[1][3] ,
         \x_mult_f_int[1][2] , \x_mult_f_int[1][1] , \x_mult_f_int[1][0] ,
         \x_mult_f_int[0][15] , \x_mult_f_int[0][14] , \x_mult_f_int[0][13] ,
         \x_mult_f_int[0][12] , \x_mult_f_int[0][11] , \x_mult_f_int[0][10] ,
         \x_mult_f_int[0][9] , \x_mult_f_int[0][8] , \x_mult_f_int[0][7] ,
         \x_mult_f_int[0][6] , \x_mult_f_int[0][5] , \x_mult_f_int[0][4] ,
         \x_mult_f_int[0][3] , \x_mult_f_int[0][2] , \x_mult_f_int[0][1] ,
         \x_mult_f_int[0][0] , \x_mult_f[31][15] , \x_mult_f[31][14] ,
         \x_mult_f[31][13] , \x_mult_f[31][12] , \x_mult_f[31][11] ,
         \x_mult_f[31][10] , \x_mult_f[31][9] , \x_mult_f[31][8] ,
         \x_mult_f[31][7] , \x_mult_f[31][6] , \x_mult_f[31][5] ,
         \x_mult_f[31][4] , \x_mult_f[31][3] , \x_mult_f[31][2] ,
         \x_mult_f[31][1] , \x_mult_f[31][0] , \x_mult_f[30][15] ,
         \x_mult_f[30][14] , \x_mult_f[30][13] , \x_mult_f[30][12] ,
         \x_mult_f[30][11] , \x_mult_f[30][10] , \x_mult_f[30][9] ,
         \x_mult_f[30][8] , \x_mult_f[30][7] , \x_mult_f[30][6] ,
         \x_mult_f[30][5] , \x_mult_f[30][4] , \x_mult_f[30][3] ,
         \x_mult_f[30][2] , \x_mult_f[30][1] , \x_mult_f[30][0] ,
         \x_mult_f[29][15] , \x_mult_f[29][14] , \x_mult_f[29][13] ,
         \x_mult_f[29][12] , \x_mult_f[29][11] , \x_mult_f[29][10] ,
         \x_mult_f[29][9] , \x_mult_f[29][8] , \x_mult_f[29][7] ,
         \x_mult_f[29][6] , \x_mult_f[29][5] , \x_mult_f[29][4] ,
         \x_mult_f[29][3] , \x_mult_f[29][2] , \x_mult_f[29][1] ,
         \x_mult_f[29][0] , \x_mult_f[28][15] , \x_mult_f[28][14] ,
         \x_mult_f[28][13] , \x_mult_f[28][12] , \x_mult_f[28][11] ,
         \x_mult_f[28][10] , \x_mult_f[28][9] , \x_mult_f[28][8] ,
         \x_mult_f[28][7] , \x_mult_f[28][6] , \x_mult_f[28][5] ,
         \x_mult_f[28][4] , \x_mult_f[28][3] , \x_mult_f[28][2] ,
         \x_mult_f[28][1] , \x_mult_f[28][0] , \x_mult_f[27][15] ,
         \x_mult_f[27][14] , \x_mult_f[27][13] , \x_mult_f[27][12] ,
         \x_mult_f[27][11] , \x_mult_f[27][10] , \x_mult_f[27][9] ,
         \x_mult_f[27][8] , \x_mult_f[27][7] , \x_mult_f[27][6] ,
         \x_mult_f[27][5] , \x_mult_f[27][4] , \x_mult_f[27][3] ,
         \x_mult_f[27][2] , \x_mult_f[27][1] , \x_mult_f[27][0] ,
         \x_mult_f[26][15] , \x_mult_f[26][14] , \x_mult_f[26][13] ,
         \x_mult_f[26][12] , \x_mult_f[26][11] , \x_mult_f[26][10] ,
         \x_mult_f[26][9] , \x_mult_f[26][8] , \x_mult_f[26][7] ,
         \x_mult_f[26][6] , \x_mult_f[26][5] , \x_mult_f[26][4] ,
         \x_mult_f[26][3] , \x_mult_f[26][2] , \x_mult_f[26][1] ,
         \x_mult_f[26][0] , \x_mult_f[25][15] , \x_mult_f[25][14] ,
         \x_mult_f[25][13] , \x_mult_f[25][12] , \x_mult_f[25][11] ,
         \x_mult_f[25][10] , \x_mult_f[25][9] , \x_mult_f[25][8] ,
         \x_mult_f[25][7] , \x_mult_f[25][6] , \x_mult_f[25][5] ,
         \x_mult_f[25][4] , \x_mult_f[25][3] , \x_mult_f[25][2] ,
         \x_mult_f[25][1] , \x_mult_f[25][0] , \x_mult_f[24][15] ,
         \x_mult_f[24][14] , \x_mult_f[24][13] , \x_mult_f[24][12] ,
         \x_mult_f[24][11] , \x_mult_f[24][10] , \x_mult_f[24][9] ,
         \x_mult_f[24][8] , \x_mult_f[24][7] , \x_mult_f[24][6] ,
         \x_mult_f[24][5] , \x_mult_f[24][4] , \x_mult_f[24][3] ,
         \x_mult_f[24][2] , \x_mult_f[24][1] , \x_mult_f[24][0] ,
         \x_mult_f[23][15] , \x_mult_f[23][14] , \x_mult_f[23][13] ,
         \x_mult_f[23][12] , \x_mult_f[23][11] , \x_mult_f[23][10] ,
         \x_mult_f[23][9] , \x_mult_f[23][8] , \x_mult_f[23][7] ,
         \x_mult_f[23][6] , \x_mult_f[23][5] , \x_mult_f[23][4] ,
         \x_mult_f[23][3] , \x_mult_f[23][2] , \x_mult_f[23][1] ,
         \x_mult_f[23][0] , \x_mult_f[22][15] , \x_mult_f[22][14] ,
         \x_mult_f[22][13] , \x_mult_f[22][12] , \x_mult_f[22][11] ,
         \x_mult_f[22][10] , \x_mult_f[22][9] , \x_mult_f[22][8] ,
         \x_mult_f[22][7] , \x_mult_f[22][6] , \x_mult_f[22][5] ,
         \x_mult_f[22][4] , \x_mult_f[22][3] , \x_mult_f[22][2] ,
         \x_mult_f[22][1] , \x_mult_f[22][0] , \x_mult_f[21][15] ,
         \x_mult_f[21][14] , \x_mult_f[21][13] , \x_mult_f[21][12] ,
         \x_mult_f[21][11] , \x_mult_f[21][10] , \x_mult_f[21][9] ,
         \x_mult_f[21][8] , \x_mult_f[21][7] , \x_mult_f[21][6] ,
         \x_mult_f[21][5] , \x_mult_f[21][4] , \x_mult_f[21][3] ,
         \x_mult_f[21][2] , \x_mult_f[21][1] , \x_mult_f[21][0] ,
         \x_mult_f[20][15] , \x_mult_f[20][14] , \x_mult_f[20][13] ,
         \x_mult_f[20][12] , \x_mult_f[20][11] , \x_mult_f[20][10] ,
         \x_mult_f[20][9] , \x_mult_f[20][8] , \x_mult_f[20][7] ,
         \x_mult_f[20][6] , \x_mult_f[20][5] , \x_mult_f[20][4] ,
         \x_mult_f[20][3] , \x_mult_f[20][2] , \x_mult_f[20][1] ,
         \x_mult_f[20][0] , \x_mult_f[19][15] , \x_mult_f[19][14] ,
         \x_mult_f[19][13] , \x_mult_f[19][12] , \x_mult_f[19][11] ,
         \x_mult_f[19][10] , \x_mult_f[19][9] , \x_mult_f[19][8] ,
         \x_mult_f[19][7] , \x_mult_f[19][6] , \x_mult_f[19][5] ,
         \x_mult_f[19][4] , \x_mult_f[19][3] , \x_mult_f[19][2] ,
         \x_mult_f[19][1] , \x_mult_f[19][0] , \x_mult_f[18][15] ,
         \x_mult_f[18][14] , \x_mult_f[18][13] , \x_mult_f[18][12] ,
         \x_mult_f[18][11] , \x_mult_f[18][10] , \x_mult_f[18][9] ,
         \x_mult_f[18][8] , \x_mult_f[18][7] , \x_mult_f[18][6] ,
         \x_mult_f[18][5] , \x_mult_f[18][4] , \x_mult_f[18][3] ,
         \x_mult_f[18][2] , \x_mult_f[18][1] , \x_mult_f[18][0] ,
         \x_mult_f[17][15] , \x_mult_f[17][14] , \x_mult_f[17][13] ,
         \x_mult_f[17][12] , \x_mult_f[17][11] , \x_mult_f[17][10] ,
         \x_mult_f[17][9] , \x_mult_f[17][8] , \x_mult_f[17][7] ,
         \x_mult_f[17][6] , \x_mult_f[17][5] , \x_mult_f[17][4] ,
         \x_mult_f[17][3] , \x_mult_f[17][2] , \x_mult_f[17][1] ,
         \x_mult_f[17][0] , \x_mult_f[16][15] , \x_mult_f[16][14] ,
         \x_mult_f[16][13] , \x_mult_f[16][12] , \x_mult_f[16][11] ,
         \x_mult_f[16][10] , \x_mult_f[16][9] , \x_mult_f[16][8] ,
         \x_mult_f[16][7] , \x_mult_f[16][6] , \x_mult_f[16][5] ,
         \x_mult_f[16][4] , \x_mult_f[16][3] , \x_mult_f[16][2] ,
         \x_mult_f[16][1] , \x_mult_f[16][0] , \x_mult_f[15][15] ,
         \x_mult_f[15][14] , \x_mult_f[15][13] , \x_mult_f[15][12] ,
         \x_mult_f[15][11] , \x_mult_f[15][10] , \x_mult_f[15][9] ,
         \x_mult_f[15][8] , \x_mult_f[15][7] , \x_mult_f[15][6] ,
         \x_mult_f[15][5] , \x_mult_f[15][4] , \x_mult_f[15][3] ,
         \x_mult_f[15][2] , \x_mult_f[15][1] , \x_mult_f[15][0] ,
         \x_mult_f[14][15] , \x_mult_f[14][14] , \x_mult_f[14][13] ,
         \x_mult_f[14][12] , \x_mult_f[14][11] , \x_mult_f[14][10] ,
         \x_mult_f[14][9] , \x_mult_f[14][8] , \x_mult_f[14][7] ,
         \x_mult_f[14][6] , \x_mult_f[14][5] , \x_mult_f[14][4] ,
         \x_mult_f[14][3] , \x_mult_f[14][2] , \x_mult_f[14][1] ,
         \x_mult_f[14][0] , \x_mult_f[13][15] , \x_mult_f[13][14] ,
         \x_mult_f[13][13] , \x_mult_f[13][12] , \x_mult_f[13][11] ,
         \x_mult_f[13][10] , \x_mult_f[13][9] , \x_mult_f[13][8] ,
         \x_mult_f[13][7] , \x_mult_f[13][6] , \x_mult_f[13][5] ,
         \x_mult_f[13][4] , \x_mult_f[13][3] , \x_mult_f[13][2] ,
         \x_mult_f[13][1] , \x_mult_f[13][0] , \x_mult_f[12][15] ,
         \x_mult_f[12][14] , \x_mult_f[12][13] , \x_mult_f[12][12] ,
         \x_mult_f[12][11] , \x_mult_f[12][10] , \x_mult_f[12][9] ,
         \x_mult_f[12][8] , \x_mult_f[12][7] , \x_mult_f[12][6] ,
         \x_mult_f[12][5] , \x_mult_f[12][4] , \x_mult_f[12][3] ,
         \x_mult_f[12][2] , \x_mult_f[12][1] , \x_mult_f[12][0] ,
         \x_mult_f[11][15] , \x_mult_f[11][14] , \x_mult_f[11][13] ,
         \x_mult_f[11][12] , \x_mult_f[11][11] , \x_mult_f[11][10] ,
         \x_mult_f[11][9] , \x_mult_f[11][8] , \x_mult_f[11][7] ,
         \x_mult_f[11][6] , \x_mult_f[11][5] , \x_mult_f[11][4] ,
         \x_mult_f[11][3] , \x_mult_f[11][2] , \x_mult_f[11][1] ,
         \x_mult_f[11][0] , \x_mult_f[10][15] , \x_mult_f[10][14] ,
         \x_mult_f[10][13] , \x_mult_f[10][12] , \x_mult_f[10][11] ,
         \x_mult_f[10][10] , \x_mult_f[10][9] , \x_mult_f[10][8] ,
         \x_mult_f[10][7] , \x_mult_f[10][6] , \x_mult_f[10][5] ,
         \x_mult_f[10][4] , \x_mult_f[10][3] , \x_mult_f[10][2] ,
         \x_mult_f[10][1] , \x_mult_f[10][0] , \x_mult_f[9][15] ,
         \x_mult_f[9][14] , \x_mult_f[9][13] , \x_mult_f[9][12] ,
         \x_mult_f[9][11] , \x_mult_f[9][10] , \x_mult_f[9][9] ,
         \x_mult_f[9][8] , \x_mult_f[9][7] , \x_mult_f[9][6] ,
         \x_mult_f[9][5] , \x_mult_f[9][4] , \x_mult_f[9][3] ,
         \x_mult_f[9][2] , \x_mult_f[9][1] , \x_mult_f[9][0] ,
         \x_mult_f[8][15] , \x_mult_f[8][14] , \x_mult_f[8][13] ,
         \x_mult_f[8][12] , \x_mult_f[8][11] , \x_mult_f[8][10] ,
         \x_mult_f[8][9] , \x_mult_f[8][8] , \x_mult_f[8][7] ,
         \x_mult_f[8][6] , \x_mult_f[8][5] , \x_mult_f[8][4] ,
         \x_mult_f[8][3] , \x_mult_f[8][2] , \x_mult_f[8][1] ,
         \x_mult_f[8][0] , \x_mult_f[7][15] , \x_mult_f[7][14] ,
         \x_mult_f[7][13] , \x_mult_f[7][12] , \x_mult_f[7][11] ,
         \x_mult_f[7][10] , \x_mult_f[7][9] , \x_mult_f[7][8] ,
         \x_mult_f[7][7] , \x_mult_f[7][6] , \x_mult_f[7][5] ,
         \x_mult_f[7][4] , \x_mult_f[7][3] , \x_mult_f[7][2] ,
         \x_mult_f[7][1] , \x_mult_f[7][0] , \x_mult_f[6][15] ,
         \x_mult_f[6][14] , \x_mult_f[6][13] , \x_mult_f[6][12] ,
         \x_mult_f[6][11] , \x_mult_f[6][10] , \x_mult_f[6][9] ,
         \x_mult_f[6][8] , \x_mult_f[6][7] , \x_mult_f[6][6] ,
         \x_mult_f[6][5] , \x_mult_f[6][4] , \x_mult_f[6][3] ,
         \x_mult_f[6][2] , \x_mult_f[6][1] , \x_mult_f[6][0] ,
         \x_mult_f[5][15] , \x_mult_f[5][14] , \x_mult_f[5][13] ,
         \x_mult_f[5][12] , \x_mult_f[5][11] , \x_mult_f[5][10] ,
         \x_mult_f[5][9] , \x_mult_f[5][8] , \x_mult_f[5][7] ,
         \x_mult_f[5][6] , \x_mult_f[5][5] , \x_mult_f[5][4] ,
         \x_mult_f[5][3] , \x_mult_f[5][2] , \x_mult_f[5][1] ,
         \x_mult_f[5][0] , \x_mult_f[4][15] , \x_mult_f[4][14] ,
         \x_mult_f[4][13] , \x_mult_f[4][12] , \x_mult_f[4][11] ,
         \x_mult_f[4][10] , \x_mult_f[4][9] , \x_mult_f[4][8] ,
         \x_mult_f[4][7] , \x_mult_f[4][6] , \x_mult_f[4][5] ,
         \x_mult_f[4][4] , \x_mult_f[4][3] , \x_mult_f[4][2] ,
         \x_mult_f[4][1] , \x_mult_f[4][0] , \x_mult_f[3][15] ,
         \x_mult_f[3][14] , \x_mult_f[3][13] , \x_mult_f[3][12] ,
         \x_mult_f[3][11] , \x_mult_f[3][10] , \x_mult_f[3][9] ,
         \x_mult_f[3][8] , \x_mult_f[3][7] , \x_mult_f[3][6] ,
         \x_mult_f[3][5] , \x_mult_f[3][4] , \x_mult_f[3][3] ,
         \x_mult_f[3][2] , \x_mult_f[3][1] , \x_mult_f[3][0] ,
         \x_mult_f[2][15] , \x_mult_f[2][14] , \x_mult_f[2][13] ,
         \x_mult_f[2][12] , \x_mult_f[2][11] , \x_mult_f[2][10] ,
         \x_mult_f[2][9] , \x_mult_f[2][8] , \x_mult_f[2][7] ,
         \x_mult_f[2][6] , \x_mult_f[2][5] , \x_mult_f[2][4] ,
         \x_mult_f[2][3] , \x_mult_f[2][2] , \x_mult_f[2][1] ,
         \x_mult_f[2][0] , \x_mult_f[1][15] , \x_mult_f[1][14] ,
         \x_mult_f[1][13] , \x_mult_f[1][12] , \x_mult_f[1][11] ,
         \x_mult_f[1][10] , \x_mult_f[1][9] , \x_mult_f[1][8] ,
         \x_mult_f[1][7] , \x_mult_f[1][6] , \x_mult_f[1][5] ,
         \x_mult_f[1][4] , \x_mult_f[1][3] , \x_mult_f[1][2] ,
         \x_mult_f[1][1] , \x_mult_f[1][0] , \x_mult_f[0][15] ,
         \x_mult_f[0][14] , \x_mult_f[0][13] , \x_mult_f[0][12] ,
         \x_mult_f[0][11] , \x_mult_f[0][10] , \x_mult_f[0][9] ,
         \x_mult_f[0][8] , \x_mult_f[0][7] , \x_mult_f[0][6] ,
         \x_mult_f[0][5] , \x_mult_f[0][4] , \x_mult_f[0][3] ,
         \x_mult_f[0][2] , \x_mult_f[0][1] , \x_mult_f[0][0] ,
         \adder_stage1[15][20] , \adder_stage1[15][15] ,
         \adder_stage1[15][14] , \adder_stage1[15][13] ,
         \adder_stage1[15][12] , \adder_stage1[15][11] ,
         \adder_stage1[15][10] , \adder_stage1[15][9] , \adder_stage1[15][8] ,
         \adder_stage1[15][7] , \adder_stage1[15][6] , \adder_stage1[15][5] ,
         \adder_stage1[15][4] , \adder_stage1[15][3] , \adder_stage1[15][2] ,
         \adder_stage1[15][1] , \adder_stage1[15][0] , \adder_stage1[14][20] ,
         \adder_stage1[14][15] , \adder_stage1[14][14] ,
         \adder_stage1[14][13] , \adder_stage1[14][12] ,
         \adder_stage1[14][11] , \adder_stage1[14][10] , \adder_stage1[14][9] ,
         \adder_stage1[14][8] , \adder_stage1[14][7] , \adder_stage1[14][6] ,
         \adder_stage1[14][5] , \adder_stage1[14][4] , \adder_stage1[14][3] ,
         \adder_stage1[14][2] , \adder_stage1[14][1] , \adder_stage1[14][0] ,
         \adder_stage1[13][20] , \adder_stage1[13][15] ,
         \adder_stage1[13][14] , \adder_stage1[13][13] ,
         \adder_stage1[13][12] , \adder_stage1[13][11] ,
         \adder_stage1[13][10] , \adder_stage1[13][9] , \adder_stage1[13][8] ,
         \adder_stage1[13][7] , \adder_stage1[13][6] , \adder_stage1[13][5] ,
         \adder_stage1[13][4] , \adder_stage1[13][3] , \adder_stage1[13][2] ,
         \adder_stage1[13][1] , \adder_stage1[13][0] , \adder_stage1[12][20] ,
         \adder_stage1[12][15] , \adder_stage1[12][14] ,
         \adder_stage1[12][13] , \adder_stage1[12][12] ,
         \adder_stage1[12][11] , \adder_stage1[12][10] , \adder_stage1[12][9] ,
         \adder_stage1[12][8] , \adder_stage1[12][7] , \adder_stage1[12][6] ,
         \adder_stage1[12][5] , \adder_stage1[12][4] , \adder_stage1[12][3] ,
         \adder_stage1[12][2] , \adder_stage1[12][1] , \adder_stage1[12][0] ,
         \adder_stage1[11][20] , \adder_stage1[11][15] ,
         \adder_stage1[11][14] , \adder_stage1[11][13] ,
         \adder_stage1[11][12] , \adder_stage1[11][11] ,
         \adder_stage1[11][10] , \adder_stage1[11][9] , \adder_stage1[11][8] ,
         \adder_stage1[11][7] , \adder_stage1[11][6] , \adder_stage1[11][5] ,
         \adder_stage1[11][4] , \adder_stage1[11][3] , \adder_stage1[11][2] ,
         \adder_stage1[11][1] , \adder_stage1[11][0] , \adder_stage1[10][20] ,
         \adder_stage1[10][15] , \adder_stage1[10][14] ,
         \adder_stage1[10][13] , \adder_stage1[10][12] ,
         \adder_stage1[10][11] , \adder_stage1[10][10] , \adder_stage1[10][9] ,
         \adder_stage1[10][8] , \adder_stage1[10][7] , \adder_stage1[10][6] ,
         \adder_stage1[10][5] , \adder_stage1[10][4] , \adder_stage1[10][3] ,
         \adder_stage1[10][2] , \adder_stage1[10][1] , \adder_stage1[10][0] ,
         \adder_stage1[9][20] , \adder_stage1[9][15] , \adder_stage1[9][14] ,
         \adder_stage1[9][13] , \adder_stage1[9][12] , \adder_stage1[9][11] ,
         \adder_stage1[9][10] , \adder_stage1[9][9] , \adder_stage1[9][8] ,
         \adder_stage1[9][7] , \adder_stage1[9][6] , \adder_stage1[9][5] ,
         \adder_stage1[9][4] , \adder_stage1[9][3] , \adder_stage1[9][2] ,
         \adder_stage1[9][1] , \adder_stage1[9][0] , \adder_stage1[8][20] ,
         \adder_stage1[8][15] , \adder_stage1[8][14] , \adder_stage1[8][13] ,
         \adder_stage1[8][12] , \adder_stage1[8][11] , \adder_stage1[8][10] ,
         \adder_stage1[8][9] , \adder_stage1[8][8] , \adder_stage1[8][7] ,
         \adder_stage1[8][6] , \adder_stage1[8][5] , \adder_stage1[8][4] ,
         \adder_stage1[8][3] , \adder_stage1[8][2] , \adder_stage1[8][1] ,
         \adder_stage1[8][0] , \adder_stage1[7][20] , \adder_stage1[7][15] ,
         \adder_stage1[7][14] , \adder_stage1[7][13] , \adder_stage1[7][12] ,
         \adder_stage1[7][11] , \adder_stage1[7][10] , \adder_stage1[7][9] ,
         \adder_stage1[7][8] , \adder_stage1[7][7] , \adder_stage1[7][6] ,
         \adder_stage1[7][5] , \adder_stage1[7][4] , \adder_stage1[7][3] ,
         \adder_stage1[7][2] , \adder_stage1[7][1] , \adder_stage1[7][0] ,
         \adder_stage1[6][20] , \adder_stage1[6][15] , \adder_stage1[6][14] ,
         \adder_stage1[6][13] , \adder_stage1[6][12] , \adder_stage1[6][11] ,
         \adder_stage1[6][10] , \adder_stage1[6][9] , \adder_stage1[6][8] ,
         \adder_stage1[6][7] , \adder_stage1[6][6] , \adder_stage1[6][5] ,
         \adder_stage1[6][4] , \adder_stage1[6][3] , \adder_stage1[6][2] ,
         \adder_stage1[6][1] , \adder_stage1[6][0] , \adder_stage1[5][20] ,
         \adder_stage1[5][15] , \adder_stage1[5][14] , \adder_stage1[5][13] ,
         \adder_stage1[5][12] , \adder_stage1[5][11] , \adder_stage1[5][10] ,
         \adder_stage1[5][9] , \adder_stage1[5][8] , \adder_stage1[5][7] ,
         \adder_stage1[5][6] , \adder_stage1[5][5] , \adder_stage1[5][4] ,
         \adder_stage1[5][3] , \adder_stage1[5][2] , \adder_stage1[5][1] ,
         \adder_stage1[5][0] , \adder_stage1[4][20] , \adder_stage1[4][15] ,
         \adder_stage1[4][14] , \adder_stage1[4][13] , \adder_stage1[4][12] ,
         \adder_stage1[4][11] , \adder_stage1[4][10] , \adder_stage1[4][9] ,
         \adder_stage1[4][8] , \adder_stage1[4][7] , \adder_stage1[4][6] ,
         \adder_stage1[4][5] , \adder_stage1[4][4] , \adder_stage1[4][3] ,
         \adder_stage1[4][2] , \adder_stage1[4][1] , \adder_stage1[4][0] ,
         \adder_stage1[3][20] , \adder_stage1[3][15] , \adder_stage1[3][14] ,
         \adder_stage1[3][13] , \adder_stage1[3][12] , \adder_stage1[3][11] ,
         \adder_stage1[3][10] , \adder_stage1[3][9] , \adder_stage1[3][8] ,
         \adder_stage1[3][7] , \adder_stage1[3][6] , \adder_stage1[3][5] ,
         \adder_stage1[3][4] , \adder_stage1[3][3] , \adder_stage1[3][2] ,
         \adder_stage1[3][1] , \adder_stage1[3][0] , \adder_stage1[2][20] ,
         \adder_stage1[2][15] , \adder_stage1[2][14] , \adder_stage1[2][13] ,
         \adder_stage1[2][12] , \adder_stage1[2][11] , \adder_stage1[2][10] ,
         \adder_stage1[2][9] , \adder_stage1[2][8] , \adder_stage1[2][7] ,
         \adder_stage1[2][6] , \adder_stage1[2][5] , \adder_stage1[2][4] ,
         \adder_stage1[2][3] , \adder_stage1[2][2] , \adder_stage1[2][1] ,
         \adder_stage1[2][0] , \adder_stage1[1][20] , \adder_stage1[1][15] ,
         \adder_stage1[1][14] , \adder_stage1[1][13] , \adder_stage1[1][12] ,
         \adder_stage1[1][11] , \adder_stage1[1][10] , \adder_stage1[1][9] ,
         \adder_stage1[1][8] , \adder_stage1[1][7] , \adder_stage1[1][6] ,
         \adder_stage1[1][5] , \adder_stage1[1][4] , \adder_stage1[1][3] ,
         \adder_stage1[1][2] , \adder_stage1[1][1] , \adder_stage1[1][0] ,
         \adder_stage1[0][20] , \adder_stage1[0][15] , \adder_stage1[0][14] ,
         \adder_stage1[0][13] , \adder_stage1[0][12] , \adder_stage1[0][11] ,
         \adder_stage1[0][10] , \adder_stage1[0][9] , \adder_stage1[0][8] ,
         \adder_stage1[0][7] , \adder_stage1[0][6] , \adder_stage1[0][5] ,
         \adder_stage1[0][4] , \adder_stage1[0][3] , \adder_stage1[0][2] ,
         \adder_stage1[0][1] , \adder_stage1[0][0] , \adder_stage2[7][20] ,
         \adder_stage2[7][19] , \adder_stage2[7][18] , \adder_stage2[7][17] ,
         \adder_stage2[7][16] , \adder_stage2[7][15] , \adder_stage2[7][14] ,
         \adder_stage2[7][13] , \adder_stage2[7][12] , \adder_stage2[7][11] ,
         \adder_stage2[7][10] , \adder_stage2[7][9] , \adder_stage2[7][8] ,
         \adder_stage2[7][7] , \adder_stage2[7][6] , \adder_stage2[7][5] ,
         \adder_stage2[7][4] , \adder_stage2[7][3] , \adder_stage2[7][2] ,
         \adder_stage2[7][1] , \adder_stage2[7][0] , \adder_stage2[6][20] ,
         \adder_stage2[6][19] , \adder_stage2[6][18] , \adder_stage2[6][17] ,
         \adder_stage2[6][16] , \adder_stage2[6][15] , \adder_stage2[6][14] ,
         \adder_stage2[6][13] , \adder_stage2[6][12] , \adder_stage2[6][11] ,
         \adder_stage2[6][10] , \adder_stage2[6][9] , \adder_stage2[6][8] ,
         \adder_stage2[6][7] , \adder_stage2[6][6] , \adder_stage2[6][5] ,
         \adder_stage2[6][4] , \adder_stage2[6][3] , \adder_stage2[6][2] ,
         \adder_stage2[6][1] , \adder_stage2[6][0] , \adder_stage2[5][20] ,
         \adder_stage2[5][19] , \adder_stage2[5][18] , \adder_stage2[5][17] ,
         \adder_stage2[5][16] , \adder_stage2[5][15] , \adder_stage2[5][14] ,
         \adder_stage2[5][13] , \adder_stage2[5][12] , \adder_stage2[5][11] ,
         \adder_stage2[5][10] , \adder_stage2[5][9] , \adder_stage2[5][8] ,
         \adder_stage2[5][7] , \adder_stage2[5][6] , \adder_stage2[5][5] ,
         \adder_stage2[5][4] , \adder_stage2[5][3] , \adder_stage2[5][2] ,
         \adder_stage2[5][1] , \adder_stage2[5][0] , \adder_stage2[4][20] ,
         \adder_stage2[4][19] , \adder_stage2[4][18] , \adder_stage2[4][17] ,
         \adder_stage2[4][16] , \adder_stage2[4][15] , \adder_stage2[4][14] ,
         \adder_stage2[4][13] , \adder_stage2[4][12] , \adder_stage2[4][11] ,
         \adder_stage2[4][10] , \adder_stage2[4][9] , \adder_stage2[4][8] ,
         \adder_stage2[4][7] , \adder_stage2[4][6] , \adder_stage2[4][5] ,
         \adder_stage2[4][4] , \adder_stage2[4][3] , \adder_stage2[4][2] ,
         \adder_stage2[4][1] , \adder_stage2[4][0] , \adder_stage2[3][20] ,
         \adder_stage2[3][19] , \adder_stage2[3][18] , \adder_stage2[3][17] ,
         \adder_stage2[3][16] , \adder_stage2[3][15] , \adder_stage2[3][14] ,
         \adder_stage2[3][13] , \adder_stage2[3][12] , \adder_stage2[3][11] ,
         \adder_stage2[3][10] , \adder_stage2[3][9] , \adder_stage2[3][8] ,
         \adder_stage2[3][7] , \adder_stage2[3][6] , \adder_stage2[3][5] ,
         \adder_stage2[3][4] , \adder_stage2[3][3] , \adder_stage2[3][2] ,
         \adder_stage2[3][1] , \adder_stage2[3][0] , \adder_stage2[2][20] ,
         \adder_stage2[2][19] , \adder_stage2[2][18] , \adder_stage2[2][17] ,
         \adder_stage2[2][16] , \adder_stage2[2][15] , \adder_stage2[2][14] ,
         \adder_stage2[2][13] , \adder_stage2[2][12] , \adder_stage2[2][11] ,
         \adder_stage2[2][10] , \adder_stage2[2][9] , \adder_stage2[2][8] ,
         \adder_stage2[2][7] , \adder_stage2[2][6] , \adder_stage2[2][5] ,
         \adder_stage2[2][4] , \adder_stage2[2][3] , \adder_stage2[2][2] ,
         \adder_stage2[2][1] , \adder_stage2[2][0] , \adder_stage2[1][20] ,
         \adder_stage2[1][19] , \adder_stage2[1][18] , \adder_stage2[1][17] ,
         \adder_stage2[1][16] , \adder_stage2[1][15] , \adder_stage2[1][14] ,
         \adder_stage2[1][13] , \adder_stage2[1][12] , \adder_stage2[1][11] ,
         \adder_stage2[1][10] , \adder_stage2[1][9] , \adder_stage2[1][8] ,
         \adder_stage2[1][7] , \adder_stage2[1][6] , \adder_stage2[1][5] ,
         \adder_stage2[1][4] , \adder_stage2[1][3] , \adder_stage2[1][2] ,
         \adder_stage2[1][1] , \adder_stage2[1][0] , \adder_stage2[0][20] ,
         \adder_stage2[0][19] , \adder_stage2[0][18] , \adder_stage2[0][17] ,
         \adder_stage2[0][16] , \adder_stage2[0][15] , \adder_stage2[0][14] ,
         \adder_stage2[0][13] , \adder_stage2[0][12] , \adder_stage2[0][11] ,
         \adder_stage2[0][10] , \adder_stage2[0][9] , \adder_stage2[0][8] ,
         \adder_stage2[0][7] , \adder_stage2[0][6] , \adder_stage2[0][5] ,
         \adder_stage2[0][4] , \adder_stage2[0][3] , \adder_stage2[0][2] ,
         \adder_stage2[0][1] , \adder_stage2[0][0] , \adder_stage3[3][20] ,
         \adder_stage3[3][19] , \adder_stage3[3][18] , \adder_stage3[3][17] ,
         \adder_stage3[3][16] , \adder_stage3[3][15] , \adder_stage3[3][14] ,
         \adder_stage3[3][13] , \adder_stage3[3][12] , \adder_stage3[3][11] ,
         \adder_stage3[3][10] , \adder_stage3[3][9] , \adder_stage3[3][8] ,
         \adder_stage3[3][7] , \adder_stage3[3][6] , \adder_stage3[3][5] ,
         \adder_stage3[3][4] , \adder_stage3[3][3] , \adder_stage3[3][2] ,
         \adder_stage3[3][1] , \adder_stage3[3][0] , \adder_stage3[2][20] ,
         \adder_stage3[2][19] , \adder_stage3[2][18] , \adder_stage3[2][17] ,
         \adder_stage3[2][16] , \adder_stage3[2][15] , \adder_stage3[2][14] ,
         \adder_stage3[2][13] , \adder_stage3[2][12] , \adder_stage3[2][11] ,
         \adder_stage3[2][10] , \adder_stage3[2][9] , \adder_stage3[2][8] ,
         \adder_stage3[2][7] , \adder_stage3[2][6] , \adder_stage3[2][5] ,
         \adder_stage3[2][4] , \adder_stage3[2][3] , \adder_stage3[2][2] ,
         \adder_stage3[2][1] , \adder_stage3[2][0] , \adder_stage3[1][20] ,
         \adder_stage3[1][19] , \adder_stage3[1][18] , \adder_stage3[1][17] ,
         \adder_stage3[1][16] , \adder_stage3[1][15] , \adder_stage3[1][14] ,
         \adder_stage3[1][13] , \adder_stage3[1][12] , \adder_stage3[1][11] ,
         \adder_stage3[1][10] , \adder_stage3[1][9] , \adder_stage3[1][8] ,
         \adder_stage3[1][7] , \adder_stage3[1][6] , \adder_stage3[1][5] ,
         \adder_stage3[1][4] , \adder_stage3[1][3] , \adder_stage3[1][2] ,
         \adder_stage3[1][1] , \adder_stage3[1][0] , \adder_stage3[0][20] ,
         \adder_stage3[0][19] , \adder_stage3[0][18] , \adder_stage3[0][17] ,
         \adder_stage3[0][16] , \adder_stage3[0][15] , \adder_stage3[0][14] ,
         \adder_stage3[0][13] , \adder_stage3[0][12] , \adder_stage3[0][11] ,
         \adder_stage3[0][10] , \adder_stage3[0][9] , \adder_stage3[0][8] ,
         \adder_stage3[0][7] , \adder_stage3[0][6] , \adder_stage3[0][5] ,
         \adder_stage3[0][4] , \adder_stage3[0][3] , \adder_stage3[0][2] ,
         \adder_stage3[0][1] , \adder_stage3[0][0] , \adder_stage4[1][20] ,
         \adder_stage4[1][19] , \adder_stage4[1][18] , \adder_stage4[1][17] ,
         \adder_stage4[1][16] , \adder_stage4[1][15] , \adder_stage4[1][14] ,
         \adder_stage4[1][13] , \adder_stage4[1][12] , \adder_stage4[1][11] ,
         \adder_stage4[1][10] , \adder_stage4[1][9] , \adder_stage4[1][8] ,
         \adder_stage4[1][7] , \adder_stage4[1][6] , \adder_stage4[1][5] ,
         \adder_stage4[1][4] , \adder_stage4[1][3] , \adder_stage4[1][2] ,
         \adder_stage4[1][1] , \adder_stage4[1][0] , \adder_stage4[0][20] ,
         \adder_stage4[0][19] , \adder_stage4[0][18] , \adder_stage4[0][17] ,
         \adder_stage4[0][16] , \adder_stage4[0][15] , \adder_stage4[0][14] ,
         \adder_stage4[0][13] , \adder_stage4[0][12] , \adder_stage4[0][11] ,
         \adder_stage4[0][10] , \adder_stage4[0][9] , \adder_stage4[0][8] ,
         \adder_stage4[0][7] , \adder_stage4[0][6] , \adder_stage4[0][5] ,
         \adder_stage4[0][4] , \adder_stage4[0][3] , \adder_stage4[0][2] ,
         \adder_stage4[0][1] , \adder_stage4[0][0] , n1909, n1910, n1911,
         n1912, n1930, n1931, n1932, n1933, n1951, n1952, n1953, n1954, n1972,
         n1973, n1974, n1975, n1993, n1994, n1995, n1996, n2014, n2015, n2016,
         n2017, n2035, n2036, n2037, n2038, n2056, n2057, n2058, n2059, n3118,
         n3119, n3120, n3121, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321;
  wire   [4:0] fmem_addr;
  wire   [6:0] \ctrl_inst/xmem_tracker ;
  wire   [3:0] \ctrl_inst/pline_cntr ;
  wire   [2:0] \ctrl_inst/state ;

  DFF_X1 \xmem_inst/mem_reg[31][7]  ( .D(n3377), .CK(clk), .Q(
        \xmem_data[31][7] ) );
  DFF_X1 \xmem_inst/mem_reg[31][6]  ( .D(n3376), .CK(clk), .Q(
        \xmem_data[31][6] ) );
  DFF_X1 \xmem_inst/mem_reg[31][5]  ( .D(n3375), .CK(clk), .Q(
        \xmem_data[31][5] ) );
  DFF_X1 \xmem_inst/mem_reg[31][4]  ( .D(n3374), .CK(clk), .Q(
        \xmem_data[31][4] ) );
  DFF_X1 \xmem_inst/mem_reg[31][3]  ( .D(n3373), .CK(clk), .Q(
        \xmem_data[31][3] ) );
  DFF_X1 \xmem_inst/mem_reg[31][2]  ( .D(n3372), .CK(clk), .Q(
        \xmem_data[31][2] ) );
  DFF_X1 \xmem_inst/mem_reg[31][1]  ( .D(n3371), .CK(clk), .Q(
        \xmem_data[31][1] ) );
  DFF_X1 \xmem_inst/mem_reg[31][0]  ( .D(n3370), .CK(clk), .Q(
        \xmem_data[31][0] ) );
  DFF_X1 \xmem_inst/mem_reg[30][7]  ( .D(n10317), .CK(clk), .Q(
        \xmem_data[30][7] ) );
  DFF_X1 \xmem_inst/mem_reg[30][6]  ( .D(n10316), .CK(clk), .Q(
        \xmem_data[30][6] ) );
  DFF_X1 \xmem_inst/mem_reg[30][5]  ( .D(n10315), .CK(clk), .Q(
        \xmem_data[30][5] ) );
  DFF_X1 \xmem_inst/mem_reg[30][4]  ( .D(n10314), .CK(clk), .Q(
        \xmem_data[30][4] ) );
  DFF_X1 \xmem_inst/mem_reg[30][3]  ( .D(n10313), .CK(clk), .Q(
        \xmem_data[30][3] ) );
  DFF_X1 \xmem_inst/mem_reg[30][2]  ( .D(n10312), .CK(clk), .Q(
        \xmem_data[30][2] ) );
  DFF_X1 \xmem_inst/mem_reg[30][1]  ( .D(n10311), .CK(clk), .Q(
        \xmem_data[30][1] ) );
  DFF_X1 \xmem_inst/mem_reg[30][0]  ( .D(n10310), .CK(clk), .Q(
        \xmem_data[30][0] ) );
  DFF_X1 \xmem_inst/mem_reg[29][7]  ( .D(n10309), .CK(clk), .Q(
        \xmem_data[29][7] ) );
  DFF_X1 \xmem_inst/mem_reg[29][6]  ( .D(n10308), .CK(clk), .Q(
        \xmem_data[29][6] ) );
  DFF_X1 \xmem_inst/mem_reg[29][5]  ( .D(n10307), .CK(clk), .Q(
        \xmem_data[29][5] ) );
  DFF_X1 \xmem_inst/mem_reg[29][4]  ( .D(n10306), .CK(clk), .Q(
        \xmem_data[29][4] ) );
  DFF_X1 \xmem_inst/mem_reg[29][3]  ( .D(n10305), .CK(clk), .Q(
        \xmem_data[29][3] ) );
  DFF_X1 \xmem_inst/mem_reg[29][2]  ( .D(n10304), .CK(clk), .Q(
        \xmem_data[29][2] ) );
  DFF_X1 \xmem_inst/mem_reg[29][1]  ( .D(n10303), .CK(clk), .Q(
        \xmem_data[29][1] ) );
  DFF_X1 \xmem_inst/mem_reg[29][0]  ( .D(n10302), .CK(clk), .Q(
        \xmem_data[29][0] ) );
  DFF_X1 \xmem_inst/mem_reg[28][7]  ( .D(n10301), .CK(clk), .Q(
        \xmem_data[28][7] ) );
  DFF_X1 \xmem_inst/mem_reg[28][6]  ( .D(n10300), .CK(clk), .Q(
        \xmem_data[28][6] ) );
  DFF_X1 \xmem_inst/mem_reg[28][5]  ( .D(n10299), .CK(clk), .Q(
        \xmem_data[28][5] ) );
  DFF_X1 \xmem_inst/mem_reg[28][4]  ( .D(n10298), .CK(clk), .Q(
        \xmem_data[28][4] ) );
  DFF_X1 \xmem_inst/mem_reg[28][3]  ( .D(n10297), .CK(clk), .Q(
        \xmem_data[28][3] ) );
  DFF_X1 \xmem_inst/mem_reg[28][2]  ( .D(n10296), .CK(clk), .Q(
        \xmem_data[28][2] ) );
  DFF_X1 \xmem_inst/mem_reg[28][1]  ( .D(n10295), .CK(clk), .Q(
        \xmem_data[28][1] ) );
  DFF_X1 \xmem_inst/mem_reg[28][0]  ( .D(n10294), .CK(clk), .Q(
        \xmem_data[28][0] ) );
  DFF_X1 \xmem_inst/mem_reg[27][7]  ( .D(n10293), .CK(clk), .Q(
        \xmem_data[27][7] ) );
  DFF_X1 \xmem_inst/mem_reg[27][6]  ( .D(n10292), .CK(clk), .Q(
        \xmem_data[27][6] ) );
  DFF_X1 \xmem_inst/mem_reg[27][5]  ( .D(n10291), .CK(clk), .Q(
        \xmem_data[27][5] ) );
  DFF_X1 \xmem_inst/mem_reg[27][4]  ( .D(n10290), .CK(clk), .Q(
        \xmem_data[27][4] ) );
  DFF_X1 \xmem_inst/mem_reg[27][3]  ( .D(n10289), .CK(clk), .Q(
        \xmem_data[27][3] ) );
  DFF_X1 \xmem_inst/mem_reg[27][2]  ( .D(n10288), .CK(clk), .Q(
        \xmem_data[27][2] ) );
  DFF_X1 \xmem_inst/mem_reg[27][1]  ( .D(n10287), .CK(clk), .Q(
        \xmem_data[27][1] ) );
  DFF_X1 \xmem_inst/mem_reg[27][0]  ( .D(n10286), .CK(clk), .Q(
        \xmem_data[27][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][7]  ( .D(n10285), .CK(clk), .Q(
        \xmem_data[26][7] ) );
  DFF_X1 \xmem_inst/mem_reg[26][6]  ( .D(n10284), .CK(clk), .Q(
        \xmem_data[26][6] ) );
  DFF_X1 \xmem_inst/mem_reg[26][5]  ( .D(n10283), .CK(clk), .Q(
        \xmem_data[26][5] ) );
  DFF_X1 \xmem_inst/mem_reg[26][4]  ( .D(n10282), .CK(clk), .Q(
        \xmem_data[26][4] ) );
  DFF_X1 \xmem_inst/mem_reg[26][3]  ( .D(n10281), .CK(clk), .Q(
        \xmem_data[26][3] ) );
  DFF_X1 \xmem_inst/mem_reg[26][2]  ( .D(n10280), .CK(clk), .Q(
        \xmem_data[26][2] ) );
  DFF_X1 \xmem_inst/mem_reg[26][1]  ( .D(n10279), .CK(clk), .Q(
        \xmem_data[26][1] ) );
  DFF_X1 \xmem_inst/mem_reg[26][0]  ( .D(n10278), .CK(clk), .Q(
        \xmem_data[26][0] ) );
  DFF_X1 \xmem_inst/mem_reg[25][7]  ( .D(n10277), .CK(clk), .Q(
        \xmem_data[25][7] ) );
  DFF_X1 \xmem_inst/mem_reg[25][6]  ( .D(n10276), .CK(clk), .Q(
        \xmem_data[25][6] ) );
  DFF_X1 \xmem_inst/mem_reg[25][5]  ( .D(n10275), .CK(clk), .Q(
        \xmem_data[25][5] ) );
  DFF_X1 \xmem_inst/mem_reg[24][5]  ( .D(n10274), .CK(clk), .Q(
        \xmem_data[24][5] ) );
  DFF_X1 \xmem_inst/mem_reg[23][5]  ( .D(n10273), .CK(clk), .Q(
        \xmem_data[23][5] ) );
  DFF_X1 \xmem_inst/mem_reg[22][5]  ( .D(n10272), .CK(clk), .Q(
        \xmem_data[22][5] ) );
  DFF_X1 \xmem_inst/mem_reg[21][5]  ( .D(n10271), .CK(clk), .Q(
        \xmem_data[21][5] ) );
  DFF_X1 \xmem_inst/mem_reg[20][5]  ( .D(n10270), .CK(clk), .Q(
        \xmem_data[20][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n10269), .CK(clk), .Q(
        \xmem_data[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n10268), .CK(clk), .Q(
        \xmem_data[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n10267), .CK(clk), .Q(
        \xmem_data[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n10266), .CK(clk), .Q(
        \xmem_data[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n10265), .CK(clk), .Q(
        \xmem_data[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n10264), .CK(clk), .Q(
        \xmem_data[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n10263), .CK(clk), .Q(
        \xmem_data[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n10262), .CK(clk), .Q(
        \xmem_data[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n10261), .CK(clk), .Q(
        \xmem_data[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n10260), .CK(clk), .Q(
        \xmem_data[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n10259), .CK(clk), .Q(
        \xmem_data[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n10258), .CK(clk), .Q(
        \xmem_data[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n10257), .CK(clk), .Q(
        \xmem_data[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n10256), .CK(clk), .Q(
        \xmem_data[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n10255), .CK(clk), .Q(
        \xmem_data[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n10254), .CK(clk), .Q(
        \xmem_data[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n10253), .CK(clk), .Q(
        \xmem_data[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n10252), .CK(clk), .Q(
        \xmem_data[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n10251), .CK(clk), .Q(
        \xmem_data[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n10250), .CK(clk), .Q(
        \xmem_data[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[25][4]  ( .D(n10249), .CK(clk), .Q(
        \xmem_data[25][4] ) );
  DFF_X1 \xmem_inst/mem_reg[24][4]  ( .D(n10248), .CK(clk), .Q(
        \xmem_data[24][4] ) );
  DFF_X1 \xmem_inst/mem_reg[23][4]  ( .D(n10247), .CK(clk), .Q(
        \xmem_data[23][4] ) );
  DFF_X1 \xmem_inst/mem_reg[22][4]  ( .D(n10246), .CK(clk), .Q(
        \xmem_data[22][4] ) );
  DFF_X1 \xmem_inst/mem_reg[21][4]  ( .D(n10245), .CK(clk), .Q(
        \xmem_data[21][4] ) );
  DFF_X1 \xmem_inst/mem_reg[20][4]  ( .D(n10244), .CK(clk), .Q(
        \xmem_data[20][4] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n10243), .CK(clk), .Q(
        \xmem_data[19][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n10242), .CK(clk), .Q(
        \xmem_data[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n10241), .CK(clk), .Q(
        \xmem_data[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n10240), .CK(clk), .Q(
        \xmem_data[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n10239), .CK(clk), .Q(
        \xmem_data[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n10238), .CK(clk), .Q(
        \xmem_data[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n10237), .CK(clk), .Q(
        \xmem_data[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n10236), .CK(clk), .Q(
        \xmem_data[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n10235), .CK(clk), .Q(
        \xmem_data[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n10234), .CK(clk), .Q(
        \xmem_data[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n10233), .CK(clk), .Q(
        \xmem_data[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n10232), .CK(clk), .Q(
        \xmem_data[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n10231), .CK(clk), .Q(
        \xmem_data[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n10230), .CK(clk), .Q(
        \xmem_data[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n10229), .CK(clk), .Q(
        \xmem_data[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n10228), .CK(clk), .Q(
        \xmem_data[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n10227), .CK(clk), .Q(
        \xmem_data[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n10226), .CK(clk), .Q(
        \xmem_data[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n10225), .CK(clk), .Q(
        \xmem_data[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n10224), .CK(clk), .Q(
        \xmem_data[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[25][3]  ( .D(n10223), .CK(clk), .Q(
        \xmem_data[25][3] ) );
  DFF_X1 \xmem_inst/mem_reg[24][3]  ( .D(n10222), .CK(clk), .Q(
        \xmem_data[24][3] ) );
  DFF_X1 \xmem_inst/mem_reg[23][3]  ( .D(n10221), .CK(clk), .Q(
        \xmem_data[23][3] ) );
  DFF_X1 \xmem_inst/mem_reg[22][3]  ( .D(n10220), .CK(clk), .Q(
        \xmem_data[22][3] ) );
  DFF_X1 \xmem_inst/mem_reg[21][3]  ( .D(n10219), .CK(clk), .Q(
        \xmem_data[21][3] ) );
  DFF_X1 \xmem_inst/mem_reg[20][3]  ( .D(n10218), .CK(clk), .Q(
        \xmem_data[20][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n10217), .CK(clk), .Q(
        \xmem_data[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n10216), .CK(clk), .Q(
        \xmem_data[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n10215), .CK(clk), .Q(
        \xmem_data[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n10214), .CK(clk), .Q(
        \xmem_data[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n10213), .CK(clk), .Q(
        \xmem_data[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n10212), .CK(clk), .Q(
        \xmem_data[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n10211), .CK(clk), .Q(
        \xmem_data[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n10210), .CK(clk), .Q(
        \xmem_data[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n10209), .CK(clk), .Q(
        \xmem_data[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n10208), .CK(clk), .Q(
        \xmem_data[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n10207), .CK(clk), .Q(
        \xmem_data[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n10206), .CK(clk), .Q(
        \xmem_data[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n10205), .CK(clk), .Q(
        \xmem_data[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n10204), .CK(clk), .Q(
        \xmem_data[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n10203), .CK(clk), .Q(
        \xmem_data[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n10202), .CK(clk), .Q(
        \xmem_data[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n10201), .CK(clk), .Q(
        \xmem_data[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n10200), .CK(clk), .Q(
        \xmem_data[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n10199), .CK(clk), .Q(
        \xmem_data[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n10198), .CK(clk), .Q(
        \xmem_data[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[25][2]  ( .D(n10197), .CK(clk), .Q(
        \xmem_data[25][2] ) );
  DFF_X1 \xmem_inst/mem_reg[24][2]  ( .D(n10196), .CK(clk), .Q(
        \xmem_data[24][2] ) );
  DFF_X1 \xmem_inst/mem_reg[23][2]  ( .D(n10195), .CK(clk), .Q(
        \xmem_data[23][2] ) );
  DFF_X1 \xmem_inst/mem_reg[22][2]  ( .D(n10194), .CK(clk), .Q(
        \xmem_data[22][2] ) );
  DFF_X1 \xmem_inst/mem_reg[21][2]  ( .D(n10193), .CK(clk), .Q(
        \xmem_data[21][2] ) );
  DFF_X1 \xmem_inst/mem_reg[20][2]  ( .D(n10192), .CK(clk), .Q(
        \xmem_data[20][2] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n10191), .CK(clk), .Q(
        \xmem_data[19][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n10190), .CK(clk), .Q(
        \xmem_data[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n10189), .CK(clk), .Q(
        \xmem_data[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n10188), .CK(clk), .Q(
        \xmem_data[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n10187), .CK(clk), .Q(
        \xmem_data[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n10186), .CK(clk), .Q(
        \xmem_data[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n10185), .CK(clk), .Q(
        \xmem_data[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n10184), .CK(clk), .Q(
        \xmem_data[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n10183), .CK(clk), .Q(
        \xmem_data[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n10182), .CK(clk), .Q(
        \xmem_data[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n10181), .CK(clk), .Q(
        \xmem_data[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n10180), .CK(clk), .Q(
        \xmem_data[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n10179), .CK(clk), .Q(
        \xmem_data[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n10178), .CK(clk), .Q(
        \xmem_data[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n10177), .CK(clk), .Q(
        \xmem_data[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n10176), .CK(clk), .Q(
        \xmem_data[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n10175), .CK(clk), .Q(
        \xmem_data[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n10174), .CK(clk), .Q(
        \xmem_data[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n10173), .CK(clk), .Q(
        \xmem_data[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n10172), .CK(clk), .Q(
        \xmem_data[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[25][1]  ( .D(n10171), .CK(clk), .Q(
        \xmem_data[25][1] ) );
  DFF_X1 \xmem_inst/mem_reg[24][1]  ( .D(n10170), .CK(clk), .Q(
        \xmem_data[24][1] ) );
  DFF_X1 \xmem_inst/mem_reg[23][1]  ( .D(n10169), .CK(clk), .Q(
        \xmem_data[23][1] ) );
  DFF_X1 \xmem_inst/mem_reg[22][1]  ( .D(n10168), .CK(clk), .Q(
        \xmem_data[22][1] ) );
  DFF_X1 \xmem_inst/mem_reg[21][1]  ( .D(n10167), .CK(clk), .Q(
        \xmem_data[21][1] ) );
  DFF_X1 \xmem_inst/mem_reg[20][1]  ( .D(n10166), .CK(clk), .Q(
        \xmem_data[20][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n10165), .CK(clk), .Q(
        \xmem_data[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n10164), .CK(clk), .Q(
        \xmem_data[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n10163), .CK(clk), .Q(
        \xmem_data[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n10162), .CK(clk), .Q(
        \xmem_data[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n10161), .CK(clk), .Q(
        \xmem_data[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n10160), .CK(clk), .Q(
        \xmem_data[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n10159), .CK(clk), .Q(
        \xmem_data[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n10158), .CK(clk), .Q(
        \xmem_data[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n10157), .CK(clk), .Q(
        \xmem_data[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n10156), .CK(clk), .Q(
        \xmem_data[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n10155), .CK(clk), .Q(
        \xmem_data[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n10154), .CK(clk), .Q(
        \xmem_data[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n10153), .CK(clk), .Q(
        \xmem_data[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n10152), .CK(clk), .Q(
        \xmem_data[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n10151), .CK(clk), .Q(
        \xmem_data[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n10150), .CK(clk), .Q(
        \xmem_data[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n10149), .CK(clk), .Q(
        \xmem_data[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n10148), .CK(clk), .Q(
        \xmem_data[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n10147), .CK(clk), .Q(
        \xmem_data[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n10146), .CK(clk), .Q(
        \xmem_data[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[25][0]  ( .D(n10145), .CK(clk), .Q(
        \xmem_data[25][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][0]  ( .D(n10144), .CK(clk), .Q(
        \xmem_data[24][0] ) );
  DFF_X1 \xmem_inst/mem_reg[23][0]  ( .D(n10143), .CK(clk), .Q(
        \xmem_data[23][0] ) );
  DFF_X1 \xmem_inst/mem_reg[22][0]  ( .D(n10142), .CK(clk), .Q(
        \xmem_data[22][0] ) );
  DFF_X1 \xmem_inst/mem_reg[21][0]  ( .D(n10141), .CK(clk), .Q(
        \xmem_data[21][0] ) );
  DFF_X1 \xmem_inst/mem_reg[20][0]  ( .D(n10140), .CK(clk), .Q(
        \xmem_data[20][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n10139), .CK(clk), .Q(
        \xmem_data[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n10138), .CK(clk), .Q(
        \xmem_data[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n10137), .CK(clk), .Q(
        \xmem_data[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n10136), .CK(clk), .Q(
        \xmem_data[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n10135), .CK(clk), .Q(
        \xmem_data[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n10134), .CK(clk), .Q(
        \xmem_data[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n10133), .CK(clk), .Q(
        \xmem_data[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n10132), .CK(clk), .Q(
        \xmem_data[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n10131), .CK(clk), .Q(
        \xmem_data[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n10130), .CK(clk), .Q(
        \xmem_data[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n10129), .CK(clk), .Q(
        \xmem_data[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n10128), .CK(clk), .Q(
        \xmem_data[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n10127), .CK(clk), .Q(
        \xmem_data[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n10126), .CK(clk), .Q(
        \xmem_data[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n10125), .CK(clk), .Q(
        \xmem_data[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n10124), .CK(clk), .Q(
        \xmem_data[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n10123), .CK(clk), .Q(
        \xmem_data[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n10122), .CK(clk), .Q(
        \xmem_data[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n10121), .CK(clk), .Q(
        \xmem_data[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n10120), .CK(clk), .Q(
        \xmem_data[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][7]  ( .D(n10119), .CK(clk), .Q(
        \xmem_data[24][7] ) );
  DFF_X1 \xmem_inst/mem_reg[23][7]  ( .D(n10118), .CK(clk), .Q(
        \xmem_data[23][7] ) );
  DFF_X1 \xmem_inst/mem_reg[22][7]  ( .D(n10117), .CK(clk), .Q(
        \xmem_data[22][7] ) );
  DFF_X1 \xmem_inst/mem_reg[21][7]  ( .D(n10116), .CK(clk), .Q(
        \xmem_data[21][7] ) );
  DFF_X1 \xmem_inst/mem_reg[20][7]  ( .D(n10115), .CK(clk), .Q(
        \xmem_data[20][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n10114), .CK(clk), .Q(
        \xmem_data[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n10113), .CK(clk), .Q(
        \xmem_data[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n10112), .CK(clk), .Q(
        \xmem_data[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n10111), .CK(clk), .Q(
        \xmem_data[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n10110), .CK(clk), .Q(
        \xmem_data[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n10109), .CK(clk), .Q(
        \xmem_data[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n10108), .CK(clk), .Q(
        \xmem_data[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n10107), .CK(clk), .Q(
        \xmem_data[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n10106), .CK(clk), .Q(
        \xmem_data[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n10105), .CK(clk), .Q(
        \xmem_data[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n10104), .CK(clk), .Q(
        \xmem_data[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n10103), .CK(clk), .Q(
        \xmem_data[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n10102), .CK(clk), .Q(
        \xmem_data[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n10101), .CK(clk), .Q(
        \xmem_data[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n10100), .CK(clk), .Q(
        \xmem_data[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n10099), .CK(clk), .Q(
        \xmem_data[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n10098), .CK(clk), .Q(
        \xmem_data[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n10097), .CK(clk), .Q(
        \xmem_data[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n10096), .CK(clk), .Q(
        \xmem_data[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n10095), .CK(clk), .Q(
        \xmem_data[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[24][6]  ( .D(n10094), .CK(clk), .Q(
        \xmem_data[24][6] ) );
  DFF_X1 \xmem_inst/mem_reg[23][6]  ( .D(n10093), .CK(clk), .Q(
        \xmem_data[23][6] ) );
  DFF_X1 \xmem_inst/mem_reg[22][6]  ( .D(n10092), .CK(clk), .Q(
        \xmem_data[22][6] ) );
  DFF_X1 \xmem_inst/mem_reg[21][6]  ( .D(n10091), .CK(clk), .Q(
        \xmem_data[21][6] ) );
  DFF_X1 \xmem_inst/mem_reg[20][6]  ( .D(n10090), .CK(clk), .Q(
        \xmem_data[20][6] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n10089), .CK(clk), .Q(
        \xmem_data[19][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n10088), .CK(clk), .Q(
        \xmem_data[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n10087), .CK(clk), .Q(
        \xmem_data[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n10086), .CK(clk), .Q(
        \xmem_data[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n10085), .CK(clk), .Q(
        \xmem_data[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n10084), .CK(clk), .Q(
        \xmem_data[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n10083), .CK(clk), .Q(
        \xmem_data[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n10082), .CK(clk), .Q(
        \xmem_data[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n10081), .CK(clk), .Q(
        \xmem_data[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n10080), .CK(clk), .Q(
        \xmem_data[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n10079), .CK(clk), .Q(
        \xmem_data[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n10078), .CK(clk), .Q(
        \xmem_data[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n10077), .CK(clk), .Q(
        \xmem_data[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n10076), .CK(clk), .Q(
        \xmem_data[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n10075), .CK(clk), .Q(
        \xmem_data[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n10074), .CK(clk), .Q(
        \xmem_data[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n10073), .CK(clk), .Q(
        \xmem_data[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n10072), .CK(clk), .Q(
        \xmem_data[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n10071), .CK(clk), .Q(
        \xmem_data[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n10070), .CK(clk), .Q(
        \xmem_data[0][6] ) );
  DFF_X1 \ctrl_inst/conv_done_reg  ( .D(n3390), .CK(clk), .Q(conv_done), .QN(
        n8718) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[0]  ( .D(n3383), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [0]), .QN(n8911) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[1]  ( .D(n10321), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [1]), .QN(n8912) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[2]  ( .D(n10320), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [2]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[3]  ( .D(n10319), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [3]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[4]  ( .D(n10318), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [4]) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[5]  ( .D(n3378), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [5]) );
  DFF_X1 \ctrl_inst/m_valid_reg  ( .D(n3389), .CK(clk), .Q(m_valid_y), .QN(
        n3511) );
  DFF_X1 \ctrl_inst/state_reg[0]  ( .D(n3388), .CK(clk), .Q(
        \ctrl_inst/state [0]) );
  DFF_X1 \ctrl_inst/xmem_full_reg  ( .D(n3391), .CK(clk), .Q(xmem_full) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[3]  ( .D(n3396), .CK(clk), .Q(
        fmem_addr[3]), .QN(n8712) );
  DFF_X1 \fmem_inst/mem_reg[0][0]  ( .D(n9546), .CK(clk), .Q(\fmem_data[0][0] ) );
  DFF_X1 \fmem_inst/mem_reg[0][1]  ( .D(n9545), .CK(clk), .Q(\fmem_data[0][1] ) );
  DFF_X1 \fmem_inst/mem_reg[0][2]  ( .D(n9544), .CK(clk), .Q(\fmem_data[0][2] ) );
  DFF_X1 \fmem_inst/mem_reg[0][3]  ( .D(n9543), .CK(clk), .Q(\fmem_data[0][3] ) );
  DFF_X1 \fmem_inst/mem_reg[0][4]  ( .D(n9542), .CK(clk), .Q(\fmem_data[0][4] ) );
  DFF_X1 \fmem_inst/mem_reg[0][5]  ( .D(n9541), .CK(clk), .Q(\fmem_data[0][5] ) );
  DFF_X1 \fmem_inst/mem_reg[0][6]  ( .D(n9540), .CK(clk), .Q(\fmem_data[0][6] ) );
  DFF_X1 \fmem_inst/mem_reg[0][7]  ( .D(n9539), .CK(clk), .Q(\fmem_data[0][7] ) );
  DFF_X1 \fmem_inst/mem_reg[1][0]  ( .D(n9538), .CK(clk), .Q(\fmem_data[1][0] ) );
  DFF_X1 \fmem_inst/mem_reg[1][1]  ( .D(n9537), .CK(clk), .Q(\fmem_data[1][1] ) );
  DFF_X1 \fmem_inst/mem_reg[1][2]  ( .D(n9536), .CK(clk), .Q(\fmem_data[1][2] ) );
  DFF_X1 \fmem_inst/mem_reg[1][3]  ( .D(n9535), .CK(clk), .Q(\fmem_data[1][3] ) );
  DFF_X1 \fmem_inst/mem_reg[1][4]  ( .D(n9534), .CK(clk), .Q(\fmem_data[1][4] ) );
  DFF_X1 \fmem_inst/mem_reg[1][5]  ( .D(n9533), .CK(clk), .Q(\fmem_data[1][5] ) );
  DFF_X1 \fmem_inst/mem_reg[1][6]  ( .D(n9532), .CK(clk), .Q(\fmem_data[1][6] ) );
  DFF_X1 \fmem_inst/mem_reg[1][7]  ( .D(n9531), .CK(clk), .Q(\fmem_data[1][7] ) );
  DFF_X1 \fmem_inst/mem_reg[2][0]  ( .D(n9530), .CK(clk), .Q(\fmem_data[2][0] ) );
  DFF_X1 \fmem_inst/mem_reg[2][1]  ( .D(n9529), .CK(clk), .Q(\fmem_data[2][1] ) );
  DFF_X1 \fmem_inst/mem_reg[2][2]  ( .D(n9528), .CK(clk), .Q(\fmem_data[2][2] ) );
  DFF_X1 \fmem_inst/mem_reg[2][3]  ( .D(n9527), .CK(clk), .Q(\fmem_data[2][3] ) );
  DFF_X1 \fmem_inst/mem_reg[2][4]  ( .D(n9526), .CK(clk), .Q(\fmem_data[2][4] ) );
  DFF_X1 \fmem_inst/mem_reg[2][5]  ( .D(n9525), .CK(clk), .Q(\fmem_data[2][5] ) );
  DFF_X1 \fmem_inst/mem_reg[2][6]  ( .D(n9524), .CK(clk), .Q(\fmem_data[2][6] ) );
  DFF_X1 \fmem_inst/mem_reg[2][7]  ( .D(n9523), .CK(clk), .Q(\fmem_data[2][7] ) );
  DFF_X1 \fmem_inst/mem_reg[3][0]  ( .D(n9522), .CK(clk), .Q(\fmem_data[3][0] ) );
  DFF_X1 \fmem_inst/mem_reg[3][1]  ( .D(n9521), .CK(clk), .Q(\fmem_data[3][1] ) );
  DFF_X1 \fmem_inst/mem_reg[3][2]  ( .D(n9520), .CK(clk), .Q(\fmem_data[3][2] ) );
  DFF_X1 \fmem_inst/mem_reg[3][3]  ( .D(n9519), .CK(clk), .Q(\fmem_data[3][3] ) );
  DFF_X1 \fmem_inst/mem_reg[3][4]  ( .D(n9518), .CK(clk), .Q(\fmem_data[3][4] ) );
  DFF_X1 \fmem_inst/mem_reg[3][5]  ( .D(n9517), .CK(clk), .Q(\fmem_data[3][5] ) );
  DFF_X1 \fmem_inst/mem_reg[3][6]  ( .D(n9516), .CK(clk), .Q(\fmem_data[3][6] ) );
  DFF_X1 \fmem_inst/mem_reg[3][7]  ( .D(n9515), .CK(clk), .Q(\fmem_data[3][7] ) );
  DFF_X1 \fmem_inst/mem_reg[4][0]  ( .D(n9514), .CK(clk), .Q(\fmem_data[4][0] ) );
  DFF_X1 \fmem_inst/mem_reg[4][1]  ( .D(n9513), .CK(clk), .Q(\fmem_data[4][1] ) );
  DFF_X1 \fmem_inst/mem_reg[4][2]  ( .D(n9512), .CK(clk), .Q(\fmem_data[4][2] ) );
  DFF_X1 \fmem_inst/mem_reg[4][3]  ( .D(n9511), .CK(clk), .Q(\fmem_data[4][3] ) );
  DFF_X1 \fmem_inst/mem_reg[4][4]  ( .D(n9510), .CK(clk), .Q(\fmem_data[4][4] ) );
  DFF_X1 \fmem_inst/mem_reg[4][5]  ( .D(n9509), .CK(clk), .Q(\fmem_data[4][5] ) );
  DFF_X1 \fmem_inst/mem_reg[4][6]  ( .D(n9508), .CK(clk), .Q(\fmem_data[4][6] ) );
  DFF_X1 \fmem_inst/mem_reg[5][0]  ( .D(n9507), .CK(clk), .Q(\fmem_data[5][0] ) );
  DFF_X1 \fmem_inst/mem_reg[5][1]  ( .D(n9506), .CK(clk), .Q(\fmem_data[5][1] ) );
  DFF_X1 \fmem_inst/mem_reg[5][2]  ( .D(n9505), .CK(clk), .Q(\fmem_data[5][2] ) );
  DFF_X1 \fmem_inst/mem_reg[5][3]  ( .D(n9504), .CK(clk), .Q(\fmem_data[5][3] ) );
  DFF_X1 \fmem_inst/mem_reg[5][4]  ( .D(n9503), .CK(clk), .Q(\fmem_data[5][4] ) );
  DFF_X1 \fmem_inst/mem_reg[5][5]  ( .D(n9502), .CK(clk), .Q(\fmem_data[5][5] ) );
  DFF_X1 \fmem_inst/mem_reg[5][6]  ( .D(n9501), .CK(clk), .Q(\fmem_data[5][6] ) );
  DFF_X1 \fmem_inst/mem_reg[5][7]  ( .D(n9500), .CK(clk), .Q(\fmem_data[5][7] ) );
  DFF_X1 \fmem_inst/mem_reg[6][0]  ( .D(n9499), .CK(clk), .Q(\fmem_data[6][0] ) );
  DFF_X1 \fmem_inst/mem_reg[6][1]  ( .D(n9498), .CK(clk), .Q(\fmem_data[6][1] ) );
  DFF_X1 \fmem_inst/mem_reg[6][2]  ( .D(n9497), .CK(clk), .Q(\fmem_data[6][2] ) );
  DFF_X1 \fmem_inst/mem_reg[6][3]  ( .D(n9496), .CK(clk), .Q(\fmem_data[6][3] ) );
  DFF_X1 \fmem_inst/mem_reg[6][4]  ( .D(n9495), .CK(clk), .Q(\fmem_data[6][4] ) );
  DFF_X1 \fmem_inst/mem_reg[6][5]  ( .D(n9494), .CK(clk), .Q(\fmem_data[6][5] ) );
  DFF_X1 \fmem_inst/mem_reg[6][6]  ( .D(n9493), .CK(clk), .Q(\fmem_data[6][6] ) );
  DFF_X1 \fmem_inst/mem_reg[6][7]  ( .D(n9492), .CK(clk), .Q(\fmem_data[6][7] ) );
  DFF_X1 \fmem_inst/mem_reg[7][0]  ( .D(n9491), .CK(clk), .Q(\fmem_data[7][0] ) );
  DFF_X1 \fmem_inst/mem_reg[7][1]  ( .D(n9490), .CK(clk), .Q(\fmem_data[7][1] ) );
  DFF_X1 \fmem_inst/mem_reg[7][2]  ( .D(n9489), .CK(clk), .Q(\fmem_data[7][2] ) );
  DFF_X1 \fmem_inst/mem_reg[7][3]  ( .D(n9488), .CK(clk), .Q(\fmem_data[7][3] ) );
  DFF_X1 \fmem_inst/mem_reg[7][4]  ( .D(n9487), .CK(clk), .Q(\fmem_data[7][4] ) );
  DFF_X1 \fmem_inst/mem_reg[7][5]  ( .D(n9486), .CK(clk), .Q(\fmem_data[7][5] ) );
  DFF_X1 \fmem_inst/mem_reg[7][6]  ( .D(n9485), .CK(clk), .Q(\fmem_data[7][6] ) );
  DFF_X1 \fmem_inst/mem_reg[7][7]  ( .D(n9484), .CK(clk), .Q(\fmem_data[7][7] ) );
  DFF_X1 \fmem_inst/mem_reg[16][0]  ( .D(n9483), .CK(clk), .Q(
        \fmem_data[16][0] ) );
  DFF_X1 \fmem_inst/mem_reg[16][1]  ( .D(n9482), .CK(clk), .Q(
        \fmem_data[16][1] ) );
  DFF_X1 \fmem_inst/mem_reg[16][2]  ( .D(n9481), .CK(clk), .Q(
        \fmem_data[16][2] ) );
  DFF_X1 \fmem_inst/mem_reg[16][3]  ( .D(n9480), .CK(clk), .Q(
        \fmem_data[16][3] ) );
  DFF_X1 \fmem_inst/mem_reg[16][4]  ( .D(n9479), .CK(clk), .Q(
        \fmem_data[16][4] ) );
  DFF_X1 \fmem_inst/mem_reg[16][5]  ( .D(n9478), .CK(clk), .Q(
        \fmem_data[16][5] ) );
  DFF_X1 \fmem_inst/mem_reg[16][6]  ( .D(n9477), .CK(clk), .Q(
        \fmem_data[16][6] ) );
  DFF_X1 \fmem_inst/mem_reg[16][7]  ( .D(n9476), .CK(clk), .Q(
        \fmem_data[16][7] ) );
  DFF_X1 \fmem_inst/mem_reg[17][0]  ( .D(n9475), .CK(clk), .Q(
        \fmem_data[17][0] ) );
  DFF_X1 \fmem_inst/mem_reg[17][1]  ( .D(n9474), .CK(clk), .Q(
        \fmem_data[17][1] ) );
  DFF_X1 \fmem_inst/mem_reg[17][2]  ( .D(n9473), .CK(clk), .Q(
        \fmem_data[17][2] ) );
  DFF_X1 \fmem_inst/mem_reg[17][3]  ( .D(n9472), .CK(clk), .Q(
        \fmem_data[17][3] ) );
  DFF_X1 \fmem_inst/mem_reg[17][4]  ( .D(n9471), .CK(clk), .Q(
        \fmem_data[17][4] ) );
  DFF_X1 \fmem_inst/mem_reg[17][5]  ( .D(n9470), .CK(clk), .Q(
        \fmem_data[17][5] ) );
  DFF_X1 \fmem_inst/mem_reg[17][6]  ( .D(n9469), .CK(clk), .Q(
        \fmem_data[17][6] ) );
  DFF_X1 \fmem_inst/mem_reg[17][7]  ( .D(n9468), .CK(clk), .Q(
        \fmem_data[17][7] ) );
  DFF_X1 \fmem_inst/mem_reg[18][0]  ( .D(n9467), .CK(clk), .Q(
        \fmem_data[18][0] ) );
  DFF_X1 \fmem_inst/mem_reg[18][1]  ( .D(n9466), .CK(clk), .Q(
        \fmem_data[18][1] ) );
  DFF_X1 \fmem_inst/mem_reg[18][2]  ( .D(n9465), .CK(clk), .Q(
        \fmem_data[18][2] ) );
  DFF_X1 \fmem_inst/mem_reg[18][3]  ( .D(n9464), .CK(clk), .Q(
        \fmem_data[18][3] ) );
  DFF_X1 \fmem_inst/mem_reg[18][4]  ( .D(n9463), .CK(clk), .Q(
        \fmem_data[18][4] ) );
  DFF_X1 \fmem_inst/mem_reg[18][5]  ( .D(n9462), .CK(clk), .Q(
        \fmem_data[18][5] ) );
  DFF_X1 \fmem_inst/mem_reg[18][6]  ( .D(n9461), .CK(clk), .Q(
        \fmem_data[18][6] ) );
  DFF_X1 \fmem_inst/mem_reg[18][7]  ( .D(n9460), .CK(clk), .Q(
        \fmem_data[18][7] ) );
  DFF_X1 \fmem_inst/mem_reg[19][0]  ( .D(n9459), .CK(clk), .Q(
        \fmem_data[19][0] ) );
  DFF_X1 \fmem_inst/mem_reg[19][1]  ( .D(n9458), .CK(clk), .Q(
        \fmem_data[19][1] ) );
  DFF_X1 \fmem_inst/mem_reg[19][2]  ( .D(n9457), .CK(clk), .Q(
        \fmem_data[19][2] ) );
  DFF_X1 \fmem_inst/mem_reg[19][3]  ( .D(n9456), .CK(clk), .Q(
        \fmem_data[19][3] ) );
  DFF_X1 \fmem_inst/mem_reg[19][4]  ( .D(n9455), .CK(clk), .Q(
        \fmem_data[19][4] ) );
  DFF_X1 \fmem_inst/mem_reg[19][5]  ( .D(n9454), .CK(clk), .Q(
        \fmem_data[19][5] ) );
  DFF_X1 \fmem_inst/mem_reg[19][6]  ( .D(n9453), .CK(clk), .Q(
        \fmem_data[19][6] ) );
  DFF_X1 \fmem_inst/mem_reg[19][7]  ( .D(n9452), .CK(clk), .Q(
        \fmem_data[19][7] ) );
  DFF_X1 \fmem_inst/mem_reg[20][0]  ( .D(n9451), .CK(clk), .Q(
        \fmem_data[20][0] ) );
  DFF_X1 \fmem_inst/mem_reg[20][1]  ( .D(n9450), .CK(clk), .Q(
        \fmem_data[20][1] ) );
  DFF_X1 \fmem_inst/mem_reg[20][2]  ( .D(n9449), .CK(clk), .Q(
        \fmem_data[20][2] ) );
  DFF_X1 \fmem_inst/mem_reg[20][3]  ( .D(n9448), .CK(clk), .Q(
        \fmem_data[20][3] ) );
  DFF_X1 \fmem_inst/mem_reg[20][4]  ( .D(n9447), .CK(clk), .Q(
        \fmem_data[20][4] ) );
  DFF_X1 \fmem_inst/mem_reg[20][5]  ( .D(n9446), .CK(clk), .Q(
        \fmem_data[20][5] ) );
  DFF_X1 \fmem_inst/mem_reg[20][6]  ( .D(n9445), .CK(clk), .Q(
        \fmem_data[20][6] ) );
  DFF_X1 \fmem_inst/mem_reg[20][7]  ( .D(n9444), .CK(clk), .Q(
        \fmem_data[20][7] ) );
  DFF_X1 \fmem_inst/mem_reg[21][0]  ( .D(n9443), .CK(clk), .Q(
        \fmem_data[21][0] ) );
  DFF_X1 \fmem_inst/mem_reg[21][1]  ( .D(n9442), .CK(clk), .Q(
        \fmem_data[21][1] ) );
  DFF_X1 \fmem_inst/mem_reg[21][2]  ( .D(n9441), .CK(clk), .Q(
        \fmem_data[21][2] ) );
  DFF_X1 \fmem_inst/mem_reg[21][3]  ( .D(n9440), .CK(clk), .Q(
        \fmem_data[21][3] ) );
  DFF_X1 \fmem_inst/mem_reg[21][4]  ( .D(n9439), .CK(clk), .Q(
        \fmem_data[21][4] ) );
  DFF_X1 \fmem_inst/mem_reg[21][5]  ( .D(n9438), .CK(clk), .Q(
        \fmem_data[21][5] ) );
  DFF_X1 \fmem_inst/mem_reg[21][6]  ( .D(n9437), .CK(clk), .Q(
        \fmem_data[21][6] ) );
  DFF_X1 \fmem_inst/mem_reg[21][7]  ( .D(n9436), .CK(clk), .Q(
        \fmem_data[21][7] ) );
  DFF_X1 \fmem_inst/mem_reg[22][0]  ( .D(n9435), .CK(clk), .Q(
        \fmem_data[22][0] ) );
  DFF_X1 \fmem_inst/mem_reg[22][1]  ( .D(n9434), .CK(clk), .Q(
        \fmem_data[22][1] ) );
  DFF_X1 \fmem_inst/mem_reg[22][2]  ( .D(n9433), .CK(clk), .Q(
        \fmem_data[22][2] ) );
  DFF_X1 \fmem_inst/mem_reg[22][3]  ( .D(n9432), .CK(clk), .Q(
        \fmem_data[22][3] ) );
  DFF_X1 \fmem_inst/mem_reg[22][4]  ( .D(n9431), .CK(clk), .Q(
        \fmem_data[22][4] ) );
  DFF_X1 \fmem_inst/mem_reg[22][5]  ( .D(n9430), .CK(clk), .Q(
        \fmem_data[22][5] ) );
  DFF_X1 \fmem_inst/mem_reg[22][6]  ( .D(n9429), .CK(clk), .Q(
        \fmem_data[22][6] ) );
  DFF_X1 \fmem_inst/mem_reg[22][7]  ( .D(n9428), .CK(clk), .Q(
        \fmem_data[22][7] ) );
  DFF_X1 \fmem_inst/mem_reg[23][0]  ( .D(n9427), .CK(clk), .Q(
        \fmem_data[23][0] ) );
  DFF_X1 \fmem_inst/mem_reg[23][1]  ( .D(n9426), .CK(clk), .Q(
        \fmem_data[23][1] ) );
  DFF_X1 \fmem_inst/mem_reg[23][2]  ( .D(n9425), .CK(clk), .Q(
        \fmem_data[23][2] ) );
  DFF_X1 \fmem_inst/mem_reg[23][3]  ( .D(n9424), .CK(clk), .Q(
        \fmem_data[23][3] ) );
  DFF_X1 \fmem_inst/mem_reg[23][4]  ( .D(n9423), .CK(clk), .Q(
        \fmem_data[23][4] ) );
  DFF_X1 \fmem_inst/mem_reg[23][5]  ( .D(n9422), .CK(clk), .Q(
        \fmem_data[23][5] ) );
  DFF_X1 \fmem_inst/mem_reg[23][6]  ( .D(n9421), .CK(clk), .Q(
        \fmem_data[23][6] ) );
  DFF_X1 \fmem_inst/mem_reg[23][7]  ( .D(n9420), .CK(clk), .Q(
        \fmem_data[23][7] ) );
  DFF_X1 \fmem_inst/mem_reg[24][0]  ( .D(n9419), .CK(clk), .Q(
        \fmem_data[24][0] ) );
  DFF_X1 \fmem_inst/mem_reg[24][1]  ( .D(n9418), .CK(clk), .Q(
        \fmem_data[24][1] ) );
  DFF_X1 \fmem_inst/mem_reg[24][2]  ( .D(n9417), .CK(clk), .Q(
        \fmem_data[24][2] ) );
  DFF_X1 \fmem_inst/mem_reg[24][3]  ( .D(n9416), .CK(clk), .Q(
        \fmem_data[24][3] ) );
  DFF_X1 \fmem_inst/mem_reg[24][4]  ( .D(n9415), .CK(clk), .Q(
        \fmem_data[24][4] ) );
  DFF_X1 \fmem_inst/mem_reg[24][5]  ( .D(n9414), .CK(clk), .Q(
        \fmem_data[24][5] ) );
  DFF_X1 \fmem_inst/mem_reg[24][6]  ( .D(n9413), .CK(clk), .Q(
        \fmem_data[24][6] ) );
  DFF_X1 \fmem_inst/mem_reg[24][7]  ( .D(n9412), .CK(clk), .Q(
        \fmem_data[24][7] ) );
  DFF_X1 \fmem_inst/mem_reg[25][0]  ( .D(n9411), .CK(clk), .Q(
        \fmem_data[25][0] ) );
  DFF_X1 \fmem_inst/mem_reg[25][1]  ( .D(n9410), .CK(clk), .Q(
        \fmem_data[25][1] ) );
  DFF_X1 \fmem_inst/mem_reg[25][2]  ( .D(n9409), .CK(clk), .Q(
        \fmem_data[25][2] ) );
  DFF_X1 \fmem_inst/mem_reg[25][3]  ( .D(n9408), .CK(clk), .Q(
        \fmem_data[25][3] ) );
  DFF_X1 \fmem_inst/mem_reg[25][4]  ( .D(n9407), .CK(clk), .Q(
        \fmem_data[25][4] ) );
  DFF_X1 \fmem_inst/mem_reg[25][5]  ( .D(n9406), .CK(clk), .Q(
        \fmem_data[25][5] ) );
  DFF_X1 \fmem_inst/mem_reg[25][6]  ( .D(n9405), .CK(clk), .Q(
        \fmem_data[25][6] ) );
  DFF_X1 \fmem_inst/mem_reg[25][7]  ( .D(n9404), .CK(clk), .Q(
        \fmem_data[25][7] ) );
  DFF_X1 \fmem_inst/mem_reg[26][0]  ( .D(n9403), .CK(clk), .Q(
        \fmem_data[26][0] ) );
  DFF_X1 \fmem_inst/mem_reg[26][1]  ( .D(n9402), .CK(clk), .Q(
        \fmem_data[26][1] ) );
  DFF_X1 \fmem_inst/mem_reg[26][2]  ( .D(n9401), .CK(clk), .Q(
        \fmem_data[26][2] ) );
  DFF_X1 \fmem_inst/mem_reg[26][3]  ( .D(n9400), .CK(clk), .Q(
        \fmem_data[26][3] ) );
  DFF_X1 \fmem_inst/mem_reg[26][4]  ( .D(n9399), .CK(clk), .Q(
        \fmem_data[26][4] ) );
  DFF_X1 \fmem_inst/mem_reg[26][5]  ( .D(n9398), .CK(clk), .Q(
        \fmem_data[26][5] ) );
  DFF_X1 \fmem_inst/mem_reg[26][6]  ( .D(n9397), .CK(clk), .Q(
        \fmem_data[26][6] ) );
  DFF_X1 \fmem_inst/mem_reg[26][7]  ( .D(n9396), .CK(clk), .Q(
        \fmem_data[26][7] ) );
  DFF_X1 \fmem_inst/mem_reg[27][0]  ( .D(n9395), .CK(clk), .Q(
        \fmem_data[27][0] ) );
  DFF_X1 \fmem_inst/mem_reg[27][1]  ( .D(n9394), .CK(clk), .Q(
        \fmem_data[27][1] ) );
  DFF_X1 \fmem_inst/mem_reg[27][2]  ( .D(n9393), .CK(clk), .Q(
        \fmem_data[27][2] ) );
  DFF_X1 \fmem_inst/mem_reg[27][3]  ( .D(n9392), .CK(clk), .Q(
        \fmem_data[27][3] ) );
  DFF_X1 \fmem_inst/mem_reg[27][4]  ( .D(n9391), .CK(clk), .Q(
        \fmem_data[27][4] ) );
  DFF_X1 \fmem_inst/mem_reg[27][5]  ( .D(n9390), .CK(clk), .Q(
        \fmem_data[27][5] ) );
  DFF_X1 \fmem_inst/mem_reg[27][6]  ( .D(n9389), .CK(clk), .Q(
        \fmem_data[27][6] ) );
  DFF_X1 \fmem_inst/mem_reg[27][7]  ( .D(n9388), .CK(clk), .Q(
        \fmem_data[27][7] ) );
  DFF_X1 \fmem_inst/mem_reg[28][0]  ( .D(n9387), .CK(clk), .Q(
        \fmem_data[28][0] ) );
  DFF_X1 \fmem_inst/mem_reg[28][1]  ( .D(n9386), .CK(clk), .Q(
        \fmem_data[28][1] ) );
  DFF_X1 \fmem_inst/mem_reg[28][2]  ( .D(n9385), .CK(clk), .Q(
        \fmem_data[28][2] ) );
  DFF_X1 \fmem_inst/mem_reg[28][3]  ( .D(n9384), .CK(clk), .Q(
        \fmem_data[28][3] ) );
  DFF_X1 \fmem_inst/mem_reg[28][4]  ( .D(n9383), .CK(clk), .Q(
        \fmem_data[28][4] ) );
  DFF_X1 \fmem_inst/mem_reg[28][5]  ( .D(n9382), .CK(clk), .Q(
        \fmem_data[28][5] ) );
  DFF_X1 \fmem_inst/mem_reg[28][6]  ( .D(n9381), .CK(clk), .Q(
        \fmem_data[28][6] ) );
  DFF_X1 \fmem_inst/mem_reg[28][7]  ( .D(n9380), .CK(clk), .Q(
        \fmem_data[28][7] ) );
  DFF_X1 \fmem_inst/mem_reg[29][0]  ( .D(n9379), .CK(clk), .Q(
        \fmem_data[29][0] ) );
  DFF_X1 \fmem_inst/mem_reg[29][1]  ( .D(n9378), .CK(clk), .Q(
        \fmem_data[29][1] ) );
  DFF_X1 \fmem_inst/mem_reg[29][2]  ( .D(n9377), .CK(clk), .Q(
        \fmem_data[29][2] ) );
  DFF_X1 \fmem_inst/mem_reg[29][3]  ( .D(n9376), .CK(clk), .Q(
        \fmem_data[29][3] ) );
  DFF_X1 \fmem_inst/mem_reg[29][4]  ( .D(n9375), .CK(clk), .Q(
        \fmem_data[29][4] ) );
  DFF_X1 \fmem_inst/mem_reg[29][5]  ( .D(n9374), .CK(clk), .Q(
        \fmem_data[29][5] ) );
  DFF_X1 \fmem_inst/mem_reg[29][6]  ( .D(n9373), .CK(clk), .Q(
        \fmem_data[29][6] ) );
  DFF_X1 \fmem_inst/mem_reg[29][7]  ( .D(n9372), .CK(clk), .Q(
        \fmem_data[29][7] ) );
  DFF_X1 \fmem_inst/mem_reg[30][0]  ( .D(n9371), .CK(clk), .Q(
        \fmem_data[30][0] ) );
  DFF_X1 \fmem_inst/mem_reg[30][1]  ( .D(n9370), .CK(clk), .Q(
        \fmem_data[30][1] ) );
  DFF_X1 \fmem_inst/mem_reg[30][2]  ( .D(n9369), .CK(clk), .Q(
        \fmem_data[30][2] ) );
  DFF_X1 \fmem_inst/mem_reg[30][3]  ( .D(n9368), .CK(clk), .Q(
        \fmem_data[30][3] ) );
  DFF_X1 \fmem_inst/mem_reg[30][4]  ( .D(n9367), .CK(clk), .Q(
        \fmem_data[30][4] ) );
  DFF_X1 \fmem_inst/mem_reg[30][5]  ( .D(n9366), .CK(clk), .Q(
        \fmem_data[30][5] ) );
  DFF_X1 \fmem_inst/mem_reg[30][6]  ( .D(n9365), .CK(clk), .Q(
        \fmem_data[30][6] ) );
  DFF_X1 \fmem_inst/mem_reg[30][7]  ( .D(n9364), .CK(clk), .Q(
        \fmem_data[30][7] ) );
  DFF_X1 \fmem_inst/mem_reg[31][0]  ( .D(n9363), .CK(clk), .Q(
        \fmem_data[31][0] ) );
  DFF_X1 \fmem_inst/mem_reg[31][1]  ( .D(n9362), .CK(clk), .Q(
        \fmem_data[31][1] ) );
  DFF_X1 \fmem_inst/mem_reg[31][2]  ( .D(n9361), .CK(clk), .Q(
        \fmem_data[31][2] ) );
  DFF_X1 \fmem_inst/mem_reg[31][3]  ( .D(n9360), .CK(clk), .Q(
        \fmem_data[31][3] ) );
  DFF_X1 \fmem_inst/mem_reg[31][4]  ( .D(n9359), .CK(clk), .Q(
        \fmem_data[31][4] ) );
  DFF_X1 \fmem_inst/mem_reg[31][5]  ( .D(n9358), .CK(clk), .Q(
        \fmem_data[31][5] ) );
  DFF_X1 \fmem_inst/mem_reg[31][6]  ( .D(n9357), .CK(clk), .Q(
        \fmem_data[31][6] ) );
  DFF_X1 \fmem_inst/mem_reg[31][7]  ( .D(n9356), .CK(clk), .Q(
        \fmem_data[31][7] ) );
  DFF_X1 \x_mult_f_reg[0][0]  ( .D(n9293), .CK(clk), .Q(\x_mult_f[0][0] ) );
  DFF_X1 \x_mult_f_reg[0][1]  ( .D(n9292), .CK(clk), .Q(\x_mult_f[0][1] ) );
  DFF_X1 \x_mult_f_reg[0][4]  ( .D(n8934), .CK(clk), .Q(\x_mult_f[0][4] ) );
  DFF_X1 \x_mult_f_reg[0][6]  ( .D(n8933), .CK(clk), .Q(\x_mult_f[0][6] ) );
  DFF_X1 \x_mult_f_reg[0][7]  ( .D(n8932), .CK(clk), .Q(\x_mult_f[0][7] ) );
  DFF_X1 \x_mult_f_reg[0][9]  ( .D(n8931), .CK(clk), .Q(\x_mult_f[0][9] ) );
  DFF_X1 \x_mult_f_reg[0][10]  ( .D(n8930), .CK(clk), .Q(\x_mult_f[0][10] ) );
  DFF_X1 \x_mult_f_reg[0][11]  ( .D(n8929), .CK(clk), .Q(\x_mult_f[0][11] ) );
  DFF_X1 \x_mult_f_reg[0][12]  ( .D(n8928), .CK(clk), .Q(\x_mult_f[0][12] ) );
  DFF_X1 \x_mult_f_reg[0][13]  ( .D(n8927), .CK(clk), .Q(\x_mult_f[0][13] ) );
  DFF_X1 \x_mult_f_reg[0][14]  ( .D(n8926), .CK(clk), .Q(\x_mult_f[0][14] ) );
  DFF_X1 \x_mult_f_reg[0][15]  ( .D(n8925), .CK(clk), .Q(\x_mult_f[0][15] ), 
        .QN(n3463) );
  DFF_X1 \x_mult_f_reg[1][0]  ( .D(n9295), .CK(clk), .Q(\x_mult_f[1][0] ) );
  DFF_X1 \x_mult_f_reg[1][1]  ( .D(n9294), .CK(clk), .Q(\x_mult_f[1][1] ) );
  DFF_X1 \x_mult_f_reg[1][2]  ( .D(n8946), .CK(clk), .Q(\x_mult_f[1][2] ) );
  DFF_X1 \x_mult_f_reg[1][3]  ( .D(n8945), .CK(clk), .Q(\x_mult_f[1][3] ) );
  DFF_X1 \x_mult_f_reg[1][4]  ( .D(n8944), .CK(clk), .Q(\x_mult_f[1][4] ) );
  DFF_X1 \x_mult_f_reg[1][6]  ( .D(n8943), .CK(clk), .Q(\x_mult_f[1][6] ) );
  DFF_X1 \x_mult_f_reg[1][7]  ( .D(n8942), .CK(clk), .Q(\x_mult_f[1][7] ) );
  DFF_X1 \x_mult_f_reg[1][9]  ( .D(n8941), .CK(clk), .Q(\x_mult_f[1][9] ) );
  DFF_X1 \x_mult_f_reg[1][10]  ( .D(n8940), .CK(clk), .Q(\x_mult_f[1][10] ) );
  DFF_X1 \x_mult_f_reg[1][11]  ( .D(n8939), .CK(clk), .Q(\x_mult_f[1][11] ) );
  DFF_X1 \x_mult_f_reg[1][12]  ( .D(n8938), .CK(clk), .Q(\x_mult_f[1][12] ) );
  DFF_X1 \x_mult_f_reg[1][13]  ( .D(n8937), .CK(clk), .Q(\x_mult_f[1][13] ) );
  DFF_X1 \x_mult_f_reg[1][14]  ( .D(n8936), .CK(clk), .Q(\x_mult_f[1][14] ) );
  DFF_X1 \x_mult_f_reg[1][15]  ( .D(n8935), .CK(clk), .Q(\x_mult_f[1][15] ), 
        .QN(n3497) );
  DFF_X1 \x_mult_f_reg[2][0]  ( .D(n9297), .CK(clk), .Q(\x_mult_f[2][0] ) );
  DFF_X1 \x_mult_f_reg[2][1]  ( .D(n9296), .CK(clk), .Q(\x_mult_f[2][1] ) );
  DFF_X1 \x_mult_f_reg[2][2]  ( .D(n8960), .CK(clk), .Q(\x_mult_f[2][2] ) );
  DFF_X1 \x_mult_f_reg[2][3]  ( .D(n8959), .CK(clk), .Q(\x_mult_f[2][3] ) );
  DFF_X1 \x_mult_f_reg[2][4]  ( .D(n8958), .CK(clk), .Q(\x_mult_f[2][4] ) );
  DFF_X1 \x_mult_f_reg[2][5]  ( .D(n8957), .CK(clk), .Q(\x_mult_f[2][5] ) );
  DFF_X1 \x_mult_f_reg[2][6]  ( .D(n8956), .CK(clk), .Q(\x_mult_f[2][6] ) );
  DFF_X1 \x_mult_f_reg[2][7]  ( .D(n8955), .CK(clk), .Q(\x_mult_f[2][7] ) );
  DFF_X1 \x_mult_f_reg[2][8]  ( .D(n8954), .CK(clk), .Q(\x_mult_f[2][8] ) );
  DFF_X1 \x_mult_f_reg[2][9]  ( .D(n8953), .CK(clk), .Q(\x_mult_f[2][9] ) );
  DFF_X1 \x_mult_f_reg[2][10]  ( .D(n8952), .CK(clk), .Q(\x_mult_f[2][10] ) );
  DFF_X1 \x_mult_f_reg[2][11]  ( .D(n8951), .CK(clk), .Q(\x_mult_f[2][11] ) );
  DFF_X1 \x_mult_f_reg[2][12]  ( .D(n8950), .CK(clk), .Q(\x_mult_f[2][12] ) );
  DFF_X1 \x_mult_f_reg[2][13]  ( .D(n8949), .CK(clk), .Q(\x_mult_f[2][13] ) );
  DFF_X1 \x_mult_f_reg[2][14]  ( .D(n8948), .CK(clk), .Q(\x_mult_f[2][14] ), 
        .QN(n3473) );
  DFF_X1 \x_mult_f_reg[2][15]  ( .D(n8947), .CK(clk), .Q(\x_mult_f[2][15] ), 
        .QN(n3476) );
  DFF_X1 \x_mult_f_reg[3][0]  ( .D(n9299), .CK(clk), .Q(\x_mult_f[3][0] ) );
  DFF_X1 \x_mult_f_reg[3][1]  ( .D(n9298), .CK(clk), .Q(\x_mult_f[3][1] ) );
  DFF_X1 \x_mult_f_reg[3][2]  ( .D(n8973), .CK(clk), .Q(\x_mult_f[3][2] ) );
  DFF_X1 \x_mult_f_reg[3][3]  ( .D(n8972), .CK(clk), .Q(\x_mult_f[3][3] ) );
  DFF_X1 \x_mult_f_reg[3][4]  ( .D(n8971), .CK(clk), .Q(\x_mult_f[3][4] ) );
  DFF_X1 \x_mult_f_reg[3][5]  ( .D(n8970), .CK(clk), .Q(\x_mult_f[3][5] ) );
  DFF_X1 \x_mult_f_reg[3][6]  ( .D(n8969), .CK(clk), .Q(\x_mult_f[3][6] ) );
  DFF_X1 \x_mult_f_reg[3][8]  ( .D(n8968), .CK(clk), .Q(\x_mult_f[3][8] ) );
  DFF_X1 \x_mult_f_reg[3][9]  ( .D(n8967), .CK(clk), .Q(\x_mult_f[3][9] ) );
  DFF_X1 \x_mult_f_reg[3][10]  ( .D(n8966), .CK(clk), .Q(\x_mult_f[3][10] ) );
  DFF_X1 \x_mult_f_reg[3][11]  ( .D(n8965), .CK(clk), .Q(\x_mult_f[3][11] ) );
  DFF_X1 \x_mult_f_reg[3][12]  ( .D(n8964), .CK(clk), .Q(\x_mult_f[3][12] ) );
  DFF_X1 \x_mult_f_reg[3][13]  ( .D(n8963), .CK(clk), .Q(\x_mult_f[3][13] ) );
  DFF_X1 \x_mult_f_reg[3][14]  ( .D(n8962), .CK(clk), .Q(\x_mult_f[3][14] ), 
        .QN(n3509) );
  DFF_X1 \x_mult_f_reg[3][15]  ( .D(n8961), .CK(clk), .Q(\x_mult_f[3][15] ), 
        .QN(n3451) );
  DFF_X1 \x_mult_f_reg[4][0]  ( .D(n9301), .CK(clk), .Q(\x_mult_f[4][0] ) );
  DFF_X1 \x_mult_f_reg[4][1]  ( .D(n9300), .CK(clk), .Q(\x_mult_f[4][1] ) );
  DFF_X1 \x_mult_f_reg[4][2]  ( .D(n8987), .CK(clk), .Q(\x_mult_f[4][2] ) );
  DFF_X1 \x_mult_f_reg[4][3]  ( .D(n8986), .CK(clk), .Q(\x_mult_f[4][3] ) );
  DFF_X1 \x_mult_f_reg[4][4]  ( .D(n8985), .CK(clk), .Q(\x_mult_f[4][4] ) );
  DFF_X1 \x_mult_f_reg[4][5]  ( .D(n8984), .CK(clk), .Q(\x_mult_f[4][5] ) );
  DFF_X1 \x_mult_f_reg[4][6]  ( .D(n8983), .CK(clk), .Q(\x_mult_f[4][6] ) );
  DFF_X1 \x_mult_f_reg[4][7]  ( .D(n8982), .CK(clk), .Q(\x_mult_f[4][7] ) );
  DFF_X1 \x_mult_f_reg[4][8]  ( .D(n8981), .CK(clk), .Q(\x_mult_f[4][8] ) );
  DFF_X1 \x_mult_f_reg[4][9]  ( .D(n8980), .CK(clk), .Q(\x_mult_f[4][9] ) );
  DFF_X1 \x_mult_f_reg[4][10]  ( .D(n8979), .CK(clk), .Q(\x_mult_f[4][10] ) );
  DFF_X1 \x_mult_f_reg[4][11]  ( .D(n8978), .CK(clk), .Q(\x_mult_f[4][11] ) );
  DFF_X1 \x_mult_f_reg[4][12]  ( .D(n8977), .CK(clk), .Q(\x_mult_f[4][12] ) );
  DFF_X1 \x_mult_f_reg[4][13]  ( .D(n8976), .CK(clk), .Q(\x_mult_f[4][13] ) );
  DFF_X1 \x_mult_f_reg[4][14]  ( .D(n8975), .CK(clk), .Q(\x_mult_f[4][14] ) );
  DFF_X1 \x_mult_f_reg[4][15]  ( .D(n8974), .CK(clk), .Q(\x_mult_f[4][15] ), 
        .QN(n3478) );
  DFF_X1 \x_mult_f_reg[5][0]  ( .D(n9303), .CK(clk), .Q(\x_mult_f[5][0] ) );
  DFF_X1 \x_mult_f_reg[5][1]  ( .D(n9302), .CK(clk), .Q(\x_mult_f[5][1] ) );
  DFF_X1 \x_mult_f_reg[5][2]  ( .D(n8998), .CK(clk), .Q(\x_mult_f[5][2] ) );
  DFF_X1 \x_mult_f_reg[5][3]  ( .D(n8997), .CK(clk), .Q(\x_mult_f[5][3] ) );
  DFF_X1 \x_mult_f_reg[5][4]  ( .D(n8996), .CK(clk), .Q(\x_mult_f[5][4] ) );
  DFF_X1 \x_mult_f_reg[5][5]  ( .D(n8995), .CK(clk), .Q(\x_mult_f[5][5] ) );
  DFF_X1 \x_mult_f_reg[5][6]  ( .D(n8994), .CK(clk), .Q(\x_mult_f[5][6] ) );
  DFF_X1 \x_mult_f_reg[5][7]  ( .D(n8993), .CK(clk), .Q(\x_mult_f[5][7] ) );
  DFF_X1 \x_mult_f_reg[5][8]  ( .D(n8992), .CK(clk), .Q(\x_mult_f[5][8] ) );
  DFF_X1 \x_mult_f_reg[5][9]  ( .D(n8991), .CK(clk), .Q(\x_mult_f[5][9] ) );
  DFF_X1 \x_mult_f_reg[5][10]  ( .D(n8990), .CK(clk), .Q(\x_mult_f[5][10] ) );
  DFF_X1 \x_mult_f_reg[5][11]  ( .D(n8989), .CK(clk), .Q(\x_mult_f[5][11] ) );
  DFF_X1 \x_mult_f_reg[5][12]  ( .D(n8988), .CK(clk), .Q(\x_mult_f[5][12] ) );
  DFF_X1 \x_mult_f_reg[6][0]  ( .D(n9305), .CK(clk), .Q(\x_mult_f[6][0] ) );
  DFF_X1 \x_mult_f_reg[6][1]  ( .D(n9304), .CK(clk), .Q(\x_mult_f[6][1] ) );
  DFF_X1 \x_mult_f_reg[6][2]  ( .D(n9012), .CK(clk), .Q(\x_mult_f[6][2] ) );
  DFF_X1 \x_mult_f_reg[6][3]  ( .D(n9011), .CK(clk), .Q(\x_mult_f[6][3] ) );
  DFF_X1 \x_mult_f_reg[6][4]  ( .D(n9010), .CK(clk), .Q(\x_mult_f[6][4] ) );
  DFF_X1 \x_mult_f_reg[6][5]  ( .D(n9009), .CK(clk), .Q(\x_mult_f[6][5] ) );
  DFF_X1 \x_mult_f_reg[6][6]  ( .D(n9008), .CK(clk), .Q(\x_mult_f[6][6] ) );
  DFF_X1 \x_mult_f_reg[6][7]  ( .D(n9007), .CK(clk), .Q(\x_mult_f[6][7] ) );
  DFF_X1 \x_mult_f_reg[6][8]  ( .D(n9006), .CK(clk), .Q(\x_mult_f[6][8] ) );
  DFF_X1 \x_mult_f_reg[6][9]  ( .D(n9005), .CK(clk), .Q(\x_mult_f[6][9] ) );
  DFF_X1 \x_mult_f_reg[6][10]  ( .D(n9004), .CK(clk), .Q(\x_mult_f[6][10] ) );
  DFF_X1 \x_mult_f_reg[6][11]  ( .D(n9003), .CK(clk), .Q(\x_mult_f[6][11] ) );
  DFF_X1 \x_mult_f_reg[6][12]  ( .D(n9002), .CK(clk), .Q(\x_mult_f[6][12] ) );
  DFF_X1 \x_mult_f_reg[6][13]  ( .D(n9001), .CK(clk), .Q(\x_mult_f[6][13] ) );
  DFF_X1 \x_mult_f_reg[6][14]  ( .D(n9000), .CK(clk), .Q(\x_mult_f[6][14] ) );
  DFF_X1 \x_mult_f_reg[6][15]  ( .D(n8999), .CK(clk), .Q(\x_mult_f[6][15] ), 
        .QN(n3459) );
  DFF_X1 \x_mult_f_reg[7][0]  ( .D(n9307), .CK(clk), .Q(\x_mult_f[7][0] ) );
  DFF_X1 \x_mult_f_reg[7][1]  ( .D(n9306), .CK(clk), .Q(\x_mult_f[7][1] ) );
  DFF_X1 \x_mult_f_reg[7][2]  ( .D(n9026), .CK(clk), .Q(\x_mult_f[7][2] ) );
  DFF_X1 \x_mult_f_reg[7][3]  ( .D(n9025), .CK(clk), .Q(\x_mult_f[7][3] ) );
  DFF_X1 \x_mult_f_reg[7][4]  ( .D(n9024), .CK(clk), .Q(\x_mult_f[7][4] ) );
  DFF_X1 \x_mult_f_reg[7][5]  ( .D(n9023), .CK(clk), .Q(\x_mult_f[7][5] ) );
  DFF_X1 \x_mult_f_reg[7][6]  ( .D(n9022), .CK(clk), .Q(\x_mult_f[7][6] ) );
  DFF_X1 \x_mult_f_reg[7][7]  ( .D(n9021), .CK(clk), .Q(\x_mult_f[7][7] ) );
  DFF_X1 \x_mult_f_reg[7][8]  ( .D(n9020), .CK(clk), .Q(\x_mult_f[7][8] ) );
  DFF_X1 \x_mult_f_reg[7][9]  ( .D(n9019), .CK(clk), .Q(\x_mult_f[7][9] ) );
  DFF_X1 \x_mult_f_reg[7][10]  ( .D(n9018), .CK(clk), .Q(\x_mult_f[7][10] ) );
  DFF_X1 \x_mult_f_reg[7][11]  ( .D(n9017), .CK(clk), .Q(\x_mult_f[7][11] ) );
  DFF_X1 \x_mult_f_reg[7][12]  ( .D(n9016), .CK(clk), .Q(\x_mult_f[7][12] ) );
  DFF_X1 \x_mult_f_reg[7][13]  ( .D(n9015), .CK(clk), .Q(\x_mult_f[7][13] ) );
  DFF_X1 \x_mult_f_reg[7][14]  ( .D(n9014), .CK(clk), .Q(\x_mult_f[7][14] ) );
  DFF_X1 \x_mult_f_reg[7][15]  ( .D(n9013), .CK(clk), .Q(\x_mult_f[7][15] ), 
        .QN(n3489) );
  DFF_X1 \x_mult_f_reg[8][0]  ( .D(n9309), .CK(clk), .Q(\x_mult_f[8][0] ) );
  DFF_X1 \x_mult_f_reg[8][1]  ( .D(n9308), .CK(clk), .Q(\x_mult_f[8][1] ) );
  DFF_X1 \x_mult_f_reg[8][2]  ( .D(n9040), .CK(clk), .Q(\x_mult_f[8][2] ) );
  DFF_X1 \x_mult_f_reg[8][3]  ( .D(n9039), .CK(clk), .Q(\x_mult_f[8][3] ) );
  DFF_X1 \x_mult_f_reg[8][4]  ( .D(n9038), .CK(clk), .Q(\x_mult_f[8][4] ) );
  DFF_X1 \x_mult_f_reg[8][5]  ( .D(n9037), .CK(clk), .Q(\x_mult_f[8][5] ) );
  DFF_X1 \x_mult_f_reg[8][6]  ( .D(n9036), .CK(clk), .Q(\x_mult_f[8][6] ) );
  DFF_X1 \x_mult_f_reg[8][7]  ( .D(n9035), .CK(clk), .Q(\x_mult_f[8][7] ) );
  DFF_X1 \x_mult_f_reg[8][8]  ( .D(n9034), .CK(clk), .Q(\x_mult_f[8][8] ) );
  DFF_X1 \x_mult_f_reg[8][9]  ( .D(n9033), .CK(clk), .Q(\x_mult_f[8][9] ) );
  DFF_X1 \x_mult_f_reg[8][10]  ( .D(n9032), .CK(clk), .Q(\x_mult_f[8][10] ) );
  DFF_X1 \x_mult_f_reg[8][11]  ( .D(n9031), .CK(clk), .Q(\x_mult_f[8][11] ) );
  DFF_X1 \x_mult_f_reg[8][12]  ( .D(n9030), .CK(clk), .Q(\x_mult_f[8][12] ) );
  DFF_X1 \x_mult_f_reg[8][13]  ( .D(n9029), .CK(clk), .Q(\x_mult_f[8][13] ) );
  DFF_X1 \x_mult_f_reg[8][14]  ( .D(n9028), .CK(clk), .Q(\x_mult_f[8][14] ) );
  DFF_X1 \x_mult_f_reg[8][15]  ( .D(n9027), .CK(clk), .Q(\x_mult_f[8][15] ), 
        .QN(n3481) );
  DFF_X1 \x_mult_f_reg[9][0]  ( .D(n9311), .CK(clk), .Q(\x_mult_f[9][0] ) );
  DFF_X1 \x_mult_f_reg[9][1]  ( .D(n9310), .CK(clk), .Q(\x_mult_f[9][1] ) );
  DFF_X1 \x_mult_f_reg[9][2]  ( .D(n9045), .CK(clk), .Q(\x_mult_f[9][2] ) );
  DFF_X1 \x_mult_f_reg[9][3]  ( .D(n9044), .CK(clk), .Q(\x_mult_f[9][3] ) );
  DFF_X1 \x_mult_f_reg[9][4]  ( .D(n9043), .CK(clk), .Q(\x_mult_f[9][4] ) );
  DFF_X1 \x_mult_f_reg[9][5]  ( .D(n9042), .CK(clk), .Q(\x_mult_f[9][5] ) );
  DFF_X1 \x_mult_f_reg[9][7]  ( .D(n9041), .CK(clk), .Q(\x_mult_f[9][7] ) );
  DFF_X1 \x_mult_f_reg[10][0]  ( .D(n9313), .CK(clk), .Q(\x_mult_f[10][0] ) );
  DFF_X1 \x_mult_f_reg[10][1]  ( .D(n9312), .CK(clk), .Q(\x_mult_f[10][1] ) );
  DFF_X1 \x_mult_f_reg[10][3]  ( .D(n9057), .CK(clk), .Q(\x_mult_f[10][3] ) );
  DFF_X1 \x_mult_f_reg[10][5]  ( .D(n9056), .CK(clk), .Q(\x_mult_f[10][5] ) );
  DFF_X1 \x_mult_f_reg[10][6]  ( .D(n9055), .CK(clk), .Q(\x_mult_f[10][6] ) );
  DFF_X1 \x_mult_f_reg[10][7]  ( .D(n9054), .CK(clk), .Q(\x_mult_f[10][7] ) );
  DFF_X1 \x_mult_f_reg[10][8]  ( .D(n9053), .CK(clk), .Q(\x_mult_f[10][8] ) );
  DFF_X1 \x_mult_f_reg[10][9]  ( .D(n9052), .CK(clk), .Q(\x_mult_f[10][9] ) );
  DFF_X1 \x_mult_f_reg[10][10]  ( .D(n9051), .CK(clk), .Q(\x_mult_f[10][10] )
         );
  DFF_X1 \x_mult_f_reg[10][11]  ( .D(n9050), .CK(clk), .Q(\x_mult_f[10][11] )
         );
  DFF_X1 \x_mult_f_reg[10][12]  ( .D(n9049), .CK(clk), .Q(\x_mult_f[10][12] )
         );
  DFF_X1 \x_mult_f_reg[10][13]  ( .D(n9048), .CK(clk), .Q(\x_mult_f[10][13] )
         );
  DFF_X1 \x_mult_f_reg[10][14]  ( .D(n9047), .CK(clk), .Q(\x_mult_f[10][14] )
         );
  DFF_X1 \x_mult_f_reg[10][15]  ( .D(n9046), .CK(clk), .Q(\x_mult_f[10][15] ), 
        .QN(n3454) );
  DFF_X1 \x_mult_f_reg[11][0]  ( .D(n9315), .CK(clk), .Q(\x_mult_f[11][0] ) );
  DFF_X1 \x_mult_f_reg[11][1]  ( .D(n9314), .CK(clk), .Q(\x_mult_f[11][1] ) );
  DFF_X1 \x_mult_f_reg[11][2]  ( .D(n9071), .CK(clk), .Q(\x_mult_f[11][2] ) );
  DFF_X1 \x_mult_f_reg[11][3]  ( .D(n9070), .CK(clk), .Q(\x_mult_f[11][3] ) );
  DFF_X1 \x_mult_f_reg[11][4]  ( .D(n9069), .CK(clk), .Q(\x_mult_f[11][4] ) );
  DFF_X1 \x_mult_f_reg[11][5]  ( .D(n9068), .CK(clk), .Q(\x_mult_f[11][5] ) );
  DFF_X1 \x_mult_f_reg[11][6]  ( .D(n9067), .CK(clk), .Q(\x_mult_f[11][6] ) );
  DFF_X1 \x_mult_f_reg[11][7]  ( .D(n9066), .CK(clk), .Q(\x_mult_f[11][7] ) );
  DFF_X1 \x_mult_f_reg[11][8]  ( .D(n9065), .CK(clk), .Q(\x_mult_f[11][8] ) );
  DFF_X1 \x_mult_f_reg[11][9]  ( .D(n9064), .CK(clk), .Q(\x_mult_f[11][9] ) );
  DFF_X1 \x_mult_f_reg[11][10]  ( .D(n9063), .CK(clk), .Q(\x_mult_f[11][10] )
         );
  DFF_X1 \x_mult_f_reg[11][11]  ( .D(n9062), .CK(clk), .Q(\x_mult_f[11][11] )
         );
  DFF_X1 \x_mult_f_reg[11][12]  ( .D(n9061), .CK(clk), .Q(\x_mult_f[11][12] )
         );
  DFF_X1 \x_mult_f_reg[11][13]  ( .D(n9060), .CK(clk), .Q(\x_mult_f[11][13] )
         );
  DFF_X1 \x_mult_f_reg[11][14]  ( .D(n9059), .CK(clk), .Q(\x_mult_f[11][14] )
         );
  DFF_X1 \x_mult_f_reg[11][15]  ( .D(n9058), .CK(clk), .Q(\x_mult_f[11][15] ), 
        .QN(n3484) );
  DFF_X1 \x_mult_f_reg[12][0]  ( .D(n9317), .CK(clk), .Q(\x_mult_f[12][0] ) );
  DFF_X1 \x_mult_f_reg[12][1]  ( .D(n9316), .CK(clk), .Q(\x_mult_f[12][1] ) );
  DFF_X1 \x_mult_f_reg[12][2]  ( .D(n9084), .CK(clk), .Q(\x_mult_f[12][2] ) );
  DFF_X1 \x_mult_f_reg[12][3]  ( .D(n9083), .CK(clk), .Q(\x_mult_f[12][3] ) );
  DFF_X1 \x_mult_f_reg[12][5]  ( .D(n9082), .CK(clk), .Q(\x_mult_f[12][5] ) );
  DFF_X1 \x_mult_f_reg[12][6]  ( .D(n9081), .CK(clk), .Q(\x_mult_f[12][6] ) );
  DFF_X1 \x_mult_f_reg[12][7]  ( .D(n9080), .CK(clk), .Q(\x_mult_f[12][7] ) );
  DFF_X1 \x_mult_f_reg[12][8]  ( .D(n9079), .CK(clk), .Q(\x_mult_f[12][8] ) );
  DFF_X1 \x_mult_f_reg[12][9]  ( .D(n9078), .CK(clk), .Q(\x_mult_f[12][9] ) );
  DFF_X1 \x_mult_f_reg[12][10]  ( .D(n9077), .CK(clk), .Q(\x_mult_f[12][10] )
         );
  DFF_X1 \x_mult_f_reg[12][11]  ( .D(n9076), .CK(clk), .Q(\x_mult_f[12][11] )
         );
  DFF_X1 \x_mult_f_reg[12][12]  ( .D(n9075), .CK(clk), .Q(\x_mult_f[12][12] )
         );
  DFF_X1 \x_mult_f_reg[12][13]  ( .D(n9074), .CK(clk), .Q(\x_mult_f[12][13] )
         );
  DFF_X1 \x_mult_f_reg[12][14]  ( .D(n9073), .CK(clk), .Q(\x_mult_f[12][14] )
         );
  DFF_X1 \x_mult_f_reg[12][15]  ( .D(n9072), .CK(clk), .Q(\x_mult_f[12][15] ), 
        .QN(n3457) );
  DFF_X1 \x_mult_f_reg[13][0]  ( .D(n9319), .CK(clk), .Q(\x_mult_f[13][0] ) );
  DFF_X1 \x_mult_f_reg[13][1]  ( .D(n9318), .CK(clk), .Q(\x_mult_f[13][1] ) );
  DFF_X1 \x_mult_f_reg[13][2]  ( .D(n9098), .CK(clk), .Q(\x_mult_f[13][2] ) );
  DFF_X1 \x_mult_f_reg[13][3]  ( .D(n9097), .CK(clk), .Q(\x_mult_f[13][3] ) );
  DFF_X1 \x_mult_f_reg[13][4]  ( .D(n9096), .CK(clk), .Q(\x_mult_f[13][4] ) );
  DFF_X1 \x_mult_f_reg[13][5]  ( .D(n9095), .CK(clk), .Q(\x_mult_f[13][5] ) );
  DFF_X1 \x_mult_f_reg[13][6]  ( .D(n9094), .CK(clk), .Q(\x_mult_f[13][6] ) );
  DFF_X1 \x_mult_f_reg[13][7]  ( .D(n9093), .CK(clk), .Q(\x_mult_f[13][7] ) );
  DFF_X1 \x_mult_f_reg[13][8]  ( .D(n9092), .CK(clk), .Q(\x_mult_f[13][8] ) );
  DFF_X1 \x_mult_f_reg[13][9]  ( .D(n9091), .CK(clk), .Q(\x_mult_f[13][9] ) );
  DFF_X1 \x_mult_f_reg[13][10]  ( .D(n9090), .CK(clk), .Q(\x_mult_f[13][10] )
         );
  DFF_X1 \x_mult_f_reg[13][11]  ( .D(n9089), .CK(clk), .Q(\x_mult_f[13][11] )
         );
  DFF_X1 \x_mult_f_reg[13][12]  ( .D(n9088), .CK(clk), .Q(\x_mult_f[13][12] )
         );
  DFF_X1 \x_mult_f_reg[13][13]  ( .D(n9087), .CK(clk), .Q(\x_mult_f[13][13] )
         );
  DFF_X1 \x_mult_f_reg[13][14]  ( .D(n9086), .CK(clk), .Q(\x_mult_f[13][14] )
         );
  DFF_X1 \x_mult_f_reg[13][15]  ( .D(n9085), .CK(clk), .Q(\x_mult_f[13][15] ), 
        .QN(n3487) );
  DFF_X1 \x_mult_f_reg[14][0]  ( .D(n9321), .CK(clk), .Q(\x_mult_f[14][0] ) );
  DFF_X1 \x_mult_f_reg[14][1]  ( .D(n9320), .CK(clk), .Q(\x_mult_f[14][1] ) );
  DFF_X1 \x_mult_f_reg[14][2]  ( .D(n9112), .CK(clk), .Q(\x_mult_f[14][2] ) );
  DFF_X1 \x_mult_f_reg[14][3]  ( .D(n9111), .CK(clk), .Q(\x_mult_f[14][3] ) );
  DFF_X1 \x_mult_f_reg[14][4]  ( .D(n9110), .CK(clk), .Q(\x_mult_f[14][4] ) );
  DFF_X1 \x_mult_f_reg[14][5]  ( .D(n9109), .CK(clk), .Q(\x_mult_f[14][5] ) );
  DFF_X1 \x_mult_f_reg[14][6]  ( .D(n9108), .CK(clk), .Q(\x_mult_f[14][6] ) );
  DFF_X1 \x_mult_f_reg[14][7]  ( .D(n9107), .CK(clk), .Q(\x_mult_f[14][7] ) );
  DFF_X1 \x_mult_f_reg[14][8]  ( .D(n9106), .CK(clk), .Q(\x_mult_f[14][8] ) );
  DFF_X1 \x_mult_f_reg[14][9]  ( .D(n9105), .CK(clk), .Q(\x_mult_f[14][9] ) );
  DFF_X1 \x_mult_f_reg[14][10]  ( .D(n9104), .CK(clk), .Q(\x_mult_f[14][10] )
         );
  DFF_X1 \x_mult_f_reg[14][11]  ( .D(n9103), .CK(clk), .Q(\x_mult_f[14][11] )
         );
  DFF_X1 \x_mult_f_reg[14][12]  ( .D(n9102), .CK(clk), .Q(\x_mult_f[14][12] )
         );
  DFF_X1 \x_mult_f_reg[14][13]  ( .D(n9101), .CK(clk), .Q(\x_mult_f[14][13] )
         );
  DFF_X1 \x_mult_f_reg[14][14]  ( .D(n9100), .CK(clk), .Q(\x_mult_f[14][14] )
         );
  DFF_X1 \x_mult_f_reg[14][15]  ( .D(n9099), .CK(clk), .Q(\x_mult_f[14][15] ), 
        .QN(n3453) );
  DFF_X1 \x_mult_f_reg[15][1]  ( .D(n9322), .CK(clk), .Q(\x_mult_f[15][1] ) );
  DFF_X1 \x_mult_f_reg[15][2]  ( .D(n9126), .CK(clk), .Q(\x_mult_f[15][2] ) );
  DFF_X1 \x_mult_f_reg[15][3]  ( .D(n9125), .CK(clk), .Q(\x_mult_f[15][3] ) );
  DFF_X1 \x_mult_f_reg[15][4]  ( .D(n9124), .CK(clk), .Q(\x_mult_f[15][4] ) );
  DFF_X1 \x_mult_f_reg[15][5]  ( .D(n9123), .CK(clk), .Q(\x_mult_f[15][5] ) );
  DFF_X1 \x_mult_f_reg[15][6]  ( .D(n9122), .CK(clk), .Q(\x_mult_f[15][6] ) );
  DFF_X1 \x_mult_f_reg[15][7]  ( .D(n9121), .CK(clk), .Q(\x_mult_f[15][7] ) );
  DFF_X1 \x_mult_f_reg[15][8]  ( .D(n9120), .CK(clk), .Q(\x_mult_f[15][8] ) );
  DFF_X1 \x_mult_f_reg[15][9]  ( .D(n9119), .CK(clk), .Q(\x_mult_f[15][9] ) );
  DFF_X1 \x_mult_f_reg[15][10]  ( .D(n9118), .CK(clk), .Q(\x_mult_f[15][10] )
         );
  DFF_X1 \x_mult_f_reg[15][11]  ( .D(n9117), .CK(clk), .Q(\x_mult_f[15][11] )
         );
  DFF_X1 \x_mult_f_reg[15][12]  ( .D(n9116), .CK(clk), .Q(\x_mult_f[15][12] )
         );
  DFF_X1 \x_mult_f_reg[15][13]  ( .D(n9115), .CK(clk), .Q(\x_mult_f[15][13] )
         );
  DFF_X1 \x_mult_f_reg[15][14]  ( .D(n9114), .CK(clk), .Q(\x_mult_f[15][14] )
         );
  DFF_X1 \x_mult_f_reg[15][15]  ( .D(n9113), .CK(clk), .Q(\x_mult_f[15][15] ), 
        .QN(n3483) );
  DFF_X1 \x_mult_f_reg[16][0]  ( .D(n9325), .CK(clk), .Q(\x_mult_f[16][0] ) );
  DFF_X1 \x_mult_f_reg[16][1]  ( .D(n9324), .CK(clk), .Q(\x_mult_f[16][1] ) );
  DFF_X1 \x_mult_f_reg[16][2]  ( .D(n9139), .CK(clk), .Q(\x_mult_f[16][2] ) );
  DFF_X1 \x_mult_f_reg[16][4]  ( .D(n9138), .CK(clk), .Q(\x_mult_f[16][4] ) );
  DFF_X1 \x_mult_f_reg[16][5]  ( .D(n9137), .CK(clk), .Q(\x_mult_f[16][5] ) );
  DFF_X1 \x_mult_f_reg[16][6]  ( .D(n9136), .CK(clk), .Q(\x_mult_f[16][6] ) );
  DFF_X1 \x_mult_f_reg[16][7]  ( .D(n9135), .CK(clk), .Q(\x_mult_f[16][7] ) );
  DFF_X1 \x_mult_f_reg[16][8]  ( .D(n9134), .CK(clk), .Q(\x_mult_f[16][8] ) );
  DFF_X1 \x_mult_f_reg[16][9]  ( .D(n9133), .CK(clk), .Q(\x_mult_f[16][9] ) );
  DFF_X1 \x_mult_f_reg[16][10]  ( .D(n9132), .CK(clk), .Q(\x_mult_f[16][10] )
         );
  DFF_X1 \x_mult_f_reg[16][11]  ( .D(n9131), .CK(clk), .Q(\x_mult_f[16][11] )
         );
  DFF_X1 \x_mult_f_reg[16][12]  ( .D(n9130), .CK(clk), .Q(\x_mult_f[16][12] )
         );
  DFF_X1 \x_mult_f_reg[16][13]  ( .D(n9129), .CK(clk), .Q(\x_mult_f[16][13] )
         );
  DFF_X1 \x_mult_f_reg[16][14]  ( .D(n9128), .CK(clk), .Q(\x_mult_f[16][14] )
         );
  DFF_X1 \x_mult_f_reg[16][15]  ( .D(n9127), .CK(clk), .Q(\x_mult_f[16][15] ), 
        .QN(n3460) );
  DFF_X1 \x_mult_f_reg[17][0]  ( .D(n9327), .CK(clk), .Q(\x_mult_f[17][0] ) );
  DFF_X1 \x_mult_f_reg[17][1]  ( .D(n9326), .CK(clk), .Q(\x_mult_f[17][1] ) );
  DFF_X1 \x_mult_f_reg[17][2]  ( .D(n9153), .CK(clk), .Q(\x_mult_f[17][2] ) );
  DFF_X1 \x_mult_f_reg[17][3]  ( .D(n9152), .CK(clk), .Q(\x_mult_f[17][3] ) );
  DFF_X1 \x_mult_f_reg[17][4]  ( .D(n9151), .CK(clk), .Q(\x_mult_f[17][4] ) );
  DFF_X1 \x_mult_f_reg[17][5]  ( .D(n9150), .CK(clk), .Q(\x_mult_f[17][5] ) );
  DFF_X1 \x_mult_f_reg[17][6]  ( .D(n9149), .CK(clk), .Q(\x_mult_f[17][6] ) );
  DFF_X1 \x_mult_f_reg[17][7]  ( .D(n9148), .CK(clk), .Q(\x_mult_f[17][7] ) );
  DFF_X1 \x_mult_f_reg[17][8]  ( .D(n9147), .CK(clk), .Q(\x_mult_f[17][8] ) );
  DFF_X1 \x_mult_f_reg[17][9]  ( .D(n9146), .CK(clk), .Q(\x_mult_f[17][9] ) );
  DFF_X1 \x_mult_f_reg[17][10]  ( .D(n9145), .CK(clk), .Q(\x_mult_f[17][10] )
         );
  DFF_X1 \x_mult_f_reg[17][11]  ( .D(n9144), .CK(clk), .Q(\x_mult_f[17][11] )
         );
  DFF_X1 \x_mult_f_reg[17][12]  ( .D(n9143), .CK(clk), .Q(\x_mult_f[17][12] )
         );
  DFF_X1 \x_mult_f_reg[17][13]  ( .D(n9142), .CK(clk), .Q(\x_mult_f[17][13] )
         );
  DFF_X1 \x_mult_f_reg[17][14]  ( .D(n9141), .CK(clk), .Q(\x_mult_f[17][14] )
         );
  DFF_X1 \x_mult_f_reg[17][15]  ( .D(n9140), .CK(clk), .Q(\x_mult_f[17][15] ), 
        .QN(n3490) );
  DFF_X1 \x_mult_f_reg[18][0]  ( .D(n9329), .CK(clk), .Q(\x_mult_f[18][0] ) );
  DFF_X1 \x_mult_f_reg[18][1]  ( .D(n9328), .CK(clk), .Q(\x_mult_f[18][1] ) );
  DFF_X1 \x_mult_f_reg[18][2]  ( .D(n9167), .CK(clk), .Q(\x_mult_f[18][2] ) );
  DFF_X1 \x_mult_f_reg[18][3]  ( .D(n9166), .CK(clk), .Q(\x_mult_f[18][3] ) );
  DFF_X1 \x_mult_f_reg[18][4]  ( .D(n9165), .CK(clk), .Q(\x_mult_f[18][4] ) );
  DFF_X1 \x_mult_f_reg[18][5]  ( .D(n9164), .CK(clk), .Q(\x_mult_f[18][5] ) );
  DFF_X1 \x_mult_f_reg[18][6]  ( .D(n9163), .CK(clk), .Q(\x_mult_f[18][6] ) );
  DFF_X1 \x_mult_f_reg[18][7]  ( .D(n9162), .CK(clk), .Q(\x_mult_f[18][7] ) );
  DFF_X1 \x_mult_f_reg[18][8]  ( .D(n9161), .CK(clk), .Q(\x_mult_f[18][8] ) );
  DFF_X1 \x_mult_f_reg[18][9]  ( .D(n9160), .CK(clk), .Q(\x_mult_f[18][9] ) );
  DFF_X1 \x_mult_f_reg[18][10]  ( .D(n9159), .CK(clk), .Q(\x_mult_f[18][10] )
         );
  DFF_X1 \x_mult_f_reg[18][11]  ( .D(n9158), .CK(clk), .Q(\x_mult_f[18][11] )
         );
  DFF_X1 \x_mult_f_reg[18][12]  ( .D(n9157), .CK(clk), .Q(\x_mult_f[18][12] )
         );
  DFF_X1 \x_mult_f_reg[18][13]  ( .D(n9156), .CK(clk), .Q(\x_mult_f[18][13] )
         );
  DFF_X1 \x_mult_f_reg[18][14]  ( .D(n9155), .CK(clk), .Q(\x_mult_f[18][14] )
         );
  DFF_X1 \x_mult_f_reg[18][15]  ( .D(n9154), .CK(clk), .Q(\x_mult_f[18][15] ), 
        .QN(n3456) );
  DFF_X1 \x_mult_f_reg[19][0]  ( .D(n9331), .CK(clk), .Q(\x_mult_f[19][0] ) );
  DFF_X1 \x_mult_f_reg[19][1]  ( .D(n9330), .CK(clk), .Q(\x_mult_f[19][1] ) );
  DFF_X1 \x_mult_f_reg[19][2]  ( .D(n9181), .CK(clk), .Q(\x_mult_f[19][2] ) );
  DFF_X1 \x_mult_f_reg[19][3]  ( .D(n9180), .CK(clk), .Q(\x_mult_f[19][3] ) );
  DFF_X1 \x_mult_f_reg[19][4]  ( .D(n9179), .CK(clk), .Q(\x_mult_f[19][4] ) );
  DFF_X1 \x_mult_f_reg[19][6]  ( .D(n9177), .CK(clk), .Q(\x_mult_f[19][6] ) );
  DFF_X1 \x_mult_f_reg[19][7]  ( .D(n9176), .CK(clk), .Q(\x_mult_f[19][7] ) );
  DFF_X1 \x_mult_f_reg[19][8]  ( .D(n9175), .CK(clk), .Q(\x_mult_f[19][8] ) );
  DFF_X1 \x_mult_f_reg[19][9]  ( .D(n9174), .CK(clk), .Q(\x_mult_f[19][9] ) );
  DFF_X1 \x_mult_f_reg[19][10]  ( .D(n9173), .CK(clk), .Q(\x_mult_f[19][10] )
         );
  DFF_X1 \x_mult_f_reg[19][11]  ( .D(n9172), .CK(clk), .Q(\x_mult_f[19][11] )
         );
  DFF_X1 \x_mult_f_reg[19][12]  ( .D(n9171), .CK(clk), .Q(\x_mult_f[19][12] )
         );
  DFF_X1 \x_mult_f_reg[19][13]  ( .D(n9170), .CK(clk), .Q(\x_mult_f[19][13] )
         );
  DFF_X1 \x_mult_f_reg[19][14]  ( .D(n9169), .CK(clk), .Q(\x_mult_f[19][14] )
         );
  DFF_X1 \x_mult_f_reg[19][15]  ( .D(n9168), .CK(clk), .Q(\x_mult_f[19][15] ), 
        .QN(n3486) );
  DFF_X1 \x_mult_f_reg[20][0]  ( .D(n9333), .CK(clk), .Q(\x_mult_f[20][0] ) );
  DFF_X1 \x_mult_f_reg[20][1]  ( .D(n9332), .CK(clk), .Q(\x_mult_f[20][1] ) );
  DFF_X1 \x_mult_f_reg[20][2]  ( .D(n9187), .CK(clk), .Q(\x_mult_f[20][2] ) );
  DFF_X1 \x_mult_f_reg[20][3]  ( .D(n9186), .CK(clk), .Q(\x_mult_f[20][3] ) );
  DFF_X1 \x_mult_f_reg[20][4]  ( .D(n9185), .CK(clk), .Q(\x_mult_f[20][4] ) );
  DFF_X1 \x_mult_f_reg[20][5]  ( .D(n9184), .CK(clk), .Q(\x_mult_f[20][5] ) );
  DFF_X1 \x_mult_f_reg[20][6]  ( .D(n9183), .CK(clk), .Q(\x_mult_f[20][6] ) );
  DFF_X1 \x_mult_f_reg[20][7]  ( .D(n9182), .CK(clk), .Q(\x_mult_f[20][7] ) );
  DFF_X1 \x_mult_f_reg[21][0]  ( .D(n9335), .CK(clk), .Q(\x_mult_f[21][0] ) );
  DFF_X1 \x_mult_f_reg[21][1]  ( .D(n9334), .CK(clk), .Q(\x_mult_f[21][1] ) );
  DFF_X1 \x_mult_f_reg[21][2]  ( .D(n9195), .CK(clk), .Q(\x_mult_f[21][2] ) );
  DFF_X1 \x_mult_f_reg[21][3]  ( .D(n9194), .CK(clk), .Q(\x_mult_f[21][3] ) );
  DFF_X1 \x_mult_f_reg[21][4]  ( .D(n9193), .CK(clk), .Q(\x_mult_f[21][4] ) );
  DFF_X1 \x_mult_f_reg[21][11]  ( .D(n9192), .CK(clk), .Q(\x_mult_f[21][11] )
         );
  DFF_X1 \x_mult_f_reg[21][12]  ( .D(n9191), .CK(clk), .Q(\x_mult_f[21][12] )
         );
  DFF_X1 \x_mult_f_reg[21][13]  ( .D(n9190), .CK(clk), .Q(\x_mult_f[21][13] )
         );
  DFF_X1 \x_mult_f_reg[21][14]  ( .D(n9189), .CK(clk), .Q(\x_mult_f[21][14] )
         );
  DFF_X1 \x_mult_f_reg[21][15]  ( .D(n9188), .CK(clk), .Q(\x_mult_f[21][15] ), 
        .QN(n3498) );
  DFF_X1 \x_mult_f_reg[22][1]  ( .D(n9336), .CK(clk), .Q(\x_mult_f[22][1] ) );
  DFF_X1 \x_mult_f_reg[22][2]  ( .D(n9204), .CK(clk), .Q(\x_mult_f[22][2] ) );
  DFF_X1 \x_mult_f_reg[22][3]  ( .D(n9203), .CK(clk), .Q(\x_mult_f[22][3] ) );
  DFF_X1 \x_mult_f_reg[22][4]  ( .D(n9202), .CK(clk), .Q(\x_mult_f[22][4] ) );
  DFF_X1 \x_mult_f_reg[22][5]  ( .D(n9201), .CK(clk), .Q(\x_mult_f[22][5] ) );
  DFF_X1 \x_mult_f_reg[22][7]  ( .D(n9200), .CK(clk), .Q(\x_mult_f[22][7] ) );
  DFF_X1 \x_mult_f_reg[22][8]  ( .D(n9199), .CK(clk), .Q(\x_mult_f[22][8] ) );
  DFF_X1 \x_mult_f_reg[22][9]  ( .D(n9198), .CK(clk), .Q(\x_mult_f[22][9] ) );
  DFF_X1 \x_mult_f_reg[22][10]  ( .D(n9197), .CK(clk), .Q(\x_mult_f[22][10] )
         );
  DFF_X1 \x_mult_f_reg[22][11]  ( .D(n9196), .CK(clk), .Q(\x_mult_f[22][11] )
         );
  DFF_X1 \x_mult_f_reg[23][0]  ( .D(n9339), .CK(clk), .Q(\x_mult_f[23][0] ) );
  DFF_X1 \x_mult_f_reg[23][1]  ( .D(n9338), .CK(clk), .Q(\x_mult_f[23][1] ) );
  DFF_X1 \x_mult_f_reg[23][2]  ( .D(n9215), .CK(clk), .Q(\x_mult_f[23][2] ) );
  DFF_X1 \x_mult_f_reg[23][3]  ( .D(n9214), .CK(clk), .Q(\x_mult_f[23][3] ) );
  DFF_X1 \x_mult_f_reg[23][4]  ( .D(n9213), .CK(clk), .Q(\x_mult_f[23][4] ) );
  DFF_X1 \x_mult_f_reg[23][5]  ( .D(n9212), .CK(clk), .Q(\x_mult_f[23][5] ) );
  DFF_X1 \x_mult_f_reg[23][6]  ( .D(n9211), .CK(clk), .Q(\x_mult_f[23][6] ) );
  DFF_X1 \x_mult_f_reg[23][7]  ( .D(n9210), .CK(clk), .Q(\x_mult_f[23][7] ) );
  DFF_X1 \x_mult_f_reg[23][8]  ( .D(n9209), .CK(clk), .Q(\x_mult_f[23][8] ) );
  DFF_X1 \x_mult_f_reg[23][9]  ( .D(n9208), .CK(clk), .Q(\x_mult_f[23][9] ) );
  DFF_X1 \x_mult_f_reg[23][10]  ( .D(n9207), .CK(clk), .Q(\x_mult_f[23][10] )
         );
  DFF_X1 \x_mult_f_reg[23][11]  ( .D(n9206), .CK(clk), .Q(\x_mult_f[23][11] )
         );
  DFF_X1 \x_mult_f_reg[23][12]  ( .D(n9205), .CK(clk), .Q(\x_mult_f[23][12] )
         );
  DFF_X1 \x_mult_f_reg[24][0]  ( .D(n9341), .CK(clk), .Q(\x_mult_f[24][0] ) );
  DFF_X1 \x_mult_f_reg[24][1]  ( .D(n9340), .CK(clk), .Q(\x_mult_f[24][1] ) );
  DFF_X1 \x_mult_f_reg[24][2]  ( .D(n9226), .CK(clk), .Q(\x_mult_f[24][2] ) );
  DFF_X1 \x_mult_f_reg[24][3]  ( .D(n9225), .CK(clk), .Q(\x_mult_f[24][3] ) );
  DFF_X1 \x_mult_f_reg[24][4]  ( .D(n9224), .CK(clk), .Q(\x_mult_f[24][4] ) );
  DFF_X1 \x_mult_f_reg[24][6]  ( .D(n9223), .CK(clk), .Q(\x_mult_f[24][6] ) );
  DFF_X1 \x_mult_f_reg[24][8]  ( .D(n9222), .CK(clk), .Q(\x_mult_f[24][8] ) );
  DFF_X1 \x_mult_f_reg[24][9]  ( .D(n9221), .CK(clk), .Q(\x_mult_f[24][9] ) );
  DFF_X1 \x_mult_f_reg[24][10]  ( .D(n9220), .CK(clk), .Q(\x_mult_f[24][10] )
         );
  DFF_X1 \x_mult_f_reg[24][11]  ( .D(n9219), .CK(clk), .Q(\x_mult_f[24][11] )
         );
  DFF_X1 \x_mult_f_reg[24][13]  ( .D(n9218), .CK(clk), .Q(\x_mult_f[24][13] )
         );
  DFF_X1 \x_mult_f_reg[24][14]  ( .D(n9217), .CK(clk), .Q(\x_mult_f[24][14] )
         );
  DFF_X1 \x_mult_f_reg[24][15]  ( .D(n9216), .CK(clk), .Q(\x_mult_f[24][15] ), 
        .QN(n3480) );
  DFF_X1 \x_mult_f_reg[25][0]  ( .D(n9343), .CK(clk), .Q(\x_mult_f[25][0] ) );
  DFF_X1 \x_mult_f_reg[25][1]  ( .D(n9342), .CK(clk), .Q(\x_mult_f[25][1] ) );
  DFF_X1 \x_mult_f_reg[25][2]  ( .D(n9229), .CK(clk), .Q(\x_mult_f[25][2] ) );
  DFF_X1 \x_mult_f_reg[25][3]  ( .D(n9228), .CK(clk), .Q(\x_mult_f[25][3] ) );
  DFF_X1 \x_mult_f_reg[25][4]  ( .D(n9227), .CK(clk), .Q(\x_mult_f[25][4] ) );
  DFF_X1 \x_mult_f_reg[26][0]  ( .D(n9345), .CK(clk), .Q(\x_mult_f[26][0] ) );
  DFF_X1 \x_mult_f_reg[26][1]  ( .D(n9344), .CK(clk), .Q(\x_mult_f[26][1] ) );
  DFF_X1 \x_mult_f_reg[26][2]  ( .D(n9233), .CK(clk), .Q(\x_mult_f[26][2] ) );
  DFF_X1 \x_mult_f_reg[26][3]  ( .D(n9232), .CK(clk), .Q(\x_mult_f[26][3] ) );
  DFF_X1 \x_mult_f_reg[26][4]  ( .D(n9231), .CK(clk), .Q(\x_mult_f[26][4] ) );
  DFF_X1 \x_mult_f_reg[26][7]  ( .D(n9230), .CK(clk), .Q(\x_mult_f[26][7] ) );
  DFF_X1 \x_mult_f_reg[27][0]  ( .D(n9347), .CK(clk), .Q(\x_mult_f[27][0] ) );
  DFF_X1 \x_mult_f_reg[27][1]  ( .D(n9346), .CK(clk), .Q(\x_mult_f[27][1] ) );
  DFF_X1 \x_mult_f_reg[27][2]  ( .D(n9246), .CK(clk), .Q(\x_mult_f[27][2] ) );
  DFF_X1 \x_mult_f_reg[27][3]  ( .D(n9245), .CK(clk), .Q(\x_mult_f[27][3] ) );
  DFF_X1 \x_mult_f_reg[27][4]  ( .D(n9244), .CK(clk), .Q(\x_mult_f[27][4] ) );
  DFF_X1 \x_mult_f_reg[27][5]  ( .D(n9243), .CK(clk), .Q(\x_mult_f[27][5] ) );
  DFF_X1 \x_mult_f_reg[27][6]  ( .D(n9242), .CK(clk), .Q(\x_mult_f[27][6] ) );
  DFF_X1 \x_mult_f_reg[27][7]  ( .D(n9241), .CK(clk), .Q(\x_mult_f[27][7] ) );
  DFF_X1 \x_mult_f_reg[27][9]  ( .D(n9240), .CK(clk), .Q(\x_mult_f[27][9] ) );
  DFF_X1 \x_mult_f_reg[27][10]  ( .D(n9239), .CK(clk), .Q(\x_mult_f[27][10] )
         );
  DFF_X1 \x_mult_f_reg[27][11]  ( .D(n9238), .CK(clk), .Q(\x_mult_f[27][11] )
         );
  DFF_X1 \x_mult_f_reg[27][12]  ( .D(n9237), .CK(clk), .Q(\x_mult_f[27][12] )
         );
  DFF_X1 \x_mult_f_reg[27][13]  ( .D(n9236), .CK(clk), .Q(\x_mult_f[27][13] )
         );
  DFF_X1 \x_mult_f_reg[27][14]  ( .D(n9235), .CK(clk), .Q(\x_mult_f[27][14] )
         );
  DFF_X1 \x_mult_f_reg[27][15]  ( .D(n9234), .CK(clk), .Q(\x_mult_f[27][15] ), 
        .QN(n3482) );
  DFF_X1 \x_mult_f_reg[28][0]  ( .D(n9349), .CK(clk), .Q(\x_mult_f[28][0] ) );
  DFF_X1 \x_mult_f_reg[28][1]  ( .D(n9348), .CK(clk), .Q(\x_mult_f[28][1] ) );
  DFF_X1 \x_mult_f_reg[28][2]  ( .D(n9252), .CK(clk), .Q(\x_mult_f[28][2] ) );
  DFF_X1 \x_mult_f_reg[28][3]  ( .D(n9251), .CK(clk), .Q(\x_mult_f[28][3] ) );
  DFF_X1 \x_mult_f_reg[28][4]  ( .D(n9250), .CK(clk), .Q(\x_mult_f[28][4] ) );
  DFF_X1 \x_mult_f_reg[28][5]  ( .D(n9249), .CK(clk), .Q(\x_mult_f[28][5] ) );
  DFF_X1 \x_mult_f_reg[28][14]  ( .D(n9248), .CK(clk), .Q(\x_mult_f[28][14] )
         );
  DFF_X1 \x_mult_f_reg[28][15]  ( .D(n9247), .CK(clk), .Q(\x_mult_f[28][15] ), 
        .QN(n3477) );
  DFF_X1 \x_mult_f_reg[29][0]  ( .D(n9351), .CK(clk), .Q(\x_mult_f[29][0] ) );
  DFF_X1 \x_mult_f_reg[29][1]  ( .D(n9350), .CK(clk), .Q(\x_mult_f[29][1] ) );
  DFF_X1 \x_mult_f_reg[29][2]  ( .D(n9263), .CK(clk), .Q(\x_mult_f[29][2] ) );
  DFF_X1 \x_mult_f_reg[29][3]  ( .D(n9262), .CK(clk), .Q(\x_mult_f[29][3] ) );
  DFF_X1 \x_mult_f_reg[29][4]  ( .D(n9261), .CK(clk), .Q(\x_mult_f[29][4] ) );
  DFF_X1 \x_mult_f_reg[29][5]  ( .D(n9260), .CK(clk), .Q(\x_mult_f[29][5] ) );
  DFF_X1 \x_mult_f_reg[29][6]  ( .D(n9259), .CK(clk), .Q(\x_mult_f[29][6] ) );
  DFF_X1 \x_mult_f_reg[29][8]  ( .D(n9257), .CK(clk), .Q(\x_mult_f[29][8] ) );
  DFF_X1 \x_mult_f_reg[29][9]  ( .D(n9256), .CK(clk), .Q(\x_mult_f[29][9] ) );
  DFF_X1 \x_mult_f_reg[29][10]  ( .D(n9255), .CK(clk), .Q(\x_mult_f[29][10] )
         );
  DFF_X1 \x_mult_f_reg[29][11]  ( .D(n9254), .CK(clk), .Q(\x_mult_f[29][11] )
         );
  DFF_X1 \x_mult_f_reg[29][12]  ( .D(n9253), .CK(clk), .Q(\x_mult_f[29][12] )
         );
  DFF_X1 \x_mult_f_reg[30][0]  ( .D(n9353), .CK(clk), .Q(\x_mult_f[30][0] ) );
  DFF_X1 \x_mult_f_reg[30][1]  ( .D(n9352), .CK(clk), .Q(\x_mult_f[30][1] ) );
  DFF_X1 \x_mult_f_reg[30][2]  ( .D(n9277), .CK(clk), .Q(\x_mult_f[30][2] ) );
  DFF_X1 \x_mult_f_reg[30][3]  ( .D(n9276), .CK(clk), .Q(\x_mult_f[30][3] ) );
  DFF_X1 \x_mult_f_reg[30][4]  ( .D(n9275), .CK(clk), .Q(\x_mult_f[30][4] ) );
  DFF_X1 \x_mult_f_reg[30][5]  ( .D(n9274), .CK(clk), .Q(\x_mult_f[30][5] ) );
  DFF_X1 \x_mult_f_reg[30][6]  ( .D(n9273), .CK(clk), .Q(\x_mult_f[30][6] ) );
  DFF_X1 \x_mult_f_reg[30][7]  ( .D(n9272), .CK(clk), .Q(\x_mult_f[30][7] ) );
  DFF_X1 \x_mult_f_reg[30][8]  ( .D(n9271), .CK(clk), .Q(\x_mult_f[30][8] ) );
  DFF_X1 \x_mult_f_reg[30][9]  ( .D(n9270), .CK(clk), .Q(\x_mult_f[30][9] ) );
  DFF_X1 \x_mult_f_reg[30][10]  ( .D(n9269), .CK(clk), .Q(\x_mult_f[30][10] )
         );
  DFF_X1 \x_mult_f_reg[30][11]  ( .D(n9268), .CK(clk), .Q(\x_mult_f[30][11] )
         );
  DFF_X1 \x_mult_f_reg[30][12]  ( .D(n9267), .CK(clk), .Q(\x_mult_f[30][12] )
         );
  DFF_X1 \x_mult_f_reg[30][13]  ( .D(n9266), .CK(clk), .Q(\x_mult_f[30][13] )
         );
  DFF_X1 \x_mult_f_reg[30][14]  ( .D(n9265), .CK(clk), .Q(\x_mult_f[30][14] )
         );
  DFF_X1 \x_mult_f_reg[30][15]  ( .D(n9264), .CK(clk), .Q(\x_mult_f[30][15] ), 
        .QN(n3458) );
  DFF_X1 \x_mult_f_reg[31][1]  ( .D(n9354), .CK(clk), .Q(\x_mult_f[31][1] ) );
  DFF_X1 \x_mult_f_reg[31][2]  ( .D(n9291), .CK(clk), .Q(\x_mult_f[31][2] ) );
  DFF_X1 \x_mult_f_reg[31][3]  ( .D(n9290), .CK(clk), .Q(\x_mult_f[31][3] ) );
  DFF_X1 \x_mult_f_reg[31][4]  ( .D(n9289), .CK(clk), .Q(\x_mult_f[31][4] ) );
  DFF_X1 \x_mult_f_reg[31][5]  ( .D(n9288), .CK(clk), .Q(\x_mult_f[31][5] ) );
  DFF_X1 \x_mult_f_reg[31][6]  ( .D(n9287), .CK(clk), .Q(\x_mult_f[31][6] ) );
  DFF_X1 \x_mult_f_reg[31][7]  ( .D(n9286), .CK(clk), .Q(\x_mult_f[31][7] ) );
  DFF_X1 \x_mult_f_reg[31][8]  ( .D(n9285), .CK(clk), .Q(\x_mult_f[31][8] ) );
  DFF_X1 \x_mult_f_reg[31][9]  ( .D(n9284), .CK(clk), .Q(\x_mult_f[31][9] ) );
  DFF_X1 \x_mult_f_reg[31][10]  ( .D(n9283), .CK(clk), .Q(\x_mult_f[31][10] )
         );
  DFF_X1 \x_mult_f_reg[31][11]  ( .D(n9282), .CK(clk), .Q(\x_mult_f[31][11] )
         );
  DFF_X1 \x_mult_f_reg[31][12]  ( .D(n9281), .CK(clk), .Q(\x_mult_f[31][12] )
         );
  DFF_X1 \x_mult_f_reg[31][13]  ( .D(n9280), .CK(clk), .Q(\x_mult_f[31][13] )
         );
  DFF_X1 \x_mult_f_reg[31][14]  ( .D(n9279), .CK(clk), .Q(\x_mult_f[31][14] )
         );
  DFF_X1 \x_mult_f_reg[31][15]  ( .D(n9278), .CK(clk), .Q(\x_mult_f[31][15] ), 
        .QN(n3488) );
  DFF_X1 \adder_stage1_reg[0][0]  ( .D(n10069), .CK(clk), .Q(
        \adder_stage1[0][0] ) );
  DFF_X1 \adder_stage1_reg[0][1]  ( .D(n10068), .CK(clk), .Q(
        \adder_stage1[0][1] ) );
  DFF_X1 \adder_stage1_reg[0][3]  ( .D(n10067), .CK(clk), .Q(
        \adder_stage1[0][3] ) );
  DFF_X1 \adder_stage1_reg[0][4]  ( .D(n10066), .CK(clk), .Q(
        \adder_stage1[0][4] ) );
  DFF_X1 \adder_stage1_reg[0][5]  ( .D(n10065), .CK(clk), .Q(
        \adder_stage1[0][5] ) );
  DFF_X1 \adder_stage1_reg[0][6]  ( .D(n10064), .CK(clk), .Q(
        \adder_stage1[0][6] ) );
  DFF_X1 \adder_stage1_reg[0][7]  ( .D(n10063), .CK(clk), .Q(
        \adder_stage1[0][7] ) );
  DFF_X1 \adder_stage1_reg[0][8]  ( .D(n10062), .CK(clk), .Q(
        \adder_stage1[0][8] ) );
  DFF_X1 \adder_stage1_reg[0][9]  ( .D(n10061), .CK(clk), .Q(
        \adder_stage1[0][9] ) );
  DFF_X1 \adder_stage1_reg[0][10]  ( .D(n10060), .CK(clk), .Q(
        \adder_stage1[0][10] ) );
  DFF_X1 \adder_stage1_reg[0][11]  ( .D(n10059), .CK(clk), .Q(
        \adder_stage1[0][11] ) );
  DFF_X1 \adder_stage1_reg[0][12]  ( .D(n10058), .CK(clk), .Q(
        \adder_stage1[0][12] ) );
  DFF_X1 \adder_stage1_reg[0][13]  ( .D(n10057), .CK(clk), .Q(
        \adder_stage1[0][13] ) );
  DFF_X1 \adder_stage1_reg[0][14]  ( .D(n10056), .CK(clk), .Q(
        \adder_stage1[0][14] ) );
  DFF_X1 \adder_stage1_reg[0][15]  ( .D(n10055), .CK(clk), .Q(
        \adder_stage1[0][15] ) );
  DFF_X1 \adder_stage1_reg[0][20]  ( .D(n10054), .CK(clk), .Q(
        \adder_stage1[0][20] ), .QN(n3479) );
  DFF_X1 \adder_stage1_reg[1][0]  ( .D(n10053), .CK(clk), .Q(
        \adder_stage1[1][0] ) );
  DFF_X1 \adder_stage1_reg[1][1]  ( .D(n10052), .CK(clk), .Q(
        \adder_stage1[1][1] ) );
  DFF_X1 \adder_stage1_reg[1][2]  ( .D(n10051), .CK(clk), .Q(
        \adder_stage1[1][2] ) );
  DFF_X1 \adder_stage1_reg[1][3]  ( .D(n10050), .CK(clk), .Q(
        \adder_stage1[1][3] ) );
  DFF_X1 \adder_stage1_reg[1][4]  ( .D(n10049), .CK(clk), .Q(
        \adder_stage1[1][4] ) );
  DFF_X1 \adder_stage1_reg[1][5]  ( .D(n10048), .CK(clk), .Q(
        \adder_stage1[1][5] ) );
  DFF_X1 \adder_stage1_reg[1][6]  ( .D(n10047), .CK(clk), .Q(
        \adder_stage1[1][6] ) );
  DFF_X1 \adder_stage1_reg[1][7]  ( .D(n10046), .CK(clk), .Q(
        \adder_stage1[1][7] ) );
  DFF_X1 \adder_stage1_reg[1][8]  ( .D(n10045), .CK(clk), .Q(
        \adder_stage1[1][8] ) );
  DFF_X1 \adder_stage1_reg[1][9]  ( .D(n10044), .CK(clk), .Q(
        \adder_stage1[1][9] ) );
  DFF_X1 \adder_stage1_reg[1][10]  ( .D(n10043), .CK(clk), .Q(
        \adder_stage1[1][10] ) );
  DFF_X1 \adder_stage1_reg[1][11]  ( .D(n10042), .CK(clk), .Q(
        \adder_stage1[1][11] ) );
  DFF_X1 \adder_stage1_reg[1][12]  ( .D(n10041), .CK(clk), .Q(
        \adder_stage1[1][12] ) );
  DFF_X1 \adder_stage1_reg[1][13]  ( .D(n10040), .CK(clk), .Q(
        \adder_stage1[1][13] ) );
  DFF_X1 \adder_stage1_reg[1][14]  ( .D(n10039), .CK(clk), .Q(
        \adder_stage1[1][14] ) );
  DFF_X1 \adder_stage1_reg[1][15]  ( .D(n10038), .CK(clk), .Q(
        \adder_stage1[1][15] ) );
  DFF_X1 \adder_stage1_reg[1][20]  ( .D(n10037), .CK(clk), .Q(
        \adder_stage1[1][20] ), .QN(n8706) );
  DFF_X1 \adder_stage1_reg[2][0]  ( .D(n10036), .CK(clk), .Q(
        \adder_stage1[2][0] ) );
  DFF_X1 \adder_stage1_reg[2][1]  ( .D(n10035), .CK(clk), .Q(
        \adder_stage1[2][1] ) );
  DFF_X1 \adder_stage1_reg[2][2]  ( .D(n10034), .CK(clk), .Q(
        \adder_stage1[2][2] ) );
  DFF_X1 \adder_stage1_reg[2][3]  ( .D(n10033), .CK(clk), .Q(
        \adder_stage1[2][3] ) );
  DFF_X1 \adder_stage1_reg[2][4]  ( .D(n10032), .CK(clk), .Q(
        \adder_stage1[2][4] ) );
  DFF_X1 \adder_stage1_reg[2][5]  ( .D(n10031), .CK(clk), .Q(
        \adder_stage1[2][5] ) );
  DFF_X1 \adder_stage1_reg[2][6]  ( .D(n10030), .CK(clk), .Q(
        \adder_stage1[2][6] ) );
  DFF_X1 \adder_stage1_reg[2][7]  ( .D(n10029), .CK(clk), .Q(
        \adder_stage1[2][7] ), .QN(n3513) );
  DFF_X1 \adder_stage1_reg[2][8]  ( .D(n10028), .CK(clk), .Q(
        \adder_stage1[2][8] ) );
  DFF_X1 \adder_stage1_reg[2][9]  ( .D(n10027), .CK(clk), .Q(
        \adder_stage1[2][9] ) );
  DFF_X1 \adder_stage1_reg[2][10]  ( .D(n10026), .CK(clk), .Q(
        \adder_stage1[2][10] ) );
  DFF_X1 \adder_stage1_reg[2][11]  ( .D(n10025), .CK(clk), .Q(
        \adder_stage1[2][11] ) );
  DFF_X1 \adder_stage1_reg[2][12]  ( .D(n10024), .CK(clk), .Q(
        \adder_stage1[2][12] ) );
  DFF_X1 \adder_stage1_reg[2][13]  ( .D(n10023), .CK(clk), .Q(
        \adder_stage1[2][13] ) );
  DFF_X1 \adder_stage1_reg[2][15]  ( .D(n10022), .CK(clk), .Q(
        \adder_stage1[2][15] ) );
  DFF_X1 \adder_stage1_reg[2][20]  ( .D(n10021), .CK(clk), .Q(
        \adder_stage1[2][20] ), .QN(n3461) );
  DFF_X1 \adder_stage1_reg[3][0]  ( .D(n10020), .CK(clk), .Q(
        \adder_stage1[3][0] ) );
  DFF_X1 \adder_stage1_reg[3][1]  ( .D(n10019), .CK(clk), .Q(
        \adder_stage1[3][1] ) );
  DFF_X1 \adder_stage1_reg[3][2]  ( .D(n10018), .CK(clk), .Q(
        \adder_stage1[3][2] ) );
  DFF_X1 \adder_stage1_reg[3][3]  ( .D(n10017), .CK(clk), .Q(
        \adder_stage1[3][3] ) );
  DFF_X1 \adder_stage1_reg[3][4]  ( .D(n10016), .CK(clk), .Q(
        \adder_stage1[3][4] ) );
  DFF_X1 \adder_stage1_reg[3][5]  ( .D(n10015), .CK(clk), .Q(
        \adder_stage1[3][5] ) );
  DFF_X1 \adder_stage1_reg[3][6]  ( .D(n10014), .CK(clk), .Q(
        \adder_stage1[3][6] ) );
  DFF_X1 \adder_stage1_reg[3][7]  ( .D(n10013), .CK(clk), .Q(
        \adder_stage1[3][7] ), .QN(n3475) );
  DFF_X1 \adder_stage1_reg[3][8]  ( .D(n10012), .CK(clk), .Q(
        \adder_stage1[3][8] ) );
  DFF_X1 \adder_stage1_reg[3][9]  ( .D(n10011), .CK(clk), .Q(
        \adder_stage1[3][9] ) );
  DFF_X1 \adder_stage1_reg[3][10]  ( .D(n10010), .CK(clk), .Q(
        \adder_stage1[3][10] ) );
  DFF_X1 \adder_stage1_reg[3][11]  ( .D(n10009), .CK(clk), .Q(
        \adder_stage1[3][11] ) );
  DFF_X1 \adder_stage1_reg[3][12]  ( .D(n10008), .CK(clk), .Q(
        \adder_stage1[3][12] ) );
  DFF_X1 \adder_stage1_reg[3][13]  ( .D(n10007), .CK(clk), .Q(
        \adder_stage1[3][13] ) );
  DFF_X1 \adder_stage1_reg[3][14]  ( .D(n10006), .CK(clk), .Q(
        \adder_stage1[3][14] ) );
  DFF_X1 \adder_stage1_reg[3][15]  ( .D(n10005), .CK(clk), .Q(
        \adder_stage1[3][15] ) );
  DFF_X1 \adder_stage1_reg[3][20]  ( .D(n10004), .CK(clk), .Q(
        \adder_stage1[3][20] ), .QN(n3492) );
  DFF_X1 \adder_stage1_reg[4][0]  ( .D(n10003), .CK(clk), .Q(
        \adder_stage1[4][0] ) );
  DFF_X1 \adder_stage1_reg[4][1]  ( .D(n10002), .CK(clk), .Q(
        \adder_stage1[4][1] ) );
  DFF_X1 \adder_stage1_reg[4][2]  ( .D(n10001), .CK(clk), .Q(
        \adder_stage1[4][2] ) );
  DFF_X1 \adder_stage1_reg[4][3]  ( .D(n10000), .CK(clk), .Q(
        \adder_stage1[4][3] ) );
  DFF_X1 \adder_stage1_reg[4][4]  ( .D(n9999), .CK(clk), .Q(
        \adder_stage1[4][4] ) );
  DFF_X1 \adder_stage1_reg[4][5]  ( .D(n9998), .CK(clk), .Q(
        \adder_stage1[4][5] ) );
  DFF_X1 \adder_stage1_reg[4][6]  ( .D(n9997), .CK(clk), .Q(
        \adder_stage1[4][6] ) );
  DFF_X1 \adder_stage1_reg[4][7]  ( .D(n9996), .CK(clk), .Q(
        \adder_stage1[4][7] ) );
  DFF_X1 \adder_stage1_reg[4][8]  ( .D(n9995), .CK(clk), .Q(
        \adder_stage1[4][8] ) );
  DFF_X1 \adder_stage1_reg[4][9]  ( .D(n9994), .CK(clk), .Q(
        \adder_stage1[4][9] ) );
  DFF_X1 \adder_stage1_reg[4][10]  ( .D(n9993), .CK(clk), .Q(
        \adder_stage1[4][10] ) );
  DFF_X1 \adder_stage1_reg[4][11]  ( .D(n9992), .CK(clk), .Q(
        \adder_stage1[4][11] ) );
  DFF_X1 \adder_stage1_reg[4][12]  ( .D(n9991), .CK(clk), .Q(
        \adder_stage1[4][12] ) );
  DFF_X1 \adder_stage1_reg[4][15]  ( .D(n9990), .CK(clk), .Q(
        \adder_stage1[4][15] ) );
  DFF_X1 \adder_stage1_reg[5][0]  ( .D(n9989), .CK(clk), .Q(
        \adder_stage1[5][0] ) );
  DFF_X1 \adder_stage1_reg[5][1]  ( .D(n9988), .CK(clk), .Q(
        \adder_stage1[5][1] ) );
  DFF_X1 \adder_stage1_reg[5][2]  ( .D(n9987), .CK(clk), .Q(
        \adder_stage1[5][2] ) );
  DFF_X1 \adder_stage1_reg[5][3]  ( .D(n9986), .CK(clk), .Q(
        \adder_stage1[5][3] ) );
  DFF_X1 \adder_stage1_reg[5][4]  ( .D(n9985), .CK(clk), .Q(
        \adder_stage1[5][4] ) );
  DFF_X1 \adder_stage1_reg[5][5]  ( .D(n9984), .CK(clk), .Q(
        \adder_stage1[5][5] ) );
  DFF_X1 \adder_stage1_reg[5][6]  ( .D(n9983), .CK(clk), .Q(
        \adder_stage1[5][6] ) );
  DFF_X1 \adder_stage1_reg[5][7]  ( .D(n9982), .CK(clk), .Q(
        \adder_stage1[5][7] ) );
  DFF_X1 \adder_stage1_reg[5][8]  ( .D(n9981), .CK(clk), .Q(
        \adder_stage1[5][8] ) );
  DFF_X1 \adder_stage1_reg[5][9]  ( .D(n9980), .CK(clk), .Q(
        \adder_stage1[5][9] ) );
  DFF_X1 \adder_stage1_reg[5][10]  ( .D(n9979), .CK(clk), .Q(
        \adder_stage1[5][10] ) );
  DFF_X1 \adder_stage1_reg[5][11]  ( .D(n9978), .CK(clk), .Q(
        \adder_stage1[5][11] ) );
  DFF_X1 \adder_stage1_reg[5][12]  ( .D(n9977), .CK(clk), .Q(
        \adder_stage1[5][12] ) );
  DFF_X1 \adder_stage1_reg[5][13]  ( .D(n9976), .CK(clk), .Q(
        \adder_stage1[5][13] ) );
  DFF_X1 \adder_stage1_reg[5][14]  ( .D(n9975), .CK(clk), .Q(
        \adder_stage1[5][14] ) );
  DFF_X1 \adder_stage1_reg[5][15]  ( .D(n9974), .CK(clk), .Q(
        \adder_stage1[5][15] ) );
  DFF_X1 \adder_stage1_reg[5][20]  ( .D(n9973), .CK(clk), .Q(
        \adder_stage1[5][20] ), .QN(n3491) );
  DFF_X1 \adder_stage1_reg[6][0]  ( .D(n9972), .CK(clk), .Q(
        \adder_stage1[6][0] ) );
  DFF_X1 \adder_stage1_reg[6][1]  ( .D(n9971), .CK(clk), .Q(
        \adder_stage1[6][1] ) );
  DFF_X1 \adder_stage1_reg[6][2]  ( .D(n9970), .CK(clk), .Q(
        \adder_stage1[6][2] ) );
  DFF_X1 \adder_stage1_reg[6][3]  ( .D(n9969), .CK(clk), .Q(
        \adder_stage1[6][3] ) );
  DFF_X1 \adder_stage1_reg[6][4]  ( .D(n9968), .CK(clk), .Q(
        \adder_stage1[6][4] ) );
  DFF_X1 \adder_stage1_reg[6][5]  ( .D(n9967), .CK(clk), .Q(
        \adder_stage1[6][5] ) );
  DFF_X1 \adder_stage1_reg[6][6]  ( .D(n9966), .CK(clk), .Q(
        \adder_stage1[6][6] ) );
  DFF_X1 \adder_stage1_reg[6][7]  ( .D(n9965), .CK(clk), .Q(
        \adder_stage1[6][7] ) );
  DFF_X1 \adder_stage1_reg[6][8]  ( .D(n9964), .CK(clk), .Q(
        \adder_stage1[6][8] ) );
  DFF_X1 \adder_stage1_reg[6][9]  ( .D(n9963), .CK(clk), .Q(
        \adder_stage1[6][9] ), .QN(n3474) );
  DFF_X1 \adder_stage1_reg[6][10]  ( .D(n9962), .CK(clk), .Q(
        \adder_stage1[6][10] ) );
  DFF_X1 \adder_stage1_reg[6][11]  ( .D(n9961), .CK(clk), .Q(
        \adder_stage1[6][11] ) );
  DFF_X1 \adder_stage1_reg[6][12]  ( .D(n9960), .CK(clk), .Q(
        \adder_stage1[6][12] ) );
  DFF_X1 \adder_stage1_reg[6][13]  ( .D(n9959), .CK(clk), .Q(
        \adder_stage1[6][13] ) );
  DFF_X1 \adder_stage1_reg[6][14]  ( .D(n9958), .CK(clk), .Q(
        \adder_stage1[6][14] ) );
  DFF_X1 \adder_stage1_reg[6][15]  ( .D(n9957), .CK(clk), .Q(
        \adder_stage1[6][15] ) );
  DFF_X1 \adder_stage1_reg[6][20]  ( .D(n9956), .CK(clk), .Q(
        \adder_stage1[6][20] ), .QN(n3464) );
  DFF_X1 \adder_stage1_reg[7][0]  ( .D(n9955), .CK(clk), .Q(
        \adder_stage1[7][0] ) );
  DFF_X1 \adder_stage1_reg[7][1]  ( .D(n9954), .CK(clk), .Q(
        \adder_stage1[7][1] ) );
  DFF_X1 \adder_stage1_reg[7][2]  ( .D(n9953), .CK(clk), .Q(
        \adder_stage1[7][2] ) );
  DFF_X1 \adder_stage1_reg[7][3]  ( .D(n9952), .CK(clk), .Q(
        \adder_stage1[7][3] ) );
  DFF_X1 \adder_stage1_reg[7][4]  ( .D(n9951), .CK(clk), .Q(
        \adder_stage1[7][4] ) );
  DFF_X1 \adder_stage1_reg[7][5]  ( .D(n9950), .CK(clk), .Q(
        \adder_stage1[7][5] ) );
  DFF_X1 \adder_stage1_reg[7][6]  ( .D(n9949), .CK(clk), .Q(
        \adder_stage1[7][6] ) );
  DFF_X1 \adder_stage1_reg[7][8]  ( .D(n9947), .CK(clk), .Q(
        \adder_stage1[7][8] ) );
  DFF_X1 \adder_stage1_reg[7][9]  ( .D(n9946), .CK(clk), .Q(
        \adder_stage1[7][9] ), .QN(n3512) );
  DFF_X1 \adder_stage1_reg[7][10]  ( .D(n9945), .CK(clk), .Q(
        \adder_stage1[7][10] ) );
  DFF_X1 \adder_stage1_reg[7][11]  ( .D(n9944), .CK(clk), .Q(
        \adder_stage1[7][11] ) );
  DFF_X1 \adder_stage1_reg[7][12]  ( .D(n9943), .CK(clk), .Q(
        \adder_stage1[7][12] ) );
  DFF_X1 \adder_stage1_reg[7][13]  ( .D(n9942), .CK(clk), .Q(
        \adder_stage1[7][13] ) );
  DFF_X1 \adder_stage1_reg[7][14]  ( .D(n9941), .CK(clk), .Q(
        \adder_stage1[7][14] ) );
  DFF_X1 \adder_stage1_reg[7][15]  ( .D(n9940), .CK(clk), .Q(
        \adder_stage1[7][15] ) );
  DFF_X1 \adder_stage1_reg[7][20]  ( .D(n9939), .CK(clk), .Q(
        \adder_stage1[7][20] ), .QN(n3493) );
  DFF_X1 \adder_stage1_reg[8][0]  ( .D(n9938), .CK(clk), .Q(
        \adder_stage1[8][0] ) );
  DFF_X1 \adder_stage1_reg[8][1]  ( .D(n9937), .CK(clk), .Q(
        \adder_stage1[8][1] ) );
  DFF_X1 \adder_stage1_reg[8][2]  ( .D(n9936), .CK(clk), .Q(
        \adder_stage1[8][2] ) );
  DFF_X1 \adder_stage1_reg[8][3]  ( .D(n9935), .CK(clk), .Q(
        \adder_stage1[8][3] ) );
  DFF_X1 \adder_stage1_reg[8][4]  ( .D(n9934), .CK(clk), .Q(
        \adder_stage1[8][4] ) );
  DFF_X1 \adder_stage1_reg[8][5]  ( .D(n9933), .CK(clk), .Q(
        \adder_stage1[8][5] ) );
  DFF_X1 \adder_stage1_reg[8][6]  ( .D(n9932), .CK(clk), .Q(
        \adder_stage1[8][6] ) );
  DFF_X1 \adder_stage1_reg[8][7]  ( .D(n9931), .CK(clk), .Q(
        \adder_stage1[8][7] ) );
  DFF_X1 \adder_stage1_reg[8][8]  ( .D(n9930), .CK(clk), .Q(
        \adder_stage1[8][8] ) );
  DFF_X1 \adder_stage1_reg[8][9]  ( .D(n9929), .CK(clk), .Q(
        \adder_stage1[8][9] ) );
  DFF_X1 \adder_stage1_reg[8][10]  ( .D(n9928), .CK(clk), .Q(
        \adder_stage1[8][10] ) );
  DFF_X1 \adder_stage1_reg[8][11]  ( .D(n9927), .CK(clk), .Q(
        \adder_stage1[8][11] ) );
  DFF_X1 \adder_stage1_reg[8][12]  ( .D(n9926), .CK(clk), .Q(
        \adder_stage1[8][12] ) );
  DFF_X1 \adder_stage1_reg[8][13]  ( .D(n9925), .CK(clk), .Q(
        \adder_stage1[8][13] ) );
  DFF_X1 \adder_stage1_reg[8][14]  ( .D(n9924), .CK(clk), .Q(
        \adder_stage1[8][14] ) );
  DFF_X1 \adder_stage1_reg[8][15]  ( .D(n9923), .CK(clk), .Q(
        \adder_stage1[8][15] ) );
  DFF_X1 \adder_stage1_reg[8][20]  ( .D(n9922), .CK(clk), .Q(
        \adder_stage1[8][20] ), .QN(n3465) );
  DFF_X1 \adder_stage1_reg[9][0]  ( .D(n9921), .CK(clk), .Q(
        \adder_stage1[9][0] ) );
  DFF_X1 \adder_stage1_reg[9][1]  ( .D(n9920), .CK(clk), .Q(
        \adder_stage1[9][1] ) );
  DFF_X1 \adder_stage1_reg[9][2]  ( .D(n9919), .CK(clk), .Q(
        \adder_stage1[9][2] ) );
  DFF_X1 \adder_stage1_reg[9][3]  ( .D(n9918), .CK(clk), .Q(
        \adder_stage1[9][3] ) );
  DFF_X1 \adder_stage1_reg[9][4]  ( .D(n9917), .CK(clk), .Q(
        \adder_stage1[9][4] ) );
  DFF_X1 \adder_stage1_reg[9][6]  ( .D(n9915), .CK(clk), .Q(
        \adder_stage1[9][6] ) );
  DFF_X1 \adder_stage1_reg[9][7]  ( .D(n9914), .CK(clk), .Q(
        \adder_stage1[9][7] ) );
  DFF_X1 \adder_stage1_reg[9][8]  ( .D(n9913), .CK(clk), .Q(
        \adder_stage1[9][8] ) );
  DFF_X1 \adder_stage1_reg[9][9]  ( .D(n9912), .CK(clk), .Q(
        \adder_stage1[9][9] ) );
  DFF_X1 \adder_stage1_reg[9][10]  ( .D(n9911), .CK(clk), .Q(
        \adder_stage1[9][10] ) );
  DFF_X1 \adder_stage1_reg[9][11]  ( .D(n9910), .CK(clk), .Q(
        \adder_stage1[9][11] ) );
  DFF_X1 \adder_stage1_reg[9][12]  ( .D(n9909), .CK(clk), .Q(
        \adder_stage1[9][12] ) );
  DFF_X1 \adder_stage1_reg[9][13]  ( .D(n9908), .CK(clk), .Q(
        \adder_stage1[9][13] ) );
  DFF_X1 \adder_stage1_reg[9][14]  ( .D(n9907), .CK(clk), .Q(
        \adder_stage1[9][14] ) );
  DFF_X1 \adder_stage1_reg[9][15]  ( .D(n9906), .CK(clk), .Q(
        \adder_stage1[9][15] ) );
  DFF_X1 \adder_stage1_reg[9][20]  ( .D(n9905), .CK(clk), .Q(
        \adder_stage1[9][20] ), .QN(n3494) );
  DFF_X1 \adder_stage1_reg[10][0]  ( .D(n9904), .CK(clk), .Q(
        \adder_stage1[10][0] ) );
  DFF_X1 \adder_stage1_reg[10][1]  ( .D(n9903), .CK(clk), .Q(
        \adder_stage1[10][1] ) );
  DFF_X1 \adder_stage1_reg[10][3]  ( .D(n9902), .CK(clk), .Q(
        \adder_stage1[10][3] ) );
  DFF_X1 \adder_stage1_reg[10][4]  ( .D(n9901), .CK(clk), .Q(
        \adder_stage1[10][4] ) );
  DFF_X1 \adder_stage1_reg[10][5]  ( .D(n9900), .CK(clk), .Q(
        \adder_stage1[10][5] ) );
  DFF_X1 \adder_stage1_reg[10][6]  ( .D(n9899), .CK(clk), .Q(
        \adder_stage1[10][6] ) );
  DFF_X1 \adder_stage1_reg[10][7]  ( .D(n9898), .CK(clk), .Q(
        \adder_stage1[10][7] ) );
  DFF_X1 \adder_stage1_reg[10][8]  ( .D(n9897), .CK(clk), .Q(
        \adder_stage1[10][8] ) );
  DFF_X1 \adder_stage1_reg[10][9]  ( .D(n9896), .CK(clk), .Q(
        \adder_stage1[10][9] ) );
  DFF_X1 \adder_stage1_reg[10][10]  ( .D(n9895), .CK(clk), .Q(
        \adder_stage1[10][10] ) );
  DFF_X1 \adder_stage1_reg[10][11]  ( .D(n9894), .CK(clk), .Q(
        \adder_stage1[10][11] ) );
  DFF_X1 \adder_stage1_reg[10][12]  ( .D(n9893), .CK(clk), .Q(
        \adder_stage1[10][12] ) );
  DFF_X1 \adder_stage1_reg[10][14]  ( .D(n9892), .CK(clk), .Q(
        \adder_stage1[10][14] ) );
  DFF_X1 \adder_stage1_reg[10][15]  ( .D(n9891), .CK(clk), .Q(
        \adder_stage1[10][15] ) );
  DFF_X1 \adder_stage1_reg[11][0]  ( .D(n9890), .CK(clk), .Q(
        \adder_stage1[11][0] ) );
  DFF_X1 \adder_stage1_reg[11][1]  ( .D(n9889), .CK(clk), .Q(
        \adder_stage1[11][1] ) );
  DFF_X1 \adder_stage1_reg[11][2]  ( .D(n9888), .CK(clk), .Q(
        \adder_stage1[11][2] ) );
  DFF_X1 \adder_stage1_reg[11][3]  ( .D(n9887), .CK(clk), .Q(
        \adder_stage1[11][3] ) );
  DFF_X1 \adder_stage1_reg[11][4]  ( .D(n9886), .CK(clk), .Q(
        \adder_stage1[11][4] ) );
  DFF_X1 \adder_stage1_reg[11][5]  ( .D(n9885), .CK(clk), .Q(
        \adder_stage1[11][5] ) );
  DFF_X1 \adder_stage1_reg[11][6]  ( .D(n9884), .CK(clk), .Q(
        \adder_stage1[11][6] ) );
  DFF_X1 \adder_stage1_reg[11][8]  ( .D(n9882), .CK(clk), .Q(
        \adder_stage1[11][8] ) );
  DFF_X1 \adder_stage1_reg[11][9]  ( .D(n9881), .CK(clk), .Q(
        \adder_stage1[11][9] ) );
  DFF_X1 \adder_stage1_reg[11][10]  ( .D(n9880), .CK(clk), .Q(
        \adder_stage1[11][10] ) );
  DFF_X1 \adder_stage1_reg[11][11]  ( .D(n9879), .CK(clk), .Q(
        \adder_stage1[11][11] ) );
  DFF_X1 \adder_stage1_reg[11][12]  ( .D(n9878), .CK(clk), .Q(
        \adder_stage1[11][12] ) );
  DFF_X1 \adder_stage1_reg[11][13]  ( .D(n9877), .CK(clk), .Q(
        \adder_stage1[11][13] ) );
  DFF_X1 \adder_stage1_reg[11][14]  ( .D(n9876), .CK(clk), .Q(
        \adder_stage1[11][14] ) );
  DFF_X1 \adder_stage1_reg[11][15]  ( .D(n9875), .CK(clk), .Q(
        \adder_stage1[11][15] ) );
  DFF_X1 \adder_stage1_reg[11][20]  ( .D(n9874), .CK(clk), .Q(
        \adder_stage1[11][20] ), .QN(n3495) );
  DFF_X1 \adder_stage1_reg[12][0]  ( .D(n9873), .CK(clk), .Q(
        \adder_stage1[12][0] ) );
  DFF_X1 \adder_stage1_reg[12][1]  ( .D(n9872), .CK(clk), .Q(
        \adder_stage1[12][1] ) );
  DFF_X1 \adder_stage1_reg[12][2]  ( .D(n9871), .CK(clk), .Q(
        \adder_stage1[12][2] ) );
  DFF_X1 \adder_stage1_reg[12][3]  ( .D(n9870), .CK(clk), .Q(
        \adder_stage1[12][3] ) );
  DFF_X1 \adder_stage1_reg[12][4]  ( .D(n9869), .CK(clk), .Q(
        \adder_stage1[12][4] ) );
  DFF_X1 \adder_stage1_reg[12][5]  ( .D(n9868), .CK(clk), .Q(
        \adder_stage1[12][5] ) );
  DFF_X1 \adder_stage1_reg[12][6]  ( .D(n9867), .CK(clk), .Q(
        \adder_stage1[12][6] ) );
  DFF_X1 \adder_stage1_reg[12][7]  ( .D(n9866), .CK(clk), .Q(
        \adder_stage1[12][7] ) );
  DFF_X1 \adder_stage1_reg[12][8]  ( .D(n9865), .CK(clk), .Q(
        \adder_stage1[12][8] ) );
  DFF_X1 \adder_stage1_reg[12][9]  ( .D(n9864), .CK(clk), .Q(
        \adder_stage1[12][9] ) );
  DFF_X1 \adder_stage1_reg[12][10]  ( .D(n9863), .CK(clk), .Q(
        \adder_stage1[12][10] ) );
  DFF_X1 \adder_stage1_reg[12][11]  ( .D(n9862), .CK(clk), .Q(
        \adder_stage1[12][11] ) );
  DFF_X1 \adder_stage1_reg[12][12]  ( .D(n9861), .CK(clk), .Q(
        \adder_stage1[12][12] ) );
  DFF_X1 \adder_stage1_reg[12][13]  ( .D(n9860), .CK(clk), .Q(
        \adder_stage1[12][13] ) );
  DFF_X1 \adder_stage1_reg[12][14]  ( .D(n9859), .CK(clk), .Q(
        \adder_stage1[12][14] ) );
  DFF_X1 \adder_stage1_reg[12][15]  ( .D(n9858), .CK(clk), .Q(
        \adder_stage1[12][15] ) );
  DFF_X1 \adder_stage1_reg[12][20]  ( .D(n9857), .CK(clk), .Q(
        \adder_stage1[12][20] ), .QN(n3462) );
  DFF_X1 \adder_stage1_reg[13][0]  ( .D(n9856), .CK(clk), .Q(
        \adder_stage1[13][0] ) );
  DFF_X1 \adder_stage1_reg[13][1]  ( .D(n9855), .CK(clk), .Q(
        \adder_stage1[13][1] ) );
  DFF_X1 \adder_stage1_reg[13][2]  ( .D(n9854), .CK(clk), .Q(
        \adder_stage1[13][2] ) );
  DFF_X1 \adder_stage1_reg[13][4]  ( .D(n9852), .CK(clk), .Q(
        \adder_stage1[13][4] ) );
  DFF_X1 \adder_stage1_reg[13][5]  ( .D(n9851), .CK(clk), .Q(
        \adder_stage1[13][5] ) );
  DFF_X1 \adder_stage1_reg[13][6]  ( .D(n9850), .CK(clk), .Q(
        \adder_stage1[13][6] ) );
  DFF_X1 \adder_stage1_reg[13][7]  ( .D(n9849), .CK(clk), .Q(
        \adder_stage1[13][7] ) );
  DFF_X1 \adder_stage1_reg[13][8]  ( .D(n9848), .CK(clk), .Q(
        \adder_stage1[13][8] ) );
  DFF_X1 \adder_stage1_reg[13][9]  ( .D(n9847), .CK(clk), .Q(
        \adder_stage1[13][9] ) );
  DFF_X1 \adder_stage1_reg[13][10]  ( .D(n9846), .CK(clk), .Q(
        \adder_stage1[13][10] ) );
  DFF_X1 \adder_stage1_reg[13][11]  ( .D(n9845), .CK(clk), .Q(
        \adder_stage1[13][11] ) );
  DFF_X1 \adder_stage1_reg[13][12]  ( .D(n9844), .CK(clk), .Q(
        \adder_stage1[13][12] ) );
  DFF_X1 \adder_stage1_reg[13][13]  ( .D(n9843), .CK(clk), .Q(
        \adder_stage1[13][13] ) );
  DFF_X1 \adder_stage1_reg[13][14]  ( .D(n9842), .CK(clk), .Q(
        \adder_stage1[13][14] ) );
  DFF_X1 \adder_stage1_reg[13][15]  ( .D(n9841), .CK(clk), .Q(
        \adder_stage1[13][15] ) );
  DFF_X1 \adder_stage1_reg[13][20]  ( .D(n9840), .CK(clk), .Q(
        \adder_stage1[13][20] ), .QN(n3496) );
  DFF_X1 \adder_stage1_reg[14][0]  ( .D(n9839), .CK(clk), .Q(
        \adder_stage1[14][0] ) );
  DFF_X1 \adder_stage1_reg[14][1]  ( .D(n9838), .CK(clk), .Q(
        \adder_stage1[14][1] ) );
  DFF_X1 \adder_stage1_reg[14][2]  ( .D(n9837), .CK(clk), .Q(
        \adder_stage1[14][2] ) );
  DFF_X1 \adder_stage1_reg[14][3]  ( .D(n9836), .CK(clk), .Q(
        \adder_stage1[14][3] ) );
  DFF_X1 \adder_stage1_reg[14][4]  ( .D(n9835), .CK(clk), .Q(
        \adder_stage1[14][4] ) );
  DFF_X1 \adder_stage1_reg[14][5]  ( .D(n9834), .CK(clk), .Q(
        \adder_stage1[14][5] ) );
  DFF_X1 \adder_stage1_reg[14][6]  ( .D(n9833), .CK(clk), .Q(
        \adder_stage1[14][6] ) );
  DFF_X1 \adder_stage1_reg[14][7]  ( .D(n9832), .CK(clk), .Q(
        \adder_stage1[14][7] ) );
  DFF_X1 \adder_stage1_reg[14][8]  ( .D(n9831), .CK(clk), .Q(
        \adder_stage1[14][8] ) );
  DFF_X1 \adder_stage1_reg[14][9]  ( .D(n9830), .CK(clk), .Q(
        \adder_stage1[14][9] ) );
  DFF_X1 \adder_stage1_reg[14][10]  ( .D(n9829), .CK(clk), .Q(
        \adder_stage1[14][10] ) );
  DFF_X1 \adder_stage1_reg[14][11]  ( .D(n9828), .CK(clk), .Q(
        \adder_stage1[14][11] ) );
  DFF_X1 \adder_stage1_reg[14][12]  ( .D(n9827), .CK(clk), .Q(
        \adder_stage1[14][12] ) );
  DFF_X1 \adder_stage1_reg[14][13]  ( .D(n9826), .CK(clk), .Q(
        \adder_stage1[14][13] ) );
  DFF_X1 \adder_stage1_reg[14][14]  ( .D(n9825), .CK(clk), .Q(
        \adder_stage1[14][14] ) );
  DFF_X1 \adder_stage1_reg[14][15]  ( .D(n9824), .CK(clk), .Q(
        \adder_stage1[14][15] ) );
  DFF_X1 \adder_stage1_reg[14][20]  ( .D(n9823), .CK(clk), .Q(
        \adder_stage1[14][20] ), .QN(n3455) );
  DFF_X1 \adder_stage1_reg[15][0]  ( .D(n9822), .CK(clk), .Q(
        \adder_stage1[15][0] ) );
  DFF_X1 \adder_stage1_reg[15][1]  ( .D(n9821), .CK(clk), .Q(
        \adder_stage1[15][1] ) );
  DFF_X1 \adder_stage1_reg[15][2]  ( .D(n9820), .CK(clk), .Q(
        \adder_stage1[15][2] ) );
  DFF_X1 \adder_stage1_reg[15][3]  ( .D(n9819), .CK(clk), .Q(
        \adder_stage1[15][3] ) );
  DFF_X1 \adder_stage1_reg[15][4]  ( .D(n9818), .CK(clk), .Q(
        \adder_stage1[15][4] ) );
  DFF_X1 \adder_stage1_reg[15][5]  ( .D(n9817), .CK(clk), .Q(
        \adder_stage1[15][5] ) );
  DFF_X1 \adder_stage1_reg[15][6]  ( .D(n9816), .CK(clk), .Q(
        \adder_stage1[15][6] ) );
  DFF_X1 \adder_stage1_reg[15][7]  ( .D(n9815), .CK(clk), .Q(
        \adder_stage1[15][7] ) );
  DFF_X1 \adder_stage1_reg[15][8]  ( .D(n9814), .CK(clk), .Q(
        \adder_stage1[15][8] ) );
  DFF_X1 \adder_stage1_reg[15][9]  ( .D(n9813), .CK(clk), .Q(
        \adder_stage1[15][9] ) );
  DFF_X1 \adder_stage1_reg[15][10]  ( .D(n9812), .CK(clk), .Q(
        \adder_stage1[15][10] ) );
  DFF_X1 \adder_stage1_reg[15][11]  ( .D(n9811), .CK(clk), .Q(
        \adder_stage1[15][11] ) );
  DFF_X1 \adder_stage1_reg[15][12]  ( .D(n9810), .CK(clk), .Q(
        \adder_stage1[15][12] ) );
  DFF_X1 \adder_stage1_reg[15][13]  ( .D(n9809), .CK(clk), .Q(
        \adder_stage1[15][13] ) );
  DFF_X1 \adder_stage1_reg[15][14]  ( .D(n9808), .CK(clk), .Q(
        \adder_stage1[15][14] ) );
  DFF_X1 \adder_stage1_reg[15][15]  ( .D(n9807), .CK(clk), .Q(
        \adder_stage1[15][15] ) );
  DFF_X1 \adder_stage1_reg[15][20]  ( .D(n9806), .CK(clk), .Q(
        \adder_stage1[15][20] ), .QN(n3485) );
  DFF_X1 \adder_stage2_reg[0][0]  ( .D(n9805), .CK(clk), .Q(
        \adder_stage2[0][0] ) );
  DFF_X1 \adder_stage2_reg[0][1]  ( .D(n9804), .CK(clk), .Q(
        \adder_stage2[0][1] ) );
  DFF_X1 \adder_stage2_reg[0][2]  ( .D(n9803), .CK(clk), .Q(
        \adder_stage2[0][2] ) );
  DFF_X1 \adder_stage2_reg[0][3]  ( .D(n9802), .CK(clk), .Q(
        \adder_stage2[0][3] ) );
  DFF_X1 \adder_stage2_reg[0][4]  ( .D(n9801), .CK(clk), .Q(
        \adder_stage2[0][4] ) );
  DFF_X1 \adder_stage2_reg[0][5]  ( .D(n9800), .CK(clk), .Q(
        \adder_stage2[0][5] ) );
  DFF_X1 \adder_stage2_reg[0][6]  ( .D(n9799), .CK(clk), .Q(
        \adder_stage2[0][6] ) );
  DFF_X1 \adder_stage2_reg[0][7]  ( .D(n9798), .CK(clk), .Q(
        \adder_stage2[0][7] ) );
  DFF_X1 \adder_stage2_reg[0][8]  ( .D(n9797), .CK(clk), .Q(
        \adder_stage2[0][8] ) );
  DFF_X1 \adder_stage2_reg[0][9]  ( .D(n9796), .CK(clk), .Q(
        \adder_stage2[0][9] ) );
  DFF_X1 \adder_stage2_reg[0][10]  ( .D(n9795), .CK(clk), .Q(
        \adder_stage2[0][10] ) );
  DFF_X1 \adder_stage2_reg[0][11]  ( .D(n9794), .CK(clk), .Q(
        \adder_stage2[0][11] ) );
  DFF_X1 \adder_stage2_reg[0][12]  ( .D(n9793), .CK(clk), .Q(
        \adder_stage2[0][12] ) );
  DFF_X1 \adder_stage2_reg[0][13]  ( .D(n9792), .CK(clk), .Q(
        \adder_stage2[0][13] ) );
  DFF_X1 \adder_stage2_reg[0][14]  ( .D(n9791), .CK(clk), .Q(
        \adder_stage2[0][14] ) );
  DFF_X1 \adder_stage2_reg[0][15]  ( .D(n9790), .CK(clk), .Q(
        \adder_stage2[0][15] ) );
  DFF_X1 \adder_stage2_reg[0][16]  ( .D(n9789), .CK(clk), .Q(
        \adder_stage2[0][16] ) );
  DFF_X1 \adder_stage2_reg[0][17]  ( .D(n2059), .CK(clk), .Q(
        \adder_stage2[0][17] ), .QN(n8735) );
  DFF_X1 \adder_stage2_reg[0][18]  ( .D(n2058), .CK(clk), .Q(
        \adder_stage2[0][18] ), .QN(n8736) );
  DFF_X1 \adder_stage2_reg[0][19]  ( .D(n2057), .CK(clk), .Q(
        \adder_stage2[0][19] ), .QN(n8737) );
  DFF_X1 \adder_stage2_reg[0][20]  ( .D(n2056), .CK(clk), .Q(
        \adder_stage2[0][20] ), .QN(n8748) );
  DFF_X1 \adder_stage2_reg[1][0]  ( .D(n9788), .CK(clk), .Q(
        \adder_stage2[1][0] ) );
  DFF_X1 \adder_stage2_reg[1][1]  ( .D(n9787), .CK(clk), .Q(
        \adder_stage2[1][1] ) );
  DFF_X1 \adder_stage2_reg[1][2]  ( .D(n9786), .CK(clk), .Q(
        \adder_stage2[1][2] ) );
  DFF_X1 \adder_stage2_reg[1][3]  ( .D(n9785), .CK(clk), .Q(
        \adder_stage2[1][3] ) );
  DFF_X1 \adder_stage2_reg[1][4]  ( .D(n9784), .CK(clk), .Q(
        \adder_stage2[1][4] ) );
  DFF_X1 \adder_stage2_reg[1][5]  ( .D(n9783), .CK(clk), .Q(
        \adder_stage2[1][5] ) );
  DFF_X1 \adder_stage2_reg[1][6]  ( .D(n9782), .CK(clk), .Q(
        \adder_stage2[1][6] ) );
  DFF_X1 \adder_stage2_reg[1][7]  ( .D(n9781), .CK(clk), .Q(
        \adder_stage2[1][7] ) );
  DFF_X1 \adder_stage2_reg[1][8]  ( .D(n9780), .CK(clk), .Q(
        \adder_stage2[1][8] ) );
  DFF_X1 \adder_stage2_reg[1][9]  ( .D(n9779), .CK(clk), .Q(
        \adder_stage2[1][9] ) );
  DFF_X1 \adder_stage2_reg[1][10]  ( .D(n9778), .CK(clk), .Q(
        \adder_stage2[1][10] ) );
  DFF_X1 \adder_stage2_reg[1][11]  ( .D(n9777), .CK(clk), .Q(
        \adder_stage2[1][11] ) );
  DFF_X1 \adder_stage2_reg[1][12]  ( .D(n9776), .CK(clk), .Q(
        \adder_stage2[1][12] ) );
  DFF_X1 \adder_stage2_reg[1][13]  ( .D(n9775), .CK(clk), .Q(
        \adder_stage2[1][13] ) );
  DFF_X1 \adder_stage2_reg[1][14]  ( .D(n9774), .CK(clk), .Q(
        \adder_stage2[1][14] ) );
  DFF_X1 \adder_stage2_reg[1][15]  ( .D(n9773), .CK(clk), .Q(
        \adder_stage2[1][15] ) );
  DFF_X1 \adder_stage2_reg[1][16]  ( .D(n9772), .CK(clk), .Q(
        \adder_stage2[1][16] ) );
  DFF_X1 \adder_stage2_reg[1][17]  ( .D(n2038), .CK(clk), .Q(
        \adder_stage2[1][17] ), .QN(n8723) );
  DFF_X1 \adder_stage2_reg[1][18]  ( .D(n2037), .CK(clk), .Q(
        \adder_stage2[1][18] ), .QN(n8724) );
  DFF_X1 \adder_stage2_reg[1][19]  ( .D(n2036), .CK(clk), .Q(
        \adder_stage2[1][19] ), .QN(n8725) );
  DFF_X1 \adder_stage2_reg[1][20]  ( .D(n2035), .CK(clk), .Q(
        \adder_stage2[1][20] ), .QN(n8752) );
  DFF_X1 \adder_stage2_reg[2][0]  ( .D(n9771), .CK(clk), .Q(
        \adder_stage2[2][0] ) );
  DFF_X1 \adder_stage2_reg[2][1]  ( .D(n9770), .CK(clk), .Q(
        \adder_stage2[2][1] ) );
  DFF_X1 \adder_stage2_reg[2][2]  ( .D(n9769), .CK(clk), .Q(
        \adder_stage2[2][2] ) );
  DFF_X1 \adder_stage2_reg[2][3]  ( .D(n9768), .CK(clk), .Q(
        \adder_stage2[2][3] ) );
  DFF_X1 \adder_stage2_reg[2][4]  ( .D(n9767), .CK(clk), .Q(
        \adder_stage2[2][4] ) );
  DFF_X1 \adder_stage2_reg[2][5]  ( .D(n9766), .CK(clk), .Q(
        \adder_stage2[2][5] ) );
  DFF_X1 \adder_stage2_reg[2][6]  ( .D(n9765), .CK(clk), .Q(
        \adder_stage2[2][6] ) );
  DFF_X1 \adder_stage2_reg[2][7]  ( .D(n9764), .CK(clk), .Q(
        \adder_stage2[2][7] ) );
  DFF_X1 \adder_stage2_reg[2][8]  ( .D(n9763), .CK(clk), .Q(
        \adder_stage2[2][8] ) );
  DFF_X1 \adder_stage2_reg[2][9]  ( .D(n9762), .CK(clk), .Q(
        \adder_stage2[2][9] ) );
  DFF_X1 \adder_stage2_reg[2][10]  ( .D(n9761), .CK(clk), .Q(
        \adder_stage2[2][10] ) );
  DFF_X1 \adder_stage2_reg[2][11]  ( .D(n9760), .CK(clk), .Q(
        \adder_stage2[2][11] ) );
  DFF_X1 \adder_stage2_reg[2][12]  ( .D(n9759), .CK(clk), .Q(
        \adder_stage2[2][12] ) );
  DFF_X1 \adder_stage2_reg[2][13]  ( .D(n9758), .CK(clk), .Q(
        \adder_stage2[2][13] ) );
  DFF_X1 \adder_stage2_reg[2][14]  ( .D(n9757), .CK(clk), .Q(
        \adder_stage2[2][14] ) );
  DFF_X1 \adder_stage2_reg[2][15]  ( .D(n9756), .CK(clk), .Q(
        \adder_stage2[2][15] ) );
  DFF_X1 \adder_stage2_reg[2][16]  ( .D(n9755), .CK(clk), .Q(
        \adder_stage2[2][16] ) );
  DFF_X1 \adder_stage2_reg[2][17]  ( .D(n2017), .CK(clk), .Q(
        \adder_stage2[2][17] ), .QN(n8732) );
  DFF_X1 \adder_stage2_reg[2][18]  ( .D(n2016), .CK(clk), .Q(
        \adder_stage2[2][18] ), .QN(n8733) );
  DFF_X1 \adder_stage2_reg[2][19]  ( .D(n2015), .CK(clk), .Q(
        \adder_stage2[2][19] ), .QN(n8734) );
  DFF_X1 \adder_stage2_reg[2][20]  ( .D(n2014), .CK(clk), .Q(
        \adder_stage2[2][20] ), .QN(n8747) );
  DFF_X1 \adder_stage2_reg[3][0]  ( .D(n9754), .CK(clk), .Q(
        \adder_stage2[3][0] ) );
  DFF_X1 \adder_stage2_reg[3][1]  ( .D(n9753), .CK(clk), .Q(
        \adder_stage2[3][1] ) );
  DFF_X1 \adder_stage2_reg[3][2]  ( .D(n9752), .CK(clk), .Q(
        \adder_stage2[3][2] ) );
  DFF_X1 \adder_stage2_reg[3][3]  ( .D(n9751), .CK(clk), .Q(
        \adder_stage2[3][3] ) );
  DFF_X1 \adder_stage2_reg[3][4]  ( .D(n9750), .CK(clk), .Q(
        \adder_stage2[3][4] ) );
  DFF_X1 \adder_stage2_reg[3][5]  ( .D(n9749), .CK(clk), .Q(
        \adder_stage2[3][5] ) );
  DFF_X1 \adder_stage2_reg[3][6]  ( .D(n9748), .CK(clk), .Q(
        \adder_stage2[3][6] ) );
  DFF_X1 \adder_stage2_reg[3][7]  ( .D(n9747), .CK(clk), .Q(
        \adder_stage2[3][7] ) );
  DFF_X1 \adder_stage2_reg[3][8]  ( .D(n9746), .CK(clk), .Q(
        \adder_stage2[3][8] ) );
  DFF_X1 \adder_stage2_reg[3][9]  ( .D(n9745), .CK(clk), .Q(
        \adder_stage2[3][9] ) );
  DFF_X1 \adder_stage2_reg[3][10]  ( .D(n9744), .CK(clk), .Q(
        \adder_stage2[3][10] ) );
  DFF_X1 \adder_stage2_reg[3][12]  ( .D(n9742), .CK(clk), .Q(
        \adder_stage2[3][12] ) );
  DFF_X1 \adder_stage2_reg[3][13]  ( .D(n9741), .CK(clk), .Q(
        \adder_stage2[3][13] ) );
  DFF_X1 \adder_stage2_reg[3][14]  ( .D(n9740), .CK(clk), .Q(
        \adder_stage2[3][14] ) );
  DFF_X1 \adder_stage2_reg[3][15]  ( .D(n9739), .CK(clk), .Q(
        \adder_stage2[3][15] ) );
  DFF_X1 \adder_stage2_reg[3][16]  ( .D(n9738), .CK(clk), .Q(
        \adder_stage2[3][16] ) );
  DFF_X1 \adder_stage2_reg[3][17]  ( .D(n1996), .CK(clk), .Q(
        \adder_stage2[3][17] ), .QN(n8726) );
  DFF_X1 \adder_stage2_reg[3][18]  ( .D(n1995), .CK(clk), .Q(
        \adder_stage2[3][18] ), .QN(n8727) );
  DFF_X1 \adder_stage2_reg[3][19]  ( .D(n1994), .CK(clk), .Q(
        \adder_stage2[3][19] ), .QN(n8728) );
  DFF_X1 \adder_stage2_reg[3][20]  ( .D(n1993), .CK(clk), .Q(
        \adder_stage2[3][20] ), .QN(n8753) );
  DFF_X1 \adder_stage2_reg[4][0]  ( .D(n9737), .CK(clk), .Q(
        \adder_stage2[4][0] ) );
  DFF_X1 \adder_stage2_reg[4][1]  ( .D(n9736), .CK(clk), .Q(
        \adder_stage2[4][1] ) );
  DFF_X1 \adder_stage2_reg[4][2]  ( .D(n9735), .CK(clk), .Q(
        \adder_stage2[4][2] ) );
  DFF_X1 \adder_stage2_reg[4][3]  ( .D(n9734), .CK(clk), .Q(
        \adder_stage2[4][3] ) );
  DFF_X1 \adder_stage2_reg[4][4]  ( .D(n9733), .CK(clk), .Q(
        \adder_stage2[4][4] ) );
  DFF_X1 \adder_stage2_reg[4][5]  ( .D(n9732), .CK(clk), .Q(
        \adder_stage2[4][5] ) );
  DFF_X1 \adder_stage2_reg[4][6]  ( .D(n9731), .CK(clk), .Q(
        \adder_stage2[4][6] ) );
  DFF_X1 \adder_stage2_reg[4][7]  ( .D(n9730), .CK(clk), .Q(
        \adder_stage2[4][7] ) );
  DFF_X1 \adder_stage2_reg[4][8]  ( .D(n9729), .CK(clk), .Q(
        \adder_stage2[4][8] ) );
  DFF_X1 \adder_stage2_reg[4][9]  ( .D(n9728), .CK(clk), .Q(
        \adder_stage2[4][9] ) );
  DFF_X1 \adder_stage2_reg[4][10]  ( .D(n9727), .CK(clk), .Q(
        \adder_stage2[4][10] ) );
  DFF_X1 \adder_stage2_reg[4][11]  ( .D(n9726), .CK(clk), .Q(
        \adder_stage2[4][11] ) );
  DFF_X1 \adder_stage2_reg[4][12]  ( .D(n9725), .CK(clk), .Q(
        \adder_stage2[4][12] ) );
  DFF_X1 \adder_stage2_reg[4][13]  ( .D(n9724), .CK(clk), .Q(
        \adder_stage2[4][13] ) );
  DFF_X1 \adder_stage2_reg[4][14]  ( .D(n9723), .CK(clk), .Q(
        \adder_stage2[4][14] ) );
  DFF_X1 \adder_stage2_reg[4][15]  ( .D(n9722), .CK(clk), .Q(
        \adder_stage2[4][15] ) );
  DFF_X1 \adder_stage2_reg[4][16]  ( .D(n9721), .CK(clk), .Q(
        \adder_stage2[4][16] ) );
  DFF_X1 \adder_stage2_reg[4][17]  ( .D(n1975), .CK(clk), .Q(
        \adder_stage2[4][17] ), .QN(n8738) );
  DFF_X1 \adder_stage2_reg[4][18]  ( .D(n1974), .CK(clk), .Q(
        \adder_stage2[4][18] ), .QN(n8739) );
  DFF_X1 \adder_stage2_reg[4][19]  ( .D(n1973), .CK(clk), .Q(
        \adder_stage2[4][19] ), .QN(n8740) );
  DFF_X1 \adder_stage2_reg[4][20]  ( .D(n1972), .CK(clk), .Q(
        \adder_stage2[4][20] ), .QN(n8749) );
  DFF_X1 \adder_stage2_reg[5][0]  ( .D(n9720), .CK(clk), .Q(
        \adder_stage2[5][0] ) );
  DFF_X1 \adder_stage2_reg[5][1]  ( .D(n9719), .CK(clk), .Q(
        \adder_stage2[5][1] ) );
  DFF_X1 \adder_stage2_reg[5][2]  ( .D(n9718), .CK(clk), .Q(
        \adder_stage2[5][2] ) );
  DFF_X1 \adder_stage2_reg[5][3]  ( .D(n9717), .CK(clk), .Q(
        \adder_stage2[5][3] ) );
  DFF_X1 \adder_stage2_reg[5][4]  ( .D(n9716), .CK(clk), .Q(
        \adder_stage2[5][4] ) );
  DFF_X1 \adder_stage2_reg[5][5]  ( .D(n9715), .CK(clk), .Q(
        \adder_stage2[5][5] ) );
  DFF_X1 \adder_stage2_reg[5][6]  ( .D(n9714), .CK(clk), .Q(
        \adder_stage2[5][6] ) );
  DFF_X1 \adder_stage2_reg[5][8]  ( .D(n9712), .CK(clk), .Q(
        \adder_stage2[5][8] ) );
  DFF_X1 \adder_stage2_reg[5][9]  ( .D(n9711), .CK(clk), .Q(
        \adder_stage2[5][9] ) );
  DFF_X1 \adder_stage2_reg[5][10]  ( .D(n9710), .CK(clk), .Q(
        \adder_stage2[5][10] ) );
  DFF_X1 \adder_stage2_reg[5][12]  ( .D(n9708), .CK(clk), .Q(
        \adder_stage2[5][12] ) );
  DFF_X1 \adder_stage2_reg[5][13]  ( .D(n9707), .CK(clk), .Q(
        \adder_stage2[5][13] ) );
  DFF_X1 \adder_stage2_reg[5][14]  ( .D(n9706), .CK(clk), .Q(
        \adder_stage2[5][14] ) );
  DFF_X1 \adder_stage2_reg[5][15]  ( .D(n9705), .CK(clk), .Q(
        \adder_stage2[5][15] ) );
  DFF_X1 \adder_stage2_reg[5][16]  ( .D(n9704), .CK(clk), .Q(
        \adder_stage2[5][16] ) );
  DFF_X1 \adder_stage2_reg[5][17]  ( .D(n1954), .CK(clk), .Q(
        \adder_stage2[5][17] ), .QN(n8729) );
  DFF_X1 \adder_stage2_reg[5][18]  ( .D(n1953), .CK(clk), .Q(
        \adder_stage2[5][18] ), .QN(n8730) );
  DFF_X1 \adder_stage2_reg[5][19]  ( .D(n1952), .CK(clk), .Q(
        \adder_stage2[5][19] ), .QN(n8731) );
  DFF_X1 \adder_stage2_reg[5][20]  ( .D(n1951), .CK(clk), .Q(
        \adder_stage2[5][20] ), .QN(n8754) );
  DFF_X1 \adder_stage2_reg[6][0]  ( .D(n9703), .CK(clk), .Q(
        \adder_stage2[6][0] ) );
  DFF_X1 \adder_stage2_reg[6][1]  ( .D(n9702), .CK(clk), .Q(
        \adder_stage2[6][1] ) );
  DFF_X1 \adder_stage2_reg[6][2]  ( .D(n9701), .CK(clk), .Q(
        \adder_stage2[6][2] ) );
  DFF_X1 \adder_stage2_reg[6][3]  ( .D(n9700), .CK(clk), .Q(
        \adder_stage2[6][3] ), .QN(n3439) );
  DFF_X1 \adder_stage2_reg[6][4]  ( .D(n9699), .CK(clk), .Q(
        \adder_stage2[6][4] ) );
  DFF_X1 \adder_stage2_reg[6][5]  ( .D(n9698), .CK(clk), .Q(
        \adder_stage2[6][5] ) );
  DFF_X1 \adder_stage2_reg[6][6]  ( .D(n9697), .CK(clk), .Q(
        \adder_stage2[6][6] ) );
  DFF_X1 \adder_stage2_reg[6][7]  ( .D(n9696), .CK(clk), .Q(
        \adder_stage2[6][7] ) );
  DFF_X1 \adder_stage2_reg[6][8]  ( .D(n9695), .CK(clk), .Q(
        \adder_stage2[6][8] ) );
  DFF_X1 \adder_stage2_reg[6][9]  ( .D(n9694), .CK(clk), .Q(
        \adder_stage2[6][9] ), .QN(n3441) );
  DFF_X1 \adder_stage2_reg[6][10]  ( .D(n9693), .CK(clk), .Q(
        \adder_stage2[6][10] ) );
  DFF_X1 \adder_stage2_reg[6][11]  ( .D(n9692), .CK(clk), .Q(
        \adder_stage2[6][11] ), .QN(n3444) );
  DFF_X1 \adder_stage2_reg[6][12]  ( .D(n9691), .CK(clk), .Q(
        \adder_stage2[6][12] ) );
  DFF_X1 \adder_stage2_reg[6][13]  ( .D(n9690), .CK(clk), .Q(
        \adder_stage2[6][13] ) );
  DFF_X1 \adder_stage2_reg[6][14]  ( .D(n9689), .CK(clk), .Q(
        \adder_stage2[6][14] ) );
  DFF_X1 \adder_stage2_reg[6][15]  ( .D(n9688), .CK(clk), .Q(
        \adder_stage2[6][15] ) );
  DFF_X1 \adder_stage2_reg[6][16]  ( .D(n9687), .CK(clk), .Q(
        \adder_stage2[6][16] ) );
  DFF_X1 \adder_stage2_reg[6][17]  ( .D(n1933), .CK(clk), .Q(
        \adder_stage2[6][17] ), .QN(n8741) );
  DFF_X1 \adder_stage2_reg[6][18]  ( .D(n1932), .CK(clk), .Q(
        \adder_stage2[6][18] ), .QN(n8742) );
  DFF_X1 \adder_stage2_reg[6][19]  ( .D(n1931), .CK(clk), .Q(
        \adder_stage2[6][19] ), .QN(n8743) );
  DFF_X1 \adder_stage2_reg[6][20]  ( .D(n1930), .CK(clk), .Q(
        \adder_stage2[6][20] ), .QN(n8750) );
  DFF_X1 \adder_stage2_reg[7][0]  ( .D(n9686), .CK(clk), .Q(
        \adder_stage2[7][0] ) );
  DFF_X1 \adder_stage2_reg[7][1]  ( .D(n9685), .CK(clk), .Q(
        \adder_stage2[7][1] ) );
  DFF_X1 \adder_stage2_reg[7][2]  ( .D(n9684), .CK(clk), .Q(
        \adder_stage2[7][2] ) );
  DFF_X1 \adder_stage2_reg[7][4]  ( .D(n9682), .CK(clk), .Q(
        \adder_stage2[7][4] ) );
  DFF_X1 \adder_stage2_reg[7][5]  ( .D(n9681), .CK(clk), .Q(
        \adder_stage2[7][5] ) );
  DFF_X1 \adder_stage2_reg[7][6]  ( .D(n9680), .CK(clk), .Q(
        \adder_stage2[7][6] ) );
  DFF_X1 \adder_stage2_reg[7][7]  ( .D(n9679), .CK(clk), .Q(
        \adder_stage2[7][7] ) );
  DFF_X1 \adder_stage2_reg[7][8]  ( .D(n9678), .CK(clk), .Q(
        \adder_stage2[7][8] ) );
  DFF_X1 \adder_stage2_reg[7][9]  ( .D(n9677), .CK(clk), .Q(
        \adder_stage2[7][9] ), .QN(n3442) );
  DFF_X1 \adder_stage2_reg[7][10]  ( .D(n9676), .CK(clk), .Q(
        \adder_stage2[7][10] ) );
  DFF_X1 \adder_stage2_reg[7][11]  ( .D(n9675), .CK(clk), .Q(
        \adder_stage2[7][11] ), .QN(n3445) );
  DFF_X1 \adder_stage2_reg[7][12]  ( .D(n9674), .CK(clk), .Q(
        \adder_stage2[7][12] ) );
  DFF_X1 \adder_stage2_reg[7][13]  ( .D(n9673), .CK(clk), .Q(
        \adder_stage2[7][13] ) );
  DFF_X1 \adder_stage2_reg[7][14]  ( .D(n9672), .CK(clk), .Q(
        \adder_stage2[7][14] ) );
  DFF_X1 \adder_stage2_reg[7][15]  ( .D(n9671), .CK(clk), .Q(
        \adder_stage2[7][15] ) );
  DFF_X1 \adder_stage2_reg[7][16]  ( .D(n9670), .CK(clk), .Q(
        \adder_stage2[7][16] ) );
  DFF_X1 \adder_stage2_reg[7][17]  ( .D(n1912), .CK(clk), .Q(
        \adder_stage2[7][17] ), .QN(n8720) );
  DFF_X1 \adder_stage2_reg[7][18]  ( .D(n1911), .CK(clk), .Q(
        \adder_stage2[7][18] ), .QN(n8721) );
  DFF_X1 \adder_stage2_reg[7][19]  ( .D(n1910), .CK(clk), .Q(
        \adder_stage2[7][19] ), .QN(n8722) );
  DFF_X1 \adder_stage3_reg[0][0]  ( .D(n9669), .CK(clk), .Q(
        \adder_stage3[0][0] ) );
  DFF_X1 \adder_stage3_reg[0][1]  ( .D(n9668), .CK(clk), .Q(
        \adder_stage3[0][1] ) );
  DFF_X1 \adder_stage3_reg[0][2]  ( .D(n9667), .CK(clk), .Q(
        \adder_stage3[0][2] ) );
  DFF_X1 \adder_stage3_reg[0][3]  ( .D(n9666), .CK(clk), .Q(
        \adder_stage3[0][3] ) );
  DFF_X1 \adder_stage3_reg[0][4]  ( .D(n9665), .CK(clk), .Q(
        \adder_stage3[0][4] ) );
  DFF_X1 \adder_stage3_reg[0][5]  ( .D(n9664), .CK(clk), .Q(
        \adder_stage3[0][5] ) );
  DFF_X1 \adder_stage3_reg[0][6]  ( .D(n9663), .CK(clk), .Q(
        \adder_stage3[0][6] ) );
  DFF_X1 \adder_stage3_reg[0][7]  ( .D(n9662), .CK(clk), .Q(
        \adder_stage3[0][7] ) );
  DFF_X1 \adder_stage3_reg[0][8]  ( .D(n9661), .CK(clk), .Q(
        \adder_stage3[0][8] ) );
  DFF_X1 \adder_stage3_reg[0][9]  ( .D(n9660), .CK(clk), .Q(
        \adder_stage3[0][9] ) );
  DFF_X1 \adder_stage3_reg[0][10]  ( .D(n9659), .CK(clk), .Q(
        \adder_stage3[0][10] ) );
  DFF_X1 \adder_stage3_reg[0][11]  ( .D(n9658), .CK(clk), .Q(
        \adder_stage3[0][11] ) );
  DFF_X1 \adder_stage3_reg[0][12]  ( .D(n9657), .CK(clk), .Q(
        \adder_stage3[0][12] ) );
  DFF_X1 \adder_stage3_reg[0][13]  ( .D(n9656), .CK(clk), .Q(
        \adder_stage3[0][13] ) );
  DFF_X1 \adder_stage3_reg[0][14]  ( .D(n9655), .CK(clk), .Q(
        \adder_stage3[0][14] ) );
  DFF_X1 \adder_stage3_reg[0][15]  ( .D(n9654), .CK(clk), .Q(
        \adder_stage3[0][15] ) );
  DFF_X1 \adder_stage3_reg[0][16]  ( .D(n9653), .CK(clk), .Q(
        \adder_stage3[0][16] ) );
  DFF_X1 \adder_stage3_reg[0][17]  ( .D(n9652), .CK(clk), .Q(
        \adder_stage3[0][17] ) );
  DFF_X1 \adder_stage3_reg[0][20]  ( .D(n9651), .CK(clk), .Q(
        \adder_stage3[0][20] ) );
  DFF_X1 \adder_stage3_reg[1][0]  ( .D(n9650), .CK(clk), .Q(
        \adder_stage3[1][0] ) );
  DFF_X1 \adder_stage3_reg[1][1]  ( .D(n9649), .CK(clk), .Q(
        \adder_stage3[1][1] ) );
  DFF_X1 \adder_stage3_reg[1][2]  ( .D(n9648), .CK(clk), .Q(
        \adder_stage3[1][2] ) );
  DFF_X1 \adder_stage3_reg[1][3]  ( .D(n9647), .CK(clk), .Q(
        \adder_stage3[1][3] ) );
  DFF_X1 \adder_stage3_reg[1][4]  ( .D(n9646), .CK(clk), .Q(
        \adder_stage3[1][4] ) );
  DFF_X1 \adder_stage3_reg[1][5]  ( .D(n9645), .CK(clk), .Q(
        \adder_stage3[1][5] ) );
  DFF_X1 \adder_stage3_reg[1][6]  ( .D(n9644), .CK(clk), .Q(
        \adder_stage3[1][6] ) );
  DFF_X1 \adder_stage3_reg[1][7]  ( .D(n9643), .CK(clk), .Q(
        \adder_stage3[1][7] ) );
  DFF_X1 \adder_stage3_reg[1][8]  ( .D(n9642), .CK(clk), .Q(
        \adder_stage3[1][8] ) );
  DFF_X1 \adder_stage3_reg[1][9]  ( .D(n9641), .CK(clk), .Q(
        \adder_stage3[1][9] ) );
  DFF_X1 \adder_stage3_reg[1][10]  ( .D(n9640), .CK(clk), .Q(
        \adder_stage3[1][10] ) );
  DFF_X1 \adder_stage3_reg[1][12]  ( .D(n9638), .CK(clk), .Q(
        \adder_stage3[1][12] ) );
  DFF_X1 \adder_stage3_reg[1][13]  ( .D(n9637), .CK(clk), .Q(
        \adder_stage3[1][13] ) );
  DFF_X1 \adder_stage3_reg[1][14]  ( .D(n9636), .CK(clk), .Q(
        \adder_stage3[1][14] ) );
  DFF_X1 \adder_stage3_reg[1][15]  ( .D(n9635), .CK(clk), .Q(
        \adder_stage3[1][15] ) );
  DFF_X1 \adder_stage3_reg[1][16]  ( .D(n9634), .CK(clk), .Q(
        \adder_stage3[1][16] ) );
  DFF_X1 \adder_stage3_reg[1][17]  ( .D(n9633), .CK(clk), .Q(
        \adder_stage3[1][17] ) );
  DFF_X1 \adder_stage3_reg[1][18]  ( .D(n9632), .CK(clk), .Q(
        \adder_stage3[1][18] ) );
  DFF_X1 \adder_stage3_reg[1][19]  ( .D(n9631), .CK(clk), .Q(
        \adder_stage3[1][19] ) );
  DFF_X1 \adder_stage3_reg[1][20]  ( .D(n9630), .CK(clk), .Q(
        \adder_stage3[1][20] ) );
  DFF_X1 \adder_stage3_reg[2][0]  ( .D(n9629), .CK(clk), .Q(
        \adder_stage3[2][0] ) );
  DFF_X1 \adder_stage3_reg[2][1]  ( .D(n9628), .CK(clk), .Q(
        \adder_stage3[2][1] ) );
  DFF_X1 \adder_stage3_reg[2][2]  ( .D(n9627), .CK(clk), .Q(
        \adder_stage3[2][2] ) );
  DFF_X1 \adder_stage3_reg[2][3]  ( .D(n9626), .CK(clk), .Q(
        \adder_stage3[2][3] ) );
  DFF_X1 \adder_stage3_reg[2][4]  ( .D(n9625), .CK(clk), .Q(
        \adder_stage3[2][4] ) );
  DFF_X1 \adder_stage3_reg[2][5]  ( .D(n9624), .CK(clk), .Q(
        \adder_stage3[2][5] ) );
  DFF_X1 \adder_stage3_reg[2][6]  ( .D(n9623), .CK(clk), .Q(
        \adder_stage3[2][6] ) );
  DFF_X1 \adder_stage3_reg[2][7]  ( .D(n9622), .CK(clk), .Q(
        \adder_stage3[2][7] ) );
  DFF_X1 \adder_stage3_reg[2][8]  ( .D(n9621), .CK(clk), .Q(
        \adder_stage3[2][8] ) );
  DFF_X1 \adder_stage3_reg[2][9]  ( .D(n9620), .CK(clk), .Q(
        \adder_stage3[2][9] ) );
  DFF_X1 \adder_stage3_reg[2][10]  ( .D(n9619), .CK(clk), .Q(
        \adder_stage3[2][10] ) );
  DFF_X1 \adder_stage3_reg[2][11]  ( .D(n9618), .CK(clk), .Q(
        \adder_stage3[2][11] ) );
  DFF_X1 \adder_stage3_reg[2][12]  ( .D(n9617), .CK(clk), .Q(
        \adder_stage3[2][12] ) );
  DFF_X1 \adder_stage3_reg[2][13]  ( .D(n9616), .CK(clk), .Q(
        \adder_stage3[2][13] ) );
  DFF_X1 \adder_stage3_reg[2][14]  ( .D(n9615), .CK(clk), .Q(
        \adder_stage3[2][14] ) );
  DFF_X1 \adder_stage3_reg[2][15]  ( .D(n9614), .CK(clk), .Q(
        \adder_stage3[2][15] ) );
  DFF_X1 \adder_stage3_reg[2][16]  ( .D(n9613), .CK(clk), .Q(
        \adder_stage3[2][16] ) );
  DFF_X1 \adder_stage3_reg[2][17]  ( .D(n9612), .CK(clk), .Q(
        \adder_stage3[2][17] ) );
  DFF_X1 \adder_stage3_reg[2][18]  ( .D(n9611), .CK(clk), .Q(
        \adder_stage3[2][18] ) );
  DFF_X1 \adder_stage3_reg[2][19]  ( .D(n9610), .CK(clk), .Q(
        \adder_stage3[2][19] ) );
  DFF_X1 \adder_stage3_reg[2][20]  ( .D(n8182), .CK(clk), .Q(
        \adder_stage3[2][20] ) );
  DFF_X1 \adder_stage3_reg[3][0]  ( .D(n9609), .CK(clk), .Q(
        \adder_stage3[3][0] ) );
  DFF_X1 \adder_stage3_reg[3][1]  ( .D(n9608), .CK(clk), .Q(
        \adder_stage3[3][1] ) );
  DFF_X1 \adder_stage3_reg[3][2]  ( .D(n9607), .CK(clk), .Q(
        \adder_stage3[3][2] ) );
  DFF_X1 \adder_stage3_reg[3][3]  ( .D(n9606), .CK(clk), .Q(
        \adder_stage3[3][3] ) );
  DFF_X1 \adder_stage3_reg[3][4]  ( .D(n9605), .CK(clk), .Q(
        \adder_stage3[3][4] ) );
  DFF_X1 \adder_stage3_reg[3][5]  ( .D(n9604), .CK(clk), .Q(
        \adder_stage3[3][5] ) );
  DFF_X1 \adder_stage3_reg[3][6]  ( .D(n9603), .CK(clk), .Q(
        \adder_stage3[3][6] ) );
  DFF_X1 \adder_stage3_reg[3][7]  ( .D(n9602), .CK(clk), .Q(
        \adder_stage3[3][7] ) );
  DFF_X1 \adder_stage3_reg[3][8]  ( .D(n9601), .CK(clk), .Q(
        \adder_stage3[3][8] ) );
  DFF_X1 \adder_stage3_reg[3][9]  ( .D(n9600), .CK(clk), .Q(
        \adder_stage3[3][9] ) );
  DFF_X1 \adder_stage3_reg[3][10]  ( .D(n9599), .CK(clk), .Q(
        \adder_stage3[3][10] ) );
  DFF_X1 \adder_stage3_reg[3][11]  ( .D(n9598), .CK(clk), .Q(
        \adder_stage3[3][11] ) );
  DFF_X1 \adder_stage3_reg[3][12]  ( .D(n9597), .CK(clk), .Q(
        \adder_stage3[3][12] ) );
  DFF_X1 \adder_stage3_reg[3][13]  ( .D(n9596), .CK(clk), .Q(
        \adder_stage3[3][13] ) );
  DFF_X1 \adder_stage3_reg[3][14]  ( .D(n9595), .CK(clk), .Q(
        \adder_stage3[3][14] ) );
  DFF_X1 \adder_stage3_reg[3][15]  ( .D(n9594), .CK(clk), .Q(
        \adder_stage3[3][15] ) );
  DFF_X1 \adder_stage3_reg[3][16]  ( .D(n9593), .CK(clk), .Q(
        \adder_stage3[3][16] ) );
  DFF_X1 \adder_stage3_reg[3][17]  ( .D(n9592), .CK(clk), .Q(
        \adder_stage3[3][17] ) );
  DFF_X1 \adder_stage3_reg[3][18]  ( .D(n9591), .CK(clk), .Q(
        \adder_stage3[3][18] ) );
  DFF_X1 \adder_stage3_reg[3][19]  ( .D(n9590), .CK(clk), .Q(
        \adder_stage3[3][19] ) );
  DFF_X1 \adder_stage3_reg[3][20]  ( .D(n9589), .CK(clk), .Q(
        \adder_stage3[3][20] ) );
  DFF_X1 \adder_stage4_reg[0][0]  ( .D(n9588), .CK(clk), .Q(
        \adder_stage4[0][0] ) );
  DFF_X1 \adder_stage4_reg[0][1]  ( .D(n9587), .CK(clk), .Q(
        \adder_stage4[0][1] ) );
  DFF_X1 \adder_stage4_reg[0][2]  ( .D(n9586), .CK(clk), .Q(
        \adder_stage4[0][2] ) );
  DFF_X1 \adder_stage4_reg[0][3]  ( .D(n9585), .CK(clk), .Q(
        \adder_stage4[0][3] ) );
  DFF_X1 \adder_stage4_reg[0][4]  ( .D(n9584), .CK(clk), .Q(
        \adder_stage4[0][4] ) );
  DFF_X1 \adder_stage4_reg[0][5]  ( .D(n9583), .CK(clk), .Q(
        \adder_stage4[0][5] ) );
  DFF_X1 \adder_stage4_reg[0][6]  ( .D(n9582), .CK(clk), .Q(
        \adder_stage4[0][6] ) );
  DFF_X1 \adder_stage4_reg[0][7]  ( .D(n9581), .CK(clk), .Q(
        \adder_stage4[0][7] ) );
  DFF_X1 \adder_stage4_reg[0][8]  ( .D(n9580), .CK(clk), .Q(
        \adder_stage4[0][8] ) );
  DFF_X1 \adder_stage4_reg[0][9]  ( .D(n9579), .CK(clk), .Q(
        \adder_stage4[0][9] ) );
  DFF_X1 \adder_stage4_reg[0][10]  ( .D(n9578), .CK(clk), .Q(
        \adder_stage4[0][10] ) );
  DFF_X1 \adder_stage4_reg[0][11]  ( .D(n9577), .CK(clk), .Q(
        \adder_stage4[0][11] ) );
  DFF_X1 \adder_stage4_reg[0][12]  ( .D(n9576), .CK(clk), .Q(
        \adder_stage4[0][12] ) );
  DFF_X1 \adder_stage4_reg[0][13]  ( .D(n9575), .CK(clk), .Q(
        \adder_stage4[0][13] ) );
  DFF_X1 \adder_stage4_reg[0][14]  ( .D(n9574), .CK(clk), .Q(
        \adder_stage4[0][14] ) );
  DFF_X1 \adder_stage4_reg[0][15]  ( .D(n9573), .CK(clk), .Q(
        \adder_stage4[0][15] ) );
  DFF_X1 \adder_stage4_reg[0][16]  ( .D(n9572), .CK(clk), .Q(
        \adder_stage4[0][16] ) );
  DFF_X1 \adder_stage4_reg[0][17]  ( .D(n9571), .CK(clk), .Q(
        \adder_stage4[0][17] ) );
  DFF_X1 \adder_stage4_reg[0][18]  ( .D(n9570), .CK(clk), .Q(
        \adder_stage4[0][18] ) );
  DFF_X1 \adder_stage4_reg[0][19]  ( .D(n9569), .CK(clk), .Q(
        \adder_stage4[0][19] ) );
  DFF_X1 \adder_stage4_reg[0][20]  ( .D(n9568), .CK(clk), .Q(
        \adder_stage4[0][20] ) );
  DFF_X1 \adder_stage4_reg[1][0]  ( .D(n9567), .CK(clk), .Q(
        \adder_stage4[1][0] ) );
  DFF_X1 \adder_stage4_reg[1][1]  ( .D(n9566), .CK(clk), .Q(
        \adder_stage4[1][1] ) );
  DFF_X1 \adder_stage4_reg[1][2]  ( .D(n9565), .CK(clk), .Q(
        \adder_stage4[1][2] ) );
  DFF_X1 \adder_stage4_reg[1][3]  ( .D(n9564), .CK(clk), .Q(
        \adder_stage4[1][3] ) );
  DFF_X1 \adder_stage4_reg[1][4]  ( .D(n9563), .CK(clk), .Q(
        \adder_stage4[1][4] ) );
  DFF_X1 \adder_stage4_reg[1][5]  ( .D(n9562), .CK(clk), .Q(
        \adder_stage4[1][5] ) );
  DFF_X1 \adder_stage4_reg[1][6]  ( .D(n9561), .CK(clk), .Q(
        \adder_stage4[1][6] ) );
  DFF_X1 \adder_stage4_reg[1][7]  ( .D(n9560), .CK(clk), .Q(
        \adder_stage4[1][7] ) );
  DFF_X1 \adder_stage4_reg[1][8]  ( .D(n9559), .CK(clk), .Q(
        \adder_stage4[1][8] ) );
  DFF_X1 \adder_stage4_reg[1][9]  ( .D(n9558), .CK(clk), .Q(
        \adder_stage4[1][9] ) );
  DFF_X1 \adder_stage4_reg[1][10]  ( .D(n9557), .CK(clk), .Q(
        \adder_stage4[1][10] ) );
  DFF_X1 \adder_stage4_reg[1][11]  ( .D(n9556), .CK(clk), .Q(
        \adder_stage4[1][11] ) );
  DFF_X1 \adder_stage4_reg[1][12]  ( .D(n9555), .CK(clk), .Q(
        \adder_stage4[1][12] ) );
  DFF_X1 \adder_stage4_reg[1][13]  ( .D(n9554), .CK(clk), .Q(
        \adder_stage4[1][13] ) );
  DFF_X1 \adder_stage4_reg[1][14]  ( .D(n9553), .CK(clk), .Q(
        \adder_stage4[1][14] ) );
  DFF_X1 \adder_stage4_reg[1][15]  ( .D(n9552), .CK(clk), .Q(
        \adder_stage4[1][15] ) );
  DFF_X1 \adder_stage4_reg[1][16]  ( .D(n9551), .CK(clk), .Q(
        \adder_stage4[1][16] ) );
  DFF_X1 \adder_stage4_reg[1][17]  ( .D(n9550), .CK(clk), .Q(
        \adder_stage4[1][17] ) );
  DFF_X1 \adder_stage4_reg[1][18]  ( .D(n9549), .CK(clk), .Q(
        \adder_stage4[1][18] ) );
  DFF_X1 \adder_stage4_reg[1][19]  ( .D(n9548), .CK(clk), .Q(
        \adder_stage4[1][19] ) );
  DFF_X1 \adder_stage4_reg[1][20]  ( .D(n9547), .CK(clk), .Q(
        \adder_stage4[1][20] ) );
  conv_128_32_DW_mult_pipe_J1_0 \multiplier[31].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8913), .tc(1'b1), .a({\xmem_data[31][7] , 
        \xmem_data[31][6] , \xmem_data[31][5] , \xmem_data[31][4] , 
        \xmem_data[31][3] , \xmem_data[31][2] , \xmem_data[31][1] , 
        \xmem_data[31][0] }), .b({\fmem_data[31][7] , \fmem_data[31][6] , 
        \fmem_data[31][5] , \fmem_data[31][4] , \fmem_data[31][3] , 
        \fmem_data[31][2] , \fmem_data[31][1] , \fmem_data[31][0] }), 
        .product({\x_mult_f_int[31][15] , \x_mult_f_int[31][14] , 
        \x_mult_f_int[31][13] , \x_mult_f_int[31][12] , \x_mult_f_int[31][11] , 
        \x_mult_f_int[31][10] , \x_mult_f_int[31][9] , \x_mult_f_int[31][8] , 
        \x_mult_f_int[31][7] , \x_mult_f_int[31][6] , \x_mult_f_int[31][5] , 
        \x_mult_f_int[31][4] , \x_mult_f_int[31][3] , \x_mult_f_int[31][2] , 
        \x_mult_f_int[31][1] , \x_mult_f_int[31][0] }) );
  conv_128_32_DW_mult_pipe_J1_1 \multiplier[30].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n3443), .tc(1'b1), .a({\xmem_data[30][7] , 
        \xmem_data[30][6] , \xmem_data[30][5] , \xmem_data[30][4] , 
        \xmem_data[30][3] , \xmem_data[30][2] , \xmem_data[30][1] , 
        \xmem_data[30][0] }), .b({\fmem_data[30][7] , \fmem_data[30][6] , 
        \fmem_data[30][5] , \fmem_data[30][4] , \fmem_data[30][3] , 
        \fmem_data[30][2] , \fmem_data[30][1] , \fmem_data[30][0] }), 
        .product({\x_mult_f_int[30][15] , \x_mult_f_int[30][14] , 
        \x_mult_f_int[30][13] , \x_mult_f_int[30][12] , \x_mult_f_int[30][11] , 
        \x_mult_f_int[30][10] , \x_mult_f_int[30][9] , \x_mult_f_int[30][8] , 
        \x_mult_f_int[30][7] , \x_mult_f_int[30][6] , \x_mult_f_int[30][5] , 
        \x_mult_f_int[30][4] , \x_mult_f_int[30][3] , \x_mult_f_int[30][2] , 
        \x_mult_f_int[30][1] , \x_mult_f_int[30][0] }) );
  conv_128_32_DW_mult_pipe_J1_2 \multiplier[29].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8915), .tc(1'b1), .a({\xmem_data[29][7] , 
        \xmem_data[29][6] , \xmem_data[29][5] , \xmem_data[29][4] , 
        \xmem_data[29][3] , \xmem_data[29][2] , \xmem_data[29][1] , 
        \xmem_data[29][0] }), .b({\fmem_data[29][7] , \fmem_data[29][6] , 
        \fmem_data[29][5] , \fmem_data[29][4] , \fmem_data[29][3] , 
        \fmem_data[29][2] , \fmem_data[29][1] , \fmem_data[29][0] }), 
        .product({\x_mult_f_int[29][15] , \x_mult_f_int[29][14] , 
        \x_mult_f_int[29][13] , \x_mult_f_int[29][12] , \x_mult_f_int[29][11] , 
        \x_mult_f_int[29][10] , \x_mult_f_int[29][9] , \x_mult_f_int[29][8] , 
        \x_mult_f_int[29][7] , \x_mult_f_int[29][6] , \x_mult_f_int[29][5] , 
        \x_mult_f_int[29][4] , \x_mult_f_int[29][3] , \x_mult_f_int[29][2] , 
        \x_mult_f_int[29][1] , \x_mult_f_int[29][0] }) );
  conv_128_32_DW_mult_pipe_J1_3 \multiplier[28].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8917), .tc(1'b1), .a({\xmem_data[28][7] , 
        \xmem_data[28][6] , \xmem_data[28][5] , \xmem_data[28][4] , 
        \xmem_data[28][3] , \xmem_data[28][2] , \xmem_data[28][1] , 
        \xmem_data[28][0] }), .b({\fmem_data[28][7] , \fmem_data[28][6] , 
        \fmem_data[28][5] , \fmem_data[28][4] , \fmem_data[28][3] , 
        \fmem_data[28][2] , \fmem_data[28][1] , \fmem_data[28][0] }), 
        .product({\x_mult_f_int[28][15] , \x_mult_f_int[28][14] , 
        \x_mult_f_int[28][13] , \x_mult_f_int[28][12] , \x_mult_f_int[28][11] , 
        \x_mult_f_int[28][10] , \x_mult_f_int[28][9] , \x_mult_f_int[28][8] , 
        \x_mult_f_int[28][7] , \x_mult_f_int[28][6] , \x_mult_f_int[28][5] , 
        \x_mult_f_int[28][4] , \x_mult_f_int[28][3] , \x_mult_f_int[28][2] , 
        \x_mult_f_int[28][1] , \x_mult_f_int[28][0] }) );
  conv_128_32_DW_mult_pipe_J1_4 \multiplier[27].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8913), .tc(1'b1), .a({\xmem_data[27][7] , 
        \xmem_data[27][6] , \xmem_data[27][5] , \xmem_data[27][4] , 
        \xmem_data[27][3] , \xmem_data[27][2] , \xmem_data[27][1] , 
        \xmem_data[27][0] }), .b({\fmem_data[27][7] , \fmem_data[27][6] , 
        \fmem_data[27][5] , \fmem_data[27][4] , \fmem_data[27][3] , 
        \fmem_data[27][2] , \fmem_data[27][1] , \fmem_data[27][0] }), 
        .product({\x_mult_f_int[27][15] , \x_mult_f_int[27][14] , 
        \x_mult_f_int[27][13] , \x_mult_f_int[27][12] , \x_mult_f_int[27][11] , 
        \x_mult_f_int[27][10] , \x_mult_f_int[27][9] , \x_mult_f_int[27][8] , 
        \x_mult_f_int[27][7] , \x_mult_f_int[27][6] , \x_mult_f_int[27][5] , 
        \x_mult_f_int[27][4] , \x_mult_f_int[27][3] , \x_mult_f_int[27][2] , 
        \x_mult_f_int[27][1] , \x_mult_f_int[27][0] }) );
  conv_128_32_DW_mult_pipe_J1_5 \multiplier[26].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8923), .tc(1'b1), .a({\xmem_data[26][7] , 
        \xmem_data[26][6] , \xmem_data[26][5] , \xmem_data[26][4] , 
        \xmem_data[26][3] , \xmem_data[26][2] , \xmem_data[26][1] , 
        \xmem_data[26][0] }), .b({\fmem_data[26][7] , \fmem_data[26][6] , 
        \fmem_data[26][5] , \fmem_data[26][4] , \fmem_data[26][3] , 
        \fmem_data[26][2] , \fmem_data[26][1] , \fmem_data[26][0] }), 
        .product({\x_mult_f_int[26][15] , \x_mult_f_int[26][14] , 
        \x_mult_f_int[26][13] , \x_mult_f_int[26][12] , \x_mult_f_int[26][11] , 
        \x_mult_f_int[26][10] , \x_mult_f_int[26][9] , \x_mult_f_int[26][8] , 
        \x_mult_f_int[26][7] , \x_mult_f_int[26][6] , \x_mult_f_int[26][5] , 
        \x_mult_f_int[26][4] , \x_mult_f_int[26][3] , \x_mult_f_int[26][2] , 
        \x_mult_f_int[26][1] , \x_mult_f_int[26][0] }) );
  conv_128_32_DW_mult_pipe_J1_6 \multiplier[25].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3449), .en(n8913), .tc(1'b1), .a({\xmem_data[25][7] , 
        \xmem_data[25][6] , \xmem_data[25][5] , \xmem_data[25][4] , 
        \xmem_data[25][3] , \xmem_data[25][2] , \xmem_data[25][1] , 
        \xmem_data[25][0] }), .b({\fmem_data[25][7] , \fmem_data[25][6] , 
        \fmem_data[25][5] , \fmem_data[25][4] , \fmem_data[25][3] , 
        \fmem_data[25][2] , \fmem_data[25][1] , \fmem_data[25][0] }), 
        .product({\x_mult_f_int[25][15] , \x_mult_f_int[25][14] , 
        \x_mult_f_int[25][13] , \x_mult_f_int[25][12] , \x_mult_f_int[25][11] , 
        \x_mult_f_int[25][10] , \x_mult_f_int[25][9] , \x_mult_f_int[25][8] , 
        \x_mult_f_int[25][7] , \x_mult_f_int[25][6] , \x_mult_f_int[25][5] , 
        \x_mult_f_int[25][4] , \x_mult_f_int[25][3] , \x_mult_f_int[25][2] , 
        \x_mult_f_int[25][1] , \x_mult_f_int[25][0] }) );
  conv_128_32_DW_mult_pipe_J1_7 \multiplier[24].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8915), .tc(1'b1), .a({\xmem_data[24][7] , 
        \xmem_data[24][6] , \xmem_data[24][5] , \xmem_data[24][4] , 
        \xmem_data[24][3] , \xmem_data[24][2] , \xmem_data[24][1] , 
        \xmem_data[24][0] }), .b({\fmem_data[24][7] , \fmem_data[24][6] , 
        \fmem_data[24][5] , \fmem_data[24][4] , \fmem_data[24][3] , 
        \fmem_data[24][2] , \fmem_data[24][1] , \fmem_data[24][0] }), 
        .product({\x_mult_f_int[24][15] , \x_mult_f_int[24][14] , 
        \x_mult_f_int[24][13] , \x_mult_f_int[24][12] , \x_mult_f_int[24][11] , 
        \x_mult_f_int[24][10] , \x_mult_f_int[24][9] , \x_mult_f_int[24][8] , 
        \x_mult_f_int[24][7] , \x_mult_f_int[24][6] , \x_mult_f_int[24][5] , 
        \x_mult_f_int[24][4] , \x_mult_f_int[24][3] , \x_mult_f_int[24][2] , 
        \x_mult_f_int[24][1] , \x_mult_f_int[24][0] }) );
  conv_128_32_DW_mult_pipe_J1_8 \multiplier[23].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8922), .tc(1'b1), .a({\xmem_data[23][7] , 
        \xmem_data[23][6] , \xmem_data[23][5] , \xmem_data[23][4] , 
        \xmem_data[23][3] , \xmem_data[23][2] , \xmem_data[23][1] , 
        \xmem_data[23][0] }), .b({\fmem_data[23][7] , \fmem_data[23][6] , 
        \fmem_data[23][5] , \fmem_data[23][4] , \fmem_data[23][3] , 
        \fmem_data[23][2] , \fmem_data[23][1] , \fmem_data[23][0] }), 
        .product({\x_mult_f_int[23][15] , \x_mult_f_int[23][14] , 
        \x_mult_f_int[23][13] , \x_mult_f_int[23][12] , \x_mult_f_int[23][11] , 
        \x_mult_f_int[23][10] , \x_mult_f_int[23][9] , \x_mult_f_int[23][8] , 
        \x_mult_f_int[23][7] , \x_mult_f_int[23][6] , \x_mult_f_int[23][5] , 
        \x_mult_f_int[23][4] , \x_mult_f_int[23][3] , \x_mult_f_int[23][2] , 
        \x_mult_f_int[23][1] , \x_mult_f_int[23][0] }) );
  conv_128_32_DW_mult_pipe_J1_9 \multiplier[22].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8916), .tc(1'b1), .a({\xmem_data[22][7] , 
        \xmem_data[22][6] , \xmem_data[22][5] , \xmem_data[22][4] , 
        \xmem_data[22][3] , \xmem_data[22][2] , \xmem_data[22][1] , 
        \xmem_data[22][0] }), .b({\fmem_data[22][7] , \fmem_data[22][6] , 
        \fmem_data[22][5] , \fmem_data[22][4] , \fmem_data[22][3] , 
        \fmem_data[22][2] , \fmem_data[22][1] , \fmem_data[22][0] }), 
        .product({\x_mult_f_int[22][15] , \x_mult_f_int[22][14] , 
        \x_mult_f_int[22][13] , \x_mult_f_int[22][12] , \x_mult_f_int[22][11] , 
        \x_mult_f_int[22][10] , \x_mult_f_int[22][9] , \x_mult_f_int[22][8] , 
        \x_mult_f_int[22][7] , \x_mult_f_int[22][6] , \x_mult_f_int[22][5] , 
        \x_mult_f_int[22][4] , \x_mult_f_int[22][3] , \x_mult_f_int[22][2] , 
        \x_mult_f_int[22][1] , \x_mult_f_int[22][0] }) );
  conv_128_32_DW_mult_pipe_J1_10 \multiplier[21].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8913), .tc(1'b1), .a({\xmem_data[21][7] , 
        \xmem_data[21][6] , \xmem_data[21][5] , \xmem_data[21][4] , 
        \xmem_data[21][3] , \xmem_data[21][2] , \xmem_data[21][1] , 
        \xmem_data[21][0] }), .b({\fmem_data[21][7] , \fmem_data[21][6] , 
        \fmem_data[21][5] , \fmem_data[21][4] , \fmem_data[21][3] , 
        \fmem_data[21][2] , \fmem_data[21][1] , \fmem_data[21][0] }), 
        .product({\x_mult_f_int[21][15] , \x_mult_f_int[21][14] , 
        \x_mult_f_int[21][13] , \x_mult_f_int[21][12] , \x_mult_f_int[21][11] , 
        \x_mult_f_int[21][10] , \x_mult_f_int[21][9] , \x_mult_f_int[21][8] , 
        \x_mult_f_int[21][7] , \x_mult_f_int[21][6] , \x_mult_f_int[21][5] , 
        \x_mult_f_int[21][4] , \x_mult_f_int[21][3] , \x_mult_f_int[21][2] , 
        \x_mult_f_int[21][1] , \x_mult_f_int[21][0] }) );
  conv_128_32_DW_mult_pipe_J1_11 \multiplier[20].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n3430), .tc(1'b1), .a({\xmem_data[20][7] , 
        \xmem_data[20][6] , \xmem_data[20][5] , \xmem_data[20][4] , 
        \xmem_data[20][3] , \xmem_data[20][2] , \xmem_data[20][1] , 
        \xmem_data[20][0] }), .b({\fmem_data[20][7] , \fmem_data[20][6] , 
        \fmem_data[20][5] , \fmem_data[20][4] , \fmem_data[20][3] , 
        \fmem_data[20][2] , \fmem_data[20][1] , \fmem_data[20][0] }), 
        .product({\x_mult_f_int[20][15] , \x_mult_f_int[20][14] , 
        \x_mult_f_int[20][13] , \x_mult_f_int[20][12] , \x_mult_f_int[20][11] , 
        \x_mult_f_int[20][10] , \x_mult_f_int[20][9] , \x_mult_f_int[20][8] , 
        \x_mult_f_int[20][7] , \x_mult_f_int[20][6] , \x_mult_f_int[20][5] , 
        \x_mult_f_int[20][4] , \x_mult_f_int[20][3] , \x_mult_f_int[20][2] , 
        \x_mult_f_int[20][1] , \x_mult_f_int[20][0] }) );
  conv_128_32_DW_mult_pipe_J1_12 \multiplier[19].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8921), .tc(1'b1), .a({\xmem_data[19][7] , 
        \xmem_data[19][6] , \xmem_data[19][5] , \xmem_data[19][4] , 
        \xmem_data[19][3] , \xmem_data[19][2] , \xmem_data[19][1] , 
        \xmem_data[19][0] }), .b({\fmem_data[19][7] , \fmem_data[19][6] , 
        \fmem_data[19][5] , \fmem_data[19][4] , \fmem_data[19][3] , 
        \fmem_data[19][2] , \fmem_data[19][1] , \fmem_data[19][0] }), 
        .product({\x_mult_f_int[19][15] , \x_mult_f_int[19][14] , 
        \x_mult_f_int[19][13] , \x_mult_f_int[19][12] , \x_mult_f_int[19][11] , 
        \x_mult_f_int[19][10] , \x_mult_f_int[19][9] , \x_mult_f_int[19][8] , 
        \x_mult_f_int[19][7] , \x_mult_f_int[19][6] , \x_mult_f_int[19][5] , 
        \x_mult_f_int[19][4] , \x_mult_f_int[19][3] , \x_mult_f_int[19][2] , 
        \x_mult_f_int[19][1] , \x_mult_f_int[19][0] }) );
  conv_128_32_DW_mult_pipe_J1_13 \multiplier[18].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8914), .tc(1'b1), .a({\xmem_data[18][7] , 
        \xmem_data[18][6] , \xmem_data[18][5] , \xmem_data[18][4] , 
        \xmem_data[18][3] , \xmem_data[18][2] , \xmem_data[18][1] , 
        \xmem_data[18][0] }), .b({\fmem_data[18][7] , \fmem_data[18][6] , 
        \fmem_data[18][5] , \fmem_data[18][4] , \fmem_data[18][3] , 
        \fmem_data[18][2] , \fmem_data[18][1] , \fmem_data[18][0] }), 
        .product({\x_mult_f_int[18][15] , \x_mult_f_int[18][14] , 
        \x_mult_f_int[18][13] , \x_mult_f_int[18][12] , \x_mult_f_int[18][11] , 
        \x_mult_f_int[18][10] , \x_mult_f_int[18][9] , \x_mult_f_int[18][8] , 
        \x_mult_f_int[18][7] , \x_mult_f_int[18][6] , \x_mult_f_int[18][5] , 
        \x_mult_f_int[18][4] , \x_mult_f_int[18][3] , \x_mult_f_int[18][2] , 
        \x_mult_f_int[18][1] , \x_mult_f_int[18][0] }) );
  conv_128_32_DW_mult_pipe_J1_14 \multiplier[17].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8921), .tc(1'b1), .a({\xmem_data[17][7] , 
        \xmem_data[17][6] , \xmem_data[17][5] , \xmem_data[17][4] , 
        \xmem_data[17][3] , \xmem_data[17][2] , \xmem_data[17][1] , 
        \xmem_data[17][0] }), .b({\fmem_data[17][7] , \fmem_data[17][6] , 
        \fmem_data[17][5] , \fmem_data[17][4] , \fmem_data[17][3] , 
        \fmem_data[17][2] , \fmem_data[17][1] , \fmem_data[17][0] }), 
        .product({\x_mult_f_int[17][15] , \x_mult_f_int[17][14] , 
        \x_mult_f_int[17][13] , \x_mult_f_int[17][12] , \x_mult_f_int[17][11] , 
        \x_mult_f_int[17][10] , \x_mult_f_int[17][9] , \x_mult_f_int[17][8] , 
        \x_mult_f_int[17][7] , \x_mult_f_int[17][6] , \x_mult_f_int[17][5] , 
        \x_mult_f_int[17][4] , \x_mult_f_int[17][3] , \x_mult_f_int[17][2] , 
        \x_mult_f_int[17][1] , \x_mult_f_int[17][0] }) );
  conv_128_32_DW_mult_pipe_J1_15 \multiplier[16].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8914), .tc(1'b1), .a({\xmem_data[16][7] , 
        \xmem_data[16][6] , \xmem_data[16][5] , \xmem_data[16][4] , 
        \xmem_data[16][3] , \xmem_data[16][2] , \xmem_data[16][1] , 
        \xmem_data[16][0] }), .b({\fmem_data[16][7] , \fmem_data[16][6] , 
        \fmem_data[16][5] , \fmem_data[16][4] , \fmem_data[16][3] , 
        \fmem_data[16][2] , \fmem_data[16][1] , \fmem_data[16][0] }), 
        .product({\x_mult_f_int[16][15] , \x_mult_f_int[16][14] , 
        \x_mult_f_int[16][13] , \x_mult_f_int[16][12] , \x_mult_f_int[16][11] , 
        \x_mult_f_int[16][10] , \x_mult_f_int[16][9] , \x_mult_f_int[16][8] , 
        \x_mult_f_int[16][7] , \x_mult_f_int[16][6] , \x_mult_f_int[16][5] , 
        \x_mult_f_int[16][4] , \x_mult_f_int[16][3] , \x_mult_f_int[16][2] , 
        \x_mult_f_int[16][1] , \x_mult_f_int[16][0] }) );
  conv_128_32_DW_mult_pipe_J1_16 \multiplier[15].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8922), .tc(1'b1), .a({\xmem_data[15][7] , 
        \xmem_data[15][6] , \xmem_data[15][5] , \xmem_data[15][4] , 
        \xmem_data[15][3] , \xmem_data[15][2] , \xmem_data[15][1] , 
        \xmem_data[15][0] }), .b({\fmem_data[15][7] , \fmem_data[15][6] , 
        \fmem_data[15][5] , \fmem_data[15][4] , \fmem_data[15][3] , 
        \fmem_data[15][2] , \fmem_data[15][1] , \fmem_data[15][0] }), 
        .product({\x_mult_f_int[15][15] , \x_mult_f_int[15][14] , 
        \x_mult_f_int[15][13] , \x_mult_f_int[15][12] , \x_mult_f_int[15][11] , 
        \x_mult_f_int[15][10] , \x_mult_f_int[15][9] , \x_mult_f_int[15][8] , 
        \x_mult_f_int[15][7] , \x_mult_f_int[15][6] , \x_mult_f_int[15][5] , 
        \x_mult_f_int[15][4] , \x_mult_f_int[15][3] , \x_mult_f_int[15][2] , 
        \x_mult_f_int[15][1] , \x_mult_f_int[15][0] }) );
  conv_128_32_DW_mult_pipe_J1_17 \multiplier[14].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3449), .en(n8917), .tc(1'b1), .a({\xmem_data[14][7] , 
        \xmem_data[14][6] , \xmem_data[14][5] , \xmem_data[14][4] , 
        \xmem_data[14][3] , \xmem_data[14][2] , \xmem_data[14][1] , 
        \xmem_data[14][0] }), .b({\fmem_data[14][7] , \fmem_data[14][6] , 
        \fmem_data[14][5] , \fmem_data[14][4] , \fmem_data[14][3] , 
        \fmem_data[14][2] , \fmem_data[14][1] , \fmem_data[14][0] }), 
        .product({\x_mult_f_int[14][15] , \x_mult_f_int[14][14] , 
        \x_mult_f_int[14][13] , \x_mult_f_int[14][12] , \x_mult_f_int[14][11] , 
        \x_mult_f_int[14][10] , \x_mult_f_int[14][9] , \x_mult_f_int[14][8] , 
        \x_mult_f_int[14][7] , \x_mult_f_int[14][6] , \x_mult_f_int[14][5] , 
        \x_mult_f_int[14][4] , \x_mult_f_int[14][3] , \x_mult_f_int[14][2] , 
        \x_mult_f_int[14][1] , \x_mult_f_int[14][0] }) );
  conv_128_32_DW_mult_pipe_J1_18 \multiplier[13].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8914), .tc(1'b1), .a({\xmem_data[13][7] , 
        \xmem_data[13][6] , \xmem_data[13][5] , \xmem_data[13][4] , 
        \xmem_data[13][3] , \xmem_data[13][2] , \xmem_data[13][1] , 
        \xmem_data[13][0] }), .b({\fmem_data[13][7] , \fmem_data[13][6] , 
        \fmem_data[13][5] , \fmem_data[13][4] , \fmem_data[13][3] , 
        \fmem_data[13][2] , \fmem_data[13][1] , \fmem_data[13][0] }), 
        .product({\x_mult_f_int[13][15] , \x_mult_f_int[13][14] , 
        \x_mult_f_int[13][13] , \x_mult_f_int[13][12] , \x_mult_f_int[13][11] , 
        \x_mult_f_int[13][10] , \x_mult_f_int[13][9] , \x_mult_f_int[13][8] , 
        \x_mult_f_int[13][7] , \x_mult_f_int[13][6] , \x_mult_f_int[13][5] , 
        \x_mult_f_int[13][4] , \x_mult_f_int[13][3] , \x_mult_f_int[13][2] , 
        \x_mult_f_int[13][1] , \x_mult_f_int[13][0] }) );
  conv_128_32_DW_mult_pipe_J1_19 \multiplier[12].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8918), .en(n8922), .tc(1'b1), .a({\xmem_data[12][7] , 
        \xmem_data[12][6] , \xmem_data[12][5] , \xmem_data[12][4] , 
        \xmem_data[12][3] , \xmem_data[12][2] , \xmem_data[12][1] , 
        \xmem_data[12][0] }), .b({\fmem_data[12][7] , \fmem_data[12][6] , 
        \fmem_data[12][5] , \fmem_data[12][4] , \fmem_data[12][3] , 
        \fmem_data[12][2] , \fmem_data[12][1] , \fmem_data[12][0] }), 
        .product({\x_mult_f_int[12][15] , \x_mult_f_int[12][14] , 
        \x_mult_f_int[12][13] , \x_mult_f_int[12][12] , \x_mult_f_int[12][11] , 
        \x_mult_f_int[12][10] , \x_mult_f_int[12][9] , \x_mult_f_int[12][8] , 
        \x_mult_f_int[12][7] , \x_mult_f_int[12][6] , \x_mult_f_int[12][5] , 
        \x_mult_f_int[12][4] , \x_mult_f_int[12][3] , \x_mult_f_int[12][2] , 
        \x_mult_f_int[12][1] , \x_mult_f_int[12][0] }) );
  conv_128_32_DW_mult_pipe_J1_20 \multiplier[11].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8915), .tc(1'b1), .a({\xmem_data[11][7] , 
        \xmem_data[11][6] , \xmem_data[11][5] , \xmem_data[11][4] , 
        \xmem_data[11][3] , \xmem_data[11][2] , \xmem_data[11][1] , 
        \xmem_data[11][0] }), .b({\fmem_data[11][7] , \fmem_data[11][6] , 
        \fmem_data[11][5] , \fmem_data[11][4] , \fmem_data[11][3] , 
        \fmem_data[11][2] , \fmem_data[11][1] , \fmem_data[11][0] }), 
        .product({\x_mult_f_int[11][15] , \x_mult_f_int[11][14] , 
        \x_mult_f_int[11][13] , \x_mult_f_int[11][12] , \x_mult_f_int[11][11] , 
        \x_mult_f_int[11][10] , \x_mult_f_int[11][9] , \x_mult_f_int[11][8] , 
        \x_mult_f_int[11][7] , \x_mult_f_int[11][6] , \x_mult_f_int[11][5] , 
        \x_mult_f_int[11][4] , \x_mult_f_int[11][3] , \x_mult_f_int[11][2] , 
        \x_mult_f_int[11][1] , \x_mult_f_int[11][0] }) );
  conv_128_32_DW_mult_pipe_J1_21 \multiplier[10].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3450), .en(n8915), .tc(1'b1), .a({\xmem_data[10][7] , 
        \xmem_data[10][6] , \xmem_data[10][5] , \xmem_data[10][4] , 
        \xmem_data[10][3] , \xmem_data[10][2] , \xmem_data[10][1] , 
        \xmem_data[10][0] }), .b({\fmem_data[10][7] , \fmem_data[10][6] , 
        \fmem_data[10][5] , \fmem_data[10][4] , \fmem_data[10][3] , 
        \fmem_data[10][2] , \fmem_data[10][1] , \fmem_data[10][0] }), 
        .product({\x_mult_f_int[10][15] , \x_mult_f_int[10][14] , 
        \x_mult_f_int[10][13] , \x_mult_f_int[10][12] , \x_mult_f_int[10][11] , 
        \x_mult_f_int[10][10] , \x_mult_f_int[10][9] , \x_mult_f_int[10][8] , 
        \x_mult_f_int[10][7] , \x_mult_f_int[10][6] , \x_mult_f_int[10][5] , 
        \x_mult_f_int[10][4] , \x_mult_f_int[10][3] , \x_mult_f_int[10][2] , 
        \x_mult_f_int[10][1] , \x_mult_f_int[10][0] }) );
  conv_128_32_DW_mult_pipe_J1_22 \multiplier[9].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8919), .en(n8920), .tc(1'b1), .a({\xmem_data[9][7] , 
        \xmem_data[9][6] , \xmem_data[9][5] , \xmem_data[9][4] , 
        \xmem_data[9][3] , \xmem_data[9][2] , \xmem_data[9][1] , 
        \xmem_data[9][0] }), .b({\fmem_data[9][7] , \fmem_data[9][6] , 
        \fmem_data[9][5] , \fmem_data[9][4] , \fmem_data[9][3] , 
        \fmem_data[9][2] , \fmem_data[9][1] , \fmem_data[9][0] }), .product({
        \x_mult_f_int[9][15] , \x_mult_f_int[9][14] , \x_mult_f_int[9][13] , 
        \x_mult_f_int[9][12] , \x_mult_f_int[9][11] , \x_mult_f_int[9][10] , 
        \x_mult_f_int[9][9] , \x_mult_f_int[9][8] , \x_mult_f_int[9][7] , 
        \x_mult_f_int[9][6] , \x_mult_f_int[9][5] , \x_mult_f_int[9][4] , 
        \x_mult_f_int[9][3] , \x_mult_f_int[9][2] , \x_mult_f_int[9][1] , 
        \x_mult_f_int[9][0] }) );
  conv_128_32_DW_mult_pipe_J1_23 \multiplier[8].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8913), .tc(1'b1), .a({\xmem_data[8][7] , 
        \xmem_data[8][6] , \xmem_data[8][5] , \xmem_data[8][4] , 
        \xmem_data[8][3] , \xmem_data[8][2] , \xmem_data[8][1] , 
        \xmem_data[8][0] }), .b({\fmem_data[8][7] , \fmem_data[8][6] , 
        \fmem_data[8][5] , \fmem_data[8][4] , \fmem_data[8][3] , 
        \fmem_data[8][2] , \fmem_data[8][1] , \fmem_data[8][0] }), .product({
        \x_mult_f_int[8][15] , \x_mult_f_int[8][14] , \x_mult_f_int[8][13] , 
        \x_mult_f_int[8][12] , \x_mult_f_int[8][11] , \x_mult_f_int[8][10] , 
        \x_mult_f_int[8][9] , \x_mult_f_int[8][8] , \x_mult_f_int[8][7] , 
        \x_mult_f_int[8][6] , \x_mult_f_int[8][5] , \x_mult_f_int[8][4] , 
        \x_mult_f_int[8][3] , \x_mult_f_int[8][2] , \x_mult_f_int[8][1] , 
        \x_mult_f_int[8][0] }) );
  conv_128_32_DW_mult_pipe_J1_24 \multiplier[7].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8920), .tc(1'b1), .a({\xmem_data[7][7] , 
        \xmem_data[7][6] , \xmem_data[7][5] , \xmem_data[7][4] , 
        \xmem_data[7][3] , \xmem_data[7][2] , \xmem_data[7][1] , 
        \xmem_data[7][0] }), .b({\fmem_data[7][7] , \fmem_data[7][6] , 
        \fmem_data[7][5] , \fmem_data[7][4] , \fmem_data[7][3] , 
        \fmem_data[7][2] , \fmem_data[7][1] , \fmem_data[7][0] }), .product({
        \x_mult_f_int[7][15] , \x_mult_f_int[7][14] , \x_mult_f_int[7][13] , 
        \x_mult_f_int[7][12] , \x_mult_f_int[7][11] , \x_mult_f_int[7][10] , 
        \x_mult_f_int[7][9] , \x_mult_f_int[7][8] , \x_mult_f_int[7][7] , 
        \x_mult_f_int[7][6] , \x_mult_f_int[7][5] , \x_mult_f_int[7][4] , 
        \x_mult_f_int[7][3] , \x_mult_f_int[7][2] , \x_mult_f_int[7][1] , 
        \x_mult_f_int[7][0] }) );
  conv_128_32_DW_mult_pipe_J1_25 \multiplier[6].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8923), .tc(1'b1), .a({\xmem_data[6][7] , 
        \xmem_data[6][6] , \xmem_data[6][5] , \xmem_data[6][4] , 
        \xmem_data[6][3] , \xmem_data[6][2] , \xmem_data[6][1] , 
        \xmem_data[6][0] }), .b({\fmem_data[6][7] , \fmem_data[6][6] , 
        \fmem_data[6][5] , \fmem_data[6][4] , \fmem_data[6][3] , 
        \fmem_data[6][2] , \fmem_data[6][1] , \fmem_data[6][0] }), .product({
        \x_mult_f_int[6][15] , \x_mult_f_int[6][14] , \x_mult_f_int[6][13] , 
        \x_mult_f_int[6][12] , \x_mult_f_int[6][11] , \x_mult_f_int[6][10] , 
        \x_mult_f_int[6][9] , \x_mult_f_int[6][8] , \x_mult_f_int[6][7] , 
        \x_mult_f_int[6][6] , \x_mult_f_int[6][5] , \x_mult_f_int[6][4] , 
        \x_mult_f_int[6][3] , \x_mult_f_int[6][2] , \x_mult_f_int[6][1] , 
        \x_mult_f_int[6][0] }) );
  conv_128_32_DW_mult_pipe_J1_26 \multiplier[5].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n8918), .en(n8916), .tc(1'b1), .a({\xmem_data[5][7] , 
        \xmem_data[5][6] , \xmem_data[5][5] , \xmem_data[5][4] , 
        \xmem_data[5][3] , \xmem_data[5][2] , \xmem_data[5][1] , 
        \xmem_data[5][0] }), .b({\fmem_data[5][7] , \fmem_data[5][6] , 
        \fmem_data[5][5] , \fmem_data[5][4] , \fmem_data[5][3] , 
        \fmem_data[5][2] , \fmem_data[5][1] , \fmem_data[5][0] }), .product({
        \x_mult_f_int[5][15] , \x_mult_f_int[5][14] , \x_mult_f_int[5][13] , 
        \x_mult_f_int[5][12] , \x_mult_f_int[5][11] , \x_mult_f_int[5][10] , 
        \x_mult_f_int[5][9] , \x_mult_f_int[5][8] , \x_mult_f_int[5][7] , 
        \x_mult_f_int[5][6] , \x_mult_f_int[5][5] , \x_mult_f_int[5][4] , 
        \x_mult_f_int[5][3] , \x_mult_f_int[5][2] , \x_mult_f_int[5][1] , 
        \x_mult_f_int[5][0] }) );
  conv_128_32_DW_mult_pipe_J1_27 \multiplier[4].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3450), .en(n8920), .tc(1'b1), .a({\xmem_data[4][7] , 
        \xmem_data[4][6] , \xmem_data[4][5] , \xmem_data[4][4] , 
        \xmem_data[4][3] , \xmem_data[4][2] , \xmem_data[4][1] , 
        \xmem_data[4][0] }), .b({\fmem_data[4][7] , \fmem_data[4][6] , 
        \fmem_data[4][5] , \fmem_data[4][4] , \fmem_data[4][3] , 
        \fmem_data[4][2] , \fmem_data[4][1] , \fmem_data[4][0] }), .product({
        \x_mult_f_int[4][15] , \x_mult_f_int[4][14] , \x_mult_f_int[4][13] , 
        \x_mult_f_int[4][12] , \x_mult_f_int[4][11] , \x_mult_f_int[4][10] , 
        \x_mult_f_int[4][9] , \x_mult_f_int[4][8] , \x_mult_f_int[4][7] , 
        \x_mult_f_int[4][6] , \x_mult_f_int[4][5] , \x_mult_f_int[4][4] , 
        \x_mult_f_int[4][3] , \x_mult_f_int[4][2] , \x_mult_f_int[4][1] , 
        \x_mult_f_int[4][0] }) );
  conv_128_32_DW_mult_pipe_J1_28 \multiplier[3].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3449), .en(n8915), .tc(1'b1), .a({\xmem_data[3][7] , 
        \xmem_data[3][6] , \xmem_data[3][5] , \xmem_data[3][4] , 
        \xmem_data[3][3] , \xmem_data[3][2] , \xmem_data[3][1] , 
        \xmem_data[3][0] }), .b({\fmem_data[3][7] , \fmem_data[3][6] , 
        \fmem_data[3][5] , \fmem_data[3][4] , \fmem_data[3][3] , 
        \fmem_data[3][2] , \fmem_data[3][1] , \fmem_data[3][0] }), .product({
        \x_mult_f_int[3][15] , \x_mult_f_int[3][14] , \x_mult_f_int[3][13] , 
        \x_mult_f_int[3][12] , \x_mult_f_int[3][11] , \x_mult_f_int[3][10] , 
        \x_mult_f_int[3][9] , \x_mult_f_int[3][8] , \x_mult_f_int[3][7] , 
        \x_mult_f_int[3][6] , \x_mult_f_int[3][5] , \x_mult_f_int[3][4] , 
        \x_mult_f_int[3][3] , \x_mult_f_int[3][2] , \x_mult_f_int[3][1] , 
        \x_mult_f_int[3][0] }) );
  conv_128_32_DW_mult_pipe_J1_29 \multiplier[2].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3449), .en(n8916), .tc(1'b1), .a({\xmem_data[2][7] , 
        \xmem_data[2][6] , \xmem_data[2][5] , \xmem_data[2][4] , 
        \xmem_data[2][3] , \xmem_data[2][2] , \xmem_data[2][1] , 
        \xmem_data[2][0] }), .b({\fmem_data[2][7] , \fmem_data[2][6] , 
        \fmem_data[2][5] , \fmem_data[2][4] , \fmem_data[2][3] , 
        \fmem_data[2][2] , \fmem_data[2][1] , \fmem_data[2][0] }), .product({
        \x_mult_f_int[2][15] , \x_mult_f_int[2][14] , \x_mult_f_int[2][13] , 
        \x_mult_f_int[2][12] , \x_mult_f_int[2][11] , \x_mult_f_int[2][10] , 
        \x_mult_f_int[2][9] , \x_mult_f_int[2][8] , \x_mult_f_int[2][7] , 
        \x_mult_f_int[2][6] , \x_mult_f_int[2][5] , \x_mult_f_int[2][4] , 
        \x_mult_f_int[2][3] , \x_mult_f_int[2][2] , \x_mult_f_int[2][1] , 
        \x_mult_f_int[2][0] }) );
  conv_128_32_DW_mult_pipe_J1_30 \multiplier[1].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8916), .tc(1'b1), .a({\xmem_data[1][7] , 
        \xmem_data[1][6] , \xmem_data[1][5] , \xmem_data[1][4] , 
        \xmem_data[1][3] , \xmem_data[1][2] , \xmem_data[1][1] , 
        \xmem_data[1][0] }), .b({\fmem_data[1][7] , \fmem_data[1][6] , 
        \fmem_data[1][5] , \fmem_data[1][4] , \fmem_data[1][3] , 
        \fmem_data[1][2] , \fmem_data[1][1] , \fmem_data[1][0] }), .product({
        \x_mult_f_int[1][15] , \x_mult_f_int[1][14] , \x_mult_f_int[1][13] , 
        \x_mult_f_int[1][12] , \x_mult_f_int[1][11] , \x_mult_f_int[1][10] , 
        \x_mult_f_int[1][9] , \x_mult_f_int[1][8] , \x_mult_f_int[1][7] , 
        \x_mult_f_int[1][6] , \x_mult_f_int[1][5] , \x_mult_f_int[1][4] , 
        \x_mult_f_int[1][3] , \x_mult_f_int[1][2] , \x_mult_f_int[1][1] , 
        \x_mult_f_int[1][0] }) );
  conv_128_32_DW_mult_pipe_J1_31 \multiplier[0].x_f_mult_inst  ( .clk(clk), 
        .rst_n(n3448), .en(n8916), .tc(1'b1), .a({\xmem_data[0][7] , 
        \xmem_data[0][6] , \xmem_data[0][5] , \xmem_data[0][4] , 
        \xmem_data[0][3] , \xmem_data[0][2] , \xmem_data[0][1] , 
        \xmem_data[0][0] }), .b({\fmem_data[0][7] , \fmem_data[0][6] , 
        \fmem_data[0][5] , \fmem_data[0][4] , \fmem_data[0][3] , 
        \fmem_data[0][2] , \fmem_data[0][1] , \fmem_data[0][0] }), .product({
        \x_mult_f_int[0][15] , \x_mult_f_int[0][14] , \x_mult_f_int[0][13] , 
        \x_mult_f_int[0][12] , \x_mult_f_int[0][11] , \x_mult_f_int[0][10] , 
        \x_mult_f_int[0][9] , \x_mult_f_int[0][8] , \x_mult_f_int[0][7] , 
        \x_mult_f_int[0][6] , \x_mult_f_int[0][5] , \x_mult_f_int[0][4] , 
        \x_mult_f_int[0][3] , \x_mult_f_int[0][2] , \x_mult_f_int[0][1] , 
        \x_mult_f_int[0][0] }) );
  DFF_X1 \x_mult_f_reg[15][0]  ( .D(n9323), .CK(clk), .Q(\x_mult_f[15][0] ) );
  DFF_X1 \x_mult_f_reg[29][7]  ( .D(n9258), .CK(clk), .Q(\x_mult_f[29][7] ) );
  DFF_X1 \adder_stage3_reg[1][11]  ( .D(n9639), .CK(clk), .Q(
        \adder_stage3[1][11] ) );
  DFF_X1 \x_mult_f_reg[31][0]  ( .D(n9355), .CK(clk), .Q(\x_mult_f[31][0] ) );
  DFF_X1 \x_mult_f_reg[22][0]  ( .D(n9337), .CK(clk), .Q(\x_mult_f[22][0] ) );
  DFF_X1 \adder_stage1_reg[11][7]  ( .D(n9883), .CK(clk), .Q(
        \adder_stage1[11][7] ) );
  DFF_X1 \adder_stage2_reg[7][3]  ( .D(n9683), .CK(clk), .Q(
        \adder_stage2[7][3] ), .QN(n3440) );
  DFF_X1 \adder_stage1_reg[7][7]  ( .D(n9948), .CK(clk), .Q(
        \adder_stage1[7][7] ) );
  DFF_X1 \x_mult_f_reg[19][5]  ( .D(n9178), .CK(clk), .Q(\x_mult_f[19][5] ) );
  DFF_X1 \adder_stage1_reg[9][5]  ( .D(n9916), .CK(clk), .Q(
        \adder_stage1[9][5] ) );
  DFF_X1 \adder_stage1_reg[13][3]  ( .D(n9853), .CK(clk), .Q(
        \adder_stage1[13][3] ) );
  DFF_X1 \adder_stage2_reg[5][7]  ( .D(n9713), .CK(clk), .Q(
        \adder_stage2[5][7] ) );
  DFF_X1 \adder_stage2_reg[3][11]  ( .D(n9743), .CK(clk), .Q(
        \adder_stage2[3][11] ) );
  DFF_X1 \adder_stage2_reg[5][11]  ( .D(n9709), .CK(clk), .Q(
        \adder_stage2[5][11] ) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[1]  ( .D(n3394), .CK(clk), .Q(
        fmem_addr[1]), .QN(n8711) );
  DFF_X1 \ctrl_fmem_write_inst/s_ready_reg  ( .D(n3392), .CK(clk), .Q(
        s_ready_f), .QN(n8716) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[0]  ( .D(n3121), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [0]), .QN(n8713) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[1]  ( .D(n3120), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [1]), .QN(n8744) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[2]  ( .D(n3119), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [2]), .QN(n8715) );
  DFF_X1 \ctrl_inst/pline_cntr_reg[3]  ( .D(n3118), .CK(clk), .Q(
        \ctrl_inst/pline_cntr [3]), .QN(n8717) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[4]  ( .D(n3397), .CK(clk), .Q(
        fmem_addr[4]), .QN(n8746) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[0]  ( .D(n3395), .CK(clk), .Q(
        fmem_addr[0]), .QN(n8710) );
  DFF_X1 \ctrl_inst/state_reg[1]  ( .D(n3387), .CK(clk), .Q(
        \ctrl_inst/state [1]), .QN(n8714) );
  DFF_X1 \ctrl_inst/state_reg[2]  ( .D(n3386), .CK(clk), .Q(
        \ctrl_inst/state [2]), .QN(n8696) );
  DFF_X1 \ctrl_inst/xmem_tracker_reg[6]  ( .D(n3384), .CK(clk), .Q(
        \ctrl_inst/xmem_tracker [6]), .QN(n8745) );
  DFF_X1 \ctrl_fmem_write_inst/mem_addr_reg[2]  ( .D(n3393), .CK(clk), .Q(
        fmem_addr[2]), .QN(n8709) );
  DFF_X1 \fmem_inst/mem_reg[12][7]  ( .D(n8870), .CK(clk), .QN(
        \fmem_data[12][7] ) );
  DFF_X1 \fmem_inst/mem_reg[12][6]  ( .D(n8871), .CK(clk), .QN(
        \fmem_data[12][6] ) );
  DFF_X1 \fmem_inst/mem_reg[12][5]  ( .D(n8872), .CK(clk), .QN(
        \fmem_data[12][5] ) );
  DFF_X1 \fmem_inst/mem_reg[12][4]  ( .D(n8873), .CK(clk), .QN(
        \fmem_data[12][4] ) );
  DFF_X1 \fmem_inst/mem_reg[12][3]  ( .D(n8874), .CK(clk), .QN(
        \fmem_data[12][3] ) );
  DFF_X1 \fmem_inst/mem_reg[12][2]  ( .D(n8875), .CK(clk), .QN(
        \fmem_data[12][2] ) );
  DFF_X1 \fmem_inst/mem_reg[12][1]  ( .D(n8876), .CK(clk), .QN(
        \fmem_data[12][1] ) );
  DFF_X1 \fmem_inst/mem_reg[12][0]  ( .D(n8877), .CK(clk), .QN(
        \fmem_data[12][0] ) );
  DFF_X1 \fmem_inst/mem_reg[14][7]  ( .D(n8854), .CK(clk), .QN(
        \fmem_data[14][7] ) );
  DFF_X1 \fmem_inst/mem_reg[14][6]  ( .D(n8855), .CK(clk), .QN(
        \fmem_data[14][6] ) );
  DFF_X1 \fmem_inst/mem_reg[14][5]  ( .D(n8856), .CK(clk), .QN(
        \fmem_data[14][5] ) );
  DFF_X1 \fmem_inst/mem_reg[14][4]  ( .D(n8857), .CK(clk), .QN(
        \fmem_data[14][4] ) );
  DFF_X1 \fmem_inst/mem_reg[14][3]  ( .D(n8858), .CK(clk), .QN(
        \fmem_data[14][3] ) );
  DFF_X1 \fmem_inst/mem_reg[14][2]  ( .D(n8859), .CK(clk), .QN(
        \fmem_data[14][2] ) );
  DFF_X1 \fmem_inst/mem_reg[14][1]  ( .D(n8860), .CK(clk), .QN(
        \fmem_data[14][1] ) );
  DFF_X1 \fmem_inst/mem_reg[14][0]  ( .D(n8861), .CK(clk), .QN(
        \fmem_data[14][0] ) );
  DFF_X1 \fmem_inst/mem_reg[10][7]  ( .D(n8886), .CK(clk), .QN(
        \fmem_data[10][7] ) );
  DFF_X1 \fmem_inst/mem_reg[10][6]  ( .D(n8887), .CK(clk), .QN(
        \fmem_data[10][6] ) );
  DFF_X1 \fmem_inst/mem_reg[10][5]  ( .D(n8888), .CK(clk), .QN(
        \fmem_data[10][5] ) );
  DFF_X1 \fmem_inst/mem_reg[10][4]  ( .D(n8889), .CK(clk), .QN(
        \fmem_data[10][4] ) );
  DFF_X1 \fmem_inst/mem_reg[10][3]  ( .D(n8890), .CK(clk), .QN(
        \fmem_data[10][3] ) );
  DFF_X1 \fmem_inst/mem_reg[10][2]  ( .D(n8891), .CK(clk), .QN(
        \fmem_data[10][2] ) );
  DFF_X1 \fmem_inst/mem_reg[10][1]  ( .D(n8892), .CK(clk), .QN(
        \fmem_data[10][1] ) );
  DFF_X1 \fmem_inst/mem_reg[10][0]  ( .D(n8893), .CK(clk), .QN(
        \fmem_data[10][0] ) );
  DFF_X1 \fmem_inst/mem_reg[8][7]  ( .D(n8902), .CK(clk), .QN(
        \fmem_data[8][7] ) );
  DFF_X1 \fmem_inst/mem_reg[8][6]  ( .D(n8903), .CK(clk), .QN(
        \fmem_data[8][6] ) );
  DFF_X1 \fmem_inst/mem_reg[8][5]  ( .D(n8904), .CK(clk), .QN(
        \fmem_data[8][5] ) );
  DFF_X1 \fmem_inst/mem_reg[8][4]  ( .D(n8905), .CK(clk), .QN(
        \fmem_data[8][4] ) );
  DFF_X1 \fmem_inst/mem_reg[8][3]  ( .D(n8906), .CK(clk), .QN(
        \fmem_data[8][3] ) );
  DFF_X1 \fmem_inst/mem_reg[8][2]  ( .D(n8907), .CK(clk), .QN(
        \fmem_data[8][2] ) );
  DFF_X1 \fmem_inst/mem_reg[8][1]  ( .D(n8908), .CK(clk), .QN(
        \fmem_data[8][1] ) );
  DFF_X1 \fmem_inst/mem_reg[8][0]  ( .D(n8909), .CK(clk), .QN(
        \fmem_data[8][0] ) );
  DFF_X1 \fmem_inst/mem_reg[13][7]  ( .D(n8862), .CK(clk), .QN(
        \fmem_data[13][7] ) );
  DFF_X1 \fmem_inst/mem_reg[13][6]  ( .D(n8863), .CK(clk), .QN(
        \fmem_data[13][6] ) );
  DFF_X1 \fmem_inst/mem_reg[13][5]  ( .D(n8864), .CK(clk), .QN(
        \fmem_data[13][5] ) );
  DFF_X1 \fmem_inst/mem_reg[13][4]  ( .D(n8865), .CK(clk), .QN(
        \fmem_data[13][4] ) );
  DFF_X1 \fmem_inst/mem_reg[13][3]  ( .D(n8866), .CK(clk), .QN(
        \fmem_data[13][3] ) );
  DFF_X1 \fmem_inst/mem_reg[13][2]  ( .D(n8867), .CK(clk), .QN(
        \fmem_data[13][2] ) );
  DFF_X1 \fmem_inst/mem_reg[13][1]  ( .D(n8868), .CK(clk), .QN(
        \fmem_data[13][1] ) );
  DFF_X1 \fmem_inst/mem_reg[13][0]  ( .D(n8869), .CK(clk), .QN(
        \fmem_data[13][0] ) );
  DFF_X1 \fmem_inst/mem_reg[9][7]  ( .D(n8894), .CK(clk), .QN(
        \fmem_data[9][7] ) );
  DFF_X1 \fmem_inst/mem_reg[9][6]  ( .D(n8895), .CK(clk), .QN(
        \fmem_data[9][6] ) );
  DFF_X1 \fmem_inst/mem_reg[9][5]  ( .D(n8896), .CK(clk), .QN(
        \fmem_data[9][5] ) );
  DFF_X1 \fmem_inst/mem_reg[9][4]  ( .D(n8897), .CK(clk), .QN(
        \fmem_data[9][4] ) );
  DFF_X1 \fmem_inst/mem_reg[9][3]  ( .D(n8898), .CK(clk), .QN(
        \fmem_data[9][3] ) );
  DFF_X1 \fmem_inst/mem_reg[9][2]  ( .D(n8899), .CK(clk), .QN(
        \fmem_data[9][2] ) );
  DFF_X1 \fmem_inst/mem_reg[9][1]  ( .D(n8900), .CK(clk), .QN(
        \fmem_data[9][1] ) );
  DFF_X1 \fmem_inst/mem_reg[9][0]  ( .D(n8901), .CK(clk), .QN(
        \fmem_data[9][0] ) );
  DFF_X1 \fmem_inst/mem_reg[11][7]  ( .D(n8878), .CK(clk), .QN(
        \fmem_data[11][7] ) );
  DFF_X1 \fmem_inst/mem_reg[11][6]  ( .D(n8879), .CK(clk), .QN(
        \fmem_data[11][6] ) );
  DFF_X1 \fmem_inst/mem_reg[11][5]  ( .D(n8880), .CK(clk), .QN(
        \fmem_data[11][5] ) );
  DFF_X1 \fmem_inst/mem_reg[11][4]  ( .D(n8881), .CK(clk), .QN(
        \fmem_data[11][4] ) );
  DFF_X1 \fmem_inst/mem_reg[11][3]  ( .D(n8882), .CK(clk), .QN(
        \fmem_data[11][3] ) );
  DFF_X1 \fmem_inst/mem_reg[11][2]  ( .D(n8883), .CK(clk), .QN(
        \fmem_data[11][2] ) );
  DFF_X1 \fmem_inst/mem_reg[11][1]  ( .D(n8884), .CK(clk), .QN(
        \fmem_data[11][1] ) );
  DFF_X1 \fmem_inst/mem_reg[11][0]  ( .D(n8885), .CK(clk), .QN(
        \fmem_data[11][0] ) );
  DFF_X1 \fmem_inst/mem_reg[15][7]  ( .D(n8846), .CK(clk), .QN(
        \fmem_data[15][7] ) );
  DFF_X1 \fmem_inst/mem_reg[15][6]  ( .D(n8847), .CK(clk), .QN(
        \fmem_data[15][6] ) );
  DFF_X1 \fmem_inst/mem_reg[15][5]  ( .D(n8848), .CK(clk), .QN(
        \fmem_data[15][5] ) );
  DFF_X1 \fmem_inst/mem_reg[15][4]  ( .D(n8849), .CK(clk), .QN(
        \fmem_data[15][4] ) );
  DFF_X1 \fmem_inst/mem_reg[15][3]  ( .D(n8850), .CK(clk), .QN(
        \fmem_data[15][3] ) );
  DFF_X1 \fmem_inst/mem_reg[15][2]  ( .D(n8851), .CK(clk), .QN(
        \fmem_data[15][2] ) );
  DFF_X1 \fmem_inst/mem_reg[15][1]  ( .D(n8852), .CK(clk), .QN(
        \fmem_data[15][1] ) );
  DFF_X1 \fmem_inst/mem_reg[15][0]  ( .D(n8853), .CK(clk), .QN(
        \fmem_data[15][0] ) );
  DFF_X1 \fmem_inst/mem_reg[4][7]  ( .D(n8910), .CK(clk), .QN(
        \fmem_data[4][7] ) );
  DFF_X1 \adder_stage1_reg[0][2]  ( .D(n8790), .CK(clk), .QN(
        \adder_stage1[0][2] ) );
  DFF_X1 \adder_stage1_reg[10][2]  ( .D(n8819), .CK(clk), .QN(
        \adder_stage1[10][2] ) );
  DFF_X1 \x_mult_f_reg[26][15]  ( .D(n8782), .CK(clk), .Q(n8704), .QN(
        \x_mult_f[26][15] ) );
  DFF_X1 \x_mult_f_reg[26][14]  ( .D(n8773), .CK(clk), .QN(\x_mult_f[26][14] )
         );
  DFF_X1 \x_mult_f_reg[26][13]  ( .D(n8765), .CK(clk), .QN(\x_mult_f[26][13] )
         );
  DFF_X1 \x_mult_f_reg[26][12]  ( .D(n8767), .CK(clk), .QN(\x_mult_f[26][12] )
         );
  DFF_X1 \x_mult_f_reg[26][11]  ( .D(n8830), .CK(clk), .QN(\x_mult_f[26][11] )
         );
  DFF_X1 \x_mult_f_reg[26][10]  ( .D(n8831), .CK(clk), .QN(\x_mult_f[26][10] )
         );
  DFF_X1 \x_mult_f_reg[26][9]  ( .D(n8832), .CK(clk), .QN(\x_mult_f[26][9] )
         );
  DFF_X1 \x_mult_f_reg[25][5]  ( .D(n8829), .CK(clk), .QN(\x_mult_f[25][5] )
         );
  DFF_X1 \x_mult_f_reg[24][12]  ( .D(n8758), .CK(clk), .QN(\x_mult_f[24][12] )
         );
  DFF_X1 \x_mult_f_reg[21][5]  ( .D(n8816), .CK(clk), .QN(\x_mult_f[21][5] )
         );
  DFF_X1 \x_mult_f_reg[5][15]  ( .D(n8781), .CK(clk), .Q(n8698), .QN(
        \x_mult_f[5][15] ) );
  DFF_X1 \x_mult_f_reg[5][14]  ( .D(n8762), .CK(clk), .QN(\x_mult_f[5][14] )
         );
  DFF_X1 \x_mult_f_reg[5][13]  ( .D(n8763), .CK(clk), .QN(\x_mult_f[5][13] )
         );
  DFF_X1 \adder_stage1_reg[10][13]  ( .D(n8818), .CK(clk), .QN(
        \adder_stage1[10][13] ) );
  DFF_X1 \x_mult_f_reg[27][8]  ( .D(n8836), .CK(clk), .QN(\x_mult_f[27][8] )
         );
  DFF_X1 \x_mult_f_reg[26][8]  ( .D(n8833), .CK(clk), .QN(\x_mult_f[26][8] )
         );
  DFF_X1 \x_mult_f_reg[26][6]  ( .D(n8834), .CK(clk), .QN(\x_mult_f[26][6] )
         );
  DFF_X1 \x_mult_f_reg[26][5]  ( .D(n8835), .CK(clk), .QN(\x_mult_f[26][5] )
         );
  DFF_X1 \x_mult_f_reg[25][15]  ( .D(n8777), .CK(clk), .Q(n8703), .QN(
        \x_mult_f[25][15] ) );
  DFF_X1 \x_mult_f_reg[25][14]  ( .D(n8775), .CK(clk), .QN(\x_mult_f[25][14] )
         );
  DFF_X1 \x_mult_f_reg[25][13]  ( .D(n8760), .CK(clk), .QN(\x_mult_f[25][13] )
         );
  DFF_X1 \x_mult_f_reg[25][12]  ( .D(n8759), .CK(clk), .QN(\x_mult_f[25][12] )
         );
  DFF_X1 \x_mult_f_reg[25][11]  ( .D(n8823), .CK(clk), .QN(\x_mult_f[25][11] )
         );
  DFF_X1 \x_mult_f_reg[25][10]  ( .D(n8824), .CK(clk), .QN(\x_mult_f[25][10] )
         );
  DFF_X1 \x_mult_f_reg[25][9]  ( .D(n8825), .CK(clk), .QN(\x_mult_f[25][9] )
         );
  DFF_X1 \x_mult_f_reg[25][8]  ( .D(n8826), .CK(clk), .QN(\x_mult_f[25][8] )
         );
  DFF_X1 \x_mult_f_reg[25][7]  ( .D(n8827), .CK(clk), .QN(\x_mult_f[25][7] )
         );
  DFF_X1 \x_mult_f_reg[25][6]  ( .D(n8828), .CK(clk), .QN(\x_mult_f[25][6] )
         );
  DFF_X1 \x_mult_f_reg[24][7]  ( .D(n8821), .CK(clk), .QN(\x_mult_f[24][7] )
         );
  DFF_X1 \x_mult_f_reg[24][5]  ( .D(n8822), .CK(clk), .QN(\x_mult_f[24][5] )
         );
  DFF_X1 \x_mult_f_reg[1][8]  ( .D(n8788), .CK(clk), .QN(\x_mult_f[1][8] ) );
  DFF_X1 \x_mult_f_reg[1][5]  ( .D(n8789), .CK(clk), .QN(\x_mult_f[1][5] ) );
  DFF_X1 \x_mult_f_reg[0][8]  ( .D(n8784), .CK(clk), .QN(\x_mult_f[0][8] ) );
  DFF_X1 \x_mult_f_reg[0][5]  ( .D(n8785), .CK(clk), .QN(\x_mult_f[0][5] ) );
  DFF_X1 \adder_stage3_reg[0][19]  ( .D(n8793), .CK(clk), .QN(
        \adder_stage3[0][19] ) );
  DFF_X1 \adder_stage3_reg[0][18]  ( .D(n8794), .CK(clk), .QN(
        \adder_stage3[0][18] ) );
  DFF_X1 \adder_stage1_reg[2][14]  ( .D(n8792), .CK(clk), .QN(
        \adder_stage1[2][14] ) );
  DFF_X1 \x_mult_f_reg[21][10]  ( .D(n8811), .CK(clk), .QN(\x_mult_f[21][10] )
         );
  DFF_X1 \x_mult_f_reg[21][9]  ( .D(n8812), .CK(clk), .QN(\x_mult_f[21][9] )
         );
  DFF_X1 \x_mult_f_reg[21][8]  ( .D(n8813), .CK(clk), .QN(\x_mult_f[21][8] )
         );
  DFF_X1 \x_mult_f_reg[21][7]  ( .D(n8814), .CK(clk), .QN(\x_mult_f[21][7] )
         );
  DFF_X1 \x_mult_f_reg[28][13]  ( .D(n8837), .CK(clk), .QN(\x_mult_f[28][13] )
         );
  DFF_X1 \x_mult_f_reg[28][12]  ( .D(n8838), .CK(clk), .QN(\x_mult_f[28][12] )
         );
  DFF_X1 \x_mult_f_reg[28][11]  ( .D(n8839), .CK(clk), .QN(\x_mult_f[28][11] )
         );
  DFF_X1 \x_mult_f_reg[28][10]  ( .D(n8840), .CK(clk), .QN(\x_mult_f[28][10] )
         );
  DFF_X1 \x_mult_f_reg[28][9]  ( .D(n8841), .CK(clk), .QN(\x_mult_f[28][9] )
         );
  DFF_X1 \x_mult_f_reg[28][8]  ( .D(n8842), .CK(clk), .QN(\x_mult_f[28][8] )
         );
  DFF_X1 \x_mult_f_reg[28][7]  ( .D(n8843), .CK(clk), .QN(\x_mult_f[28][7] )
         );
  DFF_X1 \x_mult_f_reg[28][6]  ( .D(n8844), .CK(clk), .QN(\x_mult_f[28][6] )
         );
  DFF_X1 \x_mult_f_reg[22][12]  ( .D(n8755), .CK(clk), .QN(\x_mult_f[22][12] )
         );
  DFF_X1 \x_mult_f_reg[22][15]  ( .D(n8783), .CK(clk), .Q(n8701), .QN(
        \x_mult_f[22][15] ) );
  DFF_X1 \x_mult_f_reg[22][14]  ( .D(n8778), .CK(clk), .QN(\x_mult_f[22][14] )
         );
  DFF_X1 \x_mult_f_reg[22][13]  ( .D(n8761), .CK(clk), .QN(\x_mult_f[22][13] )
         );
  DFF_X1 \x_mult_f_reg[21][6]  ( .D(n8815), .CK(clk), .QN(\x_mult_f[21][6] )
         );
  DFF_X1 \adder_stage1_reg[10][20]  ( .D(n8817), .CK(clk), .Q(n8708), .QN(
        \adder_stage1[10][20] ) );
  DFF_X1 \x_mult_f_reg[29][13]  ( .D(n8845), .CK(clk), .QN(\x_mult_f[29][13] )
         );
  DFF_X1 \adder_stage1_reg[4][14]  ( .D(n8801), .CK(clk), .QN(
        \adder_stage1[4][14] ) );
  DFF_X1 \adder_stage1_reg[4][13]  ( .D(n8802), .CK(clk), .QN(
        \adder_stage1[4][13] ) );
  DFF_X1 \x_mult_f_reg[9][13]  ( .D(n8772), .CK(clk), .QN(\x_mult_f[9][13] )
         );
  DFF_X1 \x_mult_f_reg[9][12]  ( .D(n8771), .CK(clk), .QN(\x_mult_f[9][12] )
         );
  DFF_X1 \x_mult_f_reg[9][11]  ( .D(n8795), .CK(clk), .QN(\x_mult_f[9][11] )
         );
  DFF_X1 \x_mult_f_reg[9][10]  ( .D(n8796), .CK(clk), .QN(\x_mult_f[9][10] )
         );
  DFF_X1 \x_mult_f_reg[9][9]  ( .D(n8797), .CK(clk), .QN(\x_mult_f[9][9] ) );
  DFF_X1 \x_mult_f_reg[9][8]  ( .D(n8798), .CK(clk), .QN(\x_mult_f[9][8] ) );
  DFF_X1 \x_mult_f_reg[9][6]  ( .D(n8799), .CK(clk), .QN(\x_mult_f[9][6] ) );
  DFF_X1 \x_mult_f_reg[29][15]  ( .D(n8780), .CK(clk), .Q(n8705), .QN(
        \x_mult_f[29][15] ) );
  DFF_X1 \x_mult_f_reg[29][14]  ( .D(n8770), .CK(clk), .QN(\x_mult_f[29][14] )
         );
  DFF_X1 \x_mult_f_reg[23][15]  ( .D(n8768), .CK(clk), .Q(n8702), .QN(
        \x_mult_f[23][15] ) );
  DFF_X1 \x_mult_f_reg[23][14]  ( .D(n8756), .CK(clk), .QN(\x_mult_f[23][14] )
         );
  DFF_X1 \x_mult_f_reg[23][13]  ( .D(n8757), .CK(clk), .QN(\x_mult_f[23][13] )
         );
  DFF_X1 \x_mult_f_reg[22][6]  ( .D(n8820), .CK(clk), .QN(\x_mult_f[22][6] )
         );
  DFF_X1 \x_mult_f_reg[20][15]  ( .D(n8776), .CK(clk), .Q(n8700), .QN(
        \x_mult_f[20][15] ) );
  DFF_X1 \x_mult_f_reg[20][14]  ( .D(n8774), .CK(clk), .QN(\x_mult_f[20][14] )
         );
  DFF_X1 \x_mult_f_reg[20][13]  ( .D(n8766), .CK(clk), .QN(\x_mult_f[20][13] )
         );
  DFF_X1 \x_mult_f_reg[20][12]  ( .D(n8764), .CK(clk), .QN(\x_mult_f[20][12] )
         );
  DFF_X1 \x_mult_f_reg[20][11]  ( .D(n8807), .CK(clk), .QN(\x_mult_f[20][11] )
         );
  DFF_X1 \x_mult_f_reg[20][10]  ( .D(n8808), .CK(clk), .QN(\x_mult_f[20][10] )
         );
  DFF_X1 \x_mult_f_reg[20][9]  ( .D(n8809), .CK(clk), .QN(\x_mult_f[20][9] )
         );
  DFF_X1 \x_mult_f_reg[20][8]  ( .D(n8810), .CK(clk), .QN(\x_mult_f[20][8] )
         );
  DFF_X1 \x_mult_f_reg[9][15]  ( .D(n8779), .CK(clk), .Q(n8699), .QN(
        \x_mult_f[9][15] ) );
  DFF_X1 \x_mult_f_reg[9][14]  ( .D(n8769), .CK(clk), .QN(\x_mult_f[9][14] )
         );
  DFF_X1 \adder_stage1_reg[4][20]  ( .D(n8800), .CK(clk), .Q(n8707), .QN(
        \adder_stage1[4][20] ) );
  DFF_X1 \x_mult_f_reg[10][4]  ( .D(n8803), .CK(clk), .QN(\x_mult_f[10][4] )
         );
  DFF_X1 \x_mult_f_reg[10][2]  ( .D(n8804), .CK(clk), .QN(\x_mult_f[10][2] )
         );
  DFF_X1 \x_mult_f_reg[0][3]  ( .D(n8786), .CK(clk), .QN(\x_mult_f[0][3] ) );
  DFF_X1 \x_mult_f_reg[0][2]  ( .D(n8787), .CK(clk), .QN(\x_mult_f[0][2] ) );
  DFF_X1 \x_mult_f_reg[16][3]  ( .D(n8806), .CK(clk), .QN(\x_mult_f[16][3] )
         );
  DFF_X1 \ctrl_inst/s_ready_fsm_reg  ( .D(n3385), .CK(clk), .Q(n8697), .QN(
        n8719) );
  DFF_X1 \x_mult_f_reg[12][4]  ( .D(n8805), .CK(clk), .QN(\x_mult_f[12][4] )
         );
  DFF_X1 \x_mult_f_reg[3][7]  ( .D(n8791), .CK(clk), .QN(\x_mult_f[3][7] ) );
  DFF_X1 \adder_stage2_reg[7][20]  ( .D(n1909), .CK(clk), .Q(
        \adder_stage2[7][20] ), .QN(n8751) );
  BUF_X1 U3404 ( .A(n5447), .Z(n5480) );
  INV_X1 U3405 ( .A(n3807), .ZN(n3809) );
  AND2_X1 U3406 ( .A1(\ctrl_inst/xmem_tracker [5]), .A2(
        \ctrl_inst/xmem_tracker [6]), .ZN(n3400) );
  BUF_X1 U3407 ( .A(n3950), .Z(n8318) );
  BUF_X1 U3408 ( .A(n3950), .Z(n8329) );
  CLKBUF_X2 U3409 ( .A(n6231), .Z(n8186) );
  CLKBUF_X2 U3410 ( .A(n6231), .Z(n6523) );
  BUF_X1 U3411 ( .A(n6231), .Z(n8310) );
  CLKBUF_X2 U3412 ( .A(n6231), .Z(n8229) );
  CLKBUF_X2 U3413 ( .A(n6645), .Z(n7110) );
  BUF_X1 U3414 ( .A(n6231), .Z(n7182) );
  BUF_X1 U3415 ( .A(n6645), .Z(n8398) );
  CLKBUF_X2 U3416 ( .A(n6231), .Z(n6256) );
  BUF_X1 U3417 ( .A(n6231), .Z(n7369) );
  CLKBUF_X2 U3418 ( .A(n6645), .Z(n6915) );
  CLKBUF_X2 U3419 ( .A(n6231), .Z(n8216) );
  BUF_X1 U3420 ( .A(n6231), .Z(n8291) );
  CLKBUF_X2 U3421 ( .A(n6231), .Z(n8203) );
  CLKBUF_X2 U3422 ( .A(n6645), .Z(n7356) );
  CLKBUF_X2 U3423 ( .A(n6231), .Z(n8037) );
  CLKBUF_X2 U3424 ( .A(n6645), .Z(n7454) );
  CLKBUF_X2 U3425 ( .A(n6645), .Z(n6221) );
  CLKBUF_X2 U3426 ( .A(n6645), .Z(n8194) );
  CLKBUF_X2 U3427 ( .A(n6645), .Z(n8389) );
  CLKBUF_X2 U3428 ( .A(n6231), .Z(n7511) );
  BUF_X2 U3429 ( .A(n6435), .Z(n3950) );
  INV_X1 U3430 ( .A(n3808), .ZN(n8919) );
  AND2_X1 U3431 ( .A1(m_ready_y), .A2(m_valid_y), .ZN(n3858) );
  OR2_X1 U3432 ( .A1(n8179), .A2(n3417), .ZN(n8182) );
  XNOR2_X1 U3433 ( .A(n8142), .B(n3415), .ZN(n7971) );
  INV_X1 U3434 ( .A(n6105), .ZN(n8364) );
  BUF_X2 U3435 ( .A(n5921), .Z(n8150) );
  BUF_X2 U3436 ( .A(n6435), .Z(n8282) );
  AND2_X1 U3437 ( .A1(n8919), .A2(n8917), .ZN(n6435) );
  OAI21_X1 U3438 ( .B1(n6705), .B2(n6701), .A(n6702), .ZN(n7115) );
  OAI21_X1 U3439 ( .B1(n4796), .B2(n4793), .A(n4794), .ZN(n4830) );
  AOI21_X1 U3440 ( .B1(n5140), .B2(n5102), .A(n5101), .ZN(n5298) );
  OR2_X1 U3441 ( .A1(n8712), .A2(n8481), .ZN(n8470) );
  INV_X1 U3442 ( .A(n3808), .ZN(n3448) );
  INV_X2 U3443 ( .A(n3808), .ZN(n3450) );
  INV_X2 U3444 ( .A(n3808), .ZN(n8918) );
  OR2_X1 U3445 ( .A1(fmem_addr[3]), .A2(n8481), .ZN(n8552) );
  INV_X1 U3446 ( .A(n3820), .ZN(n3408) );
  INV_X1 U3447 ( .A(n3521), .ZN(n5455) );
  INV_X1 U3448 ( .A(n8688), .ZN(n8680) );
  CLKBUF_X1 U3449 ( .A(n3858), .Z(n3425) );
  AND2_X1 U3450 ( .A1(n8696), .A2(n8714), .ZN(n3404) );
  AND2_X1 U3451 ( .A1(\ctrl_inst/state [0]), .A2(n8714), .ZN(n3521) );
  NOR2_X1 U3452 ( .A1(\x_mult_f[2][5] ), .A2(\x_mult_f[3][5] ), .ZN(n7210) );
  NOR2_X1 U3453 ( .A1(\adder_stage1[12][3] ), .A2(\adder_stage1[13][3] ), .ZN(
        n5620) );
  NOR2_X1 U3454 ( .A1(\adder_stage1[10][3] ), .A2(\adder_stage1[11][3] ), .ZN(
        n4657) );
  INV_X1 U3455 ( .A(n4793), .ZN(n3401) );
  XNOR2_X1 U3456 ( .A(n3496), .B(n3462), .ZN(n3415) );
  NAND2_X1 U3457 ( .A1(s_valid_f), .A2(s_ready_f), .ZN(n8682) );
  NOR2_X1 U3458 ( .A1(\x_mult_f[6][3] ), .A2(\x_mult_f[7][3] ), .ZN(n6654) );
  NAND2_X1 U3459 ( .A1(s_valid_x), .A2(n3402), .ZN(n3407) );
  AND2_X1 U3460 ( .A1(n3404), .A2(n3403), .ZN(n3402) );
  AND2_X1 U3461 ( .A1(n3810), .A2(\ctrl_inst/state [0]), .ZN(n3403) );
  NAND2_X1 U3462 ( .A1(n3858), .A2(n3834), .ZN(n3406) );
  NAND2_X1 U3463 ( .A1(n3400), .A2(n3405), .ZN(n3657) );
  INV_X1 U3464 ( .A(n3849), .ZN(n3405) );
  NAND4_X1 U3465 ( .A1(n3815), .A2(\ctrl_inst/xmem_tracker [2]), .A3(
        \ctrl_inst/xmem_tracker [3]), .A4(\ctrl_inst/xmem_tracker [4]), .ZN(
        n3849) );
  OAI21_X1 U3466 ( .B1(m_ready_y), .B2(n8697), .A(n3657), .ZN(n3812) );
  OAI21_X2 U3467 ( .B1(n3812), .B2(n3407), .A(n3406), .ZN(n3807) );
  NAND2_X2 U3468 ( .A1(n8688), .A2(n3408), .ZN(n3808) );
  NOR2_X2 U3469 ( .A1(conv_done), .A2(reset), .ZN(n8688) );
  INV_X1 U3470 ( .A(n3409), .ZN(n4633) );
  OAI21_X1 U3471 ( .B1(n4796), .B2(n3412), .A(n3410), .ZN(n3409) );
  AOI21_X1 U3472 ( .B1(n4828), .B2(n3411), .A(n4618), .ZN(n3410) );
  INV_X1 U3473 ( .A(n4794), .ZN(n3411) );
  NAND2_X1 U3474 ( .A1(n3401), .A2(n4828), .ZN(n3412) );
  AOI21_X1 U3475 ( .B1(n5471), .B2(n5470), .A(n5469), .ZN(n3426) );
  OAI21_X1 U3476 ( .B1(n4633), .B2(n4629), .A(n4630), .ZN(n5471) );
  AOI22_X1 U3477 ( .A1(n8142), .A2(n3414), .B1(n3496), .B2(n3462), .ZN(n3413)
         );
  NAND2_X1 U3478 ( .A1(\adder_stage1[13][20] ), .A2(\adder_stage1[12][20] ), 
        .ZN(n3414) );
  INV_X1 U3479 ( .A(n3416), .ZN(n7970) );
  AOI21_X1 U3480 ( .B1(n5304), .B2(n5305), .A(n5303), .ZN(n3416) );
  AND2_X1 U3481 ( .A1(n8181), .A2(n8180), .ZN(n3417) );
  INV_X2 U3482 ( .A(n5378), .ZN(n8178) );
  OAI21_X1 U3483 ( .B1(n7102), .B2(n7098), .A(n7099), .ZN(n7046) );
  NAND2_X1 U3484 ( .A1(n3419), .A2(n3418), .ZN(n9704) );
  NAND2_X1 U3485 ( .A1(n8094), .A2(\adder_stage2[5][16] ), .ZN(n3418) );
  NAND2_X1 U3486 ( .A1(n8095), .A2(n7909), .ZN(n3419) );
  AOI22_X1 U3487 ( .A1(n7919), .A2(n3420), .B1(\adder_stage1[1][20] ), .B2(
        n8364), .ZN(n7920) );
  AND2_X1 U3488 ( .A1(n8265), .A2(n7918), .ZN(n3420) );
  NAND2_X1 U3489 ( .A1(n3422), .A2(n3421), .ZN(n9589) );
  NAND2_X1 U3490 ( .A1(n8200), .A2(\adder_stage3[3][20] ), .ZN(n3421) );
  NAND2_X1 U3491 ( .A1(n8166), .A2(n8365), .ZN(n3422) );
  NOR2_X2 U3492 ( .A1(n8676), .A2(n8470), .ZN(n8689) );
  OAI21_X1 U3493 ( .B1(n6123), .B2(n6077), .A(n6216), .ZN(n6071) );
  NAND2_X1 U3494 ( .A1(n6149), .A2(n3423), .ZN(n6123) );
  AND2_X1 U3495 ( .A1(n6132), .A2(n6134), .ZN(n3423) );
  NAND2_X1 U3496 ( .A1(n3424), .A2(n6117), .ZN(n8107) );
  NAND2_X1 U3497 ( .A1(n6116), .A2(n6118), .ZN(n3424) );
  INV_X1 U3498 ( .A(n4998), .ZN(n3549) );
  OAI21_X1 U3499 ( .B1(n5537), .B2(n3548), .A(n5539), .ZN(n4997) );
  INV_X1 U3500 ( .A(n5540), .ZN(n3548) );
  AOI21_X1 U3501 ( .B1(n3547), .B2(n5504), .A(n3546), .ZN(n5537) );
  INV_X1 U3502 ( .A(n5507), .ZN(n3546) );
  INV_X1 U3503 ( .A(n3872), .ZN(n3651) );
  OAI21_X1 U3504 ( .B1(n5008), .B2(n3650), .A(n5010), .ZN(n3871) );
  INV_X1 U3505 ( .A(n5011), .ZN(n3650) );
  AOI21_X1 U3506 ( .B1(n3649), .B2(n5016), .A(n3648), .ZN(n5008) );
  INV_X1 U3507 ( .A(n5018), .ZN(n3648) );
  INV_X1 U3508 ( .A(n4637), .ZN(n3566) );
  OAI21_X1 U3509 ( .B1(n5203), .B2(n3565), .A(n5205), .ZN(n4636) );
  INV_X1 U3510 ( .A(n5206), .ZN(n3565) );
  AOI21_X1 U3511 ( .B1(n3564), .B2(n5245), .A(n3563), .ZN(n5203) );
  INV_X1 U3512 ( .A(n5247), .ZN(n3563) );
  INV_X1 U3513 ( .A(n6086), .ZN(n3617) );
  OAI21_X1 U3514 ( .B1(n4069), .B2(n3616), .A(n4071), .ZN(n6084) );
  INV_X1 U3515 ( .A(n4072), .ZN(n3616) );
  AOI21_X1 U3516 ( .B1(n3615), .B2(n4084), .A(n3614), .ZN(n4069) );
  INV_X1 U3517 ( .A(n4086), .ZN(n3614) );
  INV_X1 U3518 ( .A(n5464), .ZN(n3583) );
  NOR2_X1 U3519 ( .A1(n7259), .A2(n3579), .ZN(n7193) );
  INV_X1 U3520 ( .A(n7257), .ZN(n3579) );
  AOI21_X1 U3521 ( .B1(n3581), .B2(n7256), .A(n3580), .ZN(n7194) );
  INV_X1 U3522 ( .A(n7260), .ZN(n3580) );
  INV_X1 U3523 ( .A(n6100), .ZN(n3634) );
  OAI21_X1 U3524 ( .B1(n7088), .B2(n3633), .A(n7090), .ZN(n6099) );
  INV_X1 U3525 ( .A(n7091), .ZN(n3633) );
  AOI21_X1 U3526 ( .B1(n3632), .B2(n7078), .A(n3631), .ZN(n7088) );
  INV_X1 U3527 ( .A(n7080), .ZN(n3631) );
  INV_X1 U3528 ( .A(n4183), .ZN(n3600) );
  OAI21_X1 U3529 ( .B1(n6764), .B2(n3599), .A(n6766), .ZN(n4182) );
  INV_X1 U3530 ( .A(n6767), .ZN(n3599) );
  AOI21_X1 U3531 ( .B1(n3598), .B2(n6745), .A(n3597), .ZN(n6764) );
  INV_X1 U3532 ( .A(n6748), .ZN(n3597) );
  NAND2_X1 U3533 ( .A1(n3511), .A2(n8719), .ZN(n3810) );
  OAI21_X1 U3534 ( .B1(n7194), .B2(n3582), .A(n7196), .ZN(n5463) );
  INV_X1 U3535 ( .A(n7197), .ZN(n3582) );
  AOI21_X1 U3536 ( .B1(n6227), .B2(n6226), .A(n6225), .ZN(n7996) );
  NAND2_X1 U3537 ( .A1(\adder_stage1[11][15] ), .A2(\adder_stage1[10][15] ), 
        .ZN(n8091) );
  NOR2_X1 U3538 ( .A1(\adder_stage1[11][15] ), .A2(\adder_stage1[10][15] ), 
        .ZN(n8092) );
  XNOR2_X1 U3539 ( .A(n3476), .B(n3451), .ZN(n3534) );
  NAND2_X1 U3540 ( .A1(n3521), .A2(n8696), .ZN(n3834) );
  NAND2_X1 U3541 ( .A1(xmem_full), .A2(n8716), .ZN(n3820) );
  NAND2_X1 U3542 ( .A1(fmem_addr[3]), .A2(n8579), .ZN(n8576) );
  AND2_X1 U3543 ( .A1(n3439), .A2(n3440), .ZN(n4098) );
  CLKBUF_X1 U3544 ( .A(n6123), .Z(n6213) );
  NOR2_X1 U3545 ( .A1(n5506), .A2(n3545), .ZN(n5535) );
  INV_X1 U3546 ( .A(n5505), .ZN(n3545) );
  NOR2_X1 U3547 ( .A1(n5017), .A2(n3647), .ZN(n5007) );
  INV_X1 U3548 ( .A(n5044), .ZN(n3647) );
  NOR2_X1 U3549 ( .A1(n5246), .A2(n3562), .ZN(n5202) );
  INV_X1 U3550 ( .A(n5289), .ZN(n3562) );
  NOR2_X1 U3551 ( .A1(n4085), .A2(n3613), .ZN(n4068) );
  INV_X1 U3552 ( .A(n4106), .ZN(n3613) );
  NOR2_X1 U3553 ( .A1(n7079), .A2(n3630), .ZN(n7087) );
  INV_X1 U3554 ( .A(n7106), .ZN(n3630) );
  NOR2_X1 U3555 ( .A1(n6747), .A2(n3596), .ZN(n6762) );
  INV_X1 U3556 ( .A(n6746), .ZN(n3596) );
  CLKBUF_X1 U3557 ( .A(n6590), .Z(n7120) );
  BUF_X1 U3558 ( .A(n4892), .Z(n5378) );
  NAND2_X1 U3559 ( .A1(n8579), .A2(n8712), .ZN(n8654) );
  NOR2_X1 U3560 ( .A1(n8676), .A2(n8576), .ZN(n8563) );
  NOR2_X1 U3561 ( .A1(n8576), .A2(n8685), .ZN(n8570) );
  INV_X1 U3562 ( .A(n8570), .ZN(n8571) );
  NOR2_X1 U3563 ( .A1(n8576), .A2(n8643), .ZN(n8574) );
  INV_X1 U3564 ( .A(n8574), .ZN(n8575) );
  NOR2_X1 U3565 ( .A1(n8576), .A2(n8601), .ZN(n8566) );
  INV_X1 U3566 ( .A(n8566), .ZN(n8567) );
  NOR2_X1 U3567 ( .A1(n8576), .A2(n8655), .ZN(n8577) );
  INV_X1 U3568 ( .A(n8577), .ZN(n8578) );
  NOR2_X1 U3569 ( .A1(n8576), .A2(n8632), .ZN(n8572) );
  INV_X1 U3570 ( .A(n8572), .ZN(n8573) );
  NOR2_X1 U3571 ( .A1(n8576), .A2(n8590), .ZN(n8564) );
  INV_X1 U3572 ( .A(n8564), .ZN(n8565) );
  NOR2_X1 U3573 ( .A1(n8576), .A2(n8612), .ZN(n8568) );
  INV_X1 U3574 ( .A(n8568), .ZN(n8569) );
  INV_X1 U3575 ( .A(n3657), .ZN(n6360) );
  OAI21_X1 U3576 ( .B1(n8281), .B2(n8274), .A(n8273), .ZN(n8275) );
  OR2_X1 U3577 ( .A1(n8268), .A2(n8270), .ZN(n8274) );
  INV_X1 U3578 ( .A(n8272), .ZN(n8273) );
  OAI21_X1 U3579 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8272) );
  INV_X1 U3580 ( .A(n7932), .ZN(n7935) );
  OAI21_X1 U3581 ( .B1(n8281), .B2(n8268), .A(n8271), .ZN(n7932) );
  NOR2_X1 U3582 ( .A1(n3510), .A2(n3986), .ZN(n3989) );
  CLKBUF_X1 U3583 ( .A(n8250), .Z(n3447) );
  CLKBUF_X1 U3584 ( .A(n4485), .Z(n3446) );
  OAI21_X1 U3585 ( .B1(n7996), .B2(n7995), .A(n7994), .ZN(n8007) );
  NAND2_X1 U3586 ( .A1(\adder_stage1[15][15] ), .A2(\adder_stage1[14][15] ), 
        .ZN(n7994) );
  NOR2_X1 U3587 ( .A1(\adder_stage1[15][15] ), .A2(\adder_stage1[14][15] ), 
        .ZN(n7995) );
  CLKBUF_X1 U3588 ( .A(n4290), .Z(n3438) );
  AOI21_X1 U3589 ( .B1(n5471), .B2(n5470), .A(n5469), .ZN(n8093) );
  NAND2_X1 U3590 ( .A1(\adder_stage1[0][15] ), .A2(\adder_stage1[1][15] ), 
        .ZN(n7955) );
  NOR2_X1 U3591 ( .A1(\adder_stage1[1][15] ), .A2(\adder_stage1[0][15] ), .ZN(
        n7956) );
  AOI21_X1 U3592 ( .B1(n4997), .B2(n3506), .A(n3549), .ZN(n3550) );
  AOI21_X1 U3593 ( .B1(n5536), .B2(n3469), .A(n4997), .ZN(n5000) );
  NAND2_X1 U3594 ( .A1(n5538), .A2(n5537), .ZN(n5542) );
  NAND2_X1 U3595 ( .A1(n5536), .A2(n5535), .ZN(n5538) );
  AOI21_X1 U3596 ( .B1(n5536), .B2(n5505), .A(n5504), .ZN(n5509) );
  AOI21_X1 U3597 ( .B1(n3871), .B2(n3504), .A(n3651), .ZN(n3652) );
  AOI21_X1 U3598 ( .B1(n5046), .B2(n3466), .A(n3871), .ZN(n3874) );
  NAND2_X1 U3599 ( .A1(n5009), .A2(n5008), .ZN(n5013) );
  NAND2_X1 U3600 ( .A1(n5046), .A2(n5007), .ZN(n5009) );
  AOI21_X1 U3601 ( .B1(n5046), .B2(n5044), .A(n5016), .ZN(n5020) );
  AOI21_X1 U3602 ( .B1(n4636), .B2(n3502), .A(n3566), .ZN(n3567) );
  AOI21_X1 U3603 ( .B1(n5291), .B2(n3468), .A(n4636), .ZN(n4639) );
  NAND2_X1 U3604 ( .A1(n5204), .A2(n5203), .ZN(n5208) );
  NAND2_X1 U3605 ( .A1(n5291), .A2(n5202), .ZN(n5204) );
  AOI21_X1 U3606 ( .B1(n5291), .B2(n5289), .A(n5245), .ZN(n5249) );
  AOI21_X1 U3607 ( .B1(n6084), .B2(n3507), .A(n3617), .ZN(n3618) );
  AOI21_X1 U3608 ( .B1(n6085), .B2(n3471), .A(n6084), .ZN(n6088) );
  NAND2_X1 U3609 ( .A1(n4070), .A2(n4069), .ZN(n4074) );
  NAND2_X1 U3610 ( .A1(n6085), .A2(n4068), .ZN(n4070) );
  AOI21_X1 U3611 ( .B1(n6085), .B2(n4106), .A(n4084), .ZN(n4088) );
  AOI21_X1 U3612 ( .B1(n5463), .B2(n3505), .A(n3583), .ZN(n3584) );
  NAND2_X1 U3613 ( .A1(n7195), .A2(n7194), .ZN(n7199) );
  NAND2_X1 U3614 ( .A1(n7258), .A2(n7193), .ZN(n7195) );
  AOI21_X1 U3615 ( .B1(n7258), .B2(n7257), .A(n7256), .ZN(n7262) );
  AOI21_X1 U3616 ( .B1(n6099), .B2(n3503), .A(n3634), .ZN(n3635) );
  AOI21_X1 U3617 ( .B1(n7108), .B2(n3472), .A(n6099), .ZN(n6102) );
  NAND2_X1 U3618 ( .A1(n7089), .A2(n7088), .ZN(n7093) );
  NAND2_X1 U3619 ( .A1(n7108), .A2(n7087), .ZN(n7089) );
  AOI21_X1 U3620 ( .B1(n7108), .B2(n7106), .A(n7078), .ZN(n7082) );
  CLKBUF_X1 U3621 ( .A(n7772), .Z(n3429) );
  AOI21_X1 U3622 ( .B1(n4182), .B2(n3501), .A(n3600), .ZN(n3601) );
  AOI21_X1 U3623 ( .B1(n6763), .B2(n3467), .A(n4182), .ZN(n4185) );
  NAND2_X1 U3624 ( .A1(n6765), .A2(n6764), .ZN(n6769) );
  NAND2_X1 U3625 ( .A1(n6763), .A2(n6762), .ZN(n6765) );
  AOI21_X1 U3626 ( .B1(n6763), .B2(n6746), .A(n6745), .ZN(n6750) );
  CLKBUF_X1 U3627 ( .A(n6975), .Z(n6980) );
  CLKBUF_X1 U3628 ( .A(n7420), .Z(n7446) );
  INV_X1 U3629 ( .A(n8689), .ZN(n8675) );
  INV_X1 U3630 ( .A(n8417), .ZN(n8418) );
  INV_X1 U3631 ( .A(n8427), .ZN(n8428) );
  INV_X1 U3632 ( .A(n8437), .ZN(n8438) );
  INV_X1 U3633 ( .A(n8447), .ZN(n8448) );
  INV_X1 U3634 ( .A(n8457), .ZN(n8458) );
  INV_X1 U3635 ( .A(n8467), .ZN(n8468) );
  INV_X1 U3636 ( .A(n8478), .ZN(n8479) );
  NOR2_X1 U3637 ( .A1(n8676), .A2(n8552), .ZN(n8489) );
  INV_X1 U3638 ( .A(n8489), .ZN(n8490) );
  NOR2_X1 U3639 ( .A1(n8590), .A2(n8552), .ZN(n8499) );
  INV_X1 U3640 ( .A(n8499), .ZN(n8500) );
  NOR2_X1 U3641 ( .A1(n8601), .A2(n8552), .ZN(n8509) );
  INV_X1 U3642 ( .A(n8509), .ZN(n8510) );
  NOR2_X1 U3643 ( .A1(n8612), .A2(n8552), .ZN(n8519) );
  INV_X1 U3644 ( .A(n8519), .ZN(n8520) );
  NOR2_X1 U3645 ( .A1(n8685), .A2(n8552), .ZN(n8529) );
  INV_X1 U3646 ( .A(n8529), .ZN(n8530) );
  NOR2_X1 U3647 ( .A1(n8632), .A2(n8552), .ZN(n8539) );
  INV_X1 U3648 ( .A(n8539), .ZN(n8540) );
  NOR2_X1 U3649 ( .A1(n8643), .A2(n8552), .ZN(n8549) );
  INV_X1 U3650 ( .A(n8549), .ZN(n8550) );
  NOR2_X1 U3651 ( .A1(n8655), .A2(n8552), .ZN(n8560) );
  INV_X1 U3652 ( .A(n8560), .ZN(n8561) );
  NOR2_X1 U3653 ( .A1(n8676), .A2(n8654), .ZN(n8587) );
  INV_X1 U3654 ( .A(n8587), .ZN(n8588) );
  NOR2_X1 U3655 ( .A1(n8590), .A2(n8654), .ZN(n8598) );
  INV_X1 U3656 ( .A(n8598), .ZN(n8599) );
  NOR2_X1 U3657 ( .A1(n8601), .A2(n8654), .ZN(n8609) );
  INV_X1 U3658 ( .A(n8609), .ZN(n8610) );
  NOR2_X1 U3659 ( .A1(n8612), .A2(n8654), .ZN(n8619) );
  INV_X1 U3660 ( .A(n8619), .ZN(n8620) );
  NOR2_X1 U3661 ( .A1(n8685), .A2(n8654), .ZN(n8629) );
  INV_X1 U3662 ( .A(n8629), .ZN(n8630) );
  NOR2_X1 U3663 ( .A1(n8632), .A2(n8654), .ZN(n8640) );
  INV_X1 U3664 ( .A(n8640), .ZN(n8641) );
  NOR2_X1 U3665 ( .A1(n8643), .A2(n8654), .ZN(n8651) );
  INV_X1 U3666 ( .A(n8651), .ZN(n8652) );
  NOR2_X1 U3667 ( .A1(n8655), .A2(n8654), .ZN(n8663) );
  INV_X1 U3668 ( .A(n8663), .ZN(n8664) );
  INV_X1 U3669 ( .A(n8563), .ZN(n8678) );
  NOR2_X1 U3670 ( .A1(n8667), .A2(n8666), .ZN(n8674) );
  NAND3_X1 U3671 ( .A1(n3824), .A2(n8688), .A3(n3822), .ZN(n8667) );
  NAND2_X1 U3672 ( .A1(s_valid_x), .A2(n3810), .ZN(n3811) );
  AOI21_X1 U3673 ( .B1(n3658), .B2(n8719), .A(n6360), .ZN(s_ready_x) );
  INV_X1 U3674 ( .A(n3425), .ZN(n3658) );
  AOI21_X1 U3675 ( .B1(n7258), .B2(n3470), .A(n5463), .ZN(n5466) );
  XNOR2_X1 U3676 ( .A(n7996), .B(n6228), .ZN(n6229) );
  XNOR2_X1 U3677 ( .A(n7917), .B(n3534), .ZN(n3535) );
  XNOR2_X1 U3678 ( .A(\x_mult_f[3][14] ), .B(\x_mult_f[2][14] ), .ZN(n5995) );
  AOI21_X1 U3679 ( .B1(n5341), .B2(n6975), .A(n5340), .ZN(n3427) );
  AOI21_X1 U3680 ( .B1(n5426), .B2(n7772), .A(n5425), .ZN(n3428) );
  AOI21_X2 U3681 ( .B1(n7132), .B2(n7130), .A(n5788), .ZN(n7163) );
  INV_X1 U3682 ( .A(n8348), .ZN(n3430) );
  OAI21_X1 U3683 ( .B1(n5446), .B2(n5442), .A(n5443), .ZN(n3431) );
  AOI21_X2 U3684 ( .B1(n8250), .B2(n8248), .A(n4225), .ZN(n5446) );
  NAND2_X1 U3685 ( .A1(n8122), .A2(n6256), .ZN(n3432) );
  AOI21_X1 U3686 ( .B1(n7190), .B2(n7188), .A(n5319), .ZN(n3433) );
  BUF_X4 U3687 ( .A(n3807), .Z(n8913) );
  AND2_X1 U3688 ( .A1(n8688), .A2(n8681), .ZN(n3434) );
  OR2_X1 U3689 ( .A1(\x_mult_f[2][3] ), .A2(\x_mult_f[3][3] ), .ZN(n3435) );
  AOI21_X1 U3690 ( .B1(n7414), .B2(n7412), .A(n3908), .ZN(n3436) );
  AOI21_X1 U3691 ( .B1(n4670), .B2(n4668), .A(n4263), .ZN(n3437) );
  XNOR2_X1 U3692 ( .A(n5996), .B(n5995), .ZN(n5997) );
  OAI21_X1 U3693 ( .B1(n6000), .B2(n6001), .A(n6002), .ZN(n5996) );
  XNOR2_X1 U3694 ( .A(n8093), .B(n5472), .ZN(n5473) );
  OAI21_X1 U3695 ( .B1(n3426), .B2(n8092), .A(n8091), .ZN(n8137) );
  AND2_X1 U3696 ( .A1(n3441), .A2(n3442), .ZN(n4153) );
  INV_X1 U3697 ( .A(n8348), .ZN(n3443) );
  AND2_X1 U3698 ( .A1(n3444), .A2(n3445), .ZN(n8297) );
  XNOR2_X1 U3699 ( .A(n3433), .B(n5320), .ZN(n5321) );
  OAI21_X1 U3700 ( .B1(n7957), .B2(n7956), .A(n7955), .ZN(n8120) );
  AOI21_X1 U3701 ( .B1(n7190), .B2(n7188), .A(n5319), .ZN(n7957) );
  NOR2_X1 U3702 ( .A1(n8470), .A2(n8612), .ZN(n8437) );
  NOR2_X1 U3703 ( .A1(n8470), .A2(n8632), .ZN(n8457) );
  NOR2_X1 U3704 ( .A1(n8470), .A2(n8590), .ZN(n8417) );
  NOR2_X1 U3705 ( .A1(n8470), .A2(n8655), .ZN(n8478) );
  NOR2_X1 U3706 ( .A1(n8470), .A2(n8643), .ZN(n8467) );
  NOR2_X1 U3707 ( .A1(n8470), .A2(n8601), .ZN(n8427) );
  NOR2_X1 U3708 ( .A1(n8470), .A2(n8685), .ZN(n8447) );
  NOR2_X1 U3709 ( .A1(fmem_addr[4]), .A2(n8682), .ZN(n8579) );
  INV_X1 U3710 ( .A(n8682), .ZN(n8681) );
  INV_X2 U3711 ( .A(n3809), .ZN(n8922) );
  INV_X2 U3712 ( .A(n3809), .ZN(n8923) );
  INV_X4 U3713 ( .A(n3808), .ZN(n3449) );
  BUF_X1 U3714 ( .A(n5447), .Z(n6917) );
  BUF_X1 U3715 ( .A(n5628), .Z(n5811) );
  INV_X1 U3716 ( .A(n6917), .ZN(n7825) );
  INV_X1 U3717 ( .A(n6917), .ZN(n7910) );
  INV_X1 U3718 ( .A(n6917), .ZN(n7244) );
  INV_X2 U3719 ( .A(n3809), .ZN(n8920) );
  BUF_X1 U3720 ( .A(n5628), .Z(n4715) );
  BUF_X1 U3721 ( .A(n5628), .Z(n6588) );
  INV_X2 U3722 ( .A(n3809), .ZN(n8921) );
  BUF_X1 U3723 ( .A(n5628), .Z(n4526) );
  BUF_X1 U3724 ( .A(n5628), .Z(n6736) );
  INV_X1 U3725 ( .A(n5628), .ZN(n7775) );
  INV_X1 U3726 ( .A(n5480), .ZN(n7767) );
  INV_X1 U3727 ( .A(n6105), .ZN(n8215) );
  INV_X1 U3728 ( .A(n6736), .ZN(n7613) );
  INV_X1 U3729 ( .A(n5628), .ZN(n8195) );
  INV_X1 U3730 ( .A(n4651), .ZN(n7851) );
  INV_X1 U3731 ( .A(n4651), .ZN(n5626) );
  INV_X1 U3732 ( .A(n6105), .ZN(n7793) );
  INV_X1 U3733 ( .A(n8356), .ZN(n8350) );
  INV_X1 U3734 ( .A(n5378), .ZN(n8046) );
  INV_X1 U3735 ( .A(n5628), .ZN(n8200) );
  INV_X1 U3736 ( .A(n4512), .ZN(n8395) );
  INV_X1 U3737 ( .A(n4512), .ZN(n8397) );
  OR2_X2 U3738 ( .A1(n8916), .A2(n3808), .ZN(n3452) );
  BUF_X1 U3739 ( .A(n5345), .Z(n8136) );
  BUF_X1 U3740 ( .A(n5345), .Z(n8141) );
  BUF_X1 U3741 ( .A(n4892), .Z(n6368) );
  BUF_X1 U3742 ( .A(n6122), .Z(n6105) );
  BUF_X1 U3743 ( .A(n3452), .Z(n5447) );
  BUF_X1 U3744 ( .A(n5447), .Z(n4512) );
  BUF_X1 U3745 ( .A(n4892), .Z(n5410) );
  AND2_X1 U3746 ( .A1(n5007), .A2(n5011), .ZN(n3466) );
  AND2_X1 U3747 ( .A1(n6762), .A2(n6767), .ZN(n3467) );
  AND2_X1 U3748 ( .A1(n5202), .A2(n5206), .ZN(n3468) );
  AND2_X1 U3749 ( .A1(n5535), .A2(n5540), .ZN(n3469) );
  AND2_X1 U3750 ( .A1(n7193), .A2(n7197), .ZN(n3470) );
  AND2_X1 U3751 ( .A1(n4068), .A2(n4072), .ZN(n3471) );
  AND2_X1 U3752 ( .A1(n7087), .A2(n7091), .ZN(n3472) );
  BUF_X1 U3753 ( .A(n8282), .Z(n5921) );
  BUF_X2 U3754 ( .A(n3807), .Z(n8917) );
  BUF_X2 U3755 ( .A(n3835), .Z(n8355) );
  INV_X1 U3756 ( .A(n5506), .ZN(n3547) );
  INV_X1 U3757 ( .A(n5246), .ZN(n3564) );
  INV_X1 U3758 ( .A(n7259), .ZN(n3581) );
  INV_X1 U3759 ( .A(n6747), .ZN(n3598) );
  INV_X1 U3760 ( .A(n4085), .ZN(n3615) );
  INV_X1 U3761 ( .A(n7079), .ZN(n3632) );
  INV_X1 U3762 ( .A(n5017), .ZN(n3649) );
  BUF_X1 U3763 ( .A(n4892), .Z(n5345) );
  BUF_X1 U3764 ( .A(n3452), .Z(n4892) );
  BUF_X1 U3765 ( .A(n3950), .Z(n4002) );
  BUF_X1 U3766 ( .A(n6435), .Z(n6699) );
  BUF_X1 U3767 ( .A(n6435), .Z(n6955) );
  BUF_X1 U3768 ( .A(n6435), .Z(n6645) );
  BUF_X1 U3769 ( .A(n6435), .Z(n6231) );
  XNOR2_X1 U3770 ( .A(\adder_stage3[3][20] ), .B(\adder_stage3[2][20] ), .ZN(
        n3499) );
  XNOR2_X1 U3771 ( .A(\adder_stage2[7][20] ), .B(\adder_stage2[6][20] ), .ZN(
        n3500) );
  OR2_X1 U3772 ( .A1(\x_mult_f[14][13] ), .A2(\x_mult_f[15][13] ), .ZN(n3501)
         );
  OR2_X1 U3773 ( .A1(\x_mult_f[24][13] ), .A2(\x_mult_f[25][13] ), .ZN(n3502)
         );
  OR2_X1 U3774 ( .A1(\x_mult_f[18][13] ), .A2(\x_mult_f[19][13] ), .ZN(n3503)
         );
  OR2_X1 U3775 ( .A1(\x_mult_f[26][13] ), .A2(\x_mult_f[27][13] ), .ZN(n3504)
         );
  OR2_X1 U3776 ( .A1(\x_mult_f[20][13] ), .A2(\x_mult_f[21][13] ), .ZN(n3505)
         );
  OR2_X1 U3777 ( .A1(\x_mult_f[28][13] ), .A2(\x_mult_f[29][13] ), .ZN(n3506)
         );
  OR2_X1 U3778 ( .A1(\x_mult_f[22][13] ), .A2(\x_mult_f[23][13] ), .ZN(n3507)
         );
  OR2_X1 U3779 ( .A1(\adder_stage3[2][13] ), .A2(\adder_stage3[3][13] ), .ZN(
        n3508) );
  AND2_X1 U3780 ( .A1(n3985), .A2(n3984), .ZN(n3510) );
  AND2_X1 U3781 ( .A1(n3469), .A2(n3506), .ZN(n3514) );
  AND2_X1 U3782 ( .A1(n3468), .A2(n3502), .ZN(n3515) );
  AND2_X1 U3783 ( .A1(n3470), .A2(n3505), .ZN(n3516) );
  AND2_X1 U3784 ( .A1(n3467), .A2(n3501), .ZN(n3517) );
  AND2_X1 U3785 ( .A1(n3471), .A2(n3507), .ZN(n3518) );
  AND2_X1 U3786 ( .A1(n3472), .A2(n3503), .ZN(n3519) );
  AND2_X1 U3787 ( .A1(n3466), .A2(n3504), .ZN(n3520) );
  NOR2_X1 U3788 ( .A1(n8911), .A2(n8912), .ZN(n3815) );
  INV_X1 U3789 ( .A(n8916), .ZN(n8348) );
  BUF_X2 U3790 ( .A(n3807), .Z(n8914) );
  NOR2_X1 U3791 ( .A1(\x_mult_f[2][2] ), .A2(\x_mult_f[3][2] ), .ZN(n7272) );
  NOR2_X1 U3792 ( .A1(\x_mult_f[2][3] ), .A2(\x_mult_f[3][3] ), .ZN(n6693) );
  NOR2_X1 U3793 ( .A1(n7272), .A2(n6693), .ZN(n3523) );
  NOR2_X1 U3794 ( .A1(\x_mult_f[2][1] ), .A2(\x_mult_f[3][1] ), .ZN(n7265) );
  NAND2_X1 U3795 ( .A1(\x_mult_f[2][0] ), .A2(\x_mult_f[3][0] ), .ZN(n7268) );
  NAND2_X1 U3796 ( .A1(\x_mult_f[2][1] ), .A2(\x_mult_f[3][1] ), .ZN(n7266) );
  OAI21_X1 U3797 ( .B1(n7265), .B2(n7268), .A(n7266), .ZN(n6692) );
  NAND2_X1 U3798 ( .A1(\x_mult_f[2][2] ), .A2(\x_mult_f[3][2] ), .ZN(n7273) );
  NAND2_X1 U3799 ( .A1(\x_mult_f[2][3] ), .A2(\x_mult_f[3][3] ), .ZN(n6694) );
  OAI21_X1 U3800 ( .B1(n6693), .B2(n7273), .A(n6694), .ZN(n3522) );
  AOI21_X1 U3801 ( .B1(n3523), .B2(n6692), .A(n3522), .ZN(n6685) );
  NOR2_X1 U3802 ( .A1(\x_mult_f[2][4] ), .A2(\x_mult_f[3][4] ), .ZN(n7208) );
  NOR2_X1 U3803 ( .A1(n7208), .A2(n7210), .ZN(n6687) );
  NOR2_X1 U3804 ( .A1(\x_mult_f[2][6] ), .A2(\x_mult_f[3][6] ), .ZN(n6715) );
  NOR2_X1 U3805 ( .A1(\x_mult_f[2][7] ), .A2(\x_mult_f[3][7] ), .ZN(n6717) );
  NOR2_X1 U3806 ( .A1(n6715), .A2(n6717), .ZN(n3525) );
  NAND2_X1 U3807 ( .A1(n6687), .A2(n3525), .ZN(n3527) );
  NAND2_X1 U3808 ( .A1(\x_mult_f[2][4] ), .A2(\x_mult_f[3][4] ), .ZN(n7246) );
  NAND2_X1 U3809 ( .A1(\x_mult_f[2][5] ), .A2(\x_mult_f[3][5] ), .ZN(n7211) );
  OAI21_X1 U3810 ( .B1(n7210), .B2(n7246), .A(n7211), .ZN(n6686) );
  NAND2_X1 U3811 ( .A1(\x_mult_f[2][6] ), .A2(\x_mult_f[3][6] ), .ZN(n6714) );
  NAND2_X1 U3812 ( .A1(\x_mult_f[2][7] ), .A2(\x_mult_f[3][7] ), .ZN(n6718) );
  OAI21_X1 U3813 ( .B1(n6717), .B2(n6714), .A(n6718), .ZN(n3524) );
  AOI21_X1 U3814 ( .B1(n3525), .B2(n6686), .A(n3524), .ZN(n3526) );
  OAI21_X1 U3815 ( .B1(n6685), .B2(n3527), .A(n3526), .ZN(n7282) );
  OR2_X1 U3816 ( .A1(\x_mult_f[2][8] ), .A2(\x_mult_f[3][8] ), .ZN(n7280) );
  NAND2_X1 U3817 ( .A1(\x_mult_f[2][8] ), .A2(\x_mult_f[3][8] ), .ZN(n7279) );
  INV_X1 U3818 ( .A(n7279), .ZN(n3528) );
  AOI21_X1 U3819 ( .B1(n7282), .B2(n7280), .A(n3528), .ZN(n6705) );
  NOR2_X1 U3820 ( .A1(\x_mult_f[2][9] ), .A2(\x_mult_f[3][9] ), .ZN(n6701) );
  NAND2_X1 U3821 ( .A1(\x_mult_f[2][9] ), .A2(\x_mult_f[3][9] ), .ZN(n6702) );
  OR2_X1 U3822 ( .A1(\x_mult_f[2][10] ), .A2(\x_mult_f[3][10] ), .ZN(n7113) );
  NAND2_X1 U3823 ( .A1(\x_mult_f[2][10] ), .A2(\x_mult_f[3][10] ), .ZN(n7112)
         );
  INV_X1 U3824 ( .A(n7112), .ZN(n3529) );
  AOI21_X1 U3825 ( .B1(n7115), .B2(n7113), .A(n3529), .ZN(n7102) );
  NOR2_X1 U3826 ( .A1(\x_mult_f[2][11] ), .A2(\x_mult_f[3][11] ), .ZN(n7098)
         );
  NAND2_X1 U3827 ( .A1(\x_mult_f[2][11] ), .A2(\x_mult_f[3][11] ), .ZN(n7099)
         );
  OR2_X1 U3828 ( .A1(\x_mult_f[2][12] ), .A2(\x_mult_f[3][12] ), .ZN(n7044) );
  NAND2_X1 U3829 ( .A1(\x_mult_f[2][12] ), .A2(\x_mult_f[3][12] ), .ZN(n7043)
         );
  INV_X1 U3830 ( .A(n7043), .ZN(n3530) );
  AOI21_X1 U3831 ( .B1(n7046), .B2(n7044), .A(n3530), .ZN(n6000) );
  NOR2_X1 U3832 ( .A1(\x_mult_f[2][13] ), .A2(\x_mult_f[3][13] ), .ZN(n6001)
         );
  NAND2_X1 U3833 ( .A1(\x_mult_f[2][13] ), .A2(\x_mult_f[3][13] ), .ZN(n6002)
         );
  NAND2_X1 U3834 ( .A1(n3509), .A2(n3473), .ZN(n3531) );
  NAND2_X1 U3835 ( .A1(n5996), .A2(n3531), .ZN(n3533) );
  NAND2_X1 U3836 ( .A1(\x_mult_f[3][14] ), .A2(\x_mult_f[2][14] ), .ZN(n3532)
         );
  NAND2_X1 U3837 ( .A1(n3533), .A2(n3532), .ZN(n7917) );
  NAND2_X1 U3838 ( .A1(n3535), .A2(n8265), .ZN(n3537) );
  BUF_X2 U3839 ( .A(n3807), .Z(n8916) );
  NAND2_X1 U3840 ( .A1(n8364), .A2(\adder_stage1[1][15] ), .ZN(n3536) );
  NAND2_X1 U3841 ( .A1(n3537), .A2(n3536), .ZN(n10038) );
  NOR2_X1 U3842 ( .A1(\x_mult_f[28][1] ), .A2(\x_mult_f[29][1] ), .ZN(n4599)
         );
  NAND2_X1 U3843 ( .A1(\x_mult_f[28][0] ), .A2(\x_mult_f[29][0] ), .ZN(n4602)
         );
  NAND2_X1 U3844 ( .A1(\x_mult_f[28][1] ), .A2(\x_mult_f[29][1] ), .ZN(n4600)
         );
  OAI21_X1 U3845 ( .B1(n4599), .B2(n4602), .A(n4600), .ZN(n4587) );
  NOR2_X1 U3846 ( .A1(\x_mult_f[28][2] ), .A2(\x_mult_f[29][2] ), .ZN(n5076)
         );
  NOR2_X1 U3847 ( .A1(\x_mult_f[28][3] ), .A2(\x_mult_f[29][3] ), .ZN(n5078)
         );
  NOR2_X1 U3848 ( .A1(n5076), .A2(n5078), .ZN(n3539) );
  NAND2_X1 U3849 ( .A1(\x_mult_f[28][2] ), .A2(\x_mult_f[29][2] ), .ZN(n5075)
         );
  NAND2_X1 U3850 ( .A1(\x_mult_f[28][3] ), .A2(\x_mult_f[29][3] ), .ZN(n5079)
         );
  OAI21_X1 U3851 ( .B1(n5078), .B2(n5075), .A(n5079), .ZN(n3538) );
  AOI21_X1 U3852 ( .B1(n4587), .B2(n3539), .A(n3538), .ZN(n5065) );
  NOR2_X1 U3853 ( .A1(\x_mult_f[28][4] ), .A2(\x_mult_f[29][4] ), .ZN(n5066)
         );
  NOR2_X1 U3854 ( .A1(\x_mult_f[28][5] ), .A2(\x_mult_f[29][5] ), .ZN(n5068)
         );
  NOR2_X1 U3855 ( .A1(n5066), .A2(n5068), .ZN(n5498) );
  NOR2_X1 U3856 ( .A1(\x_mult_f[28][6] ), .A2(\x_mult_f[29][6] ), .ZN(n5520)
         );
  NOR2_X1 U3857 ( .A1(\x_mult_f[28][7] ), .A2(\x_mult_f[29][7] ), .ZN(n5522)
         );
  NOR2_X1 U3858 ( .A1(n5520), .A2(n5522), .ZN(n3541) );
  NAND2_X1 U3859 ( .A1(n5498), .A2(n3541), .ZN(n3543) );
  NAND2_X1 U3860 ( .A1(\x_mult_f[28][4] ), .A2(\x_mult_f[29][4] ), .ZN(n5085)
         );
  NAND2_X1 U3861 ( .A1(\x_mult_f[28][5] ), .A2(\x_mult_f[29][5] ), .ZN(n5069)
         );
  OAI21_X1 U3862 ( .B1(n5068), .B2(n5085), .A(n5069), .ZN(n5497) );
  NAND2_X1 U3863 ( .A1(\x_mult_f[28][6] ), .A2(\x_mult_f[29][6] ), .ZN(n5519)
         );
  NAND2_X1 U3864 ( .A1(\x_mult_f[28][7] ), .A2(\x_mult_f[29][7] ), .ZN(n5523)
         );
  OAI21_X1 U3865 ( .B1(n5522), .B2(n5519), .A(n5523), .ZN(n3540) );
  AOI21_X1 U3866 ( .B1(n3541), .B2(n5497), .A(n3540), .ZN(n3542) );
  OAI21_X1 U3867 ( .B1(n5065), .B2(n3543), .A(n3542), .ZN(n5532) );
  OR2_X1 U3868 ( .A1(\x_mult_f[28][8] ), .A2(\x_mult_f[29][8] ), .ZN(n5530) );
  NAND2_X1 U3869 ( .A1(\x_mult_f[28][8] ), .A2(\x_mult_f[29][8] ), .ZN(n5529)
         );
  INV_X1 U3870 ( .A(n5529), .ZN(n3544) );
  AOI21_X1 U3871 ( .B1(n5532), .B2(n5530), .A(n3544), .ZN(n5516) );
  NOR2_X1 U3872 ( .A1(\x_mult_f[28][9] ), .A2(\x_mult_f[29][9] ), .ZN(n5512)
         );
  NAND2_X1 U3873 ( .A1(\x_mult_f[28][9] ), .A2(\x_mult_f[29][9] ), .ZN(n5513)
         );
  OAI21_X1 U3874 ( .B1(n5516), .B2(n5512), .A(n5513), .ZN(n5536) );
  NOR2_X1 U3875 ( .A1(\x_mult_f[28][11] ), .A2(\x_mult_f[29][11] ), .ZN(n5506)
         );
  OR2_X1 U3876 ( .A1(\x_mult_f[28][10] ), .A2(\x_mult_f[29][10] ), .ZN(n5505)
         );
  OR2_X1 U3877 ( .A1(\x_mult_f[28][12] ), .A2(\x_mult_f[29][12] ), .ZN(n5540)
         );
  NAND2_X1 U3878 ( .A1(n5536), .A2(n3514), .ZN(n3551) );
  NAND2_X1 U3879 ( .A1(\x_mult_f[28][10] ), .A2(\x_mult_f[29][10] ), .ZN(n5493) );
  INV_X1 U3880 ( .A(n5493), .ZN(n5504) );
  NAND2_X1 U3881 ( .A1(\x_mult_f[28][11] ), .A2(\x_mult_f[29][11] ), .ZN(n5507) );
  NAND2_X1 U3882 ( .A1(\x_mult_f[28][12] ), .A2(\x_mult_f[29][12] ), .ZN(n5539) );
  NAND2_X1 U3883 ( .A1(\x_mult_f[28][13] ), .A2(\x_mult_f[29][13] ), .ZN(n4998) );
  NAND2_X1 U3884 ( .A1(n3551), .A2(n3550), .ZN(n5991) );
  NAND2_X1 U3885 ( .A1(n3552), .A2(n4596), .ZN(n3554) );
  INV_X2 U3886 ( .A(n6368), .ZN(n7944) );
  NAND2_X1 U3887 ( .A1(n7944), .A2(\adder_stage1[14][15] ), .ZN(n3553) );
  NAND2_X1 U3888 ( .A1(n3554), .A2(n3553), .ZN(n9824) );
  NOR2_X1 U3889 ( .A1(\x_mult_f[24][1] ), .A2(\x_mult_f[25][1] ), .ZN(n4729)
         );
  NAND2_X1 U3890 ( .A1(\x_mult_f[24][0] ), .A2(\x_mult_f[25][0] ), .ZN(n4735)
         );
  NAND2_X1 U3891 ( .A1(\x_mult_f[24][1] ), .A2(\x_mult_f[25][1] ), .ZN(n4730)
         );
  OAI21_X1 U3892 ( .B1(n4729), .B2(n4735), .A(n4730), .ZN(n5252) );
  NOR2_X1 U3893 ( .A1(\x_mult_f[24][2] ), .A2(\x_mult_f[25][2] ), .ZN(n5267)
         );
  NOR2_X1 U3894 ( .A1(\x_mult_f[24][3] ), .A2(\x_mult_f[25][3] ), .ZN(n5253)
         );
  NOR2_X1 U3895 ( .A1(n5267), .A2(n5253), .ZN(n3556) );
  NAND2_X1 U3896 ( .A1(\x_mult_f[24][2] ), .A2(\x_mult_f[25][2] ), .ZN(n5268)
         );
  NAND2_X1 U3897 ( .A1(\x_mult_f[24][3] ), .A2(\x_mult_f[25][3] ), .ZN(n5254)
         );
  OAI21_X1 U3898 ( .B1(n5253), .B2(n5268), .A(n5254), .ZN(n3555) );
  AOI21_X1 U3899 ( .B1(n5252), .B2(n3556), .A(n3555), .ZN(n5211) );
  NOR2_X1 U3900 ( .A1(\x_mult_f[24][4] ), .A2(\x_mult_f[25][4] ), .ZN(n5212)
         );
  NOR2_X1 U3901 ( .A1(\x_mult_f[24][5] ), .A2(\x_mult_f[25][5] ), .ZN(n5214)
         );
  NOR2_X1 U3902 ( .A1(n5212), .A2(n5214), .ZN(n5231) );
  NOR2_X1 U3903 ( .A1(\x_mult_f[24][6] ), .A2(\x_mult_f[25][6] ), .ZN(n5281)
         );
  NOR2_X1 U3904 ( .A1(\x_mult_f[24][7] ), .A2(\x_mult_f[25][7] ), .ZN(n5232)
         );
  NOR2_X1 U3905 ( .A1(n5281), .A2(n5232), .ZN(n3558) );
  NAND2_X1 U3906 ( .A1(n5231), .A2(n3558), .ZN(n3560) );
  NAND2_X1 U3907 ( .A1(\x_mult_f[24][4] ), .A2(\x_mult_f[25][4] ), .ZN(n5275)
         );
  NAND2_X1 U3908 ( .A1(\x_mult_f[24][5] ), .A2(\x_mult_f[25][5] ), .ZN(n5215)
         );
  OAI21_X1 U3909 ( .B1(n5214), .B2(n5275), .A(n5215), .ZN(n5230) );
  NAND2_X1 U3910 ( .A1(\x_mult_f[24][6] ), .A2(\x_mult_f[25][6] ), .ZN(n5282)
         );
  NAND2_X1 U3911 ( .A1(\x_mult_f[24][7] ), .A2(\x_mult_f[25][7] ), .ZN(n5233)
         );
  OAI21_X1 U3912 ( .B1(n5232), .B2(n5282), .A(n5233), .ZN(n3557) );
  AOI21_X1 U3913 ( .B1(n3558), .B2(n5230), .A(n3557), .ZN(n3559) );
  OAI21_X1 U3914 ( .B1(n5211), .B2(n3560), .A(n3559), .ZN(n5242) );
  OR2_X1 U3915 ( .A1(\x_mult_f[24][8] ), .A2(\x_mult_f[25][8] ), .ZN(n5240) );
  NAND2_X1 U3916 ( .A1(\x_mult_f[24][8] ), .A2(\x_mult_f[25][8] ), .ZN(n5239)
         );
  INV_X1 U3917 ( .A(n5239), .ZN(n3561) );
  AOI21_X1 U3918 ( .B1(n5242), .B2(n5240), .A(n3561), .ZN(n5264) );
  NOR2_X1 U3919 ( .A1(\x_mult_f[24][9] ), .A2(\x_mult_f[25][9] ), .ZN(n5260)
         );
  NAND2_X1 U3920 ( .A1(\x_mult_f[24][9] ), .A2(\x_mult_f[25][9] ), .ZN(n5261)
         );
  OAI21_X1 U3921 ( .B1(n5264), .B2(n5260), .A(n5261), .ZN(n5291) );
  NOR2_X1 U3922 ( .A1(\x_mult_f[24][11] ), .A2(\x_mult_f[25][11] ), .ZN(n5246)
         );
  OR2_X1 U3923 ( .A1(\x_mult_f[24][10] ), .A2(\x_mult_f[25][10] ), .ZN(n5289)
         );
  OR2_X1 U3924 ( .A1(\x_mult_f[24][12] ), .A2(\x_mult_f[25][12] ), .ZN(n5206)
         );
  NAND2_X1 U3925 ( .A1(n5291), .A2(n3515), .ZN(n3568) );
  NAND2_X1 U3926 ( .A1(\x_mult_f[24][10] ), .A2(\x_mult_f[25][10] ), .ZN(n5288) );
  INV_X1 U3927 ( .A(n5288), .ZN(n5245) );
  NAND2_X1 U3928 ( .A1(\x_mult_f[24][11] ), .A2(\x_mult_f[25][11] ), .ZN(n5247) );
  NAND2_X1 U3929 ( .A1(\x_mult_f[24][12] ), .A2(\x_mult_f[25][12] ), .ZN(n5205) );
  NAND2_X1 U3930 ( .A1(\x_mult_f[24][13] ), .A2(\x_mult_f[25][13] ), .ZN(n4637) );
  NAND2_X1 U3931 ( .A1(n3568), .A2(n3567), .ZN(n5439) );
  NAND2_X1 U3932 ( .A1(n3569), .A2(n8189), .ZN(n3571) );
  NAND2_X1 U3933 ( .A1(n7825), .A2(\adder_stage1[12][15] ), .ZN(n3570) );
  NAND2_X1 U3934 ( .A1(n3571), .A2(n3570), .ZN(n9858) );
  NOR2_X1 U3935 ( .A1(\x_mult_f[20][1] ), .A2(\x_mult_f[21][1] ), .ZN(n4875)
         );
  NAND2_X1 U3936 ( .A1(\x_mult_f[20][0] ), .A2(\x_mult_f[21][0] ), .ZN(n4881)
         );
  NAND2_X1 U3937 ( .A1(\x_mult_f[20][1] ), .A2(\x_mult_f[21][1] ), .ZN(n4876)
         );
  OAI21_X1 U3938 ( .B1(n4875), .B2(n4881), .A(n4876), .ZN(n4841) );
  NOR2_X1 U3939 ( .A1(\x_mult_f[20][2] ), .A2(\x_mult_f[21][2] ), .ZN(n4885)
         );
  NOR2_X1 U3940 ( .A1(\x_mult_f[20][3] ), .A2(\x_mult_f[21][3] ), .ZN(n4842)
         );
  NOR2_X1 U3941 ( .A1(n4885), .A2(n4842), .ZN(n3573) );
  NAND2_X1 U3942 ( .A1(\x_mult_f[20][2] ), .A2(\x_mult_f[21][2] ), .ZN(n4886)
         );
  NAND2_X1 U3943 ( .A1(\x_mult_f[20][3] ), .A2(\x_mult_f[21][3] ), .ZN(n4843)
         );
  OAI21_X1 U3944 ( .B1(n4842), .B2(n4886), .A(n4843), .ZN(n3572) );
  AOI21_X1 U3945 ( .B1(n4841), .B2(n3573), .A(n3572), .ZN(n4851) );
  NOR2_X1 U3946 ( .A1(\x_mult_f[20][4] ), .A2(\x_mult_f[21][4] ), .ZN(n4852)
         );
  NOR2_X1 U3947 ( .A1(\x_mult_f[20][5] ), .A2(\x_mult_f[21][5] ), .ZN(n4854)
         );
  NOR2_X1 U3948 ( .A1(n4852), .A2(n4854), .ZN(n4863) );
  NOR2_X1 U3949 ( .A1(\x_mult_f[20][6] ), .A2(\x_mult_f[21][6] ), .ZN(n6375)
         );
  NOR2_X1 U3950 ( .A1(\x_mult_f[20][7] ), .A2(\x_mult_f[21][7] ), .ZN(n6377)
         );
  NOR2_X1 U3951 ( .A1(n6375), .A2(n6377), .ZN(n3575) );
  NAND2_X1 U3952 ( .A1(n4863), .A2(n3575), .ZN(n3577) );
  NAND2_X1 U3953 ( .A1(\x_mult_f[20][4] ), .A2(\x_mult_f[21][4] ), .ZN(n4868)
         );
  NAND2_X1 U3954 ( .A1(\x_mult_f[20][5] ), .A2(\x_mult_f[21][5] ), .ZN(n4855)
         );
  OAI21_X1 U3955 ( .B1(n4854), .B2(n4868), .A(n4855), .ZN(n4862) );
  NAND2_X1 U3956 ( .A1(\x_mult_f[20][6] ), .A2(\x_mult_f[21][6] ), .ZN(n6374)
         );
  NAND2_X1 U3957 ( .A1(\x_mult_f[20][7] ), .A2(\x_mult_f[21][7] ), .ZN(n6378)
         );
  OAI21_X1 U3958 ( .B1(n6377), .B2(n6374), .A(n6378), .ZN(n3574) );
  AOI21_X1 U3959 ( .B1(n3575), .B2(n4862), .A(n3574), .ZN(n3576) );
  OAI21_X1 U3960 ( .B1(n4851), .B2(n3577), .A(n3576), .ZN(n7205) );
  OR2_X1 U3961 ( .A1(\x_mult_f[20][8] ), .A2(\x_mult_f[21][8] ), .ZN(n7203) );
  NAND2_X1 U3962 ( .A1(\x_mult_f[20][8] ), .A2(\x_mult_f[21][8] ), .ZN(n7202)
         );
  INV_X1 U3963 ( .A(n7202), .ZN(n3578) );
  AOI21_X1 U3964 ( .B1(n7205), .B2(n7203), .A(n3578), .ZN(n7221) );
  NOR2_X1 U3965 ( .A1(\x_mult_f[20][9] ), .A2(\x_mult_f[21][9] ), .ZN(n7217)
         );
  NAND2_X1 U3966 ( .A1(\x_mult_f[20][9] ), .A2(\x_mult_f[21][9] ), .ZN(n7218)
         );
  OAI21_X1 U3967 ( .B1(n7221), .B2(n7217), .A(n7218), .ZN(n7258) );
  NOR2_X1 U3968 ( .A1(\x_mult_f[20][11] ), .A2(\x_mult_f[21][11] ), .ZN(n7259)
         );
  OR2_X1 U3969 ( .A1(\x_mult_f[20][10] ), .A2(\x_mult_f[21][10] ), .ZN(n7257)
         );
  OR2_X1 U3970 ( .A1(\x_mult_f[20][12] ), .A2(\x_mult_f[21][12] ), .ZN(n7197)
         );
  NAND2_X1 U3971 ( .A1(n7258), .A2(n3516), .ZN(n3585) );
  NAND2_X1 U3972 ( .A1(\x_mult_f[20][10] ), .A2(\x_mult_f[21][10] ), .ZN(n7252) );
  INV_X1 U3973 ( .A(n7252), .ZN(n7256) );
  NAND2_X1 U3974 ( .A1(\x_mult_f[20][11] ), .A2(\x_mult_f[21][11] ), .ZN(n7260) );
  NAND2_X1 U3975 ( .A1(\x_mult_f[20][12] ), .A2(\x_mult_f[21][12] ), .ZN(n7196) );
  NAND2_X1 U3976 ( .A1(\x_mult_f[20][13] ), .A2(\x_mult_f[21][13] ), .ZN(n5464) );
  NAND2_X1 U3977 ( .A1(n3585), .A2(n3584), .ZN(n5949) );
  BUF_X2 U3978 ( .A(n8282), .Z(n8401) );
  NAND2_X1 U3979 ( .A1(n3586), .A2(n8401), .ZN(n3588) );
  NAND2_X1 U3980 ( .A1(n8395), .A2(\adder_stage1[10][15] ), .ZN(n3587) );
  NAND2_X1 U3981 ( .A1(n3588), .A2(n3587), .ZN(n9891) );
  NOR2_X1 U3982 ( .A1(\x_mult_f[14][1] ), .A2(\x_mult_f[15][1] ), .ZN(n5632)
         );
  NAND2_X1 U3983 ( .A1(\x_mult_f[14][0] ), .A2(\x_mult_f[15][0] ), .ZN(n5635)
         );
  NAND2_X1 U3984 ( .A1(\x_mult_f[14][1] ), .A2(\x_mult_f[15][1] ), .ZN(n5633)
         );
  OAI21_X1 U3985 ( .B1(n5632), .B2(n5635), .A(n5633), .ZN(n5649) );
  NOR2_X1 U3986 ( .A1(\x_mult_f[14][2] ), .A2(\x_mult_f[15][2] ), .ZN(n6549)
         );
  NOR2_X1 U3987 ( .A1(\x_mult_f[14][3] ), .A2(\x_mult_f[15][3] ), .ZN(n5650)
         );
  NOR2_X1 U3988 ( .A1(n6549), .A2(n5650), .ZN(n3590) );
  NAND2_X1 U3989 ( .A1(\x_mult_f[14][2] ), .A2(\x_mult_f[15][2] ), .ZN(n6550)
         );
  NAND2_X1 U3990 ( .A1(\x_mult_f[14][3] ), .A2(\x_mult_f[15][3] ), .ZN(n5651)
         );
  OAI21_X1 U3991 ( .B1(n5650), .B2(n6550), .A(n5651), .ZN(n3589) );
  AOI21_X1 U3992 ( .B1(n5649), .B2(n3590), .A(n3589), .ZN(n5639) );
  NOR2_X1 U3993 ( .A1(\x_mult_f[14][4] ), .A2(\x_mult_f[15][4] ), .ZN(n5640)
         );
  NOR2_X1 U3994 ( .A1(\x_mult_f[14][5] ), .A2(\x_mult_f[15][5] ), .ZN(n5642)
         );
  NOR2_X1 U3995 ( .A1(n5640), .A2(n5642), .ZN(n6557) );
  NOR2_X1 U3996 ( .A1(\x_mult_f[14][6] ), .A2(\x_mult_f[15][6] ), .ZN(n6635)
         );
  NOR2_X1 U3997 ( .A1(\x_mult_f[14][7] ), .A2(\x_mult_f[15][7] ), .ZN(n6637)
         );
  NOR2_X1 U3998 ( .A1(n6635), .A2(n6637), .ZN(n3592) );
  NAND2_X1 U3999 ( .A1(n6557), .A2(n3592), .ZN(n3594) );
  NAND2_X1 U4000 ( .A1(\x_mult_f[14][4] ), .A2(\x_mult_f[15][4] ), .ZN(n5657)
         );
  NAND2_X1 U4001 ( .A1(\x_mult_f[14][5] ), .A2(\x_mult_f[15][5] ), .ZN(n5643)
         );
  OAI21_X1 U4002 ( .B1(n5642), .B2(n5657), .A(n5643), .ZN(n6556) );
  NAND2_X1 U4003 ( .A1(\x_mult_f[14][6] ), .A2(\x_mult_f[15][6] ), .ZN(n6634)
         );
  NAND2_X1 U4004 ( .A1(\x_mult_f[14][7] ), .A2(\x_mult_f[15][7] ), .ZN(n6638)
         );
  OAI21_X1 U4005 ( .B1(n6637), .B2(n6634), .A(n6638), .ZN(n3591) );
  AOI21_X1 U4006 ( .B1(n3592), .B2(n6556), .A(n3591), .ZN(n3593) );
  OAI21_X1 U4007 ( .B1(n5639), .B2(n3594), .A(n3593), .ZN(n6631) );
  OR2_X1 U4008 ( .A1(\x_mult_f[14][8] ), .A2(\x_mult_f[15][8] ), .ZN(n6629) );
  NAND2_X1 U4009 ( .A1(\x_mult_f[14][8] ), .A2(\x_mult_f[15][8] ), .ZN(n6628)
         );
  INV_X1 U4010 ( .A(n6628), .ZN(n3595) );
  AOI21_X1 U4011 ( .B1(n6631), .B2(n6629), .A(n3595), .ZN(n6758) );
  NOR2_X1 U4012 ( .A1(\x_mult_f[14][9] ), .A2(\x_mult_f[15][9] ), .ZN(n6754)
         );
  NAND2_X1 U4013 ( .A1(\x_mult_f[14][9] ), .A2(\x_mult_f[15][9] ), .ZN(n6755)
         );
  OAI21_X1 U4014 ( .B1(n6758), .B2(n6754), .A(n6755), .ZN(n6763) );
  NOR2_X1 U4015 ( .A1(\x_mult_f[14][11] ), .A2(\x_mult_f[15][11] ), .ZN(n6747)
         );
  OR2_X1 U4016 ( .A1(\x_mult_f[14][10] ), .A2(\x_mult_f[15][10] ), .ZN(n6746)
         );
  OR2_X1 U4017 ( .A1(\x_mult_f[14][12] ), .A2(\x_mult_f[15][12] ), .ZN(n6767)
         );
  NAND2_X1 U4018 ( .A1(n6763), .A2(n3517), .ZN(n3602) );
  NAND2_X1 U4019 ( .A1(\x_mult_f[14][10] ), .A2(\x_mult_f[15][10] ), .ZN(n6740) );
  INV_X1 U4020 ( .A(n6740), .ZN(n6745) );
  NAND2_X1 U4021 ( .A1(\x_mult_f[14][11] ), .A2(\x_mult_f[15][11] ), .ZN(n6748) );
  NAND2_X1 U4022 ( .A1(\x_mult_f[14][12] ), .A2(\x_mult_f[15][12] ), .ZN(n6766) );
  NAND2_X1 U4023 ( .A1(\x_mult_f[14][13] ), .A2(\x_mult_f[15][13] ), .ZN(n4183) );
  NAND2_X1 U4024 ( .A1(n3602), .A2(n3601), .ZN(n5911) );
  NAND2_X1 U4025 ( .A1(n3603), .A2(n8180), .ZN(n3605) );
  INV_X2 U4026 ( .A(n5345), .ZN(n8059) );
  NAND2_X1 U4027 ( .A1(n8059), .A2(\adder_stage1[7][15] ), .ZN(n3604) );
  NAND2_X1 U4028 ( .A1(n3605), .A2(n3604), .ZN(n9940) );
  NOR2_X1 U4029 ( .A1(\x_mult_f[22][1] ), .A2(\x_mult_f[23][1] ), .ZN(n4440)
         );
  NAND2_X1 U4030 ( .A1(\x_mult_f[22][0] ), .A2(\x_mult_f[23][0] ), .ZN(n4443)
         );
  NAND2_X1 U4031 ( .A1(\x_mult_f[22][1] ), .A2(\x_mult_f[23][1] ), .ZN(n4441)
         );
  OAI21_X1 U4032 ( .B1(n4440), .B2(n4443), .A(n4441), .ZN(n4447) );
  NOR2_X1 U4033 ( .A1(\x_mult_f[22][2] ), .A2(\x_mult_f[23][2] ), .ZN(n4622)
         );
  NOR2_X1 U4034 ( .A1(\x_mult_f[22][3] ), .A2(\x_mult_f[23][3] ), .ZN(n4448)
         );
  NOR2_X1 U4035 ( .A1(n4622), .A2(n4448), .ZN(n3607) );
  NAND2_X1 U4036 ( .A1(\x_mult_f[22][2] ), .A2(\x_mult_f[23][2] ), .ZN(n4623)
         );
  NAND2_X1 U4037 ( .A1(\x_mult_f[22][3] ), .A2(\x_mult_f[23][3] ), .ZN(n4449)
         );
  OAI21_X1 U4038 ( .B1(n4448), .B2(n4623), .A(n4449), .ZN(n3606) );
  AOI21_X1 U4039 ( .B1(n4447), .B2(n3607), .A(n3606), .ZN(n3969) );
  NOR2_X1 U4040 ( .A1(\x_mult_f[22][4] ), .A2(\x_mult_f[23][4] ), .ZN(n4433)
         );
  NOR2_X1 U4041 ( .A1(\x_mult_f[22][5] ), .A2(\x_mult_f[23][5] ), .ZN(n4462)
         );
  NOR2_X1 U4042 ( .A1(n4433), .A2(n4462), .ZN(n3971) );
  NOR2_X1 U4043 ( .A1(\x_mult_f[22][6] ), .A2(\x_mult_f[23][6] ), .ZN(n4518)
         );
  NOR2_X1 U4044 ( .A1(\x_mult_f[22][7] ), .A2(\x_mult_f[23][7] ), .ZN(n3972)
         );
  NOR2_X1 U4045 ( .A1(n4518), .A2(n3972), .ZN(n3609) );
  NAND2_X1 U4046 ( .A1(n3971), .A2(n3609), .ZN(n3611) );
  NAND2_X1 U4047 ( .A1(\x_mult_f[22][4] ), .A2(\x_mult_f[23][4] ), .ZN(n4458)
         );
  NAND2_X1 U4048 ( .A1(\x_mult_f[22][5] ), .A2(\x_mult_f[23][5] ), .ZN(n4463)
         );
  OAI21_X1 U4049 ( .B1(n4462), .B2(n4458), .A(n4463), .ZN(n3970) );
  NAND2_X1 U4050 ( .A1(\x_mult_f[22][6] ), .A2(\x_mult_f[23][6] ), .ZN(n4519)
         );
  NAND2_X1 U4051 ( .A1(\x_mult_f[22][7] ), .A2(\x_mult_f[23][7] ), .ZN(n3973)
         );
  OAI21_X1 U4052 ( .B1(n3972), .B2(n4519), .A(n3973), .ZN(n3608) );
  AOI21_X1 U4053 ( .B1(n3609), .B2(n3970), .A(n3608), .ZN(n3610) );
  OAI21_X1 U4054 ( .B1(n3969), .B2(n3611), .A(n3610), .ZN(n4137) );
  OR2_X1 U4055 ( .A1(\x_mult_f[22][8] ), .A2(\x_mult_f[23][8] ), .ZN(n4135) );
  NAND2_X1 U4056 ( .A1(\x_mult_f[22][8] ), .A2(\x_mult_f[23][8] ), .ZN(n4134)
         );
  INV_X1 U4057 ( .A(n4134), .ZN(n3612) );
  AOI21_X1 U4058 ( .B1(n4137), .B2(n4135), .A(n3612), .ZN(n4114) );
  NOR2_X1 U4059 ( .A1(\x_mult_f[22][9] ), .A2(\x_mult_f[23][9] ), .ZN(n4110)
         );
  NAND2_X1 U4060 ( .A1(\x_mult_f[22][9] ), .A2(\x_mult_f[23][9] ), .ZN(n4111)
         );
  OAI21_X1 U4061 ( .B1(n4114), .B2(n4110), .A(n4111), .ZN(n6085) );
  NOR2_X1 U4062 ( .A1(\x_mult_f[22][11] ), .A2(\x_mult_f[23][11] ), .ZN(n4085)
         );
  OR2_X1 U4063 ( .A1(\x_mult_f[22][10] ), .A2(\x_mult_f[23][10] ), .ZN(n4106)
         );
  OR2_X1 U4064 ( .A1(\x_mult_f[22][12] ), .A2(\x_mult_f[23][12] ), .ZN(n4072)
         );
  NAND2_X1 U4065 ( .A1(n6085), .A2(n3518), .ZN(n3619) );
  NAND2_X1 U4066 ( .A1(\x_mult_f[22][10] ), .A2(\x_mult_f[23][10] ), .ZN(n4105) );
  INV_X1 U4067 ( .A(n4105), .ZN(n4084) );
  NAND2_X1 U4068 ( .A1(\x_mult_f[22][11] ), .A2(\x_mult_f[23][11] ), .ZN(n4086) );
  NAND2_X1 U4069 ( .A1(\x_mult_f[22][12] ), .A2(\x_mult_f[23][12] ), .ZN(n4071) );
  NAND2_X1 U4070 ( .A1(\x_mult_f[22][13] ), .A2(\x_mult_f[23][13] ), .ZN(n6086) );
  NAND2_X1 U4071 ( .A1(n3619), .A2(n3618), .ZN(n5961) );
  BUF_X2 U4072 ( .A(n8282), .Z(n5950) );
  NAND2_X1 U4073 ( .A1(n3620), .A2(n8114), .ZN(n3622) );
  INV_X2 U4074 ( .A(n5345), .ZN(n8078) );
  NAND2_X1 U4075 ( .A1(n8078), .A2(\adder_stage1[11][15] ), .ZN(n3621) );
  NAND2_X1 U4076 ( .A1(n3622), .A2(n3621), .ZN(n9875) );
  NOR2_X1 U4077 ( .A1(\x_mult_f[18][1] ), .A2(\x_mult_f[19][1] ), .ZN(n7685)
         );
  NAND2_X1 U4078 ( .A1(\x_mult_f[18][0] ), .A2(\x_mult_f[19][0] ), .ZN(n7688)
         );
  NAND2_X1 U4079 ( .A1(\x_mult_f[18][1] ), .A2(\x_mult_f[19][1] ), .ZN(n7686)
         );
  OAI21_X1 U4080 ( .B1(n7685), .B2(n7688), .A(n7686), .ZN(n6947) );
  NOR2_X1 U4081 ( .A1(\x_mult_f[18][2] ), .A2(\x_mult_f[19][2] ), .ZN(n7692)
         );
  NOR2_X1 U4082 ( .A1(\x_mult_f[18][3] ), .A2(\x_mult_f[19][3] ), .ZN(n6948)
         );
  NOR2_X1 U4083 ( .A1(n7692), .A2(n6948), .ZN(n3624) );
  NAND2_X1 U4084 ( .A1(\x_mult_f[18][2] ), .A2(\x_mult_f[19][2] ), .ZN(n7693)
         );
  NAND2_X1 U4085 ( .A1(\x_mult_f[18][3] ), .A2(\x_mult_f[19][3] ), .ZN(n6949)
         );
  OAI21_X1 U4086 ( .B1(n6948), .B2(n7693), .A(n6949), .ZN(n3623) );
  AOI21_X1 U4087 ( .B1(n6947), .B2(n3624), .A(n3623), .ZN(n6600) );
  NOR2_X1 U4088 ( .A1(\x_mult_f[18][4] ), .A2(\x_mult_f[19][4] ), .ZN(n7069)
         );
  NOR2_X1 U4089 ( .A1(\x_mult_f[18][5] ), .A2(\x_mult_f[19][5] ), .ZN(n7071)
         );
  NOR2_X1 U4090 ( .A1(n7069), .A2(n7071), .ZN(n6602) );
  NOR2_X1 U4091 ( .A1(\x_mult_f[18][6] ), .A2(\x_mult_f[19][6] ), .ZN(n7060)
         );
  NOR2_X1 U4092 ( .A1(\x_mult_f[18][7] ), .A2(\x_mult_f[19][7] ), .ZN(n7062)
         );
  NOR2_X1 U4093 ( .A1(n7060), .A2(n7062), .ZN(n3626) );
  NAND2_X1 U4094 ( .A1(n6602), .A2(n3626), .ZN(n3628) );
  NAND2_X1 U4095 ( .A1(\x_mult_f[18][4] ), .A2(\x_mult_f[19][4] ), .ZN(n7679)
         );
  NAND2_X1 U4096 ( .A1(\x_mult_f[18][5] ), .A2(\x_mult_f[19][5] ), .ZN(n7072)
         );
  OAI21_X1 U4097 ( .B1(n7071), .B2(n7679), .A(n7072), .ZN(n6601) );
  NAND2_X1 U4098 ( .A1(\x_mult_f[18][6] ), .A2(\x_mult_f[19][6] ), .ZN(n7059)
         );
  NAND2_X1 U4099 ( .A1(\x_mult_f[18][7] ), .A2(\x_mult_f[19][7] ), .ZN(n7063)
         );
  OAI21_X1 U4100 ( .B1(n7062), .B2(n7059), .A(n7063), .ZN(n3625) );
  AOI21_X1 U4101 ( .B1(n3626), .B2(n6601), .A(n3625), .ZN(n3627) );
  OAI21_X1 U4102 ( .B1(n6600), .B2(n3628), .A(n3627), .ZN(n6619) );
  OR2_X1 U4103 ( .A1(\x_mult_f[18][8] ), .A2(\x_mult_f[19][8] ), .ZN(n6617) );
  NAND2_X1 U4104 ( .A1(\x_mult_f[18][8] ), .A2(\x_mult_f[19][8] ), .ZN(n6616)
         );
  INV_X1 U4105 ( .A(n6616), .ZN(n3629) );
  AOI21_X1 U4106 ( .B1(n6619), .B2(n6617), .A(n3629), .ZN(n6611) );
  NOR2_X1 U4107 ( .A1(\x_mult_f[18][9] ), .A2(\x_mult_f[19][9] ), .ZN(n6607)
         );
  NAND2_X1 U4108 ( .A1(\x_mult_f[18][9] ), .A2(\x_mult_f[19][9] ), .ZN(n6608)
         );
  OAI21_X1 U4109 ( .B1(n6611), .B2(n6607), .A(n6608), .ZN(n7108) );
  NOR2_X1 U4110 ( .A1(\x_mult_f[18][11] ), .A2(\x_mult_f[19][11] ), .ZN(n7079)
         );
  OR2_X1 U4111 ( .A1(\x_mult_f[18][10] ), .A2(\x_mult_f[19][10] ), .ZN(n7106)
         );
  OR2_X1 U4112 ( .A1(\x_mult_f[18][12] ), .A2(\x_mult_f[19][12] ), .ZN(n7091)
         );
  NAND2_X1 U4113 ( .A1(n7108), .A2(n3519), .ZN(n3636) );
  NAND2_X1 U4114 ( .A1(\x_mult_f[18][10] ), .A2(\x_mult_f[19][10] ), .ZN(n7105) );
  INV_X1 U4115 ( .A(n7105), .ZN(n7078) );
  NAND2_X1 U4116 ( .A1(\x_mult_f[18][11] ), .A2(\x_mult_f[19][11] ), .ZN(n7080) );
  NAND2_X1 U4117 ( .A1(\x_mult_f[18][12] ), .A2(\x_mult_f[19][12] ), .ZN(n7090) );
  NAND2_X1 U4118 ( .A1(\x_mult_f[18][13] ), .A2(\x_mult_f[19][13] ), .ZN(n6100) );
  NAND2_X1 U4119 ( .A1(n3636), .A2(n3635), .ZN(n6094) );
  NAND2_X1 U4120 ( .A1(n3637), .A2(n7698), .ZN(n3639) );
  NAND2_X1 U4121 ( .A1(n7910), .A2(\adder_stage1[9][15] ), .ZN(n3638) );
  NAND2_X1 U4122 ( .A1(n3639), .A2(n3638), .ZN(n9906) );
  NOR2_X1 U4123 ( .A1(\x_mult_f[26][1] ), .A2(\x_mult_f[27][1] ), .ZN(n5163)
         );
  NAND2_X1 U4124 ( .A1(\x_mult_f[26][0] ), .A2(\x_mult_f[27][0] ), .ZN(n5166)
         );
  NAND2_X1 U4125 ( .A1(\x_mult_f[26][1] ), .A2(\x_mult_f[27][1] ), .ZN(n5164)
         );
  OAI21_X1 U4126 ( .B1(n5163), .B2(n5166), .A(n5164), .ZN(n5029) );
  NOR2_X1 U4127 ( .A1(\x_mult_f[26][2] ), .A2(\x_mult_f[27][2] ), .ZN(n5121)
         );
  NOR2_X1 U4128 ( .A1(\x_mult_f[26][3] ), .A2(\x_mult_f[27][3] ), .ZN(n5030)
         );
  NOR2_X1 U4129 ( .A1(n5121), .A2(n5030), .ZN(n3641) );
  NAND2_X1 U4130 ( .A1(\x_mult_f[26][2] ), .A2(\x_mult_f[27][2] ), .ZN(n5122)
         );
  NAND2_X1 U4131 ( .A1(\x_mult_f[26][3] ), .A2(\x_mult_f[27][3] ), .ZN(n5031)
         );
  OAI21_X1 U4132 ( .B1(n5030), .B2(n5122), .A(n5031), .ZN(n3640) );
  AOI21_X1 U4133 ( .B1(n5029), .B2(n3641), .A(n3640), .ZN(n4527) );
  NOR2_X1 U4134 ( .A1(\x_mult_f[26][4] ), .A2(\x_mult_f[27][4] ), .ZN(n4528)
         );
  NOR2_X1 U4135 ( .A1(\x_mult_f[26][5] ), .A2(\x_mult_f[27][5] ), .ZN(n4530)
         );
  NOR2_X1 U4136 ( .A1(n4528), .A2(n4530), .ZN(n5024) );
  NOR2_X1 U4137 ( .A1(\x_mult_f[26][6] ), .A2(\x_mult_f[27][6] ), .ZN(n5056)
         );
  NOR2_X1 U4138 ( .A1(\x_mult_f[26][7] ), .A2(\x_mult_f[27][7] ), .ZN(n5058)
         );
  NOR2_X1 U4139 ( .A1(n5056), .A2(n5058), .ZN(n3643) );
  NAND2_X1 U4140 ( .A1(n5024), .A2(n3643), .ZN(n3645) );
  NAND2_X1 U4141 ( .A1(\x_mult_f[26][4] ), .A2(\x_mult_f[27][4] ), .ZN(n5037)
         );
  NAND2_X1 U4142 ( .A1(\x_mult_f[26][5] ), .A2(\x_mult_f[27][5] ), .ZN(n4531)
         );
  OAI21_X1 U4143 ( .B1(n4530), .B2(n5037), .A(n4531), .ZN(n5023) );
  NAND2_X1 U4144 ( .A1(\x_mult_f[26][6] ), .A2(\x_mult_f[27][6] ), .ZN(n5055)
         );
  NAND2_X1 U4145 ( .A1(\x_mult_f[26][7] ), .A2(\x_mult_f[27][7] ), .ZN(n5059)
         );
  OAI21_X1 U4146 ( .B1(n5058), .B2(n5055), .A(n5059), .ZN(n3642) );
  AOI21_X1 U4147 ( .B1(n3643), .B2(n5023), .A(n3642), .ZN(n3644) );
  OAI21_X1 U4148 ( .B1(n4527), .B2(n3645), .A(n3644), .ZN(n5052) );
  OR2_X1 U4149 ( .A1(\x_mult_f[26][8] ), .A2(\x_mult_f[27][8] ), .ZN(n5050) );
  NAND2_X1 U4150 ( .A1(\x_mult_f[26][8] ), .A2(\x_mult_f[27][8] ), .ZN(n5049)
         );
  INV_X1 U4151 ( .A(n5049), .ZN(n3646) );
  AOI21_X1 U4152 ( .B1(n5052), .B2(n5050), .A(n3646), .ZN(n4542) );
  NOR2_X1 U4153 ( .A1(\x_mult_f[26][9] ), .A2(\x_mult_f[27][9] ), .ZN(n4538)
         );
  NAND2_X1 U4154 ( .A1(\x_mult_f[26][9] ), .A2(\x_mult_f[27][9] ), .ZN(n4539)
         );
  OAI21_X1 U4155 ( .B1(n4542), .B2(n4538), .A(n4539), .ZN(n5046) );
  NOR2_X1 U4156 ( .A1(\x_mult_f[26][11] ), .A2(\x_mult_f[27][11] ), .ZN(n5017)
         );
  OR2_X1 U4157 ( .A1(\x_mult_f[26][10] ), .A2(\x_mult_f[27][10] ), .ZN(n5044)
         );
  OR2_X1 U4158 ( .A1(\x_mult_f[26][12] ), .A2(\x_mult_f[27][12] ), .ZN(n5011)
         );
  NAND2_X1 U4159 ( .A1(n5046), .A2(n3520), .ZN(n3653) );
  NAND2_X1 U4160 ( .A1(\x_mult_f[26][10] ), .A2(\x_mult_f[27][10] ), .ZN(n5043) );
  INV_X1 U4161 ( .A(n5043), .ZN(n5016) );
  NAND2_X1 U4162 ( .A1(\x_mult_f[26][11] ), .A2(\x_mult_f[27][11] ), .ZN(n5018) );
  NAND2_X1 U4163 ( .A1(\x_mult_f[26][12] ), .A2(\x_mult_f[27][12] ), .ZN(n5010) );
  NAND2_X1 U4164 ( .A1(\x_mult_f[26][13] ), .A2(\x_mult_f[27][13] ), .ZN(n3872) );
  NAND2_X1 U4165 ( .A1(n3653), .A2(n3652), .ZN(n5323) );
  NAND2_X1 U4166 ( .A1(n3654), .A2(n7511), .ZN(n3656) );
  INV_X2 U4167 ( .A(n5628), .ZN(n8048) );
  NAND2_X1 U4168 ( .A1(n8048), .A2(\adder_stage1[13][15] ), .ZN(n3655) );
  NAND2_X1 U4169 ( .A1(n3656), .A2(n3655), .ZN(n9841) );
  NOR2_X1 U4170 ( .A1(\adder_stage4[0][2] ), .A2(\adder_stage4[1][2] ), .ZN(
        n3797) );
  NOR2_X1 U4171 ( .A1(\adder_stage4[0][3] ), .A2(\adder_stage4[1][3] ), .ZN(
        n3792) );
  NOR2_X1 U4172 ( .A1(n3797), .A2(n3792), .ZN(n3660) );
  NOR2_X1 U4173 ( .A1(\adder_stage4[0][1] ), .A2(\adder_stage4[1][1] ), .ZN(
        n3802) );
  NAND2_X1 U4174 ( .A1(\adder_stage4[0][0] ), .A2(\adder_stage4[1][0] ), .ZN(
        n3805) );
  NAND2_X1 U4175 ( .A1(\adder_stage4[0][1] ), .A2(\adder_stage4[1][1] ), .ZN(
        n3803) );
  OAI21_X1 U4176 ( .B1(n3802), .B2(n3805), .A(n3803), .ZN(n3791) );
  NAND2_X1 U4177 ( .A1(\adder_stage4[0][2] ), .A2(\adder_stage4[1][2] ), .ZN(
        n3798) );
  NAND2_X1 U4178 ( .A1(\adder_stage4[0][3] ), .A2(\adder_stage4[1][3] ), .ZN(
        n3793) );
  OAI21_X1 U4179 ( .B1(n3792), .B2(n3798), .A(n3793), .ZN(n3659) );
  AOI21_X1 U4180 ( .B1(n3660), .B2(n3791), .A(n3659), .ZN(n3757) );
  NOR2_X1 U4181 ( .A1(\adder_stage4[0][4] ), .A2(\adder_stage4[1][4] ), .ZN(
        n3780) );
  NOR2_X1 U4182 ( .A1(\adder_stage4[0][5] ), .A2(\adder_stage4[1][5] ), .ZN(
        n3782) );
  NOR2_X1 U4183 ( .A1(n3780), .A2(n3782), .ZN(n3759) );
  NOR2_X1 U4184 ( .A1(\adder_stage4[0][6] ), .A2(\adder_stage4[1][6] ), .ZN(
        n3770) );
  NOR2_X1 U4185 ( .A1(\adder_stage4[0][7] ), .A2(\adder_stage4[1][7] ), .ZN(
        n3760) );
  NOR2_X1 U4186 ( .A1(n3770), .A2(n3760), .ZN(n3662) );
  NAND2_X1 U4187 ( .A1(n3759), .A2(n3662), .ZN(n3664) );
  NAND2_X1 U4188 ( .A1(\adder_stage4[0][4] ), .A2(\adder_stage4[1][4] ), .ZN(
        n3787) );
  NAND2_X1 U4189 ( .A1(\adder_stage4[0][5] ), .A2(\adder_stage4[1][5] ), .ZN(
        n3783) );
  OAI21_X1 U4190 ( .B1(n3782), .B2(n3787), .A(n3783), .ZN(n3758) );
  NAND2_X1 U4191 ( .A1(\adder_stage4[0][6] ), .A2(\adder_stage4[1][6] ), .ZN(
        n3771) );
  NAND2_X1 U4192 ( .A1(\adder_stage4[0][7] ), .A2(\adder_stage4[1][7] ), .ZN(
        n3761) );
  OAI21_X1 U4193 ( .B1(n3760), .B2(n3771), .A(n3761), .ZN(n3661) );
  AOI21_X1 U4194 ( .B1(n3662), .B2(n3758), .A(n3661), .ZN(n3663) );
  OAI21_X1 U4195 ( .B1(n3757), .B2(n3664), .A(n3663), .ZN(n3681) );
  NOR2_X1 U4196 ( .A1(\adder_stage4[0][8] ), .A2(\adder_stage4[1][8] ), .ZN(
        n3775) );
  NOR2_X1 U4197 ( .A1(\adder_stage4[1][9] ), .A2(\adder_stage4[0][9] ), .ZN(
        n3765) );
  NOR2_X1 U4198 ( .A1(n3775), .A2(n3765), .ZN(n3715) );
  NOR2_X1 U4199 ( .A1(\adder_stage4[0][10] ), .A2(\adder_stage4[1][10] ), .ZN(
        n3719) );
  NOR2_X1 U4200 ( .A1(\adder_stage4[0][11] ), .A2(\adder_stage4[1][11] ), .ZN(
        n3721) );
  NOR2_X1 U4201 ( .A1(n3719), .A2(n3721), .ZN(n3665) );
  NAND2_X1 U4202 ( .A1(n3715), .A2(n3665), .ZN(n3683) );
  NOR2_X1 U4203 ( .A1(\adder_stage4[0][12] ), .A2(\adder_stage4[1][12] ), .ZN(
        n3726) );
  NOR2_X1 U4204 ( .A1(\adder_stage4[0][13] ), .A2(\adder_stage4[1][13] ), .ZN(
        n3729) );
  NOR2_X1 U4205 ( .A1(n3726), .A2(n3729), .ZN(n3684) );
  NOR2_X1 U4206 ( .A1(\adder_stage4[0][14] ), .A2(\adder_stage4[1][14] ), .ZN(
        n3688) );
  NOR2_X1 U4207 ( .A1(\adder_stage4[0][15] ), .A2(\adder_stage4[1][15] ), .ZN(
        n3694) );
  NOR2_X1 U4208 ( .A1(n3688), .A2(n3694), .ZN(n3669) );
  NAND2_X1 U4209 ( .A1(n3684), .A2(n3669), .ZN(n3671) );
  NOR2_X1 U4210 ( .A1(n3683), .A2(n3671), .ZN(n3673) );
  NAND2_X1 U4211 ( .A1(\adder_stage4[1][8] ), .A2(\adder_stage4[0][8] ), .ZN(
        n3776) );
  NAND2_X1 U4212 ( .A1(\adder_stage4[0][9] ), .A2(\adder_stage4[1][9] ), .ZN(
        n3766) );
  OAI21_X1 U4213 ( .B1(n3765), .B2(n3776), .A(n3766), .ZN(n3716) );
  AND2_X1 U4214 ( .A1(n3665), .A2(n3716), .ZN(n3667) );
  NAND2_X1 U4215 ( .A1(\adder_stage4[0][10] ), .A2(\adder_stage4[1][10] ), 
        .ZN(n3753) );
  NAND2_X1 U4216 ( .A1(\adder_stage4[0][11] ), .A2(\adder_stage4[1][11] ), 
        .ZN(n3722) );
  OAI21_X1 U4217 ( .B1(n3721), .B2(n3753), .A(n3722), .ZN(n3666) );
  NOR2_X1 U4218 ( .A1(n3667), .A2(n3666), .ZN(n3682) );
  NAND2_X1 U4219 ( .A1(\adder_stage4[0][12] ), .A2(\adder_stage4[1][12] ), 
        .ZN(n3734) );
  NAND2_X1 U4220 ( .A1(\adder_stage4[0][13] ), .A2(\adder_stage4[1][13] ), 
        .ZN(n3730) );
  OAI21_X1 U4221 ( .B1(n3729), .B2(n3734), .A(n3730), .ZN(n3685) );
  NAND2_X1 U4222 ( .A1(\adder_stage4[0][14] ), .A2(\adder_stage4[1][14] ), 
        .ZN(n3690) );
  NAND2_X1 U4223 ( .A1(\adder_stage4[0][15] ), .A2(\adder_stage4[1][15] ), 
        .ZN(n3695) );
  OAI21_X1 U4224 ( .B1(n3694), .B2(n3690), .A(n3695), .ZN(n3668) );
  AOI21_X1 U4225 ( .B1(n3669), .B2(n3685), .A(n3668), .ZN(n3670) );
  OAI21_X1 U4226 ( .B1(n3682), .B2(n3671), .A(n3670), .ZN(n3672) );
  AOI21_X1 U4227 ( .B1(n3681), .B2(n3673), .A(n3672), .ZN(n3747) );
  NOR2_X1 U4228 ( .A1(\adder_stage4[0][16] ), .A2(\adder_stage4[1][16] ), .ZN(
        n3700) );
  INV_X1 U4229 ( .A(n3700), .ZN(n3675) );
  NAND2_X1 U4230 ( .A1(\adder_stage4[0][16] ), .A2(\adder_stage4[1][16] ), 
        .ZN(n3699) );
  NAND2_X1 U4231 ( .A1(n3675), .A2(n3699), .ZN(n3674) );
  XOR2_X1 U4232 ( .A(n3747), .B(n3674), .Z(m_data_out_y[16]) );
  OR2_X1 U4233 ( .A1(\adder_stage4[0][17] ), .A2(\adder_stage4[1][17] ), .ZN(
        n3702) );
  NAND2_X1 U4234 ( .A1(n3702), .A2(n3675), .ZN(n3705) );
  INV_X1 U4235 ( .A(n3699), .ZN(n3677) );
  NAND2_X1 U4236 ( .A1(\adder_stage4[0][17] ), .A2(\adder_stage4[1][17] ), 
        .ZN(n3701) );
  INV_X1 U4237 ( .A(n3701), .ZN(n3676) );
  AOI21_X1 U4238 ( .B1(n3702), .B2(n3677), .A(n3676), .ZN(n3710) );
  OAI21_X1 U4239 ( .B1(n3747), .B2(n3705), .A(n3710), .ZN(n3678) );
  INV_X1 U4240 ( .A(n3678), .ZN(n3680) );
  NOR2_X1 U4241 ( .A1(\adder_stage4[0][18] ), .A2(\adder_stage4[1][18] ), .ZN(
        n3709) );
  INV_X1 U4242 ( .A(n3709), .ZN(n3706) );
  NAND2_X1 U4243 ( .A1(\adder_stage4[0][18] ), .A2(\adder_stage4[1][18] ), 
        .ZN(n3708) );
  NAND2_X1 U4244 ( .A1(n3706), .A2(n3708), .ZN(n3679) );
  XOR2_X1 U4245 ( .A(n3680), .B(n3679), .Z(m_data_out_y[18]) );
  INV_X1 U4246 ( .A(n3681), .ZN(n3779) );
  OAI21_X1 U4247 ( .B1(n3779), .B2(n3683), .A(n3682), .ZN(n3728) );
  INV_X1 U4248 ( .A(n3728), .ZN(n3737) );
  INV_X1 U4249 ( .A(n3684), .ZN(n3687) );
  INV_X1 U4250 ( .A(n3685), .ZN(n3686) );
  OAI21_X1 U4251 ( .B1(n3737), .B2(n3687), .A(n3686), .ZN(n3693) );
  INV_X1 U4252 ( .A(n3688), .ZN(n3692) );
  NAND2_X1 U4253 ( .A1(n3692), .A2(n3690), .ZN(n3689) );
  XNOR2_X1 U4254 ( .A(n3693), .B(n3689), .ZN(m_data_out_y[14]) );
  INV_X1 U4255 ( .A(n3690), .ZN(n3691) );
  AOI21_X1 U4256 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3698) );
  INV_X1 U4257 ( .A(n3694), .ZN(n3696) );
  NAND2_X1 U4258 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  XOR2_X1 U4259 ( .A(n3698), .B(n3697), .Z(m_data_out_y[15]) );
  OAI21_X1 U4260 ( .B1(n3747), .B2(n3700), .A(n3699), .ZN(n3704) );
  NAND2_X1 U4261 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  XNOR2_X1 U4262 ( .A(n3704), .B(n3703), .ZN(m_data_out_y[17]) );
  INV_X1 U4263 ( .A(n3705), .ZN(n3707) );
  NAND2_X1 U4264 ( .A1(n3707), .A2(n3706), .ZN(n3738) );
  OAI21_X1 U4265 ( .B1(n3710), .B2(n3709), .A(n3708), .ZN(n3711) );
  INV_X1 U4266 ( .A(n3711), .ZN(n3743) );
  OAI21_X1 U4267 ( .B1(n3747), .B2(n3738), .A(n3743), .ZN(n3713) );
  OR2_X1 U4268 ( .A1(\adder_stage4[0][19] ), .A2(\adder_stage4[1][19] ), .ZN(
        n3740) );
  NAND2_X1 U4269 ( .A1(\adder_stage4[0][19] ), .A2(\adder_stage4[1][19] ), 
        .ZN(n3741) );
  NAND2_X1 U4270 ( .A1(n3740), .A2(n3741), .ZN(n3712) );
  XNOR2_X1 U4271 ( .A(n3713), .B(n3712), .ZN(m_data_out_y[19]) );
  OR2_X1 U4272 ( .A1(\adder_stage4[0][0] ), .A2(\adder_stage4[1][0] ), .ZN(
        n3714) );
  AND2_X1 U4273 ( .A1(n3714), .A2(n3805), .ZN(m_data_out_y[0]) );
  INV_X1 U4274 ( .A(n3715), .ZN(n3718) );
  INV_X1 U4275 ( .A(n3716), .ZN(n3717) );
  OAI21_X1 U4276 ( .B1(n3779), .B2(n3718), .A(n3717), .ZN(n3756) );
  INV_X1 U4277 ( .A(n3719), .ZN(n3754) );
  INV_X1 U4278 ( .A(n3753), .ZN(n3720) );
  AOI21_X1 U4279 ( .B1(n3756), .B2(n3754), .A(n3720), .ZN(n3725) );
  INV_X1 U4280 ( .A(n3721), .ZN(n3723) );
  NAND2_X1 U4281 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  XOR2_X1 U4282 ( .A(n3725), .B(n3724), .Z(m_data_out_y[11]) );
  INV_X1 U4283 ( .A(n3726), .ZN(n3735) );
  INV_X1 U4284 ( .A(n3734), .ZN(n3727) );
  AOI21_X1 U4285 ( .B1(n3728), .B2(n3735), .A(n3727), .ZN(n3733) );
  INV_X1 U4286 ( .A(n3729), .ZN(n3731) );
  NAND2_X1 U4287 ( .A1(n3731), .A2(n3730), .ZN(n3732) );
  XOR2_X1 U4288 ( .A(n3733), .B(n3732), .Z(m_data_out_y[13]) );
  NAND2_X1 U4289 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  XOR2_X1 U4290 ( .A(n3737), .B(n3736), .Z(m_data_out_y[12]) );
  INV_X1 U4291 ( .A(n3738), .ZN(n3739) );
  NAND2_X1 U4292 ( .A1(n3739), .A2(n3740), .ZN(n3746) );
  INV_X1 U4293 ( .A(n3740), .ZN(n3742) );
  OAI21_X1 U4294 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(n3744) );
  INV_X1 U4295 ( .A(n3744), .ZN(n3745) );
  OAI21_X1 U4296 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(n3748) );
  INV_X1 U4297 ( .A(n3748), .ZN(n3752) );
  OR2_X1 U4298 ( .A1(\adder_stage4[0][20] ), .A2(\adder_stage4[1][20] ), .ZN(
        n3750) );
  NAND2_X1 U4299 ( .A1(\adder_stage4[0][20] ), .A2(\adder_stage4[1][20] ), 
        .ZN(n3749) );
  NAND2_X1 U4300 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  XOR2_X1 U4301 ( .A(n3752), .B(n3751), .Z(m_data_out_y[20]) );
  NAND2_X1 U4302 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  XNOR2_X1 U4303 ( .A(n3756), .B(n3755), .ZN(m_data_out_y[10]) );
  INV_X1 U4304 ( .A(n3757), .ZN(n3790) );
  AOI21_X1 U4305 ( .B1(n3790), .B2(n3759), .A(n3758), .ZN(n3774) );
  OAI21_X1 U4306 ( .B1(n3774), .B2(n3770), .A(n3771), .ZN(n3764) );
  INV_X1 U4307 ( .A(n3760), .ZN(n3762) );
  NAND2_X1 U4308 ( .A1(n3762), .A2(n3761), .ZN(n3763) );
  XNOR2_X1 U4309 ( .A(n3764), .B(n3763), .ZN(m_data_out_y[7]) );
  OAI21_X1 U4310 ( .B1(n3779), .B2(n3775), .A(n3776), .ZN(n3769) );
  INV_X1 U4311 ( .A(n3765), .ZN(n3767) );
  NAND2_X1 U4312 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  XNOR2_X1 U4313 ( .A(n3769), .B(n3768), .ZN(m_data_out_y[9]) );
  INV_X1 U4314 ( .A(n3770), .ZN(n3772) );
  NAND2_X1 U4315 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  XOR2_X1 U4316 ( .A(n3774), .B(n3773), .Z(m_data_out_y[6]) );
  INV_X1 U4317 ( .A(n3775), .ZN(n3777) );
  NAND2_X1 U4318 ( .A1(n3777), .A2(n3776), .ZN(n3778) );
  XOR2_X1 U4319 ( .A(n3779), .B(n3778), .Z(m_data_out_y[8]) );
  INV_X1 U4320 ( .A(n3780), .ZN(n3788) );
  INV_X1 U4321 ( .A(n3787), .ZN(n3781) );
  AOI21_X1 U4322 ( .B1(n3790), .B2(n3788), .A(n3781), .ZN(n3786) );
  INV_X1 U4323 ( .A(n3782), .ZN(n3784) );
  NAND2_X1 U4324 ( .A1(n3784), .A2(n3783), .ZN(n3785) );
  XOR2_X1 U4325 ( .A(n3786), .B(n3785), .Z(m_data_out_y[5]) );
  NAND2_X1 U4326 ( .A1(n3788), .A2(n3787), .ZN(n3789) );
  XNOR2_X1 U4327 ( .A(n3790), .B(n3789), .ZN(m_data_out_y[4]) );
  INV_X1 U4328 ( .A(n3791), .ZN(n3801) );
  OAI21_X1 U4329 ( .B1(n3801), .B2(n3797), .A(n3798), .ZN(n3796) );
  INV_X1 U4330 ( .A(n3792), .ZN(n3794) );
  NAND2_X1 U4331 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  XNOR2_X1 U4332 ( .A(n3796), .B(n3795), .ZN(m_data_out_y[3]) );
  INV_X1 U4333 ( .A(n3797), .ZN(n3799) );
  NAND2_X1 U4334 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  XOR2_X1 U4335 ( .A(n3801), .B(n3800), .Z(m_data_out_y[2]) );
  INV_X1 U4336 ( .A(n3802), .ZN(n3804) );
  NAND2_X1 U4337 ( .A1(n3804), .A2(n3803), .ZN(n3806) );
  XOR2_X1 U4338 ( .A(n3806), .B(n3805), .Z(m_data_out_y[1]) );
  BUF_X2 U4339 ( .A(n3807), .Z(n8915) );
  NOR2_X1 U4340 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  INV_X2 U4341 ( .A(n3813), .ZN(n3835) );
  NOR2_X1 U4342 ( .A1(\ctrl_inst/state [1]), .A2(\ctrl_inst/state [0]), .ZN(
        n6431) );
  NAND2_X1 U4343 ( .A1(n6431), .A2(n8696), .ZN(n8357) );
  NOR3_X1 U4344 ( .A1(\ctrl_inst/xmem_tracker [5]), .A2(
        \ctrl_inst/xmem_tracker [6]), .A3(n3849), .ZN(n3821) );
  INV_X1 U4345 ( .A(n3821), .ZN(n3814) );
  OR2_X1 U4346 ( .A1(n8357), .A2(n3814), .ZN(n3822) );
  AOI21_X1 U4347 ( .B1(n8350), .B2(n3822), .A(n8680), .ZN(n8332) );
  INV_X1 U4348 ( .A(n8332), .ZN(n3818) );
  INV_X1 U4349 ( .A(\ctrl_inst/xmem_tracker [1]), .ZN(n3817) );
  INV_X1 U4350 ( .A(n3815), .ZN(n8666) );
  OAI21_X1 U4351 ( .B1(\ctrl_inst/xmem_tracker [0]), .B2(
        \ctrl_inst/xmem_tracker [1]), .A(n8666), .ZN(n3816) );
  INV_X1 U4352 ( .A(n3835), .ZN(n3824) );
  OAI22_X1 U4353 ( .A1(n3818), .A2(n3817), .B1(n3816), .B2(n8667), .ZN(n10321)
         );
  NOR3_X1 U4354 ( .A1(n8714), .A2(\ctrl_inst/state [2]), .A3(
        \ctrl_inst/state [0]), .ZN(n3819) );
  AND2_X1 U4355 ( .A1(n3835), .A2(n3819), .ZN(n3827) );
  NOR2_X1 U4356 ( .A1(n3822), .A2(n3820), .ZN(n3829) );
  AOI21_X1 U4357 ( .B1(n3827), .B2(n3425), .A(n3829), .ZN(n5457) );
  NOR2_X1 U4358 ( .A1(n3821), .A2(n8357), .ZN(n3830) );
  NOR2_X1 U4359 ( .A1(reset), .A2(n3830), .ZN(n3839) );
  INV_X1 U4360 ( .A(n3822), .ZN(n3823) );
  NAND2_X1 U4361 ( .A1(n3824), .A2(n3823), .ZN(n8358) );
  NAND2_X1 U4362 ( .A1(n8715), .A2(\ctrl_inst/pline_cntr [3]), .ZN(n3825) );
  OR2_X1 U4363 ( .A1(\ctrl_inst/pline_cntr [0]), .A2(\ctrl_inst/pline_cntr [1]), .ZN(n3851) );
  NOR2_X1 U4364 ( .A1(n3825), .A2(n3851), .ZN(n3837) );
  OAI211_X1 U4365 ( .C1(n3837), .C2(\ctrl_inst/state [1]), .A(
        \ctrl_inst/state [0]), .B(n8696), .ZN(n3826) );
  OR2_X1 U4366 ( .A1(n3835), .A2(n3826), .ZN(n3856) );
  NAND4_X1 U4367 ( .A1(n5457), .A2(n3839), .A3(n8358), .A4(n3856), .ZN(n3833)
         );
  INV_X1 U4368 ( .A(n3827), .ZN(n3828) );
  NOR2_X1 U4369 ( .A1(n3828), .A2(n6360), .ZN(n5460) );
  OR3_X1 U4370 ( .A1(n3830), .A2(n3829), .A3(n5460), .ZN(n3831) );
  INV_X1 U4371 ( .A(reset), .ZN(n8359) );
  NAND3_X1 U4372 ( .A1(n3831), .A2(n8359), .A3(n3833), .ZN(n3832) );
  OAI21_X1 U4373 ( .B1(n3833), .B2(n8719), .A(n3832), .ZN(n3385) );
  OR3_X1 U4374 ( .A1(n3835), .A2(n3837), .A3(n3834), .ZN(n3838) );
  NAND3_X1 U4375 ( .A1(n8915), .A2(\ctrl_inst/state [2]), .A3(n6431), .ZN(
        n3840) );
  NAND2_X1 U4376 ( .A1(n3838), .A2(n3840), .ZN(n8693) );
  INV_X1 U4377 ( .A(n8693), .ZN(n3848) );
  NAND2_X1 U4378 ( .A1(n6431), .A2(\ctrl_inst/state [2]), .ZN(n3854) );
  NOR2_X1 U4379 ( .A1(n3854), .A2(reset), .ZN(n8342) );
  NAND2_X1 U4380 ( .A1(\ctrl_inst/state [0]), .A2(n8359), .ZN(n3836) );
  NOR2_X1 U4381 ( .A1(n3836), .A2(\ctrl_inst/state [2]), .ZN(n5461) );
  NAND3_X1 U4382 ( .A1(\ctrl_inst/pline_cntr [0]), .A2(
        \ctrl_inst/pline_cntr [1]), .A3(n5461), .ZN(n8338) );
  NOR2_X1 U4383 ( .A1(\ctrl_inst/pline_cntr [2]), .A2(n8338), .ZN(n8335) );
  AOI21_X1 U4384 ( .B1(n8342), .B2(n3837), .A(n8335), .ZN(n3847) );
  NAND3_X1 U4385 ( .A1(n3840), .A2(n3839), .A3(n3838), .ZN(n8344) );
  NAND2_X1 U4386 ( .A1(n5461), .A2(n8713), .ZN(n8343) );
  INV_X1 U4387 ( .A(n8343), .ZN(n3841) );
  AOI21_X1 U4388 ( .B1(\ctrl_inst/pline_cntr [0]), .B2(n8342), .A(n3841), .ZN(
        n3842) );
  AND2_X1 U4389 ( .A1(n8344), .A2(n3842), .ZN(n8695) );
  INV_X1 U4390 ( .A(n8342), .ZN(n8347) );
  NOR2_X1 U4391 ( .A1(n8347), .A2(n8744), .ZN(n3844) );
  AND2_X1 U4392 ( .A1(n5461), .A2(n8744), .ZN(n3843) );
  NOR2_X1 U4393 ( .A1(n3844), .A2(n3843), .ZN(n3845) );
  NAND2_X1 U4394 ( .A1(n8695), .A2(n3845), .ZN(n8337) );
  NAND2_X1 U4395 ( .A1(n8337), .A2(\ctrl_inst/pline_cntr [2]), .ZN(n3846) );
  OAI21_X1 U4396 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3119) );
  NOR2_X1 U4397 ( .A1(n8667), .A2(n3849), .ZN(n8668) );
  NAND2_X1 U4398 ( .A1(\ctrl_inst/xmem_tracker [5]), .A2(n8668), .ZN(n3850) );
  OAI21_X1 U4399 ( .B1(n8680), .B2(n8745), .A(n3850), .ZN(n3384) );
  INV_X1 U4400 ( .A(n3851), .ZN(n3853) );
  NOR2_X1 U4401 ( .A1(\ctrl_inst/pline_cntr [2]), .A2(
        \ctrl_inst/pline_cntr [3]), .ZN(n3852) );
  NAND2_X1 U4402 ( .A1(n3853), .A2(n3852), .ZN(n8349) );
  NOR2_X1 U4403 ( .A1(n8349), .A2(n3854), .ZN(n3855) );
  NAND2_X1 U4404 ( .A1(n8922), .A2(n3855), .ZN(n8360) );
  AND2_X1 U4405 ( .A1(n3856), .A2(n8359), .ZN(n3857) );
  NAND2_X1 U4406 ( .A1(n8360), .A2(n3857), .ZN(n5458) );
  AOI21_X1 U4407 ( .B1(n5460), .B2(n3425), .A(n5458), .ZN(n3859) );
  OAI22_X1 U4408 ( .A1(n3859), .A2(n5461), .B1(m_valid_y), .B2(n5458), .ZN(
        n3860) );
  INV_X1 U4409 ( .A(n3860), .ZN(n3389) );
  INV_X1 U4410 ( .A(n8668), .ZN(n3862) );
  NAND3_X1 U4411 ( .A1(n3862), .A2(n8688), .A3(\ctrl_inst/xmem_tracker [5]), 
        .ZN(n3861) );
  OAI21_X1 U4412 ( .B1(\ctrl_inst/xmem_tracker [5]), .B2(n3862), .A(n3861), 
        .ZN(n3378) );
  AOI22_X1 U4413 ( .A1(n8365), .A2(\x_mult_f_int[27][5] ), .B1(n8200), .B2(
        \x_mult_f[27][5] ), .ZN(n3863) );
  INV_X1 U4414 ( .A(n3863), .ZN(n9243) );
  INV_X2 U4415 ( .A(n6711), .ZN(n8383) );
  AOI22_X1 U4416 ( .A1(\x_mult_f_int[9][7] ), .A2(n8387), .B1(n8383), .B2(
        \x_mult_f[9][7] ), .ZN(n3864) );
  INV_X1 U4417 ( .A(n3864), .ZN(n9041) );
  AOI22_X1 U4418 ( .A1(n8203), .A2(\x_mult_f_int[9][5] ), .B1(n8383), .B2(
        \x_mult_f[9][5] ), .ZN(n3865) );
  INV_X1 U4419 ( .A(n3865), .ZN(n9042) );
  AOI22_X1 U4420 ( .A1(n8189), .A2(\x_mult_f_int[4][5] ), .B1(n8200), .B2(
        \x_mult_f[4][5] ), .ZN(n3866) );
  INV_X1 U4421 ( .A(n3866), .ZN(n8984) );
  BUF_X2 U4422 ( .A(n6645), .Z(n8114) );
  AOI22_X1 U4423 ( .A1(\x_mult_f_int[27][6] ), .A2(n8114), .B1(n8200), .B2(
        \x_mult_f[27][6] ), .ZN(n3867) );
  INV_X1 U4424 ( .A(n3867), .ZN(n9242) );
  AOI22_X1 U4425 ( .A1(\x_mult_f_int[27][7] ), .A2(n8114), .B1(n8200), .B2(
        \x_mult_f[27][7] ), .ZN(n3868) );
  INV_X1 U4426 ( .A(n3868), .ZN(n9241) );
  AOI22_X1 U4427 ( .A1(\x_mult_f_int[4][6] ), .A2(n8203), .B1(n8200), .B2(
        \x_mult_f[4][6] ), .ZN(n3869) );
  INV_X1 U4428 ( .A(n3869), .ZN(n8983) );
  BUF_X2 U4429 ( .A(n8282), .Z(n8365) );
  AOI22_X1 U4430 ( .A1(\x_mult_f_int[4][11] ), .A2(n8365), .B1(n8048), .B2(
        \x_mult_f[4][11] ), .ZN(n3870) );
  INV_X1 U4431 ( .A(n3870), .ZN(n8978) );
  NAND2_X1 U4432 ( .A1(n3504), .A2(n3872), .ZN(n3873) );
  XOR2_X1 U4433 ( .A(n3874), .B(n3873), .Z(n3875) );
  AOI22_X1 U4434 ( .A1(n3875), .A2(n8114), .B1(n8048), .B2(
        \adder_stage1[13][13] ), .ZN(n3876) );
  INV_X1 U4435 ( .A(n3876), .ZN(n9843) );
  AOI22_X1 U4436 ( .A1(\x_mult_f_int[4][10] ), .A2(n8203), .B1(n8048), .B2(
        \x_mult_f[4][10] ), .ZN(n3877) );
  INV_X1 U4437 ( .A(n3877), .ZN(n8979) );
  AOI22_X1 U4438 ( .A1(\x_mult_f_int[4][7] ), .A2(n8203), .B1(n8048), .B2(
        \x_mult_f[4][7] ), .ZN(n3878) );
  INV_X1 U4439 ( .A(n3878), .ZN(n8982) );
  AOI22_X1 U4440 ( .A1(\x_mult_f_int[4][8] ), .A2(n8203), .B1(n8048), .B2(
        \x_mult_f[4][8] ), .ZN(n3879) );
  INV_X1 U4441 ( .A(n3879), .ZN(n8981) );
  AOI22_X1 U4442 ( .A1(\x_mult_f_int[4][9] ), .A2(n8203), .B1(n8048), .B2(
        \x_mult_f[4][9] ), .ZN(n3880) );
  INV_X1 U4443 ( .A(n3880), .ZN(n8980) );
  AOI22_X1 U4444 ( .A1(\x_mult_f_int[9][10] ), .A2(n8213), .B1(n8383), .B2(
        \x_mult_f[9][10] ), .ZN(n8796) );
  AOI22_X1 U4445 ( .A1(\x_mult_f_int[9][11] ), .A2(n8365), .B1(n8383), .B2(
        \x_mult_f[9][11] ), .ZN(n8795) );
  AOI22_X1 U4446 ( .A1(\x_mult_f_int[9][9] ), .A2(n8387), .B1(n8383), .B2(
        \x_mult_f[9][9] ), .ZN(n8797) );
  AOI22_X1 U4447 ( .A1(\x_mult_f_int[9][8] ), .A2(n8401), .B1(n8383), .B2(
        \x_mult_f[9][8] ), .ZN(n8798) );
  INV_X2 U4448 ( .A(n5410), .ZN(n8386) );
  AOI22_X1 U4449 ( .A1(n8213), .A2(\x_mult_f_int[17][5] ), .B1(n8386), .B2(
        \x_mult_f[17][5] ), .ZN(n3881) );
  INV_X1 U4450 ( .A(n3881), .ZN(n9150) );
  INV_X2 U4451 ( .A(n4651), .ZN(n8088) );
  AOI22_X1 U4452 ( .A1(n4002), .A2(\x_mult_f_int[11][5] ), .B1(n8088), .B2(
        \x_mult_f[11][5] ), .ZN(n3882) );
  INV_X1 U4453 ( .A(n3882), .ZN(n9068) );
  OR2_X1 U4454 ( .A1(\x_mult_f[10][8] ), .A2(\x_mult_f[11][8] ), .ZN(n6592) );
  OR2_X1 U4455 ( .A1(\x_mult_f[10][9] ), .A2(\x_mult_f[11][9] ), .ZN(n6594) );
  AND2_X1 U4456 ( .A1(n6592), .A2(n6594), .ZN(n7119) );
  OR2_X1 U4457 ( .A1(\x_mult_f[10][10] ), .A2(\x_mult_f[11][10] ), .ZN(n7124)
         );
  AND2_X1 U4458 ( .A1(n7119), .A2(n7124), .ZN(n3892) );
  NOR2_X1 U4459 ( .A1(\x_mult_f[10][2] ), .A2(\x_mult_f[11][2] ), .ZN(n6300)
         );
  NOR2_X1 U4460 ( .A1(\x_mult_f[10][3] ), .A2(\x_mult_f[11][3] ), .ZN(n6261)
         );
  NOR2_X1 U4461 ( .A1(n6300), .A2(n6261), .ZN(n3884) );
  NOR2_X1 U4462 ( .A1(\x_mult_f[10][1] ), .A2(\x_mult_f[11][1] ), .ZN(n6311)
         );
  NAND2_X1 U4463 ( .A1(\x_mult_f[10][0] ), .A2(\x_mult_f[11][0] ), .ZN(n6323)
         );
  NAND2_X1 U4464 ( .A1(\x_mult_f[10][1] ), .A2(\x_mult_f[11][1] ), .ZN(n6312)
         );
  OAI21_X1 U4465 ( .B1(n6311), .B2(n6323), .A(n6312), .ZN(n6260) );
  NAND2_X1 U4466 ( .A1(\x_mult_f[11][2] ), .A2(\x_mult_f[10][2] ), .ZN(n6301)
         );
  NAND2_X1 U4467 ( .A1(\x_mult_f[10][3] ), .A2(\x_mult_f[11][3] ), .ZN(n6262)
         );
  OAI21_X1 U4468 ( .B1(n6261), .B2(n6301), .A(n6262), .ZN(n3883) );
  AOI21_X1 U4469 ( .B1(n3884), .B2(n6260), .A(n3883), .ZN(n6268) );
  NOR2_X1 U4470 ( .A1(\x_mult_f[10][4] ), .A2(\x_mult_f[11][4] ), .ZN(n6269)
         );
  NOR2_X1 U4471 ( .A1(\x_mult_f[10][5] ), .A2(\x_mult_f[11][5] ), .ZN(n6271)
         );
  NOR2_X1 U4472 ( .A1(n6269), .A2(n6271), .ZN(n6279) );
  NOR2_X1 U4473 ( .A1(\x_mult_f[10][6] ), .A2(\x_mult_f[11][6] ), .ZN(n6285)
         );
  NOR2_X1 U4474 ( .A1(\x_mult_f[10][7] ), .A2(\x_mult_f[11][7] ), .ZN(n6287)
         );
  NOR2_X1 U4475 ( .A1(n6285), .A2(n6287), .ZN(n3886) );
  NAND2_X1 U4476 ( .A1(n6279), .A2(n3886), .ZN(n3888) );
  NAND2_X1 U4477 ( .A1(\x_mult_f[10][4] ), .A2(\x_mult_f[11][4] ), .ZN(n6294)
         );
  NAND2_X1 U4478 ( .A1(\x_mult_f[10][5] ), .A2(\x_mult_f[11][5] ), .ZN(n6272)
         );
  OAI21_X1 U4479 ( .B1(n6271), .B2(n6294), .A(n6272), .ZN(n6278) );
  NAND2_X1 U4480 ( .A1(\x_mult_f[10][6] ), .A2(\x_mult_f[11][6] ), .ZN(n6284)
         );
  NAND2_X1 U4481 ( .A1(\x_mult_f[10][7] ), .A2(\x_mult_f[11][7] ), .ZN(n6288)
         );
  OAI21_X1 U4482 ( .B1(n6287), .B2(n6284), .A(n6288), .ZN(n3885) );
  AOI21_X1 U4483 ( .B1(n3886), .B2(n6278), .A(n3885), .ZN(n3887) );
  OAI21_X1 U4484 ( .B1(n6268), .B2(n3888), .A(n3887), .ZN(n6590) );
  NAND2_X1 U4485 ( .A1(\x_mult_f[10][8] ), .A2(\x_mult_f[11][8] ), .ZN(n6307)
         );
  INV_X1 U4486 ( .A(n6307), .ZN(n6591) );
  NAND2_X1 U4487 ( .A1(\x_mult_f[10][9] ), .A2(\x_mult_f[11][9] ), .ZN(n6593)
         );
  INV_X1 U4488 ( .A(n6593), .ZN(n3889) );
  AOI21_X1 U4489 ( .B1(n6591), .B2(n6594), .A(n3889), .ZN(n7121) );
  INV_X1 U4490 ( .A(n7124), .ZN(n3890) );
  NAND2_X1 U4491 ( .A1(\x_mult_f[10][10] ), .A2(\x_mult_f[11][10] ), .ZN(n7123) );
  OAI21_X1 U4492 ( .B1(n7121), .B2(n3890), .A(n7123), .ZN(n3891) );
  AOI21_X1 U4493 ( .B1(n3892), .B2(n6590), .A(n3891), .ZN(n7040) );
  NOR2_X1 U4494 ( .A1(\x_mult_f[10][11] ), .A2(\x_mult_f[11][11] ), .ZN(n7036)
         );
  NAND2_X1 U4495 ( .A1(\x_mult_f[10][11] ), .A2(\x_mult_f[11][11] ), .ZN(n7037) );
  OAI21_X1 U4496 ( .B1(n7040), .B2(n7036), .A(n7037), .ZN(n7052) );
  OR2_X1 U4497 ( .A1(\x_mult_f[10][12] ), .A2(\x_mult_f[11][12] ), .ZN(n7050)
         );
  NAND2_X1 U4498 ( .A1(\x_mult_f[10][12] ), .A2(\x_mult_f[11][12] ), .ZN(n7049) );
  INV_X1 U4499 ( .A(n7049), .ZN(n3893) );
  AOI21_X1 U4500 ( .B1(n7052), .B2(n7050), .A(n3893), .ZN(n4192) );
  NOR2_X1 U4501 ( .A1(\x_mult_f[10][13] ), .A2(\x_mult_f[11][13] ), .ZN(n4188)
         );
  NAND2_X1 U4502 ( .A1(\x_mult_f[10][13] ), .A2(\x_mult_f[11][13] ), .ZN(n4189) );
  OAI21_X1 U4503 ( .B1(n4192), .B2(n4188), .A(n4189), .ZN(n4159) );
  INV_X1 U4504 ( .A(n3894), .ZN(n3895) );
  AOI22_X1 U4505 ( .A1(n3895), .A2(n8186), .B1(n8088), .B2(
        \adder_stage1[5][20] ), .ZN(n3896) );
  INV_X1 U4506 ( .A(n3896), .ZN(n9973) );
  NOR2_X1 U4507 ( .A1(\x_mult_f[8][2] ), .A2(\x_mult_f[9][2] ), .ZN(n7437) );
  NOR2_X1 U4508 ( .A1(\x_mult_f[8][3] ), .A2(\x_mult_f[9][3] ), .ZN(n7430) );
  NOR2_X1 U4509 ( .A1(n7437), .A2(n7430), .ZN(n3898) );
  NOR2_X1 U4510 ( .A1(\x_mult_f[8][1] ), .A2(\x_mult_f[9][1] ), .ZN(n7387) );
  NAND2_X1 U4511 ( .A1(\x_mult_f[8][0] ), .A2(\x_mult_f[9][0] ), .ZN(n7390) );
  NAND2_X1 U4512 ( .A1(\x_mult_f[8][1] ), .A2(\x_mult_f[9][1] ), .ZN(n7388) );
  OAI21_X1 U4513 ( .B1(n7387), .B2(n7390), .A(n7388), .ZN(n7429) );
  NAND2_X1 U4514 ( .A1(\x_mult_f[8][2] ), .A2(\x_mult_f[9][2] ), .ZN(n7438) );
  NAND2_X1 U4515 ( .A1(\x_mult_f[8][3] ), .A2(\x_mult_f[9][3] ), .ZN(n7431) );
  OAI21_X1 U4516 ( .B1(n7430), .B2(n7438), .A(n7431), .ZN(n3897) );
  AOI21_X1 U4517 ( .B1(n3898), .B2(n7429), .A(n3897), .ZN(n6776) );
  NOR2_X1 U4518 ( .A1(\x_mult_f[8][4] ), .A2(\x_mult_f[9][4] ), .ZN(n7371) );
  NOR2_X1 U4519 ( .A1(\x_mult_f[8][5] ), .A2(\x_mult_f[9][5] ), .ZN(n7373) );
  NOR2_X1 U4520 ( .A1(n7371), .A2(n7373), .ZN(n6778) );
  NOR2_X1 U4521 ( .A1(\x_mult_f[8][6] ), .A2(\x_mult_f[9][6] ), .ZN(n7395) );
  NOR2_X1 U4522 ( .A1(\x_mult_f[8][7] ), .A2(\x_mult_f[9][7] ), .ZN(n7397) );
  NOR2_X1 U4523 ( .A1(n7395), .A2(n7397), .ZN(n3900) );
  NAND2_X1 U4524 ( .A1(n6778), .A2(n3900), .ZN(n3902) );
  NAND2_X1 U4525 ( .A1(\x_mult_f[8][4] ), .A2(\x_mult_f[9][4] ), .ZN(n7423) );
  NAND2_X1 U4526 ( .A1(\x_mult_f[8][5] ), .A2(\x_mult_f[9][5] ), .ZN(n7374) );
  OAI21_X1 U4527 ( .B1(n7373), .B2(n7423), .A(n7374), .ZN(n6777) );
  NAND2_X1 U4528 ( .A1(\x_mult_f[8][6] ), .A2(\x_mult_f[9][6] ), .ZN(n7394) );
  NAND2_X1 U4529 ( .A1(\x_mult_f[8][7] ), .A2(\x_mult_f[9][7] ), .ZN(n7398) );
  OAI21_X1 U4530 ( .B1(n7397), .B2(n7394), .A(n7398), .ZN(n3899) );
  AOI21_X1 U4531 ( .B1(n3900), .B2(n6777), .A(n3899), .ZN(n3901) );
  OAI21_X1 U4532 ( .B1(n6776), .B2(n3902), .A(n3901), .ZN(n7420) );
  OR2_X1 U4533 ( .A1(\x_mult_f[8][8] ), .A2(\x_mult_f[9][8] ), .ZN(n7418) );
  OR2_X1 U4534 ( .A1(\x_mult_f[8][9] ), .A2(\x_mult_f[9][9] ), .ZN(n7406) );
  AND2_X1 U4535 ( .A1(n7418), .A2(n7406), .ZN(n7445) );
  NOR2_X1 U4536 ( .A1(\x_mult_f[8][10] ), .A2(\x_mult_f[9][10] ), .ZN(n3904)
         );
  INV_X1 U4537 ( .A(n3904), .ZN(n7450) );
  NAND3_X1 U4538 ( .A1(n7420), .A2(n7445), .A3(n7450), .ZN(n3907) );
  NAND2_X1 U4539 ( .A1(\x_mult_f[8][8] ), .A2(\x_mult_f[9][8] ), .ZN(n7417) );
  INV_X1 U4540 ( .A(n7417), .ZN(n7404) );
  NAND2_X1 U4541 ( .A1(\x_mult_f[8][9] ), .A2(\x_mult_f[9][9] ), .ZN(n7405) );
  INV_X1 U4542 ( .A(n7405), .ZN(n3903) );
  AOI21_X1 U4543 ( .B1(n7404), .B2(n7406), .A(n3903), .ZN(n7447) );
  NAND2_X1 U4544 ( .A1(\x_mult_f[8][10] ), .A2(\x_mult_f[9][10] ), .ZN(n7449)
         );
  OAI21_X1 U4545 ( .B1(n7447), .B2(n3904), .A(n7449), .ZN(n3905) );
  INV_X1 U4546 ( .A(n3905), .ZN(n3906) );
  AND2_X1 U4547 ( .A1(n3907), .A2(n3906), .ZN(n7384) );
  NOR2_X1 U4548 ( .A1(\x_mult_f[8][11] ), .A2(\x_mult_f[9][11] ), .ZN(n7380)
         );
  NAND2_X1 U4549 ( .A1(\x_mult_f[8][11] ), .A2(\x_mult_f[9][11] ), .ZN(n7381)
         );
  OAI21_X1 U4550 ( .B1(n7384), .B2(n7380), .A(n7381), .ZN(n7414) );
  OR2_X1 U4551 ( .A1(\x_mult_f[8][12] ), .A2(\x_mult_f[9][12] ), .ZN(n7412) );
  NAND2_X1 U4552 ( .A1(\x_mult_f[8][12] ), .A2(\x_mult_f[9][12] ), .ZN(n7411)
         );
  INV_X1 U4553 ( .A(n7411), .ZN(n3908) );
  AOI21_X1 U4554 ( .B1(n7414), .B2(n7412), .A(n3908), .ZN(n3914) );
  NOR2_X1 U4555 ( .A1(\x_mult_f[8][13] ), .A2(\x_mult_f[9][13] ), .ZN(n3910)
         );
  NAND2_X1 U4556 ( .A1(\x_mult_f[8][13] ), .A2(\x_mult_f[9][13] ), .ZN(n3911)
         );
  OAI21_X1 U4557 ( .B1(n3436), .B2(n3910), .A(n3911), .ZN(n7947) );
  BUF_X2 U4558 ( .A(n8282), .Z(n8387) );
  AOI22_X1 U4559 ( .A1(n3909), .A2(n8387), .B1(n8386), .B2(
        \adder_stage1[4][14] ), .ZN(n8801) );
  INV_X1 U4560 ( .A(n3910), .ZN(n3912) );
  NAND2_X1 U4561 ( .A1(n3912), .A2(n3911), .ZN(n3913) );
  XOR2_X1 U4562 ( .A(n3914), .B(n3913), .Z(n3915) );
  AOI22_X1 U4563 ( .A1(n3915), .A2(n8387), .B1(n8386), .B2(
        \adder_stage1[4][13] ), .ZN(n8802) );
  BUF_X2 U4564 ( .A(n8282), .Z(n8265) );
  AOI22_X1 U4565 ( .A1(\x_mult_f_int[16][12] ), .A2(n8265), .B1(n8088), .B2(
        \x_mult_f[16][12] ), .ZN(n3916) );
  INV_X1 U4566 ( .A(n3916), .ZN(n9130) );
  AOI22_X1 U4567 ( .A1(\x_mult_f_int[10][10] ), .A2(n8216), .B1(n8154), .B2(
        \x_mult_f[10][10] ), .ZN(n3917) );
  INV_X1 U4568 ( .A(n3917), .ZN(n9051) );
  AOI22_X1 U4569 ( .A1(\x_mult_f_int[10][9] ), .A2(n8216), .B1(n8157), .B2(
        \x_mult_f[10][9] ), .ZN(n3918) );
  INV_X1 U4570 ( .A(n3918), .ZN(n9052) );
  AOI22_X1 U4571 ( .A1(\x_mult_f_int[16][13] ), .A2(n8265), .B1(n7944), .B2(
        \x_mult_f[16][13] ), .ZN(n3919) );
  INV_X1 U4572 ( .A(n3919), .ZN(n9129) );
  AOI22_X1 U4573 ( .A1(\x_mult_f_int[16][11] ), .A2(n8265), .B1(n8228), .B2(
        \x_mult_f[16][11] ), .ZN(n3920) );
  INV_X1 U4574 ( .A(n3920), .ZN(n9131) );
  AOI22_X1 U4575 ( .A1(\x_mult_f_int[10][11] ), .A2(n8216), .B1(n8397), .B2(
        \x_mult_f[10][11] ), .ZN(n3921) );
  INV_X1 U4576 ( .A(n3921), .ZN(n9050) );
  BUF_X2 U4577 ( .A(n3452), .Z(n5628) );
  NOR2_X1 U4578 ( .A1(\adder_stage3[2][8] ), .A2(\adder_stage3[3][8] ), .ZN(
        n4035) );
  NOR2_X1 U4579 ( .A1(\adder_stage3[2][9] ), .A2(\adder_stage3[3][9] ), .ZN(
        n3962) );
  NOR2_X1 U4580 ( .A1(n4035), .A2(n3962), .ZN(n3937) );
  NOR2_X1 U4581 ( .A1(\adder_stage3[2][10] ), .A2(\adder_stage3[3][10] ), .ZN(
        n3941) );
  NOR2_X1 U4582 ( .A1(\adder_stage3[2][11] ), .A2(\adder_stage3[3][11] ), .ZN(
        n3943) );
  NOR2_X1 U4583 ( .A1(n3941), .A2(n3943), .ZN(n3930) );
  NAND2_X1 U4584 ( .A1(n3937), .A2(n3930), .ZN(n4141) );
  NOR2_X1 U4585 ( .A1(\adder_stage3[2][12] ), .A2(\adder_stage3[3][12] ), .ZN(
        n4143) );
  NOR2_X1 U4586 ( .A1(n4141), .A2(n4143), .ZN(n3984) );
  AND2_X1 U4587 ( .A1(n3984), .A2(n3508), .ZN(n3928) );
  NOR2_X1 U4588 ( .A1(\adder_stage3[2][2] ), .A2(\adder_stage3[3][2] ), .ZN(
        n8321) );
  NOR2_X1 U4589 ( .A1(\adder_stage3[2][3] ), .A2(\adder_stage3[3][3] ), .ZN(
        n8323) );
  NOR2_X1 U4590 ( .A1(n8321), .A2(n8323), .ZN(n3923) );
  NOR2_X1 U4591 ( .A1(\adder_stage3[2][1] ), .A2(\adder_stage3[3][1] ), .ZN(
        n8312) );
  NAND2_X1 U4592 ( .A1(\adder_stage3[2][0] ), .A2(\adder_stage3[3][0] ), .ZN(
        n8315) );
  NAND2_X1 U4593 ( .A1(\adder_stage3[2][1] ), .A2(\adder_stage3[3][1] ), .ZN(
        n8313) );
  OAI21_X1 U4594 ( .B1(n8312), .B2(n8315), .A(n8313), .ZN(n4788) );
  NAND2_X1 U4595 ( .A1(\adder_stage3[2][2] ), .A2(\adder_stage3[3][2] ), .ZN(
        n8320) );
  NAND2_X1 U4596 ( .A1(\adder_stage3[2][3] ), .A2(\adder_stage3[3][3] ), .ZN(
        n8324) );
  OAI21_X1 U4597 ( .B1(n8323), .B2(n8320), .A(n8324), .ZN(n3922) );
  AOI21_X1 U4598 ( .B1(n3923), .B2(n4788), .A(n3922), .ZN(n3951) );
  NOR2_X1 U4599 ( .A1(\adder_stage3[2][4] ), .A2(\adder_stage3[3][4] ), .ZN(
        n3952) );
  NOR2_X1 U4600 ( .A1(\adder_stage3[2][5] ), .A2(\adder_stage3[3][5] ), .ZN(
        n3954) );
  NOR2_X1 U4601 ( .A1(n3952), .A2(n3954), .ZN(n4042) );
  NOR2_X1 U4602 ( .A1(\adder_stage3[2][6] ), .A2(\adder_stage3[3][6] ), .ZN(
        n4077) );
  NOR2_X1 U4603 ( .A1(\adder_stage3[2][7] ), .A2(\adder_stage3[3][7] ), .ZN(
        n4044) );
  NOR2_X1 U4604 ( .A1(n4077), .A2(n4044), .ZN(n3925) );
  NAND2_X1 U4605 ( .A1(n4042), .A2(n3925), .ZN(n3927) );
  NAND2_X1 U4606 ( .A1(\adder_stage3[2][4] ), .A2(\adder_stage3[3][4] ), .ZN(
        n3979) );
  NAND2_X1 U4607 ( .A1(\adder_stage3[2][5] ), .A2(\adder_stage3[3][5] ), .ZN(
        n3955) );
  OAI21_X1 U4608 ( .B1(n3954), .B2(n3979), .A(n3955), .ZN(n4041) );
  NAND2_X1 U4609 ( .A1(\adder_stage3[2][6] ), .A2(\adder_stage3[3][6] ), .ZN(
        n4078) );
  NAND2_X1 U4610 ( .A1(\adder_stage3[2][7] ), .A2(\adder_stage3[3][7] ), .ZN(
        n4045) );
  OAI21_X1 U4611 ( .B1(n4044), .B2(n4078), .A(n4045), .ZN(n3924) );
  AOI21_X1 U4612 ( .B1(n3925), .B2(n4041), .A(n3924), .ZN(n3926) );
  OAI21_X1 U4613 ( .B1(n3951), .B2(n3927), .A(n3926), .ZN(n3985) );
  NAND2_X1 U4614 ( .A1(n3928), .A2(n3985), .ZN(n3933) );
  NAND2_X1 U4615 ( .A1(\adder_stage3[2][8] ), .A2(\adder_stage3[3][8] ), .ZN(
        n4036) );
  NAND2_X1 U4616 ( .A1(\adder_stage3[2][9] ), .A2(\adder_stage3[3][9] ), .ZN(
        n3963) );
  OAI21_X1 U4617 ( .B1(n3962), .B2(n4036), .A(n3963), .ZN(n3938) );
  NAND2_X1 U4618 ( .A1(\adder_stage3[2][10] ), .A2(\adder_stage3[3][10] ), 
        .ZN(n4014) );
  NAND2_X1 U4619 ( .A1(\adder_stage3[2][11] ), .A2(\adder_stage3[3][11] ), 
        .ZN(n3944) );
  OAI21_X1 U4620 ( .B1(n3943), .B2(n4014), .A(n3944), .ZN(n3929) );
  AOI21_X1 U4621 ( .B1(n3930), .B2(n3938), .A(n3929), .ZN(n4140) );
  NAND2_X1 U4622 ( .A1(\adder_stage3[2][12] ), .A2(\adder_stage3[3][12] ), 
        .ZN(n4144) );
  OAI21_X1 U4623 ( .B1(n4140), .B2(n4143), .A(n4144), .ZN(n3986) );
  NAND2_X1 U4624 ( .A1(\adder_stage3[2][13] ), .A2(\adder_stage3[3][13] ), 
        .ZN(n3987) );
  INV_X1 U4625 ( .A(n3987), .ZN(n3931) );
  AOI21_X1 U4626 ( .B1(n3986), .B2(n3508), .A(n3931), .ZN(n3932) );
  NAND2_X1 U4627 ( .A1(n3933), .A2(n3932), .ZN(n3995) );
  OR2_X1 U4628 ( .A1(\adder_stage3[2][14] ), .A2(\adder_stage3[3][14] ), .ZN(
        n3994) );
  NAND2_X1 U4629 ( .A1(\adder_stage3[2][14] ), .A2(\adder_stage3[3][14] ), 
        .ZN(n3992) );
  NAND2_X1 U4630 ( .A1(n3994), .A2(n3992), .ZN(n3934) );
  XNOR2_X1 U4631 ( .A(n3995), .B(n3934), .ZN(n3935) );
  AOI22_X1 U4632 ( .A1(n8157), .A2(\adder_stage4[1][14] ), .B1(n7909), .B2(
        n3935), .ZN(n3936) );
  INV_X1 U4633 ( .A(n3936), .ZN(n9553) );
  INV_X1 U4634 ( .A(n3985), .ZN(n4142) );
  INV_X1 U4635 ( .A(n3937), .ZN(n3940) );
  INV_X1 U4636 ( .A(n3938), .ZN(n3939) );
  OAI21_X1 U4637 ( .B1(n4142), .B2(n3940), .A(n3939), .ZN(n4017) );
  INV_X1 U4638 ( .A(n3941), .ZN(n4015) );
  INV_X1 U4639 ( .A(n4014), .ZN(n3942) );
  AOI21_X1 U4640 ( .B1(n4017), .B2(n4015), .A(n3942), .ZN(n3947) );
  INV_X1 U4641 ( .A(n3943), .ZN(n3945) );
  NAND2_X1 U4642 ( .A1(n3945), .A2(n3944), .ZN(n3946) );
  XOR2_X1 U4643 ( .A(n3947), .B(n3946), .Z(n3948) );
  AOI22_X1 U4644 ( .A1(n5544), .A2(\adder_stage4[1][11] ), .B1(n8203), .B2(
        n3948), .ZN(n3949) );
  INV_X1 U4645 ( .A(n3949), .ZN(n9556) );
  INV_X1 U4646 ( .A(n3951), .ZN(n4043) );
  INV_X1 U4647 ( .A(n3952), .ZN(n3980) );
  INV_X1 U4648 ( .A(n3979), .ZN(n3953) );
  AOI21_X1 U4649 ( .B1(n4043), .B2(n3980), .A(n3953), .ZN(n3958) );
  INV_X1 U4650 ( .A(n3954), .ZN(n3956) );
  NAND2_X1 U4651 ( .A1(n3956), .A2(n3955), .ZN(n3957) );
  XOR2_X1 U4652 ( .A(n3958), .B(n3957), .Z(n3959) );
  AOI22_X1 U4653 ( .A1(n8383), .A2(\adder_stage4[1][5] ), .B1(n4002), .B2(
        n3959), .ZN(n3960) );
  INV_X1 U4654 ( .A(n3960), .ZN(n9562) );
  AOI22_X1 U4655 ( .A1(n7767), .A2(\x_mult_f[23][3] ), .B1(n8329), .B2(
        \x_mult_f_int[23][3] ), .ZN(n3961) );
  INV_X1 U4656 ( .A(n3961), .ZN(n9214) );
  OAI21_X1 U4657 ( .B1(n4142), .B2(n4035), .A(n4036), .ZN(n3966) );
  INV_X1 U4658 ( .A(n3962), .ZN(n3964) );
  NAND2_X1 U4659 ( .A1(n3964), .A2(n3963), .ZN(n3965) );
  XNOR2_X1 U4660 ( .A(n3966), .B(n3965), .ZN(n3967) );
  AOI22_X1 U4661 ( .A1(n6373), .A2(\adder_stage4[1][9] ), .B1(n4002), .B2(
        n3967), .ZN(n3968) );
  INV_X1 U4662 ( .A(n3968), .ZN(n9558) );
  INV_X1 U4663 ( .A(n3969), .ZN(n4461) );
  AOI21_X1 U4664 ( .B1(n4461), .B2(n3971), .A(n3970), .ZN(n4522) );
  OAI21_X1 U4665 ( .B1(n4522), .B2(n4518), .A(n4519), .ZN(n3976) );
  INV_X1 U4666 ( .A(n3972), .ZN(n3974) );
  NAND2_X1 U4667 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  XNOR2_X1 U4668 ( .A(n3976), .B(n3975), .ZN(n3977) );
  AOI22_X1 U4669 ( .A1(n6373), .A2(\adder_stage1[11][7] ), .B1(n6523), .B2(
        n3977), .ZN(n3978) );
  INV_X1 U4670 ( .A(n3978), .ZN(n9883) );
  NAND2_X1 U4671 ( .A1(n3980), .A2(n3979), .ZN(n3981) );
  XNOR2_X1 U4672 ( .A(n4043), .B(n3981), .ZN(n3982) );
  AOI22_X1 U4673 ( .A1(n8202), .A2(\adder_stage4[1][4] ), .B1(n8318), .B2(
        n3982), .ZN(n3983) );
  INV_X1 U4674 ( .A(n3983), .ZN(n9563) );
  NAND2_X1 U4675 ( .A1(n3508), .A2(n3987), .ZN(n3988) );
  XOR2_X1 U4676 ( .A(n3989), .B(n3988), .Z(n3990) );
  AOI22_X1 U4677 ( .A1(n7944), .A2(\adder_stage4[1][13] ), .B1(n7284), .B2(
        n3990), .ZN(n3991) );
  INV_X1 U4678 ( .A(n3991), .ZN(n9554) );
  INV_X1 U4679 ( .A(n3992), .ZN(n3993) );
  AOI21_X1 U4680 ( .B1(n3995), .B2(n3994), .A(n3993), .ZN(n4645) );
  NOR2_X1 U4681 ( .A1(\adder_stage3[2][15] ), .A2(\adder_stage3[3][15] ), .ZN(
        n4644) );
  INV_X1 U4682 ( .A(n4644), .ZN(n3996) );
  NAND2_X1 U4683 ( .A1(\adder_stage3[2][15] ), .A2(\adder_stage3[3][15] ), 
        .ZN(n4643) );
  NAND2_X1 U4684 ( .A1(n3996), .A2(n4643), .ZN(n3997) );
  XOR2_X1 U4685 ( .A(n4645), .B(n3997), .Z(n3998) );
  AOI22_X1 U4686 ( .A1(n8386), .A2(\adder_stage4[1][15] ), .B1(n8208), .B2(
        n3998), .ZN(n3999) );
  INV_X1 U4687 ( .A(n3999), .ZN(n9552) );
  AOI22_X1 U4688 ( .A1(n6330), .A2(\x_mult_f[23][0] ), .B1(n8329), .B2(
        \x_mult_f_int[23][0] ), .ZN(n4000) );
  INV_X1 U4689 ( .A(n4000), .ZN(n9339) );
  AOI22_X1 U4690 ( .A1(n7443), .A2(\x_mult_f[23][2] ), .B1(n8329), .B2(
        \x_mult_f_int[23][2] ), .ZN(n4001) );
  INV_X1 U4691 ( .A(n4001), .ZN(n9215) );
  NOR2_X1 U4692 ( .A1(\adder_stage2[6][2] ), .A2(\adder_stage2[7][2] ), .ZN(
        n4117) );
  NOR2_X1 U4693 ( .A1(n4117), .A2(n4098), .ZN(n4004) );
  NOR2_X1 U4694 ( .A1(\adder_stage2[6][1] ), .A2(\adder_stage2[7][1] ), .ZN(
        n4124) );
  NAND2_X1 U4695 ( .A1(\adder_stage2[6][0] ), .A2(\adder_stage2[7][0] ), .ZN(
        n4130) );
  NAND2_X1 U4696 ( .A1(\adder_stage2[6][1] ), .A2(\adder_stage2[7][1] ), .ZN(
        n4125) );
  OAI21_X1 U4697 ( .B1(n4124), .B2(n4130), .A(n4125), .ZN(n4097) );
  NAND2_X1 U4698 ( .A1(\adder_stage2[6][2] ), .A2(\adder_stage2[7][2] ), .ZN(
        n4118) );
  NAND2_X1 U4699 ( .A1(\adder_stage2[6][3] ), .A2(\adder_stage2[7][3] ), .ZN(
        n4099) );
  OAI21_X1 U4700 ( .B1(n4098), .B2(n4118), .A(n4099), .ZN(n4003) );
  AOI21_X1 U4701 ( .B1(n4004), .B2(n4097), .A(n4003), .ZN(n4024) );
  NOR2_X1 U4702 ( .A1(\adder_stage2[6][4] ), .A2(\adder_stage2[7][4] ), .ZN(
        n4059) );
  NOR2_X1 U4703 ( .A1(\adder_stage2[6][5] ), .A2(\adder_stage2[7][5] ), .ZN(
        n4061) );
  NOR2_X1 U4704 ( .A1(n4059), .A2(n4061), .ZN(n4026) );
  NOR2_X1 U4705 ( .A1(\adder_stage2[6][6] ), .A2(\adder_stage2[7][6] ), .ZN(
        n4051) );
  NOR2_X1 U4706 ( .A1(\adder_stage2[6][7] ), .A2(\adder_stage2[7][7] ), .ZN(
        n4027) );
  NOR2_X1 U4707 ( .A1(n4051), .A2(n4027), .ZN(n4006) );
  NAND2_X1 U4708 ( .A1(n4026), .A2(n4006), .ZN(n4008) );
  NAND2_X1 U4709 ( .A1(\adder_stage2[6][4] ), .A2(\adder_stage2[7][4] ), .ZN(
        n4091) );
  NAND2_X1 U4710 ( .A1(\adder_stage2[6][5] ), .A2(\adder_stage2[7][5] ), .ZN(
        n4062) );
  OAI21_X1 U4711 ( .B1(n4061), .B2(n4091), .A(n4062), .ZN(n4025) );
  NAND2_X1 U4712 ( .A1(\adder_stage2[6][6] ), .A2(\adder_stage2[7][6] ), .ZN(
        n4052) );
  NAND2_X1 U4713 ( .A1(\adder_stage2[6][7] ), .A2(\adder_stage2[7][7] ), .ZN(
        n4028) );
  OAI21_X1 U4714 ( .B1(n4027), .B2(n4052), .A(n4028), .ZN(n4005) );
  AOI21_X1 U4715 ( .B1(n4006), .B2(n4025), .A(n4005), .ZN(n4007) );
  OAI21_X1 U4716 ( .B1(n4024), .B2(n4008), .A(n4007), .ZN(n4223) );
  INV_X1 U4717 ( .A(n4223), .ZN(n4504) );
  NOR2_X1 U4718 ( .A1(\adder_stage2[6][8] ), .A2(\adder_stage2[7][8] ), .ZN(
        n4150) );
  NAND2_X1 U4719 ( .A1(\adder_stage2[6][8] ), .A2(\adder_stage2[7][8] ), .ZN(
        n4152) );
  OAI21_X1 U4720 ( .B1(n4504), .B2(n4150), .A(n4152), .ZN(n4011) );
  INV_X1 U4721 ( .A(n4153), .ZN(n4009) );
  NAND2_X1 U4722 ( .A1(\adder_stage2[6][9] ), .A2(\adder_stage2[7][9] ), .ZN(
        n4151) );
  NAND2_X1 U4723 ( .A1(n4009), .A2(n4151), .ZN(n4010) );
  XNOR2_X1 U4724 ( .A(n4011), .B(n4010), .ZN(n4012) );
  AOI22_X1 U4725 ( .A1(n8078), .A2(\adder_stage3[3][9] ), .B1(n8390), .B2(
        n4012), .ZN(n4013) );
  INV_X1 U4726 ( .A(n4013), .ZN(n9600) );
  NAND2_X1 U4727 ( .A1(n4015), .A2(n4014), .ZN(n4016) );
  XNOR2_X1 U4728 ( .A(n4017), .B(n4016), .ZN(n4018) );
  AOI22_X1 U4729 ( .A1(n8155), .A2(\adder_stage4[1][10] ), .B1(n8189), .B2(
        n4018), .ZN(n4019) );
  INV_X1 U4730 ( .A(n4019), .ZN(n9557) );
  INV_X1 U4731 ( .A(n4150), .ZN(n4020) );
  NAND2_X1 U4732 ( .A1(n4020), .A2(n4152), .ZN(n4021) );
  XOR2_X1 U4733 ( .A(n4504), .B(n4021), .Z(n4022) );
  AOI22_X1 U4734 ( .A1(n8212), .A2(\adder_stage3[3][8] ), .B1(n8329), .B2(
        n4022), .ZN(n4023) );
  INV_X1 U4735 ( .A(n4023), .ZN(n9601) );
  INV_X1 U4736 ( .A(n4024), .ZN(n4094) );
  AOI21_X1 U4737 ( .B1(n4094), .B2(n4026), .A(n4025), .ZN(n4055) );
  OAI21_X1 U4738 ( .B1(n4055), .B2(n4051), .A(n4052), .ZN(n4031) );
  INV_X1 U4739 ( .A(n4027), .ZN(n4029) );
  NAND2_X1 U4740 ( .A1(n4029), .A2(n4028), .ZN(n4030) );
  XNOR2_X1 U4741 ( .A(n4031), .B(n4030), .ZN(n4032) );
  AOI22_X1 U4742 ( .A1(n8218), .A2(\adder_stage3[3][7] ), .B1(n7110), .B2(
        n4032), .ZN(n4033) );
  INV_X1 U4743 ( .A(n4033), .ZN(n9602) );
  AOI22_X1 U4744 ( .A1(n6337), .A2(\x_mult_f[23][1] ), .B1(n8329), .B2(
        \x_mult_f_int[23][1] ), .ZN(n4034) );
  INV_X1 U4745 ( .A(n4034), .ZN(n9338) );
  INV_X1 U4746 ( .A(n4035), .ZN(n4037) );
  NAND2_X1 U4747 ( .A1(n4037), .A2(n4036), .ZN(n4038) );
  XOR2_X1 U4748 ( .A(n4142), .B(n4038), .Z(n4039) );
  AOI22_X1 U4749 ( .A1(n8059), .A2(\adder_stage4[1][8] ), .B1(n6915), .B2(
        n4039), .ZN(n4040) );
  INV_X1 U4750 ( .A(n4040), .ZN(n9559) );
  AOI21_X1 U4751 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4081) );
  OAI21_X1 U4752 ( .B1(n4081), .B2(n4077), .A(n4078), .ZN(n4048) );
  INV_X1 U4753 ( .A(n4044), .ZN(n4046) );
  NAND2_X1 U4754 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  XNOR2_X1 U4755 ( .A(n4048), .B(n4047), .ZN(n4049) );
  AOI22_X1 U4756 ( .A1(n7851), .A2(\adder_stage4[1][7] ), .B1(n8194), .B2(
        n4049), .ZN(n4050) );
  INV_X1 U4757 ( .A(n4050), .ZN(n9560) );
  INV_X1 U4758 ( .A(n4051), .ZN(n4053) );
  NAND2_X1 U4759 ( .A1(n4053), .A2(n4052), .ZN(n4054) );
  XOR2_X1 U4760 ( .A(n4055), .B(n4054), .Z(n4056) );
  AOI22_X1 U4761 ( .A1(n7793), .A2(\adder_stage3[3][6] ), .B1(n8318), .B2(
        n4056), .ZN(n4057) );
  INV_X1 U4762 ( .A(n4057), .ZN(n9603) );
  AOI22_X1 U4763 ( .A1(n8330), .A2(\x_mult_f[23][4] ), .B1(n8329), .B2(
        \x_mult_f_int[23][4] ), .ZN(n4058) );
  INV_X1 U4764 ( .A(n4058), .ZN(n9213) );
  INV_X1 U4765 ( .A(n4059), .ZN(n4092) );
  INV_X1 U4766 ( .A(n4091), .ZN(n4060) );
  AOI21_X1 U4767 ( .B1(n4094), .B2(n4092), .A(n4060), .ZN(n4065) );
  INV_X1 U4768 ( .A(n4061), .ZN(n4063) );
  NAND2_X1 U4769 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  XOR2_X1 U4770 ( .A(n4065), .B(n4064), .Z(n4066) );
  AOI22_X1 U4771 ( .A1(n7330), .A2(\adder_stage3[3][5] ), .B1(n8329), .B2(
        n4066), .ZN(n4067) );
  INV_X1 U4772 ( .A(n4067), .ZN(n9604) );
  NAND2_X1 U4773 ( .A1(n4072), .A2(n4071), .ZN(n4073) );
  XNOR2_X1 U4774 ( .A(n4074), .B(n4073), .ZN(n4075) );
  AOI22_X1 U4775 ( .A1(n8228), .A2(\adder_stage1[11][12] ), .B1(n8318), .B2(
        n4075), .ZN(n4076) );
  INV_X1 U4776 ( .A(n4076), .ZN(n9878) );
  INV_X1 U4777 ( .A(n4077), .ZN(n4079) );
  NAND2_X1 U4778 ( .A1(n4079), .A2(n4078), .ZN(n4080) );
  XOR2_X1 U4779 ( .A(n4081), .B(n4080), .Z(n4082) );
  AOI22_X1 U4780 ( .A1(n8048), .A2(\adder_stage4[1][6] ), .B1(n6221), .B2(
        n4082), .ZN(n4083) );
  INV_X1 U4781 ( .A(n4083), .ZN(n9561) );
  NAND2_X1 U4782 ( .A1(n3615), .A2(n4086), .ZN(n4087) );
  XOR2_X1 U4783 ( .A(n4088), .B(n4087), .Z(n4089) );
  AOI22_X1 U4784 ( .A1(n4689), .A2(\adder_stage1[11][11] ), .B1(n8318), .B2(
        n4089), .ZN(n4090) );
  INV_X1 U4785 ( .A(n4090), .ZN(n9879) );
  NAND2_X1 U4786 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  XNOR2_X1 U4787 ( .A(n4094), .B(n4093), .ZN(n4095) );
  AOI22_X1 U4788 ( .A1(n6330), .A2(\adder_stage3[3][4] ), .B1(n8318), .B2(
        n4095), .ZN(n4096) );
  INV_X1 U4789 ( .A(n4096), .ZN(n9605) );
  INV_X1 U4790 ( .A(n4097), .ZN(n4121) );
  OAI21_X1 U4791 ( .B1(n4121), .B2(n4117), .A(n4118), .ZN(n4102) );
  INV_X1 U4792 ( .A(n4098), .ZN(n4100) );
  NAND2_X1 U4793 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  XNOR2_X1 U4794 ( .A(n4102), .B(n4101), .ZN(n4103) );
  AOI22_X1 U4795 ( .A1(n8157), .A2(\adder_stage3[3][3] ), .B1(n7454), .B2(
        n4103), .ZN(n4104) );
  INV_X1 U4796 ( .A(n4104), .ZN(n9606) );
  NAND2_X1 U4797 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  XNOR2_X1 U4798 ( .A(n6085), .B(n4107), .ZN(n4108) );
  AOI22_X1 U4799 ( .A1(n8330), .A2(\adder_stage1[11][10] ), .B1(n8318), .B2(
        n4108), .ZN(n4109) );
  INV_X1 U4800 ( .A(n4109), .ZN(n9880) );
  INV_X1 U4801 ( .A(n4110), .ZN(n4112) );
  NAND2_X1 U4802 ( .A1(n4112), .A2(n4111), .ZN(n4113) );
  XOR2_X1 U4803 ( .A(n4114), .B(n4113), .Z(n4115) );
  AOI22_X1 U4804 ( .A1(n8202), .A2(\adder_stage1[11][9] ), .B1(n8318), .B2(
        n4115), .ZN(n4116) );
  INV_X1 U4805 ( .A(n4116), .ZN(n9881) );
  INV_X1 U4806 ( .A(n4117), .ZN(n4119) );
  NAND2_X1 U4807 ( .A1(n4119), .A2(n4118), .ZN(n4120) );
  XOR2_X1 U4808 ( .A(n4121), .B(n4120), .Z(n4122) );
  AOI22_X1 U4809 ( .A1(n8048), .A2(\adder_stage3[3][2] ), .B1(n8318), .B2(
        n4122), .ZN(n4123) );
  INV_X1 U4810 ( .A(n4123), .ZN(n9607) );
  INV_X1 U4811 ( .A(n4124), .ZN(n4126) );
  NAND2_X1 U4812 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  XOR2_X1 U4813 ( .A(n4127), .B(n4130), .Z(n4128) );
  AOI22_X1 U4814 ( .A1(n7443), .A2(\adder_stage3[3][1] ), .B1(n8329), .B2(
        n4128), .ZN(n4129) );
  INV_X1 U4815 ( .A(n4129), .ZN(n9608) );
  OR2_X1 U4816 ( .A1(\adder_stage2[6][0] ), .A2(\adder_stage2[7][0] ), .ZN(
        n4131) );
  AND2_X1 U4817 ( .A1(n4131), .A2(n4130), .ZN(n4132) );
  AOI22_X1 U4818 ( .A1(n8391), .A2(\adder_stage3[3][0] ), .B1(n8329), .B2(
        n4132), .ZN(n4133) );
  INV_X1 U4819 ( .A(n4133), .ZN(n9609) );
  NAND2_X1 U4820 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  XNOR2_X1 U4821 ( .A(n4137), .B(n4136), .ZN(n4138) );
  AOI22_X1 U4822 ( .A1(n7944), .A2(\adder_stage1[11][8] ), .B1(n8318), .B2(
        n4138), .ZN(n4139) );
  INV_X1 U4823 ( .A(n4139), .ZN(n9882) );
  OAI21_X1 U4824 ( .B1(n4142), .B2(n4141), .A(n4140), .ZN(n4147) );
  INV_X1 U4825 ( .A(n4143), .ZN(n4145) );
  NAND2_X1 U4826 ( .A1(n4145), .A2(n4144), .ZN(n4146) );
  XNOR2_X1 U4827 ( .A(n4147), .B(n4146), .ZN(n4148) );
  AOI22_X1 U4828 ( .A1(n5626), .A2(\adder_stage4[1][12] ), .B1(n8329), .B2(
        n4148), .ZN(n4149) );
  INV_X1 U4829 ( .A(n4149), .ZN(n9555) );
  NOR2_X1 U4830 ( .A1(n4150), .A2(n4153), .ZN(n4217) );
  INV_X1 U4831 ( .A(n4217), .ZN(n4155) );
  OAI21_X1 U4832 ( .B1(n4153), .B2(n4152), .A(n4151), .ZN(n4219) );
  INV_X1 U4833 ( .A(n4219), .ZN(n4154) );
  OAI21_X1 U4834 ( .B1(n4504), .B2(n4155), .A(n4154), .ZN(n8296) );
  NOR2_X1 U4835 ( .A1(\adder_stage2[6][10] ), .A2(\adder_stage2[7][10] ), .ZN(
        n4216) );
  INV_X1 U4836 ( .A(n4216), .ZN(n8295) );
  NAND2_X1 U4837 ( .A1(\adder_stage2[6][10] ), .A2(\adder_stage2[7][10] ), 
        .ZN(n8293) );
  NAND2_X1 U4838 ( .A1(n8295), .A2(n8293), .ZN(n4156) );
  XNOR2_X1 U4839 ( .A(n8296), .B(n4156), .ZN(n4157) );
  AOI22_X1 U4840 ( .A1(n5294), .A2(\adder_stage3[3][10] ), .B1(n8114), .B2(
        n4157), .ZN(n4158) );
  INV_X1 U4841 ( .A(n4158), .ZN(n9599) );
  FA_X1 U4842 ( .A(\x_mult_f[10][14] ), .B(\x_mult_f[11][14] ), .CI(n4159), 
        .CO(n7987), .S(n4160) );
  AOI22_X1 U4843 ( .A1(n4160), .A2(n8398), .B1(n8088), .B2(
        \adder_stage1[5][14] ), .ZN(n4161) );
  INV_X1 U4844 ( .A(n4161), .ZN(n9975) );
  NOR2_X1 U4845 ( .A1(\adder_stage1[4][2] ), .A2(\adder_stage1[5][2] ), .ZN(
        n7778) );
  NOR2_X1 U4846 ( .A1(\adder_stage1[4][3] ), .A2(\adder_stage1[5][3] ), .ZN(
        n7780) );
  NOR2_X1 U4847 ( .A1(n7778), .A2(n7780), .ZN(n4163) );
  NOR2_X1 U4848 ( .A1(\adder_stage1[4][1] ), .A2(\adder_stage1[5][1] ), .ZN(
        n7787) );
  NAND2_X1 U4849 ( .A1(\adder_stage1[5][0] ), .A2(\adder_stage1[4][0] ), .ZN(
        n7790) );
  NAND2_X1 U4850 ( .A1(\adder_stage1[4][1] ), .A2(\adder_stage1[5][1] ), .ZN(
        n7788) );
  OAI21_X1 U4851 ( .B1(n7787), .B2(n7790), .A(n7788), .ZN(n6926) );
  NAND2_X1 U4852 ( .A1(\adder_stage1[4][2] ), .A2(\adder_stage1[5][2] ), .ZN(
        n7777) );
  NAND2_X1 U4853 ( .A1(\adder_stage1[4][3] ), .A2(\adder_stage1[5][3] ), .ZN(
        n7781) );
  OAI21_X1 U4854 ( .B1(n7780), .B2(n7777), .A(n7781), .ZN(n4162) );
  AOI21_X1 U4855 ( .B1(n4163), .B2(n6926), .A(n4162), .ZN(n6931) );
  NOR2_X1 U4856 ( .A1(\adder_stage1[4][4] ), .A2(\adder_stage1[5][4] ), .ZN(
        n6932) );
  NOR2_X1 U4857 ( .A1(\adder_stage1[4][5] ), .A2(\adder_stage1[5][5] ), .ZN(
        n6997) );
  NOR2_X1 U4858 ( .A1(n6932), .A2(n6997), .ZN(n6937) );
  NOR2_X1 U4859 ( .A1(\adder_stage1[4][6] ), .A2(\adder_stage1[5][6] ), .ZN(
        n7803) );
  NOR2_X1 U4860 ( .A1(\adder_stage1[4][7] ), .A2(\adder_stage1[5][7] ), .ZN(
        n6938) );
  NOR2_X1 U4861 ( .A1(n7803), .A2(n6938), .ZN(n4165) );
  NAND2_X1 U4862 ( .A1(n6937), .A2(n4165), .ZN(n4167) );
  NAND2_X1 U4863 ( .A1(\adder_stage1[4][4] ), .A2(\adder_stage1[5][4] ), .ZN(
        n6993) );
  NAND2_X1 U4864 ( .A1(\adder_stage1[4][5] ), .A2(\adder_stage1[5][5] ), .ZN(
        n6998) );
  OAI21_X1 U4865 ( .B1(n6997), .B2(n6993), .A(n6998), .ZN(n6936) );
  NAND2_X1 U4866 ( .A1(\adder_stage1[4][6] ), .A2(\adder_stage1[5][6] ), .ZN(
        n7804) );
  NAND2_X1 U4867 ( .A1(\adder_stage1[4][7] ), .A2(\adder_stage1[5][7] ), .ZN(
        n6939) );
  OAI21_X1 U4868 ( .B1(n6938), .B2(n7804), .A(n6939), .ZN(n4164) );
  AOI21_X1 U4869 ( .B1(n4165), .B2(n6936), .A(n4164), .ZN(n4166) );
  OAI21_X1 U4870 ( .B1(n6931), .B2(n4167), .A(n4166), .ZN(n7795) );
  NOR2_X1 U4871 ( .A1(\adder_stage1[4][8] ), .A2(\adder_stage1[5][8] ), .ZN(
        n7796) );
  INV_X1 U4872 ( .A(n7796), .ZN(n7821) );
  OR2_X1 U4873 ( .A1(\adder_stage1[4][9] ), .A2(\adder_stage1[5][9] ), .ZN(
        n7798) );
  NAND2_X1 U4874 ( .A1(n7821), .A2(n7798), .ZN(n7811) );
  NOR2_X1 U4875 ( .A1(\adder_stage1[4][10] ), .A2(\adder_stage1[5][10] ), .ZN(
        n7812) );
  NOR2_X1 U4876 ( .A1(n7811), .A2(n7812), .ZN(n4171) );
  NAND2_X1 U4877 ( .A1(\adder_stage1[4][8] ), .A2(\adder_stage1[5][8] ), .ZN(
        n7820) );
  INV_X1 U4878 ( .A(n7820), .ZN(n4169) );
  NAND2_X1 U4879 ( .A1(\adder_stage1[4][9] ), .A2(\adder_stage1[5][9] ), .ZN(
        n7797) );
  INV_X1 U4880 ( .A(n7797), .ZN(n4168) );
  AOI21_X1 U4881 ( .B1(n7798), .B2(n4169), .A(n4168), .ZN(n7810) );
  NAND2_X1 U4882 ( .A1(\adder_stage1[4][10] ), .A2(\adder_stage1[5][10] ), 
        .ZN(n7813) );
  OAI21_X1 U4883 ( .B1(n7810), .B2(n7812), .A(n7813), .ZN(n4170) );
  AOI21_X1 U4884 ( .B1(n7795), .B2(n4171), .A(n4170), .ZN(n7843) );
  OR2_X1 U4885 ( .A1(\adder_stage1[4][12] ), .A2(\adder_stage1[5][12] ), .ZN(
        n7845) );
  NOR2_X1 U4886 ( .A1(\adder_stage1[4][11] ), .A2(\adder_stage1[5][11] ), .ZN(
        n7842) );
  INV_X1 U4887 ( .A(n7842), .ZN(n7827) );
  NAND2_X1 U4888 ( .A1(n7845), .A2(n7827), .ZN(n7831) );
  INV_X1 U4889 ( .A(n7831), .ZN(n4172) );
  NOR2_X1 U4890 ( .A1(\adder_stage1[4][13] ), .A2(\adder_stage1[5][13] ), .ZN(
        n4175) );
  INV_X1 U4891 ( .A(n4175), .ZN(n7836) );
  NAND2_X1 U4892 ( .A1(n4172), .A2(n7836), .ZN(n7145) );
  OR2_X1 U4893 ( .A1(\adder_stage1[4][14] ), .A2(\adder_stage1[5][14] ), .ZN(
        n7147) );
  INV_X1 U4894 ( .A(n7147), .ZN(n4177) );
  NOR3_X1 U4895 ( .A1(n7843), .A2(n7145), .A3(n4177), .ZN(n4179) );
  NAND2_X1 U4896 ( .A1(\adder_stage1[4][11] ), .A2(\adder_stage1[5][11] ), 
        .ZN(n7841) );
  INV_X1 U4897 ( .A(n7841), .ZN(n4174) );
  NAND2_X1 U4898 ( .A1(\adder_stage1[4][12] ), .A2(\adder_stage1[5][12] ), 
        .ZN(n7844) );
  INV_X1 U4899 ( .A(n7844), .ZN(n4173) );
  AOI21_X1 U4900 ( .B1(n7845), .B2(n4174), .A(n4173), .ZN(n7832) );
  NAND2_X1 U4901 ( .A1(\adder_stage1[4][13] ), .A2(\adder_stage1[5][13] ), 
        .ZN(n7835) );
  OAI21_X1 U4902 ( .B1(n7832), .B2(n4175), .A(n7835), .ZN(n4176) );
  INV_X1 U4903 ( .A(n4176), .ZN(n7144) );
  NAND2_X1 U4904 ( .A1(\adder_stage1[4][14] ), .A2(\adder_stage1[5][14] ), 
        .ZN(n7146) );
  OAI21_X1 U4905 ( .B1(n7144), .B2(n4177), .A(n7146), .ZN(n4178) );
  OR2_X1 U4906 ( .A1(n4179), .A2(n4178), .ZN(n7983) );
  AOI22_X1 U4907 ( .A1(n4180), .A2(n7356), .B1(n8088), .B2(
        \adder_stage2[2][15] ), .ZN(n4181) );
  INV_X1 U4908 ( .A(n4181), .ZN(n9756) );
  NAND2_X1 U4909 ( .A1(n3501), .A2(n4183), .ZN(n4184) );
  XOR2_X1 U4910 ( .A(n4185), .B(n4184), .Z(n4186) );
  AOI22_X1 U4911 ( .A1(n4186), .A2(n8208), .B1(n8088), .B2(
        \adder_stage1[7][13] ), .ZN(n4187) );
  INV_X1 U4912 ( .A(n4187), .ZN(n9942) );
  INV_X1 U4913 ( .A(n4188), .ZN(n4190) );
  NAND2_X1 U4914 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  XOR2_X1 U4915 ( .A(n4192), .B(n4191), .Z(n4193) );
  AOI22_X1 U4916 ( .A1(n4193), .A2(n6915), .B1(n8088), .B2(
        \adder_stage1[5][13] ), .ZN(n4194) );
  INV_X1 U4917 ( .A(n4194), .ZN(n9976) );
  AOI22_X1 U4918 ( .A1(\x_mult_f_int[11][6] ), .A2(n8186), .B1(n8088), .B2(
        \x_mult_f[11][6] ), .ZN(n4195) );
  INV_X1 U4919 ( .A(n4195), .ZN(n9067) );
  NOR2_X1 U4920 ( .A1(\adder_stage1[6][8] ), .A2(\adder_stage1[7][8] ), .ZN(
        n5902) );
  INV_X1 U4921 ( .A(n5902), .ZN(n5897) );
  NAND2_X1 U4922 ( .A1(n3512), .A2(n3474), .ZN(n5904) );
  NAND2_X1 U4923 ( .A1(n5897), .A2(n5904), .ZN(n6573) );
  NOR2_X1 U4924 ( .A1(\adder_stage1[6][10] ), .A2(\adder_stage1[7][10] ), .ZN(
        n6575) );
  NOR2_X1 U4925 ( .A1(n6573), .A2(n6575), .ZN(n6534) );
  NOR2_X1 U4926 ( .A1(\adder_stage1[6][2] ), .A2(\adder_stage1[7][2] ), .ZN(
        n5872) );
  NOR2_X1 U4927 ( .A1(\adder_stage1[6][3] ), .A2(\adder_stage1[7][3] ), .ZN(
        n5874) );
  NOR2_X1 U4928 ( .A1(n5872), .A2(n5874), .ZN(n4197) );
  NOR2_X1 U4929 ( .A1(\adder_stage1[6][1] ), .A2(\adder_stage1[7][1] ), .ZN(
        n5881) );
  NAND2_X1 U4930 ( .A1(\adder_stage1[6][0] ), .A2(\adder_stage1[7][0] ), .ZN(
        n5884) );
  NAND2_X1 U4931 ( .A1(\adder_stage1[6][1] ), .A2(\adder_stage1[7][1] ), .ZN(
        n5882) );
  OAI21_X1 U4932 ( .B1(n5881), .B2(n5884), .A(n5882), .ZN(n5863) );
  NAND2_X1 U4933 ( .A1(\adder_stage1[6][2] ), .A2(\adder_stage1[7][2] ), .ZN(
        n5871) );
  NAND2_X1 U4934 ( .A1(\adder_stage1[6][3] ), .A2(\adder_stage1[7][3] ), .ZN(
        n5875) );
  OAI21_X1 U4935 ( .B1(n5874), .B2(n5871), .A(n5875), .ZN(n4196) );
  AOI21_X1 U4936 ( .B1(n4197), .B2(n5863), .A(n4196), .ZN(n5831) );
  NOR2_X1 U4937 ( .A1(\adder_stage1[6][4] ), .A2(\adder_stage1[7][4] ), .ZN(
        n5832) );
  NOR2_X1 U4938 ( .A1(\adder_stage1[6][5] ), .A2(\adder_stage1[7][5] ), .ZN(
        n5856) );
  NOR2_X1 U4939 ( .A1(n5832), .A2(n5856), .ZN(n5837) );
  NOR2_X1 U4940 ( .A1(\adder_stage1[6][6] ), .A2(\adder_stage1[7][6] ), .ZN(
        n5843) );
  NOR2_X1 U4941 ( .A1(\adder_stage1[6][7] ), .A2(\adder_stage1[7][7] ), .ZN(
        n5845) );
  NOR2_X1 U4942 ( .A1(n5843), .A2(n5845), .ZN(n4199) );
  NAND2_X1 U4943 ( .A1(n5837), .A2(n4199), .ZN(n4201) );
  NAND2_X1 U4944 ( .A1(\adder_stage1[6][4] ), .A2(\adder_stage1[7][4] ), .ZN(
        n5852) );
  NAND2_X1 U4945 ( .A1(\adder_stage1[6][5] ), .A2(\adder_stage1[7][5] ), .ZN(
        n5857) );
  OAI21_X1 U4946 ( .B1(n5856), .B2(n5852), .A(n5857), .ZN(n5836) );
  NAND2_X1 U4947 ( .A1(\adder_stage1[6][6] ), .A2(\adder_stage1[7][6] ), .ZN(
        n5842) );
  NAND2_X1 U4948 ( .A1(\adder_stage1[6][7] ), .A2(\adder_stage1[7][7] ), .ZN(
        n5846) );
  OAI21_X1 U4949 ( .B1(n5845), .B2(n5842), .A(n5846), .ZN(n4198) );
  AOI21_X1 U4950 ( .B1(n4199), .B2(n5836), .A(n4198), .ZN(n4200) );
  OAI21_X1 U4951 ( .B1(n5831), .B2(n4201), .A(n4200), .ZN(n6533) );
  OR2_X1 U4952 ( .A1(\adder_stage1[6][11] ), .A2(\adder_stage1[7][11] ), .ZN(
        n6538) );
  NAND3_X1 U4953 ( .A1(n6534), .A2(n6533), .A3(n6538), .ZN(n6527) );
  OR2_X1 U4954 ( .A1(\adder_stage1[6][12] ), .A2(\adder_stage1[7][12] ), .ZN(
        n6564) );
  OR2_X1 U4955 ( .A1(\adder_stage1[6][13] ), .A2(\adder_stage1[7][13] ), .ZN(
        n6567) );
  NAND2_X1 U4956 ( .A1(n6564), .A2(n6567), .ZN(n4211) );
  NAND2_X1 U4957 ( .A1(\adder_stage1[6][11] ), .A2(\adder_stage1[7][11] ), 
        .ZN(n6537) );
  OR2_X1 U4958 ( .A1(n4211), .A2(n6537), .ZN(n4209) );
  NAND2_X1 U4959 ( .A1(\adder_stage1[7][8] ), .A2(\adder_stage1[6][8] ), .ZN(
        n5901) );
  INV_X1 U4960 ( .A(n5901), .ZN(n4203) );
  NAND2_X1 U4961 ( .A1(\adder_stage1[7][9] ), .A2(\adder_stage1[6][9] ), .ZN(
        n5903) );
  INV_X1 U4962 ( .A(n5903), .ZN(n4202) );
  AOI21_X1 U4963 ( .B1(n4203), .B2(n5904), .A(n4202), .ZN(n6572) );
  NAND2_X1 U4964 ( .A1(\adder_stage1[6][10] ), .A2(\adder_stage1[7][10] ), 
        .ZN(n6576) );
  OAI21_X1 U4965 ( .B1(n6572), .B2(n6575), .A(n6576), .ZN(n6532) );
  INV_X1 U4966 ( .A(n4211), .ZN(n4204) );
  AND2_X1 U4967 ( .A1(n4204), .A2(n6538), .ZN(n4207) );
  NAND2_X1 U4968 ( .A1(\adder_stage1[6][12] ), .A2(\adder_stage1[7][12] ), 
        .ZN(n6528) );
  INV_X1 U4969 ( .A(n6528), .ZN(n6563) );
  NAND2_X1 U4970 ( .A1(n6563), .A2(n6567), .ZN(n4205) );
  NAND2_X1 U4971 ( .A1(\adder_stage1[6][13] ), .A2(\adder_stage1[7][13] ), 
        .ZN(n6566) );
  NAND2_X1 U4972 ( .A1(n4205), .A2(n6566), .ZN(n4206) );
  AOI21_X1 U4973 ( .B1(n6532), .B2(n4207), .A(n4206), .ZN(n4208) );
  AND2_X1 U4974 ( .A1(n4209), .A2(n4208), .ZN(n4210) );
  OAI21_X1 U4975 ( .B1(n6527), .B2(n4211), .A(n4210), .ZN(n6546) );
  OR2_X1 U4976 ( .A1(\adder_stage1[6][14] ), .A2(\adder_stage1[7][14] ), .ZN(
        n6544) );
  NAND2_X1 U4977 ( .A1(\adder_stage1[6][14] ), .A2(\adder_stage1[7][14] ), 
        .ZN(n6543) );
  INV_X1 U4978 ( .A(n6543), .ZN(n4212) );
  AOI21_X1 U4979 ( .B1(n6546), .B2(n6544), .A(n4212), .ZN(n4213) );
  INV_X1 U4980 ( .A(n4213), .ZN(n8087) );
  AOI22_X1 U4981 ( .A1(n4214), .A2(n8387), .B1(n8088), .B2(
        \adder_stage2[3][15] ), .ZN(n4215) );
  INV_X1 U4982 ( .A(n4215), .ZN(n9739) );
  NOR2_X1 U4983 ( .A1(n4216), .A2(n8297), .ZN(n4220) );
  NAND2_X1 U4984 ( .A1(n4217), .A2(n4220), .ZN(n4503) );
  NOR2_X1 U4985 ( .A1(\adder_stage2[6][12] ), .A2(\adder_stage2[7][12] ), .ZN(
        n4505) );
  NOR2_X1 U4986 ( .A1(n4503), .A2(n4505), .ZN(n4222) );
  NAND2_X1 U4987 ( .A1(\adder_stage2[6][11] ), .A2(\adder_stage2[7][11] ), 
        .ZN(n8298) );
  OAI21_X1 U4988 ( .B1(n8297), .B2(n8293), .A(n8298), .ZN(n4218) );
  AOI21_X1 U4989 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n4502) );
  NAND2_X1 U4990 ( .A1(\adder_stage2[6][12] ), .A2(\adder_stage2[7][12] ), 
        .ZN(n4506) );
  OAI21_X1 U4991 ( .B1(n4502), .B2(n4505), .A(n4506), .ZN(n4221) );
  AOI21_X1 U4992 ( .B1(n4223), .B2(n4222), .A(n4221), .ZN(n4492) );
  NOR2_X1 U4993 ( .A1(\adder_stage2[6][13] ), .A2(\adder_stage2[7][13] ), .ZN(
        n4488) );
  NAND2_X1 U4994 ( .A1(\adder_stage2[6][13] ), .A2(\adder_stage2[7][13] ), 
        .ZN(n4489) );
  OAI21_X1 U4995 ( .B1(n4492), .B2(n4488), .A(n4489), .ZN(n4485) );
  OR2_X1 U4996 ( .A1(\adder_stage2[6][14] ), .A2(\adder_stage2[7][14] ), .ZN(
        n4483) );
  NAND2_X1 U4997 ( .A1(\adder_stage2[6][14] ), .A2(\adder_stage2[7][14] ), 
        .ZN(n4482) );
  INV_X1 U4998 ( .A(n4482), .ZN(n4224) );
  AOI21_X1 U4999 ( .B1(n4485), .B2(n4483), .A(n4224), .ZN(n4499) );
  NOR2_X1 U5000 ( .A1(\adder_stage2[6][15] ), .A2(\adder_stage2[7][15] ), .ZN(
        n4495) );
  NAND2_X1 U5001 ( .A1(\adder_stage2[6][15] ), .A2(\adder_stage2[7][15] ), 
        .ZN(n4496) );
  OAI21_X1 U5002 ( .B1(n4499), .B2(n4495), .A(n4496), .ZN(n8250) );
  OR2_X1 U5003 ( .A1(\adder_stage2[6][16] ), .A2(\adder_stage2[7][16] ), .ZN(
        n8248) );
  NAND2_X1 U5004 ( .A1(\adder_stage2[6][16] ), .A2(\adder_stage2[7][16] ), 
        .ZN(n8247) );
  INV_X1 U5005 ( .A(n8247), .ZN(n4225) );
  NOR2_X1 U5006 ( .A1(\adder_stage2[6][17] ), .A2(\adder_stage2[7][17] ), .ZN(
        n5442) );
  NAND2_X1 U5007 ( .A1(\adder_stage2[6][17] ), .A2(\adder_stage2[7][17] ), 
        .ZN(n5443) );
  OAI21_X1 U5008 ( .B1(n5446), .B2(n5442), .A(n5443), .ZN(n8161) );
  OR2_X1 U5009 ( .A1(\adder_stage2[6][18] ), .A2(\adder_stage2[7][18] ), .ZN(
        n8160) );
  NAND2_X1 U5010 ( .A1(\adder_stage2[6][18] ), .A2(\adder_stage2[7][18] ), 
        .ZN(n7921) );
  NAND2_X1 U5011 ( .A1(n8160), .A2(n7921), .ZN(n4226) );
  XNOR2_X1 U5012 ( .A(n3431), .B(n4226), .ZN(n4227) );
  AOI22_X1 U5013 ( .A1(n4227), .A2(n8401), .B1(n8200), .B2(
        \adder_stage3[3][18] ), .ZN(n4228) );
  INV_X1 U5014 ( .A(n4228), .ZN(n9591) );
  INV_X2 U5015 ( .A(n4715), .ZN(n4689) );
  NOR2_X1 U5016 ( .A1(\adder_stage1[14][2] ), .A2(\adder_stage1[15][2] ), .ZN(
        n4896) );
  NOR2_X1 U5017 ( .A1(\adder_stage1[14][3] ), .A2(\adder_stage1[15][3] ), .ZN(
        n4898) );
  NOR2_X1 U5018 ( .A1(n4896), .A2(n4898), .ZN(n4230) );
  NOR2_X1 U5019 ( .A1(\adder_stage1[14][1] ), .A2(\adder_stage1[15][1] ), .ZN(
        n6317) );
  NAND2_X1 U5020 ( .A1(\adder_stage1[14][0] ), .A2(\adder_stage1[15][0] ), 
        .ZN(n6327) );
  NAND2_X1 U5021 ( .A1(\adder_stage1[14][1] ), .A2(\adder_stage1[15][1] ), 
        .ZN(n6318) );
  OAI21_X1 U5022 ( .B1(n6317), .B2(n6327), .A(n6318), .ZN(n4368) );
  NAND2_X1 U5023 ( .A1(\adder_stage1[14][2] ), .A2(\adder_stage1[15][2] ), 
        .ZN(n4895) );
  NAND2_X1 U5024 ( .A1(\adder_stage1[14][3] ), .A2(\adder_stage1[15][3] ), 
        .ZN(n4899) );
  OAI21_X1 U5025 ( .B1(n4898), .B2(n4895), .A(n4899), .ZN(n4229) );
  AOI21_X1 U5026 ( .B1(n4230), .B2(n4368), .A(n4229), .ZN(n4352) );
  NOR2_X1 U5027 ( .A1(\adder_stage1[14][4] ), .A2(\adder_stage1[15][4] ), .ZN(
        n4353) );
  NOR2_X1 U5028 ( .A1(\adder_stage1[14][5] ), .A2(\adder_stage1[15][5] ), .ZN(
        n4355) );
  NOR2_X1 U5029 ( .A1(n4353), .A2(n4355), .ZN(n4363) );
  NOR2_X1 U5030 ( .A1(\adder_stage1[14][6] ), .A2(\adder_stage1[15][6] ), .ZN(
        n4374) );
  NOR2_X1 U5031 ( .A1(\adder_stage1[14][7] ), .A2(\adder_stage1[15][7] ), .ZN(
        n4376) );
  NOR2_X1 U5032 ( .A1(n4374), .A2(n4376), .ZN(n4232) );
  NAND2_X1 U5033 ( .A1(n4363), .A2(n4232), .ZN(n4234) );
  NAND2_X1 U5034 ( .A1(\adder_stage1[14][4] ), .A2(\adder_stage1[15][4] ), 
        .ZN(n4383) );
  NAND2_X1 U5035 ( .A1(\adder_stage1[14][5] ), .A2(\adder_stage1[15][5] ), 
        .ZN(n4356) );
  OAI21_X1 U5036 ( .B1(n4355), .B2(n4383), .A(n4356), .ZN(n4362) );
  NAND2_X1 U5037 ( .A1(\adder_stage1[14][6] ), .A2(\adder_stage1[15][6] ), 
        .ZN(n4373) );
  NAND2_X1 U5038 ( .A1(\adder_stage1[14][7] ), .A2(\adder_stage1[15][7] ), 
        .ZN(n4377) );
  OAI21_X1 U5039 ( .B1(n4376), .B2(n4373), .A(n4377), .ZN(n4231) );
  AOI21_X1 U5040 ( .B1(n4232), .B2(n4362), .A(n4231), .ZN(n4233) );
  OAI21_X1 U5041 ( .B1(n4352), .B2(n4234), .A(n4233), .ZN(n4262) );
  INV_X1 U5042 ( .A(n4262), .ZN(n4682) );
  NOR2_X1 U5043 ( .A1(\adder_stage1[14][8] ), .A2(\adder_stage1[15][8] ), .ZN(
        n4239) );
  NAND2_X1 U5044 ( .A1(\adder_stage1[14][8] ), .A2(\adder_stage1[15][8] ), 
        .ZN(n4255) );
  OAI21_X1 U5045 ( .B1(n4682), .B2(n4239), .A(n4255), .ZN(n4236) );
  OR2_X1 U5046 ( .A1(\adder_stage1[14][9] ), .A2(\adder_stage1[15][9] ), .ZN(
        n4259) );
  NAND2_X1 U5047 ( .A1(\adder_stage1[14][9] ), .A2(\adder_stage1[15][9] ), 
        .ZN(n4256) );
  NAND2_X1 U5048 ( .A1(n4259), .A2(n4256), .ZN(n4235) );
  XNOR2_X1 U5049 ( .A(n4236), .B(n4235), .ZN(n4237) );
  AOI22_X1 U5050 ( .A1(n4689), .A2(\adder_stage2[7][9] ), .B1(n4596), .B2(
        n4237), .ZN(n4238) );
  INV_X1 U5051 ( .A(n4238), .ZN(n9677) );
  INV_X1 U5052 ( .A(n4239), .ZN(n4254) );
  NAND2_X1 U5053 ( .A1(n4254), .A2(n4255), .ZN(n4240) );
  XOR2_X1 U5054 ( .A(n4682), .B(n4240), .Z(n4241) );
  AOI22_X1 U5055 ( .A1(n4689), .A2(\adder_stage2[7][8] ), .B1(n8365), .B2(
        n4241), .ZN(n4242) );
  INV_X1 U5056 ( .A(n4242), .ZN(n9678) );
  NOR2_X1 U5057 ( .A1(\x_mult_f[30][2] ), .A2(\x_mult_f[31][2] ), .ZN(n4293)
         );
  NOR2_X1 U5058 ( .A1(\x_mult_f[30][3] ), .A2(\x_mult_f[31][3] ), .ZN(n4268)
         );
  NOR2_X1 U5059 ( .A1(n4293), .A2(n4268), .ZN(n4244) );
  NOR2_X1 U5060 ( .A1(\x_mult_f[30][1] ), .A2(\x_mult_f[31][1] ), .ZN(n4248)
         );
  NAND2_X1 U5061 ( .A1(\x_mult_f[31][0] ), .A2(\x_mult_f[30][0] ), .ZN(n4282)
         );
  NAND2_X1 U5062 ( .A1(\x_mult_f[30][1] ), .A2(\x_mult_f[31][1] ), .ZN(n4249)
         );
  OAI21_X1 U5063 ( .B1(n4248), .B2(n4282), .A(n4249), .ZN(n4267) );
  NAND2_X1 U5064 ( .A1(\x_mult_f[30][2] ), .A2(\x_mult_f[31][2] ), .ZN(n4294)
         );
  NAND2_X1 U5065 ( .A1(\x_mult_f[30][3] ), .A2(\x_mult_f[31][3] ), .ZN(n4269)
         );
  OAI21_X1 U5066 ( .B1(n4268), .B2(n4294), .A(n4269), .ZN(n4243) );
  AOI21_X1 U5067 ( .B1(n4244), .B2(n4267), .A(n4243), .ZN(n4320) );
  INV_X1 U5068 ( .A(n4320), .ZN(n4304) );
  NOR2_X1 U5069 ( .A1(\x_mult_f[30][4] ), .A2(\x_mult_f[31][4] ), .ZN(n4300)
         );
  INV_X1 U5070 ( .A(n4300), .ZN(n4276) );
  NAND2_X1 U5071 ( .A1(\x_mult_f[30][4] ), .A2(\x_mult_f[31][4] ), .ZN(n4302)
         );
  NAND2_X1 U5072 ( .A1(n4276), .A2(n4302), .ZN(n4245) );
  XNOR2_X1 U5073 ( .A(n4304), .B(n4245), .ZN(n4246) );
  AOI22_X1 U5074 ( .A1(n4689), .A2(\adder_stage1[15][4] ), .B1(n8265), .B2(
        n4246), .ZN(n4247) );
  INV_X1 U5075 ( .A(n4247), .ZN(n9818) );
  INV_X1 U5076 ( .A(n4248), .ZN(n4250) );
  NAND2_X1 U5077 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  XOR2_X1 U5078 ( .A(n4251), .B(n4282), .Z(n4252) );
  AOI22_X1 U5079 ( .A1(n4689), .A2(\adder_stage1[15][1] ), .B1(n8387), .B2(
        n4252), .ZN(n4253) );
  INV_X1 U5080 ( .A(n4253), .ZN(n9821) );
  NAND2_X1 U5081 ( .A1(n4254), .A2(n4259), .ZN(n4681) );
  NOR2_X1 U5082 ( .A1(\adder_stage1[14][10] ), .A2(\adder_stage1[15][10] ), 
        .ZN(n4683) );
  NOR2_X1 U5083 ( .A1(n4681), .A2(n4683), .ZN(n4261) );
  INV_X1 U5084 ( .A(n4255), .ZN(n4258) );
  INV_X1 U5085 ( .A(n4256), .ZN(n4257) );
  AOI21_X1 U5086 ( .B1(n4259), .B2(n4258), .A(n4257), .ZN(n4680) );
  NAND2_X1 U5087 ( .A1(\adder_stage1[14][10] ), .A2(\adder_stage1[15][10] ), 
        .ZN(n4684) );
  OAI21_X1 U5088 ( .B1(n4680), .B2(n4683), .A(n4684), .ZN(n4260) );
  AOI21_X1 U5089 ( .B1(n4262), .B2(n4261), .A(n4260), .ZN(n4290) );
  NOR2_X1 U5090 ( .A1(\adder_stage1[14][11] ), .A2(\adder_stage1[15][11] ), 
        .ZN(n4286) );
  NAND2_X1 U5091 ( .A1(\adder_stage1[14][11] ), .A2(\adder_stage1[15][11] ), 
        .ZN(n4287) );
  OAI21_X1 U5092 ( .B1(n4290), .B2(n4286), .A(n4287), .ZN(n4670) );
  OR2_X1 U5093 ( .A1(\adder_stage1[14][12] ), .A2(\adder_stage1[15][12] ), 
        .ZN(n4668) );
  NAND2_X1 U5094 ( .A1(\adder_stage1[14][12] ), .A2(\adder_stage1[15][12] ), 
        .ZN(n4667) );
  INV_X1 U5095 ( .A(n4667), .ZN(n4263) );
  AOI21_X1 U5096 ( .B1(n4670), .B2(n4668), .A(n4263), .ZN(n4677) );
  NOR2_X1 U5097 ( .A1(\adder_stage1[14][13] ), .A2(\adder_stage1[15][13] ), 
        .ZN(n4673) );
  NAND2_X1 U5098 ( .A1(\adder_stage1[14][13] ), .A2(\adder_stage1[15][13] ), 
        .ZN(n4674) );
  OAI21_X1 U5099 ( .B1(n3437), .B2(n4673), .A(n4674), .ZN(n6227) );
  OR2_X1 U5100 ( .A1(\adder_stage1[14][14] ), .A2(\adder_stage1[15][14] ), 
        .ZN(n6226) );
  NAND2_X1 U5101 ( .A1(\adder_stage1[14][14] ), .A2(\adder_stage1[15][14] ), 
        .ZN(n6224) );
  NAND2_X1 U5102 ( .A1(n6226), .A2(n6224), .ZN(n4264) );
  XNOR2_X1 U5103 ( .A(n6227), .B(n4264), .ZN(n4265) );
  AOI22_X1 U5104 ( .A1(n4689), .A2(\adder_stage2[7][14] ), .B1(n8401), .B2(
        n4265), .ZN(n4266) );
  INV_X1 U5105 ( .A(n4266), .ZN(n9672) );
  INV_X1 U5106 ( .A(n4267), .ZN(n4297) );
  OAI21_X1 U5107 ( .B1(n4297), .B2(n4293), .A(n4294), .ZN(n4272) );
  INV_X1 U5108 ( .A(n4268), .ZN(n4270) );
  NAND2_X1 U5109 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  XNOR2_X1 U5110 ( .A(n4272), .B(n4271), .ZN(n4273) );
  AOI22_X1 U5111 ( .A1(n4689), .A2(\adder_stage1[15][3] ), .B1(n8365), .B2(
        n4273), .ZN(n4274) );
  INV_X1 U5112 ( .A(n4274), .ZN(n9819) );
  INV_X1 U5113 ( .A(n4302), .ZN(n4275) );
  AOI21_X1 U5114 ( .B1(n4304), .B2(n4276), .A(n4275), .ZN(n4279) );
  NOR2_X1 U5115 ( .A1(\x_mult_f[30][5] ), .A2(\x_mult_f[31][5] ), .ZN(n4303)
         );
  INV_X1 U5116 ( .A(n4303), .ZN(n4277) );
  NAND2_X1 U5117 ( .A1(\x_mult_f[30][5] ), .A2(\x_mult_f[31][5] ), .ZN(n4301)
         );
  NAND2_X1 U5118 ( .A1(n4277), .A2(n4301), .ZN(n4278) );
  XOR2_X1 U5119 ( .A(n4279), .B(n4278), .Z(n4280) );
  AOI22_X1 U5120 ( .A1(n8383), .A2(\adder_stage1[15][5] ), .B1(n8213), .B2(
        n4280), .ZN(n4281) );
  INV_X1 U5121 ( .A(n4281), .ZN(n9817) );
  OR2_X1 U5122 ( .A1(\x_mult_f[30][0] ), .A2(\x_mult_f[31][0] ), .ZN(n4283) );
  AND2_X1 U5123 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  AOI22_X1 U5124 ( .A1(n4689), .A2(\adder_stage1[15][0] ), .B1(n5921), .B2(
        n4284), .ZN(n4285) );
  INV_X1 U5125 ( .A(n4285), .ZN(n9822) );
  INV_X1 U5126 ( .A(n4286), .ZN(n4288) );
  NAND2_X1 U5127 ( .A1(n4288), .A2(n4287), .ZN(n4289) );
  XOR2_X1 U5128 ( .A(n3438), .B(n4289), .Z(n4291) );
  AOI22_X1 U5129 ( .A1(n4689), .A2(\adder_stage2[7][11] ), .B1(n8387), .B2(
        n4291), .ZN(n4292) );
  INV_X1 U5130 ( .A(n4292), .ZN(n9675) );
  INV_X1 U5131 ( .A(n4293), .ZN(n4295) );
  NAND2_X1 U5132 ( .A1(n4295), .A2(n4294), .ZN(n4296) );
  XOR2_X1 U5133 ( .A(n4297), .B(n4296), .Z(n4298) );
  AOI22_X1 U5134 ( .A1(n4689), .A2(\adder_stage1[15][2] ), .B1(n8216), .B2(
        n4298), .ZN(n4299) );
  INV_X1 U5135 ( .A(n4299), .ZN(n9820) );
  BUF_X2 U5136 ( .A(n8282), .Z(n4596) );
  NOR2_X1 U5137 ( .A1(n4300), .A2(n4303), .ZN(n4312) );
  OAI21_X1 U5138 ( .B1(n4303), .B2(n4302), .A(n4301), .ZN(n4316) );
  AOI21_X1 U5139 ( .B1(n4304), .B2(n4312), .A(n4316), .ZN(n4336) );
  NOR2_X1 U5140 ( .A1(\x_mult_f[30][6] ), .A2(\x_mult_f[31][6] ), .ZN(n4332)
         );
  NAND2_X1 U5141 ( .A1(\x_mult_f[30][6] ), .A2(\x_mult_f[31][6] ), .ZN(n4333)
         );
  OAI21_X1 U5142 ( .B1(n4336), .B2(n4332), .A(n4333), .ZN(n4307) );
  NOR2_X1 U5143 ( .A1(\x_mult_f[30][7] ), .A2(\x_mult_f[31][7] ), .ZN(n4314)
         );
  INV_X1 U5144 ( .A(n4314), .ZN(n4305) );
  NAND2_X1 U5145 ( .A1(\x_mult_f[30][7] ), .A2(\x_mult_f[31][7] ), .ZN(n4313)
         );
  NAND2_X1 U5146 ( .A1(n4305), .A2(n4313), .ZN(n4306) );
  XNOR2_X1 U5147 ( .A(n4307), .B(n4306), .ZN(n4308) );
  AOI22_X1 U5148 ( .A1(n8048), .A2(\adder_stage1[15][7] ), .B1(n4596), .B2(
        n4308), .ZN(n4309) );
  INV_X1 U5149 ( .A(n4309), .ZN(n9815) );
  AOI22_X1 U5150 ( .A1(n8155), .A2(\x_mult_f[31][3] ), .B1(n4596), .B2(
        \x_mult_f_int[31][3] ), .ZN(n4310) );
  INV_X1 U5151 ( .A(n4310), .ZN(n9290) );
  AOI22_X1 U5152 ( .A1(n8212), .A2(\x_mult_f[31][1] ), .B1(n4596), .B2(
        \x_mult_f_int[31][1] ), .ZN(n4311) );
  INV_X1 U5153 ( .A(n4311), .ZN(n9354) );
  NOR2_X1 U5154 ( .A1(n4332), .A2(n4314), .ZN(n4317) );
  NAND2_X1 U5155 ( .A1(n4312), .A2(n4317), .ZN(n4319) );
  OAI21_X1 U5156 ( .B1(n4314), .B2(n4333), .A(n4313), .ZN(n4315) );
  AOI21_X1 U5157 ( .B1(n4317), .B2(n4316), .A(n4315), .ZN(n4318) );
  OAI21_X1 U5158 ( .B1(n4320), .B2(n4319), .A(n4318), .ZN(n4329) );
  OR2_X1 U5159 ( .A1(\x_mult_f[30][8] ), .A2(\x_mult_f[31][8] ), .ZN(n4327) );
  NAND2_X1 U5160 ( .A1(\x_mult_f[30][8] ), .A2(\x_mult_f[31][8] ), .ZN(n4326)
         );
  INV_X1 U5161 ( .A(n4326), .ZN(n4321) );
  AOI21_X1 U5162 ( .B1(n4329), .B2(n4327), .A(n4321), .ZN(n4341) );
  NOR2_X1 U5163 ( .A1(\x_mult_f[30][9] ), .A2(\x_mult_f[31][9] ), .ZN(n4340)
         );
  INV_X1 U5164 ( .A(n4340), .ZN(n4322) );
  NAND2_X1 U5165 ( .A1(\x_mult_f[30][9] ), .A2(\x_mult_f[31][9] ), .ZN(n4339)
         );
  NAND2_X1 U5166 ( .A1(n4322), .A2(n4339), .ZN(n4323) );
  XOR2_X1 U5167 ( .A(n4341), .B(n4323), .Z(n4324) );
  AOI22_X1 U5168 ( .A1(n8059), .A2(\adder_stage1[15][9] ), .B1(n4596), .B2(
        n4324), .ZN(n4325) );
  INV_X1 U5169 ( .A(n4325), .ZN(n9813) );
  NAND2_X1 U5170 ( .A1(n4327), .A2(n4326), .ZN(n4328) );
  XNOR2_X1 U5171 ( .A(n4329), .B(n4328), .ZN(n4330) );
  AOI22_X1 U5172 ( .A1(n5544), .A2(\adder_stage1[15][8] ), .B1(n4596), .B2(
        n4330), .ZN(n4331) );
  INV_X1 U5173 ( .A(n4331), .ZN(n9814) );
  INV_X1 U5174 ( .A(n4332), .ZN(n4334) );
  NAND2_X1 U5175 ( .A1(n4334), .A2(n4333), .ZN(n4335) );
  XOR2_X1 U5176 ( .A(n4336), .B(n4335), .Z(n4337) );
  AOI22_X1 U5177 ( .A1(n8036), .A2(\adder_stage1[15][6] ), .B1(n4596), .B2(
        n4337), .ZN(n4338) );
  INV_X1 U5178 ( .A(n4338), .ZN(n9816) );
  OAI21_X1 U5179 ( .B1(n4341), .B2(n4340), .A(n4339), .ZN(n6009) );
  OR2_X1 U5180 ( .A1(\x_mult_f[30][10] ), .A2(\x_mult_f[31][10] ), .ZN(n4721)
         );
  OR2_X1 U5181 ( .A1(\x_mult_f[30][11] ), .A2(\x_mult_f[31][11] ), .ZN(n4723)
         );
  AND2_X1 U5182 ( .A1(n4721), .A2(n4723), .ZN(n5681) );
  NAND2_X1 U5183 ( .A1(n6009), .A2(n5681), .ZN(n4343) );
  NAND2_X1 U5184 ( .A1(\x_mult_f[30][10] ), .A2(\x_mult_f[31][10] ), .ZN(n4348) );
  INV_X1 U5185 ( .A(n4348), .ZN(n4720) );
  NAND2_X1 U5186 ( .A1(\x_mult_f[30][11] ), .A2(\x_mult_f[31][11] ), .ZN(n4722) );
  INV_X1 U5187 ( .A(n4722), .ZN(n4342) );
  AOI21_X1 U5188 ( .B1(n4720), .B2(n4723), .A(n4342), .ZN(n5686) );
  NAND2_X1 U5189 ( .A1(n4343), .A2(n5686), .ZN(n4345) );
  OR2_X1 U5190 ( .A1(\x_mult_f[30][12] ), .A2(\x_mult_f[31][12] ), .ZN(n5683)
         );
  NAND2_X1 U5191 ( .A1(\x_mult_f[30][12] ), .A2(\x_mult_f[31][12] ), .ZN(n5684) );
  NAND2_X1 U5192 ( .A1(n5683), .A2(n5684), .ZN(n4344) );
  XNOR2_X1 U5193 ( .A(n4345), .B(n4344), .ZN(n4346) );
  AOI22_X1 U5194 ( .A1(n6373), .A2(\adder_stage1[15][12] ), .B1(n4596), .B2(
        n4346), .ZN(n4347) );
  INV_X1 U5195 ( .A(n4347), .ZN(n9810) );
  NAND2_X1 U5196 ( .A1(n4721), .A2(n4348), .ZN(n4349) );
  XNOR2_X1 U5197 ( .A(n6009), .B(n4349), .ZN(n4350) );
  AOI22_X1 U5198 ( .A1(n6330), .A2(\adder_stage1[15][10] ), .B1(n4596), .B2(
        n4350), .ZN(n4351) );
  INV_X1 U5199 ( .A(n4351), .ZN(n9812) );
  INV_X2 U5200 ( .A(n4526), .ZN(n6330) );
  INV_X1 U5201 ( .A(n4352), .ZN(n4386) );
  INV_X1 U5202 ( .A(n4353), .ZN(n4384) );
  INV_X1 U5203 ( .A(n4383), .ZN(n4354) );
  AOI21_X1 U5204 ( .B1(n4386), .B2(n4384), .A(n4354), .ZN(n4359) );
  INV_X1 U5205 ( .A(n4355), .ZN(n4357) );
  NAND2_X1 U5206 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  XOR2_X1 U5207 ( .A(n4359), .B(n4358), .Z(n4360) );
  AOI22_X1 U5208 ( .A1(n6330), .A2(\adder_stage2[7][5] ), .B1(n8216), .B2(
        n4360), .ZN(n4361) );
  INV_X1 U5209 ( .A(n4361), .ZN(n9681) );
  AOI21_X1 U5210 ( .B1(n4386), .B2(n4363), .A(n4362), .ZN(n4375) );
  INV_X1 U5211 ( .A(n4374), .ZN(n4364) );
  NAND2_X1 U5212 ( .A1(n4364), .A2(n4373), .ZN(n4365) );
  XOR2_X1 U5213 ( .A(n4375), .B(n4365), .Z(n4366) );
  AOI22_X1 U5214 ( .A1(n6330), .A2(\adder_stage2[7][6] ), .B1(n5950), .B2(
        n4366), .ZN(n4367) );
  INV_X1 U5215 ( .A(n4367), .ZN(n9680) );
  INV_X1 U5216 ( .A(n4368), .ZN(n4897) );
  INV_X1 U5217 ( .A(n4896), .ZN(n4369) );
  NAND2_X1 U5218 ( .A1(n4369), .A2(n4895), .ZN(n4370) );
  XOR2_X1 U5219 ( .A(n4897), .B(n4370), .Z(n4371) );
  AOI22_X1 U5220 ( .A1(n6330), .A2(\adder_stage2[7][2] ), .B1(n4596), .B2(
        n4371), .ZN(n4372) );
  INV_X1 U5221 ( .A(n4372), .ZN(n9684) );
  OAI21_X1 U5222 ( .B1(n4375), .B2(n4374), .A(n4373), .ZN(n4380) );
  INV_X1 U5223 ( .A(n4376), .ZN(n4378) );
  NAND2_X1 U5224 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  XNOR2_X1 U5225 ( .A(n4380), .B(n4379), .ZN(n4381) );
  AOI22_X1 U5226 ( .A1(n6330), .A2(\adder_stage2[7][7] ), .B1(n8387), .B2(
        n4381), .ZN(n4382) );
  INV_X1 U5227 ( .A(n4382), .ZN(n9679) );
  NAND2_X1 U5228 ( .A1(n4384), .A2(n4383), .ZN(n4385) );
  XNOR2_X1 U5229 ( .A(n4386), .B(n4385), .ZN(n4387) );
  AOI22_X1 U5230 ( .A1(n6330), .A2(\adder_stage2[7][4] ), .B1(n8365), .B2(
        n4387), .ZN(n4388) );
  INV_X1 U5231 ( .A(n4388), .ZN(n9682) );
  AOI22_X1 U5232 ( .A1(n8399), .A2(\x_mult_f_int[10][5] ), .B1(n8155), .B2(
        \x_mult_f[10][5] ), .ZN(n4389) );
  INV_X1 U5233 ( .A(n4389), .ZN(n9056) );
  NOR2_X1 U5234 ( .A1(\adder_stage3[0][2] ), .A2(\adder_stage3[1][2] ), .ZN(
        n6248) );
  NOR2_X1 U5235 ( .A1(\adder_stage3[0][3] ), .A2(\adder_stage3[1][3] ), .ZN(
        n6250) );
  NOR2_X1 U5236 ( .A1(n6248), .A2(n6250), .ZN(n4391) );
  NOR2_X1 U5237 ( .A1(\adder_stage3[0][1] ), .A2(\adder_stage3[1][1] ), .ZN(
        n6241) );
  NAND2_X1 U5238 ( .A1(\adder_stage3[0][0] ), .A2(\adder_stage3[1][0] ), .ZN(
        n6505) );
  NAND2_X1 U5239 ( .A1(\adder_stage3[0][1] ), .A2(\adder_stage3[1][1] ), .ZN(
        n6242) );
  OAI21_X1 U5240 ( .B1(n6241), .B2(n6505), .A(n6242), .ZN(n6236) );
  NAND2_X1 U5241 ( .A1(\adder_stage3[0][2] ), .A2(\adder_stage3[1][2] ), .ZN(
        n6247) );
  NAND2_X1 U5242 ( .A1(\adder_stage3[0][3] ), .A2(\adder_stage3[1][3] ), .ZN(
        n6251) );
  OAI21_X1 U5243 ( .B1(n6250), .B2(n6247), .A(n6251), .ZN(n4390) );
  AOI21_X1 U5244 ( .B1(n4391), .B2(n6236), .A(n4390), .ZN(n5734) );
  NOR2_X1 U5245 ( .A1(\adder_stage3[0][4] ), .A2(\adder_stage3[1][4] ), .ZN(
        n5735) );
  NOR2_X1 U5246 ( .A1(\adder_stage3[0][5] ), .A2(\adder_stage3[1][5] ), .ZN(
        n5737) );
  NOR2_X1 U5247 ( .A1(n5735), .A2(n5737), .ZN(n5745) );
  NOR2_X1 U5248 ( .A1(\adder_stage3[0][6] ), .A2(\adder_stage3[1][6] ), .ZN(
        n5775) );
  NOR2_X1 U5249 ( .A1(\adder_stage3[0][7] ), .A2(\adder_stage3[1][7] ), .ZN(
        n5746) );
  NOR2_X1 U5250 ( .A1(n5775), .A2(n5746), .ZN(n4393) );
  NAND2_X1 U5251 ( .A1(n5745), .A2(n4393), .ZN(n4395) );
  NAND2_X1 U5252 ( .A1(\adder_stage3[0][4] ), .A2(\adder_stage3[1][4] ), .ZN(
        n5769) );
  NAND2_X1 U5253 ( .A1(\adder_stage3[0][5] ), .A2(\adder_stage3[1][5] ), .ZN(
        n5738) );
  OAI21_X1 U5254 ( .B1(n5737), .B2(n5769), .A(n5738), .ZN(n5744) );
  NAND2_X1 U5255 ( .A1(\adder_stage3[0][6] ), .A2(\adder_stage3[1][6] ), .ZN(
        n5776) );
  NAND2_X1 U5256 ( .A1(\adder_stage3[0][7] ), .A2(\adder_stage3[1][7] ), .ZN(
        n5747) );
  OAI21_X1 U5257 ( .B1(n5746), .B2(n5776), .A(n5747), .ZN(n4392) );
  AOI21_X1 U5258 ( .B1(n4393), .B2(n5744), .A(n4392), .ZN(n4394) );
  OAI21_X1 U5259 ( .B1(n5734), .B2(n4395), .A(n4394), .ZN(n5694) );
  NOR2_X1 U5260 ( .A1(\adder_stage3[0][8] ), .A2(\adder_stage3[1][8] ), .ZN(
        n5760) );
  NOR2_X1 U5261 ( .A1(\adder_stage3[0][9] ), .A2(\adder_stage3[1][9] ), .ZN(
        n5762) );
  NOR2_X1 U5262 ( .A1(n5760), .A2(n5762), .ZN(n5715) );
  NOR2_X1 U5263 ( .A1(\adder_stage3[0][10] ), .A2(\adder_stage3[1][10] ), .ZN(
        n5719) );
  NOR2_X1 U5264 ( .A1(\adder_stage3[0][11] ), .A2(\adder_stage3[1][11] ), .ZN(
        n5721) );
  NOR2_X1 U5265 ( .A1(n5719), .A2(n5721), .ZN(n4397) );
  NAND2_X1 U5266 ( .A1(n5715), .A2(n4397), .ZN(n5696) );
  NOR2_X1 U5267 ( .A1(\adder_stage3[0][12] ), .A2(\adder_stage3[1][12] ), .ZN(
        n5697) );
  NOR2_X1 U5268 ( .A1(n5696), .A2(n5697), .ZN(n4399) );
  NAND2_X1 U5269 ( .A1(\adder_stage3[0][8] ), .A2(\adder_stage3[1][8] ), .ZN(
        n5759) );
  NAND2_X1 U5270 ( .A1(\adder_stage3[0][9] ), .A2(\adder_stage3[1][9] ), .ZN(
        n5763) );
  OAI21_X1 U5271 ( .B1(n5762), .B2(n5759), .A(n5763), .ZN(n5716) );
  NAND2_X1 U5272 ( .A1(\adder_stage3[0][10] ), .A2(\adder_stage3[1][10] ), 
        .ZN(n5728) );
  NAND2_X1 U5273 ( .A1(\adder_stage3[0][11] ), .A2(\adder_stage3[1][11] ), 
        .ZN(n5722) );
  OAI21_X1 U5274 ( .B1(n5721), .B2(n5728), .A(n5722), .ZN(n4396) );
  AOI21_X1 U5275 ( .B1(n4397), .B2(n5716), .A(n4396), .ZN(n5695) );
  NAND2_X1 U5276 ( .A1(\adder_stage3[0][12] ), .A2(\adder_stage3[1][12] ), 
        .ZN(n5698) );
  OAI21_X1 U5277 ( .B1(n5695), .B2(n5697), .A(n5698), .ZN(n4398) );
  AOI21_X1 U5278 ( .B1(n5694), .B2(n4399), .A(n4398), .ZN(n5712) );
  NOR2_X1 U5279 ( .A1(\adder_stage3[0][13] ), .A2(\adder_stage3[1][13] ), .ZN(
        n5708) );
  NAND2_X1 U5280 ( .A1(\adder_stage3[0][13] ), .A2(\adder_stage3[1][13] ), 
        .ZN(n5709) );
  OAI21_X1 U5281 ( .B1(n5712), .B2(n5708), .A(n5709), .ZN(n5756) );
  OR2_X1 U5282 ( .A1(\adder_stage3[0][14] ), .A2(\adder_stage3[1][14] ), .ZN(
        n5754) );
  NAND2_X1 U5283 ( .A1(\adder_stage3[0][14] ), .A2(\adder_stage3[1][14] ), 
        .ZN(n5753) );
  INV_X1 U5284 ( .A(n5753), .ZN(n4400) );
  AOI21_X1 U5285 ( .B1(n5756), .B2(n5754), .A(n4400), .ZN(n8308) );
  NOR2_X1 U5286 ( .A1(\adder_stage3[0][15] ), .A2(\adder_stage3[1][15] ), .ZN(
        n8304) );
  NAND2_X1 U5287 ( .A1(\adder_stage3[0][15] ), .A2(\adder_stage3[1][15] ), 
        .ZN(n8305) );
  OAI21_X1 U5288 ( .B1(n8308), .B2(n8304), .A(n8305), .ZN(n8255) );
  OR2_X1 U5289 ( .A1(\adder_stage3[0][16] ), .A2(\adder_stage3[1][16] ), .ZN(
        n4418) );
  OR2_X1 U5290 ( .A1(\adder_stage3[0][17] ), .A2(\adder_stage3[1][17] ), .ZN(
        n4409) );
  AND2_X1 U5291 ( .A1(n4418), .A2(n4409), .ZN(n4423) );
  NAND2_X1 U5292 ( .A1(n8255), .A2(n4423), .ZN(n4402) );
  NAND2_X1 U5293 ( .A1(\adder_stage3[0][16] ), .A2(\adder_stage3[1][16] ), 
        .ZN(n4417) );
  INV_X1 U5294 ( .A(n4417), .ZN(n4407) );
  NAND2_X1 U5295 ( .A1(\adder_stage3[0][17] ), .A2(\adder_stage3[1][17] ), 
        .ZN(n4408) );
  INV_X1 U5296 ( .A(n4408), .ZN(n4401) );
  AOI21_X1 U5297 ( .B1(n4407), .B2(n4409), .A(n4401), .ZN(n4427) );
  NAND2_X1 U5298 ( .A1(n4402), .A2(n4427), .ZN(n4404) );
  OR2_X1 U5299 ( .A1(\adder_stage3[0][18] ), .A2(\adder_stage3[1][18] ), .ZN(
        n4424) );
  NAND2_X1 U5300 ( .A1(\adder_stage3[0][18] ), .A2(\adder_stage3[1][18] ), 
        .ZN(n4425) );
  NAND2_X1 U5301 ( .A1(n4424), .A2(n4425), .ZN(n4403) );
  XNOR2_X1 U5302 ( .A(n4404), .B(n4403), .ZN(n4405) );
  AOI22_X1 U5303 ( .A1(n4405), .A2(n8265), .B1(n8078), .B2(
        \adder_stage4[0][18] ), .ZN(n4406) );
  INV_X1 U5304 ( .A(n4406), .ZN(n9570) );
  AOI21_X1 U5305 ( .B1(n8255), .B2(n4418), .A(n4407), .ZN(n4411) );
  NAND2_X1 U5306 ( .A1(n4409), .A2(n4408), .ZN(n4410) );
  XOR2_X1 U5307 ( .A(n4411), .B(n4410), .Z(n4412) );
  AOI22_X1 U5308 ( .A1(n4412), .A2(n8265), .B1(n8059), .B2(
        \adder_stage4[0][17] ), .ZN(n4413) );
  INV_X1 U5309 ( .A(n4413), .ZN(n9571) );
  AOI22_X1 U5310 ( .A1(\x_mult_f_int[10][7] ), .A2(n8216), .B1(n8212), .B2(
        \x_mult_f[10][7] ), .ZN(n4414) );
  INV_X1 U5311 ( .A(n4414), .ZN(n9054) );
  AOI22_X1 U5312 ( .A1(\x_mult_f_int[10][8] ), .A2(n8216), .B1(n8157), .B2(
        \x_mult_f[10][8] ), .ZN(n4415) );
  INV_X1 U5313 ( .A(n4415), .ZN(n9053) );
  AOI22_X1 U5314 ( .A1(\x_mult_f_int[11][13] ), .A2(n8186), .B1(n8078), .B2(
        \x_mult_f[11][13] ), .ZN(n4416) );
  INV_X1 U5315 ( .A(n4416), .ZN(n9060) );
  NAND2_X1 U5316 ( .A1(n4418), .A2(n4417), .ZN(n4419) );
  XNOR2_X1 U5317 ( .A(n8255), .B(n4419), .ZN(n4420) );
  AOI22_X1 U5318 ( .A1(n8229), .A2(n4420), .B1(n8059), .B2(
        \adder_stage4[0][16] ), .ZN(n4421) );
  INV_X1 U5319 ( .A(n4421), .ZN(n9572) );
  AOI22_X1 U5320 ( .A1(\x_mult_f_int[10][6] ), .A2(n8216), .B1(n8155), .B2(
        \x_mult_f[10][6] ), .ZN(n4422) );
  INV_X1 U5321 ( .A(n4422), .ZN(n9055) );
  AND2_X1 U5322 ( .A1(n4423), .A2(n4424), .ZN(n8253) );
  INV_X1 U5323 ( .A(n4424), .ZN(n4426) );
  OAI21_X1 U5324 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n8259) );
  AOI21_X1 U5325 ( .B1(n8255), .B2(n8253), .A(n8259), .ZN(n4429) );
  OR2_X1 U5326 ( .A1(\adder_stage3[0][19] ), .A2(\adder_stage3[1][19] ), .ZN(
        n8258) );
  NAND2_X1 U5327 ( .A1(\adder_stage3[0][19] ), .A2(\adder_stage3[1][19] ), 
        .ZN(n8256) );
  NAND2_X1 U5328 ( .A1(n8258), .A2(n8256), .ZN(n4428) );
  XOR2_X1 U5329 ( .A(n4429), .B(n4428), .Z(n4430) );
  AOI22_X1 U5330 ( .A1(n4430), .A2(n8265), .B1(n8212), .B2(
        \adder_stage4[0][19] ), .ZN(n4431) );
  INV_X1 U5331 ( .A(n4431), .ZN(n9569) );
  INV_X2 U5332 ( .A(n4651), .ZN(n4713) );
  AOI22_X1 U5333 ( .A1(n4713), .A2(\x_mult_f[25][3] ), .B1(n8203), .B2(
        \x_mult_f_int[25][3] ), .ZN(n4432) );
  INV_X1 U5334 ( .A(n4432), .ZN(n9228) );
  INV_X2 U5335 ( .A(n6588), .ZN(n7443) );
  INV_X1 U5336 ( .A(n4433), .ZN(n4460) );
  NAND2_X1 U5337 ( .A1(n4460), .A2(n4458), .ZN(n4434) );
  XNOR2_X1 U5338 ( .A(n4461), .B(n4434), .ZN(n4435) );
  AOI22_X1 U5339 ( .A1(n7443), .A2(\adder_stage1[11][4] ), .B1(n8318), .B2(
        n4435), .ZN(n4436) );
  INV_X1 U5340 ( .A(n4436), .ZN(n9886) );
  OR2_X1 U5341 ( .A1(\x_mult_f[22][0] ), .A2(\x_mult_f[23][0] ), .ZN(n4437) );
  AND2_X1 U5342 ( .A1(n4437), .A2(n4443), .ZN(n4438) );
  AOI22_X1 U5343 ( .A1(n7443), .A2(\adder_stage1[11][0] ), .B1(n8389), .B2(
        n4438), .ZN(n4439) );
  INV_X1 U5344 ( .A(n4439), .ZN(n9890) );
  INV_X1 U5345 ( .A(n4440), .ZN(n4442) );
  NAND2_X1 U5346 ( .A1(n4442), .A2(n4441), .ZN(n4444) );
  XOR2_X1 U5347 ( .A(n4444), .B(n4443), .Z(n4445) );
  AOI22_X1 U5348 ( .A1(n7443), .A2(\adder_stage1[11][1] ), .B1(n7356), .B2(
        n4445), .ZN(n4446) );
  INV_X1 U5349 ( .A(n4446), .ZN(n9889) );
  INV_X1 U5350 ( .A(n4447), .ZN(n4626) );
  OAI21_X1 U5351 ( .B1(n4626), .B2(n4622), .A(n4623), .ZN(n4452) );
  INV_X1 U5352 ( .A(n4448), .ZN(n4450) );
  NAND2_X1 U5353 ( .A1(n4450), .A2(n4449), .ZN(n4451) );
  XNOR2_X1 U5354 ( .A(n4452), .B(n4451), .ZN(n4453) );
  AOI22_X1 U5355 ( .A1(n7443), .A2(\adder_stage1[11][3] ), .B1(n8318), .B2(
        n4453), .ZN(n4454) );
  INV_X1 U5356 ( .A(n4454), .ZN(n9887) );
  OR2_X1 U5357 ( .A1(\adder_stage2[4][0] ), .A2(\adder_stage2[5][0] ), .ZN(
        n4455) );
  NAND2_X1 U5358 ( .A1(\adder_stage2[4][0] ), .A2(\adder_stage2[5][0] ), .ZN(
        n4709) );
  AND2_X1 U5359 ( .A1(n4455), .A2(n4709), .ZN(n4456) );
  AOI22_X1 U5360 ( .A1(n4713), .A2(\adder_stage3[2][0] ), .B1(n8401), .B2(
        n4456), .ZN(n4457) );
  INV_X1 U5361 ( .A(n4457), .ZN(n9629) );
  INV_X1 U5362 ( .A(n4458), .ZN(n4459) );
  AOI21_X1 U5363 ( .B1(n4461), .B2(n4460), .A(n4459), .ZN(n4466) );
  INV_X1 U5364 ( .A(n4462), .ZN(n4464) );
  NAND2_X1 U5365 ( .A1(n4464), .A2(n4463), .ZN(n4465) );
  XOR2_X1 U5366 ( .A(n4466), .B(n4465), .Z(n4467) );
  AOI22_X1 U5367 ( .A1(n7443), .A2(\adder_stage1[11][5] ), .B1(n8318), .B2(
        n4467), .ZN(n4468) );
  INV_X1 U5368 ( .A(n4468), .ZN(n9885) );
  AOI22_X1 U5369 ( .A1(n4713), .A2(\x_mult_f[24][0] ), .B1(n8365), .B2(
        \x_mult_f_int[24][0] ), .ZN(n4469) );
  INV_X1 U5370 ( .A(n4469), .ZN(n9341) );
  NOR2_X1 U5371 ( .A1(\adder_stage2[4][1] ), .A2(\adder_stage2[5][1] ), .ZN(
        n4706) );
  NAND2_X1 U5372 ( .A1(\adder_stage2[4][1] ), .A2(\adder_stage2[5][1] ), .ZN(
        n4707) );
  OAI21_X1 U5373 ( .B1(n4706), .B2(n4709), .A(n4707), .ZN(n4475) );
  INV_X1 U5374 ( .A(n4475), .ZN(n4697) );
  NOR2_X1 U5375 ( .A1(\adder_stage2[4][2] ), .A2(\adder_stage2[5][2] ), .ZN(
        n4696) );
  INV_X1 U5376 ( .A(n4696), .ZN(n4470) );
  NAND2_X1 U5377 ( .A1(\adder_stage2[5][2] ), .A2(\adder_stage2[4][2] ), .ZN(
        n4695) );
  NAND2_X1 U5378 ( .A1(n4470), .A2(n4695), .ZN(n4471) );
  XOR2_X1 U5379 ( .A(n4697), .B(n4471), .Z(n4472) );
  AOI22_X1 U5380 ( .A1(n4713), .A2(\adder_stage3[2][2] ), .B1(n8213), .B2(
        n4472), .ZN(n4473) );
  INV_X1 U5381 ( .A(n4473), .ZN(n9627) );
  NOR2_X1 U5382 ( .A1(\adder_stage2[4][3] ), .A2(\adder_stage2[5][3] ), .ZN(
        n4698) );
  NOR2_X1 U5383 ( .A1(n4696), .A2(n4698), .ZN(n4476) );
  NAND2_X1 U5384 ( .A1(\adder_stage2[4][3] ), .A2(\adder_stage2[5][3] ), .ZN(
        n4699) );
  OAI21_X1 U5385 ( .B1(n4698), .B2(n4695), .A(n4699), .ZN(n4474) );
  AOI21_X1 U5386 ( .B1(n4476), .B2(n4475), .A(n4474), .ZN(n4915) );
  INV_X1 U5387 ( .A(n4915), .ZN(n4557) );
  NOR2_X1 U5388 ( .A1(\adder_stage2[4][4] ), .A2(\adder_stage2[5][4] ), .ZN(
        n4553) );
  INV_X1 U5389 ( .A(n4553), .ZN(n4547) );
  NAND2_X1 U5390 ( .A1(\adder_stage2[4][4] ), .A2(\adder_stage2[5][4] ), .ZN(
        n4555) );
  NAND2_X1 U5391 ( .A1(n4547), .A2(n4555), .ZN(n4477) );
  XNOR2_X1 U5392 ( .A(n4557), .B(n4477), .ZN(n4478) );
  AOI22_X1 U5393 ( .A1(n4713), .A2(\adder_stage3[2][4] ), .B1(n4596), .B2(
        n4478), .ZN(n4479) );
  INV_X1 U5394 ( .A(n4479), .ZN(n9625) );
  AOI22_X1 U5395 ( .A1(\x_mult_f_int[17][6] ), .A2(n8213), .B1(n8386), .B2(
        \x_mult_f[17][6] ), .ZN(n4480) );
  INV_X1 U5396 ( .A(n4480), .ZN(n9149) );
  AOI22_X1 U5397 ( .A1(\x_mult_f_int[17][7] ), .A2(n8401), .B1(n8386), .B2(
        \x_mult_f[17][7] ), .ZN(n4481) );
  INV_X1 U5398 ( .A(n4481), .ZN(n9148) );
  NAND2_X1 U5399 ( .A1(n4483), .A2(n4482), .ZN(n4484) );
  XNOR2_X1 U5400 ( .A(n3446), .B(n4484), .ZN(n4486) );
  AOI22_X1 U5401 ( .A1(n6330), .A2(\adder_stage3[3][14] ), .B1(n7029), .B2(
        n4486), .ZN(n4487) );
  INV_X1 U5402 ( .A(n4487), .ZN(n9595) );
  INV_X1 U5403 ( .A(n4488), .ZN(n4490) );
  NAND2_X1 U5404 ( .A1(n4490), .A2(n4489), .ZN(n4491) );
  XOR2_X1 U5405 ( .A(n4492), .B(n4491), .Z(n4493) );
  AOI22_X1 U5406 ( .A1(n6330), .A2(\adder_stage3[3][13] ), .B1(n8399), .B2(
        n4493), .ZN(n4494) );
  INV_X1 U5407 ( .A(n4494), .ZN(n9596) );
  INV_X1 U5408 ( .A(n4495), .ZN(n4497) );
  NAND2_X1 U5409 ( .A1(n4497), .A2(n4496), .ZN(n4498) );
  XOR2_X1 U5410 ( .A(n4499), .B(n4498), .Z(n4500) );
  AOI22_X1 U5411 ( .A1(n6330), .A2(\adder_stage3[3][15] ), .B1(n7117), .B2(
        n4500), .ZN(n4501) );
  INV_X1 U5412 ( .A(n4501), .ZN(n9594) );
  OAI21_X1 U5413 ( .B1(n4504), .B2(n4503), .A(n4502), .ZN(n4509) );
  INV_X1 U5414 ( .A(n4505), .ZN(n4507) );
  NAND2_X1 U5415 ( .A1(n4507), .A2(n4506), .ZN(n4508) );
  XNOR2_X1 U5416 ( .A(n4509), .B(n4508), .ZN(n4510) );
  AOI22_X1 U5417 ( .A1(n6330), .A2(\adder_stage3[3][12] ), .B1(n8390), .B2(
        n4510), .ZN(n4511) );
  INV_X1 U5418 ( .A(n4511), .ZN(n9597) );
  INV_X2 U5419 ( .A(n4512), .ZN(n8392) );
  AOI22_X1 U5420 ( .A1(\x_mult_f_int[21][12] ), .A2(n8265), .B1(n8392), .B2(
        \x_mult_f[21][12] ), .ZN(n4513) );
  INV_X1 U5421 ( .A(n4513), .ZN(n9191) );
  AOI22_X1 U5422 ( .A1(\x_mult_f_int[21][11] ), .A2(n8401), .B1(n8392), .B2(
        \x_mult_f[21][11] ), .ZN(n4514) );
  INV_X1 U5423 ( .A(n4514), .ZN(n9192) );
  AOI22_X1 U5424 ( .A1(n6643), .A2(\x_mult_f_int[20][5] ), .B1(n8392), .B2(
        \x_mult_f[20][5] ), .ZN(n4515) );
  INV_X1 U5425 ( .A(n4515), .ZN(n9184) );
  AOI22_X1 U5426 ( .A1(\x_mult_f_int[20][6] ), .A2(n8203), .B1(n8392), .B2(
        \x_mult_f[20][6] ), .ZN(n4516) );
  INV_X1 U5427 ( .A(n4516), .ZN(n9183) );
  BUF_X2 U5428 ( .A(n6122), .Z(n4651) );
  INV_X2 U5429 ( .A(n4651), .ZN(n5544) );
  AOI22_X1 U5430 ( .A1(n5544), .A2(\x_mult_f[29][3] ), .B1(n8363), .B2(
        \x_mult_f_int[29][3] ), .ZN(n4517) );
  INV_X1 U5431 ( .A(n4517), .ZN(n9262) );
  INV_X1 U5432 ( .A(n4518), .ZN(n4520) );
  NAND2_X1 U5433 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  XOR2_X1 U5434 ( .A(n4522), .B(n4521), .Z(n4523) );
  AOI22_X1 U5435 ( .A1(n7775), .A2(\adder_stage1[11][6] ), .B1(n8329), .B2(
        n4523), .ZN(n4524) );
  INV_X1 U5436 ( .A(n4524), .ZN(n9884) );
  AOI22_X1 U5437 ( .A1(n5544), .A2(\x_mult_f[29][4] ), .B1(n7698), .B2(
        \x_mult_f_int[29][4] ), .ZN(n4525) );
  INV_X1 U5438 ( .A(n4525), .ZN(n9261) );
  INV_X1 U5439 ( .A(n4527), .ZN(n5040) );
  INV_X1 U5440 ( .A(n4528), .ZN(n5038) );
  INV_X1 U5441 ( .A(n5037), .ZN(n4529) );
  AOI21_X1 U5442 ( .B1(n5040), .B2(n5038), .A(n4529), .ZN(n4534) );
  INV_X1 U5443 ( .A(n4530), .ZN(n4532) );
  NAND2_X1 U5444 ( .A1(n4532), .A2(n4531), .ZN(n4533) );
  XOR2_X1 U5445 ( .A(n4534), .B(n4533), .Z(n4535) );
  AOI22_X1 U5446 ( .A1(n8218), .A2(\adder_stage1[13][5] ), .B1(n7117), .B2(
        n4535), .ZN(n4536) );
  INV_X1 U5447 ( .A(n4536), .ZN(n9851) );
  AOI22_X1 U5448 ( .A1(n5544), .A2(\x_mult_f[29][0] ), .B1(n8390), .B2(
        \x_mult_f_int[29][0] ), .ZN(n4537) );
  INV_X1 U5449 ( .A(n4537), .ZN(n9351) );
  INV_X1 U5450 ( .A(n4538), .ZN(n4540) );
  NAND2_X1 U5451 ( .A1(n4540), .A2(n4539), .ZN(n4541) );
  XOR2_X1 U5452 ( .A(n4542), .B(n4541), .Z(n4543) );
  AOI22_X1 U5453 ( .A1(n8157), .A2(\adder_stage1[13][9] ), .B1(n8282), .B2(
        n4543), .ZN(n4544) );
  INV_X1 U5454 ( .A(n4544), .ZN(n9847) );
  AOI22_X1 U5455 ( .A1(n5294), .A2(\x_mult_f[27][0] ), .B1(n7110), .B2(
        \x_mult_f_int[27][0] ), .ZN(n4545) );
  INV_X1 U5456 ( .A(n4545), .ZN(n9347) );
  INV_X1 U5457 ( .A(n4555), .ZN(n4546) );
  AOI21_X1 U5458 ( .B1(n4557), .B2(n4547), .A(n4546), .ZN(n4550) );
  NOR2_X1 U5459 ( .A1(\adder_stage2[4][5] ), .A2(\adder_stage2[5][5] ), .ZN(
        n4556) );
  INV_X1 U5460 ( .A(n4556), .ZN(n4548) );
  NAND2_X1 U5461 ( .A1(\adder_stage2[4][5] ), .A2(\adder_stage2[5][5] ), .ZN(
        n4554) );
  NAND2_X1 U5462 ( .A1(n4548), .A2(n4554), .ZN(n4549) );
  XOR2_X1 U5463 ( .A(n4550), .B(n4549), .Z(n4551) );
  AOI22_X1 U5464 ( .A1(n8157), .A2(\adder_stage3[2][5] ), .B1(n5950), .B2(
        n4551), .ZN(n4552) );
  INV_X1 U5465 ( .A(n4552), .ZN(n9624) );
  NOR2_X1 U5466 ( .A1(n4553), .A2(n4556), .ZN(n4906) );
  OAI21_X1 U5467 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n4911) );
  AOI21_X1 U5468 ( .B1(n4557), .B2(n4906), .A(n4911), .ZN(n4564) );
  NOR2_X1 U5469 ( .A1(\adder_stage2[4][6] ), .A2(\adder_stage2[5][6] ), .ZN(
        n4905) );
  INV_X1 U5470 ( .A(n4905), .ZN(n4558) );
  NAND2_X1 U5471 ( .A1(\adder_stage2[4][6] ), .A2(\adder_stage2[5][6] ), .ZN(
        n4908) );
  NAND2_X1 U5472 ( .A1(n4558), .A2(n4908), .ZN(n4559) );
  XOR2_X1 U5473 ( .A(n4564), .B(n4559), .Z(n4560) );
  AOI22_X1 U5474 ( .A1(n5273), .A2(\adder_stage3[2][6] ), .B1(n8401), .B2(
        n4560), .ZN(n4561) );
  INV_X1 U5475 ( .A(n4561), .ZN(n9623) );
  AOI22_X1 U5476 ( .A1(n5544), .A2(\x_mult_f[29][1] ), .B1(n8401), .B2(
        \x_mult_f_int[29][1] ), .ZN(n4562) );
  INV_X1 U5477 ( .A(n4562), .ZN(n9350) );
  AOI22_X1 U5478 ( .A1(n5544), .A2(\x_mult_f[27][1] ), .B1(n8389), .B2(
        \x_mult_f_int[27][1] ), .ZN(n4563) );
  INV_X1 U5479 ( .A(n4563), .ZN(n9346) );
  OAI21_X1 U5480 ( .B1(n4564), .B2(n4905), .A(n4908), .ZN(n4567) );
  NOR2_X1 U5481 ( .A1(\adder_stage2[4][7] ), .A2(\adder_stage2[5][7] ), .ZN(
        n4909) );
  INV_X1 U5482 ( .A(n4909), .ZN(n4565) );
  NAND2_X1 U5483 ( .A1(\adder_stage2[4][7] ), .A2(\adder_stage2[5][7] ), .ZN(
        n4907) );
  NAND2_X1 U5484 ( .A1(n4565), .A2(n4907), .ZN(n4566) );
  XNOR2_X1 U5485 ( .A(n4567), .B(n4566), .ZN(n4568) );
  AOI22_X1 U5486 ( .A1(n7775), .A2(\adder_stage3[2][7] ), .B1(n5921), .B2(
        n4568), .ZN(n4569) );
  INV_X1 U5487 ( .A(n4569), .ZN(n9622) );
  NOR2_X1 U5488 ( .A1(\x_mult_f[0][2] ), .A2(\x_mult_f[1][2] ), .ZN(n7587) );
  NOR2_X1 U5489 ( .A1(\x_mult_f[0][3] ), .A2(\x_mult_f[1][3] ), .ZN(n7566) );
  NOR2_X1 U5490 ( .A1(n7587), .A2(n7566), .ZN(n4571) );
  NOR2_X1 U5491 ( .A1(\x_mult_f[0][1] ), .A2(\x_mult_f[1][1] ), .ZN(n7672) );
  NAND2_X1 U5492 ( .A1(\x_mult_f[0][0] ), .A2(\x_mult_f[1][0] ), .ZN(n7675) );
  NAND2_X1 U5493 ( .A1(\x_mult_f[0][1] ), .A2(\x_mult_f[1][1] ), .ZN(n7673) );
  OAI21_X1 U5494 ( .B1(n7672), .B2(n7675), .A(n7673), .ZN(n7565) );
  NAND2_X1 U5495 ( .A1(\x_mult_f[0][2] ), .A2(\x_mult_f[1][2] ), .ZN(n7588) );
  NAND2_X1 U5496 ( .A1(\x_mult_f[0][3] ), .A2(\x_mult_f[1][3] ), .ZN(n7567) );
  OAI21_X1 U5497 ( .B1(n7566), .B2(n7588), .A(n7567), .ZN(n4570) );
  AOI21_X1 U5498 ( .B1(n4571), .B2(n7565), .A(n4570), .ZN(n7514) );
  NOR2_X1 U5499 ( .A1(\x_mult_f[0][4] ), .A2(\x_mult_f[1][4] ), .ZN(n7515) );
  NOR2_X1 U5500 ( .A1(\x_mult_f[0][5] ), .A2(\x_mult_f[1][5] ), .ZN(n7517) );
  NOR2_X1 U5501 ( .A1(n7515), .A2(n7517), .ZN(n7541) );
  NOR2_X1 U5502 ( .A1(\x_mult_f[0][6] ), .A2(\x_mult_f[1][6] ), .ZN(n7579) );
  NOR2_X1 U5503 ( .A1(\x_mult_f[0][7] ), .A2(\x_mult_f[1][7] ), .ZN(n7542) );
  NOR2_X1 U5504 ( .A1(n7579), .A2(n7542), .ZN(n4573) );
  NAND2_X1 U5505 ( .A1(n7541), .A2(n4573), .ZN(n4575) );
  NAND2_X1 U5506 ( .A1(\x_mult_f[1][4] ), .A2(\x_mult_f[0][4] ), .ZN(n7559) );
  NAND2_X1 U5507 ( .A1(\x_mult_f[0][5] ), .A2(\x_mult_f[1][5] ), .ZN(n7518) );
  OAI21_X1 U5508 ( .B1(n7517), .B2(n7559), .A(n7518), .ZN(n7540) );
  NAND2_X1 U5509 ( .A1(\x_mult_f[0][6] ), .A2(\x_mult_f[1][6] ), .ZN(n7580) );
  NAND2_X1 U5510 ( .A1(\x_mult_f[0][7] ), .A2(\x_mult_f[1][7] ), .ZN(n7543) );
  OAI21_X1 U5511 ( .B1(n7542), .B2(n7580), .A(n7543), .ZN(n4572) );
  AOI21_X1 U5512 ( .B1(n4573), .B2(n7540), .A(n4572), .ZN(n4574) );
  OAI21_X1 U5513 ( .B1(n7514), .B2(n4575), .A(n4574), .ZN(n7664) );
  OR2_X1 U5514 ( .A1(\x_mult_f[0][11] ), .A2(\x_mult_f[1][11] ), .ZN(n7667) );
  NAND2_X1 U5515 ( .A1(n7664), .A2(n7667), .ZN(n4582) );
  OR2_X1 U5516 ( .A1(\x_mult_f[0][8] ), .A2(\x_mult_f[1][8] ), .ZN(n7632) );
  OR2_X1 U5517 ( .A1(\x_mult_f[0][9] ), .A2(\x_mult_f[1][9] ), .ZN(n7529) );
  AND2_X1 U5518 ( .A1(n7632), .A2(n7529), .ZN(n7600) );
  OR2_X1 U5519 ( .A1(\x_mult_f[0][10] ), .A2(\x_mult_f[1][10] ), .ZN(n7602) );
  NAND2_X1 U5520 ( .A1(n7600), .A2(n7602), .ZN(n7659) );
  NAND2_X1 U5521 ( .A1(\x_mult_f[0][8] ), .A2(\x_mult_f[1][8] ), .ZN(n7631) );
  INV_X1 U5522 ( .A(n7631), .ZN(n7527) );
  NAND2_X1 U5523 ( .A1(\x_mult_f[0][9] ), .A2(\x_mult_f[1][9] ), .ZN(n7528) );
  INV_X1 U5524 ( .A(n7528), .ZN(n4576) );
  AOI21_X1 U5525 ( .B1(n7527), .B2(n7529), .A(n4576), .ZN(n7662) );
  INV_X1 U5526 ( .A(n7662), .ZN(n4580) );
  INV_X1 U5527 ( .A(n7602), .ZN(n7661) );
  INV_X1 U5528 ( .A(n7667), .ZN(n4577) );
  NOR2_X1 U5529 ( .A1(n7661), .A2(n4577), .ZN(n4579) );
  NAND2_X1 U5530 ( .A1(\x_mult_f[0][10] ), .A2(\x_mult_f[1][10] ), .ZN(n7660)
         );
  NAND2_X1 U5531 ( .A1(\x_mult_f[0][11] ), .A2(\x_mult_f[1][11] ), .ZN(n7666)
         );
  OAI21_X1 U5532 ( .B1(n7660), .B2(n4577), .A(n7666), .ZN(n4578) );
  AOI21_X1 U5533 ( .B1(n4580), .B2(n4579), .A(n4578), .ZN(n4581) );
  OAI21_X1 U5534 ( .B1(n4582), .B2(n7659), .A(n4581), .ZN(n7576) );
  OR2_X1 U5535 ( .A1(\x_mult_f[0][12] ), .A2(\x_mult_f[1][12] ), .ZN(n7574) );
  NAND2_X1 U5536 ( .A1(\x_mult_f[0][12] ), .A2(\x_mult_f[1][12] ), .ZN(n7573)
         );
  INV_X1 U5537 ( .A(n7573), .ZN(n4583) );
  AOI21_X1 U5538 ( .B1(n7576), .B2(n7574), .A(n4583), .ZN(n4743) );
  NOR2_X1 U5539 ( .A1(\x_mult_f[0][13] ), .A2(\x_mult_f[1][13] ), .ZN(n4739)
         );
  NAND2_X1 U5540 ( .A1(\x_mult_f[0][13] ), .A2(\x_mult_f[1][13] ), .ZN(n4740)
         );
  OAI21_X1 U5541 ( .B1(n4743), .B2(n4739), .A(n4740), .ZN(n4746) );
  INV_X1 U5542 ( .A(n4584), .ZN(n4585) );
  AOI22_X1 U5543 ( .A1(n4585), .A2(n6643), .B1(n8200), .B2(
        \adder_stage1[0][20] ), .ZN(n4586) );
  INV_X1 U5544 ( .A(n4586), .ZN(n10054) );
  INV_X2 U5545 ( .A(n4651), .ZN(n5294) );
  INV_X1 U5546 ( .A(n4587), .ZN(n5077) );
  INV_X1 U5547 ( .A(n5076), .ZN(n4588) );
  NAND2_X1 U5548 ( .A1(n4588), .A2(n5075), .ZN(n4589) );
  XOR2_X1 U5549 ( .A(n5077), .B(n4589), .Z(n4590) );
  AOI22_X1 U5550 ( .A1(n5294), .A2(\adder_stage1[14][2] ), .B1(n4596), .B2(
        n4590), .ZN(n4591) );
  INV_X1 U5551 ( .A(n4591), .ZN(n9837) );
  OR2_X1 U5552 ( .A1(\x_mult_f[28][0] ), .A2(\x_mult_f[29][0] ), .ZN(n4592) );
  AND2_X1 U5553 ( .A1(n4592), .A2(n4602), .ZN(n4593) );
  AOI22_X1 U5554 ( .A1(n5294), .A2(\adder_stage1[14][0] ), .B1(n4596), .B2(
        n4593), .ZN(n4594) );
  INV_X1 U5555 ( .A(n4594), .ZN(n9839) );
  INV_X2 U5556 ( .A(n4715), .ZN(n5273) );
  AOI22_X1 U5557 ( .A1(n5273), .A2(\x_mult_f[27][3] ), .B1(n5950), .B2(
        \x_mult_f_int[27][3] ), .ZN(n4595) );
  INV_X1 U5558 ( .A(n4595), .ZN(n9245) );
  AOI22_X1 U5559 ( .A1(n7775), .A2(\x_mult_f[25][0] ), .B1(n7698), .B2(
        \x_mult_f_int[25][0] ), .ZN(n4597) );
  INV_X1 U5560 ( .A(n4597), .ZN(n9343) );
  AOI22_X1 U5561 ( .A1(n5273), .A2(\x_mult_f[27][2] ), .B1(n5950), .B2(
        \x_mult_f_int[27][2] ), .ZN(n4598) );
  INV_X1 U5562 ( .A(n4598), .ZN(n9246) );
  INV_X1 U5563 ( .A(n4599), .ZN(n4601) );
  NAND2_X1 U5564 ( .A1(n4601), .A2(n4600), .ZN(n4603) );
  XOR2_X1 U5565 ( .A(n4603), .B(n4602), .Z(n4604) );
  AOI22_X1 U5566 ( .A1(n5294), .A2(\adder_stage1[14][1] ), .B1(n4596), .B2(
        n4604), .ZN(n4605) );
  INV_X1 U5567 ( .A(n4605), .ZN(n9838) );
  AOI22_X1 U5568 ( .A1(n5273), .A2(\x_mult_f[27][4] ), .B1(n5950), .B2(
        \x_mult_f_int[27][4] ), .ZN(n4606) );
  INV_X1 U5569 ( .A(n4606), .ZN(n9244) );
  AOI22_X1 U5570 ( .A1(n6337), .A2(\x_mult_f[25][1] ), .B1(n7284), .B2(
        \x_mult_f_int[25][1] ), .ZN(n4607) );
  INV_X1 U5571 ( .A(n4607), .ZN(n9342) );
  NOR2_X1 U5572 ( .A1(\adder_stage1[10][2] ), .A2(\adder_stage1[11][2] ), .ZN(
        n4773) );
  NOR2_X1 U5573 ( .A1(n4773), .A2(n4657), .ZN(n4609) );
  NOR2_X1 U5574 ( .A1(\adder_stage1[10][1] ), .A2(\adder_stage1[11][1] ), .ZN(
        n6332) );
  NAND2_X1 U5575 ( .A1(\adder_stage1[10][0] ), .A2(\adder_stage1[11][0] ), 
        .ZN(n6339) );
  NAND2_X1 U5576 ( .A1(\adder_stage1[10][1] ), .A2(\adder_stage1[11][1] ), 
        .ZN(n6333) );
  OAI21_X1 U5577 ( .B1(n6332), .B2(n6339), .A(n6333), .ZN(n4656) );
  NAND2_X1 U5578 ( .A1(\adder_stage1[10][2] ), .A2(\adder_stage1[11][2] ), 
        .ZN(n4774) );
  NAND2_X1 U5579 ( .A1(\adder_stage1[10][3] ), .A2(\adder_stage1[11][3] ), 
        .ZN(n4658) );
  OAI21_X1 U5580 ( .B1(n4657), .B2(n4774), .A(n4658), .ZN(n4608) );
  AOI21_X1 U5581 ( .B1(n4609), .B2(n4656), .A(n4608), .ZN(n4751) );
  NOR2_X1 U5582 ( .A1(\adder_stage1[10][4] ), .A2(\adder_stage1[11][4] ), .ZN(
        n4752) );
  NOR2_X1 U5583 ( .A1(\adder_stage1[10][5] ), .A2(\adder_stage1[11][5] ), .ZN(
        n4754) );
  NOR2_X1 U5584 ( .A1(n4752), .A2(n4754), .ZN(n4765) );
  NOR2_X1 U5585 ( .A1(\adder_stage1[10][6] ), .A2(\adder_stage1[11][6] ), .ZN(
        n4814) );
  NOR2_X1 U5586 ( .A1(\adder_stage1[10][7] ), .A2(\adder_stage1[11][7] ), .ZN(
        n4766) );
  NOR2_X1 U5587 ( .A1(n4814), .A2(n4766), .ZN(n4611) );
  NAND2_X1 U5588 ( .A1(n4765), .A2(n4611), .ZN(n4613) );
  NAND2_X1 U5589 ( .A1(\adder_stage1[10][4] ), .A2(\adder_stage1[11][4] ), 
        .ZN(n4799) );
  NAND2_X1 U5590 ( .A1(\adder_stage1[10][5] ), .A2(\adder_stage1[11][5] ), 
        .ZN(n4755) );
  OAI21_X1 U5591 ( .B1(n4754), .B2(n4799), .A(n4755), .ZN(n4764) );
  NAND2_X1 U5592 ( .A1(\adder_stage1[10][6] ), .A2(\adder_stage1[11][6] ), 
        .ZN(n4815) );
  NAND2_X1 U5593 ( .A1(\adder_stage1[10][7] ), .A2(\adder_stage1[11][7] ), 
        .ZN(n4767) );
  OAI21_X1 U5594 ( .B1(n4766), .B2(n4815), .A(n4767), .ZN(n4610) );
  AOI21_X1 U5595 ( .B1(n4611), .B2(n4764), .A(n4610), .ZN(n4612) );
  OAI21_X1 U5596 ( .B1(n4751), .B2(n4613), .A(n4612), .ZN(n4780) );
  NOR2_X1 U5597 ( .A1(\adder_stage1[10][8] ), .A2(\adder_stage1[11][8] ), .ZN(
        n4781) );
  INV_X1 U5598 ( .A(n4781), .ZN(n4822) );
  OR2_X1 U5599 ( .A1(\adder_stage1[10][9] ), .A2(\adder_stage1[11][9] ), .ZN(
        n4783) );
  NAND2_X1 U5600 ( .A1(n4822), .A2(n4783), .ZN(n4806) );
  NOR2_X1 U5601 ( .A1(\adder_stage1[10][10] ), .A2(\adder_stage1[11][10] ), 
        .ZN(n4807) );
  NOR2_X1 U5602 ( .A1(n4806), .A2(n4807), .ZN(n4617) );
  NAND2_X1 U5603 ( .A1(\adder_stage1[10][8] ), .A2(\adder_stage1[11][8] ), 
        .ZN(n4821) );
  INV_X1 U5604 ( .A(n4821), .ZN(n4615) );
  NAND2_X1 U5605 ( .A1(\adder_stage1[10][9] ), .A2(\adder_stage1[11][9] ), 
        .ZN(n4782) );
  INV_X1 U5606 ( .A(n4782), .ZN(n4614) );
  AOI21_X1 U5607 ( .B1(n4783), .B2(n4615), .A(n4614), .ZN(n4805) );
  NAND2_X1 U5608 ( .A1(\adder_stage1[10][10] ), .A2(\adder_stage1[11][10] ), 
        .ZN(n4808) );
  OAI21_X1 U5609 ( .B1(n4805), .B2(n4807), .A(n4808), .ZN(n4616) );
  AOI21_X1 U5610 ( .B1(n4780), .B2(n4617), .A(n4616), .ZN(n4796) );
  NOR2_X1 U5611 ( .A1(\adder_stage1[10][11] ), .A2(\adder_stage1[11][11] ), 
        .ZN(n4793) );
  NAND2_X1 U5612 ( .A1(\adder_stage1[10][11] ), .A2(\adder_stage1[11][11] ), 
        .ZN(n4794) );
  OR2_X1 U5613 ( .A1(\adder_stage1[10][12] ), .A2(\adder_stage1[11][12] ), 
        .ZN(n4828) );
  NAND2_X1 U5614 ( .A1(\adder_stage1[10][12] ), .A2(\adder_stage1[11][12] ), 
        .ZN(n4827) );
  INV_X1 U5615 ( .A(n4827), .ZN(n4618) );
  NOR2_X1 U5616 ( .A1(\adder_stage1[10][13] ), .A2(\adder_stage1[11][13] ), 
        .ZN(n4629) );
  NAND2_X1 U5617 ( .A1(\adder_stage1[10][13] ), .A2(\adder_stage1[11][13] ), 
        .ZN(n4630) );
  OR2_X1 U5618 ( .A1(\adder_stage1[10][14] ), .A2(\adder_stage1[11][14] ), 
        .ZN(n5470) );
  NAND2_X1 U5619 ( .A1(\adder_stage1[10][14] ), .A2(\adder_stage1[11][14] ), 
        .ZN(n5468) );
  NAND2_X1 U5620 ( .A1(n5470), .A2(n5468), .ZN(n4619) );
  XNOR2_X1 U5621 ( .A(n5471), .B(n4619), .ZN(n4620) );
  AOI22_X1 U5622 ( .A1(n7443), .A2(\adder_stage2[5][14] ), .B1(n7698), .B2(
        n4620), .ZN(n4621) );
  INV_X1 U5623 ( .A(n4621), .ZN(n9706) );
  INV_X1 U5624 ( .A(n4622), .ZN(n4624) );
  NAND2_X1 U5625 ( .A1(n4624), .A2(n4623), .ZN(n4625) );
  XOR2_X1 U5626 ( .A(n4626), .B(n4625), .Z(n4627) );
  AOI22_X1 U5627 ( .A1(n7443), .A2(\adder_stage1[11][2] ), .B1(n8329), .B2(
        n4627), .ZN(n4628) );
  INV_X1 U5628 ( .A(n4628), .ZN(n9888) );
  INV_X1 U5629 ( .A(n4629), .ZN(n4631) );
  NAND2_X1 U5630 ( .A1(n4631), .A2(n4630), .ZN(n4632) );
  XOR2_X1 U5631 ( .A(n4633), .B(n4632), .Z(n4634) );
  AOI22_X1 U5632 ( .A1(n7443), .A2(\adder_stage2[5][13] ), .B1(n8037), .B2(
        n4634), .ZN(n4635) );
  INV_X1 U5633 ( .A(n4635), .ZN(n9707) );
  NAND2_X1 U5634 ( .A1(n3502), .A2(n4637), .ZN(n4638) );
  XOR2_X1 U5635 ( .A(n4639), .B(n4638), .Z(n4640) );
  AOI22_X1 U5636 ( .A1(n4640), .A2(n8399), .B1(n6373), .B2(
        \adder_stage1[12][13] ), .ZN(n4641) );
  INV_X1 U5637 ( .A(n4641), .ZN(n9860) );
  AOI22_X1 U5638 ( .A1(\x_mult_f_int[1][14] ), .A2(n7110), .B1(n8202), .B2(
        \x_mult_f[1][14] ), .ZN(n4642) );
  INV_X1 U5639 ( .A(n4642), .ZN(n8936) );
  OAI21_X1 U5640 ( .B1(n4645), .B2(n4644), .A(n4643), .ZN(n5934) );
  OR2_X1 U5641 ( .A1(\adder_stage3[2][16] ), .A2(\adder_stage3[3][16] ), .ZN(
        n5932) );
  NAND2_X1 U5642 ( .A1(\adder_stage3[2][16] ), .A2(\adder_stage3[3][16] ), 
        .ZN(n5931) );
  INV_X1 U5643 ( .A(n5931), .ZN(n4646) );
  AOI21_X1 U5644 ( .B1(n5934), .B2(n5932), .A(n4646), .ZN(n8281) );
  NOR2_X1 U5645 ( .A1(\adder_stage3[2][17] ), .A2(\adder_stage3[3][17] ), .ZN(
        n8278) );
  NAND2_X1 U5646 ( .A1(\adder_stage3[2][17] ), .A2(\adder_stage3[3][17] ), 
        .ZN(n8279) );
  OAI21_X1 U5647 ( .B1(n8281), .B2(n8278), .A(n8279), .ZN(n4648) );
  OR2_X1 U5648 ( .A1(\adder_stage3[2][18] ), .A2(\adder_stage3[3][18] ), .ZN(
        n7931) );
  NAND2_X1 U5649 ( .A1(\adder_stage3[2][18] ), .A2(\adder_stage3[3][18] ), 
        .ZN(n7928) );
  NAND2_X1 U5650 ( .A1(n7931), .A2(n7928), .ZN(n4647) );
  XNOR2_X1 U5651 ( .A(n4648), .B(n4647), .ZN(n4649) );
  AOI22_X1 U5652 ( .A1(n4649), .A2(n5908), .B1(n6373), .B2(
        \adder_stage4[1][18] ), .ZN(n4650) );
  INV_X1 U5653 ( .A(n4650), .ZN(n9549) );
  NOR2_X1 U5654 ( .A1(\adder_stage1[12][1] ), .A2(\adder_stage1[13][1] ), .ZN(
        n5092) );
  INV_X1 U5655 ( .A(n5092), .ZN(n4652) );
  NAND2_X1 U5656 ( .A1(\adder_stage1[12][1] ), .A2(\adder_stage1[13][1] ), 
        .ZN(n5090) );
  NAND2_X1 U5657 ( .A1(n4652), .A2(n5090), .ZN(n4653) );
  NAND2_X1 U5658 ( .A1(\adder_stage1[12][0] ), .A2(\adder_stage1[13][0] ), 
        .ZN(n5091) );
  XOR2_X1 U5659 ( .A(n4653), .B(n5091), .Z(n4654) );
  AOI22_X1 U5660 ( .A1(n5626), .A2(\adder_stage2[6][1] ), .B1(n6523), .B2(
        n4654), .ZN(n4655) );
  INV_X1 U5661 ( .A(n4655), .ZN(n9702) );
  INV_X2 U5662 ( .A(n6588), .ZN(n6337) );
  INV_X1 U5663 ( .A(n4656), .ZN(n4777) );
  OAI21_X1 U5664 ( .B1(n4777), .B2(n4773), .A(n4774), .ZN(n4661) );
  INV_X1 U5665 ( .A(n4657), .ZN(n4659) );
  NAND2_X1 U5666 ( .A1(n4659), .A2(n4658), .ZN(n4660) );
  XNOR2_X1 U5667 ( .A(n4661), .B(n4660), .ZN(n4662) );
  AOI22_X1 U5668 ( .A1(n6337), .A2(\adder_stage2[5][3] ), .B1(n8189), .B2(
        n4662), .ZN(n4663) );
  INV_X1 U5669 ( .A(n4663), .ZN(n9717) );
  OR2_X1 U5670 ( .A1(\adder_stage1[12][0] ), .A2(\adder_stage1[13][0] ), .ZN(
        n4664) );
  AND2_X1 U5671 ( .A1(n4664), .A2(n5091), .ZN(n4665) );
  AOI22_X1 U5672 ( .A1(n5626), .A2(\adder_stage2[6][0] ), .B1(n7992), .B2(
        n4665), .ZN(n4666) );
  INV_X1 U5673 ( .A(n4666), .ZN(n9703) );
  NAND2_X1 U5674 ( .A1(n4668), .A2(n4667), .ZN(n4669) );
  XNOR2_X1 U5675 ( .A(n4670), .B(n4669), .ZN(n4671) );
  AOI22_X1 U5676 ( .A1(n4689), .A2(\adder_stage2[7][12] ), .B1(n8387), .B2(
        n4671), .ZN(n4672) );
  INV_X1 U5677 ( .A(n4672), .ZN(n9674) );
  INV_X1 U5678 ( .A(n4673), .ZN(n4675) );
  NAND2_X1 U5679 ( .A1(n4675), .A2(n4674), .ZN(n4676) );
  XOR2_X1 U5680 ( .A(n4677), .B(n4676), .Z(n4678) );
  AOI22_X1 U5681 ( .A1(n4689), .A2(\adder_stage2[7][13] ), .B1(n8401), .B2(
        n4678), .ZN(n4679) );
  INV_X1 U5682 ( .A(n4679), .ZN(n9673) );
  OAI21_X1 U5683 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4687) );
  INV_X1 U5684 ( .A(n4683), .ZN(n4685) );
  NAND2_X1 U5685 ( .A1(n4685), .A2(n4684), .ZN(n4686) );
  XNOR2_X1 U5686 ( .A(n4687), .B(n4686), .ZN(n4688) );
  AOI22_X1 U5687 ( .A1(n4689), .A2(\adder_stage2[7][10] ), .B1(n7284), .B2(
        n4688), .ZN(n4690) );
  INV_X1 U5688 ( .A(n4690), .ZN(n9676) );
  AOI22_X1 U5689 ( .A1(n5544), .A2(\x_mult_f[29][2] ), .B1(n8213), .B2(
        \x_mult_f_int[29][2] ), .ZN(n4691) );
  INV_X1 U5690 ( .A(n4691), .ZN(n9263) );
  AOI22_X1 U5691 ( .A1(n4713), .A2(\x_mult_f[24][3] ), .B1(n8318), .B2(
        \x_mult_f_int[24][3] ), .ZN(n4692) );
  INV_X1 U5692 ( .A(n4692), .ZN(n9225) );
  AOI22_X1 U5693 ( .A1(n4713), .A2(\x_mult_f[24][4] ), .B1(n7698), .B2(
        \x_mult_f_int[24][4] ), .ZN(n4693) );
  INV_X1 U5694 ( .A(n4693), .ZN(n9224) );
  AOI22_X1 U5695 ( .A1(n4713), .A2(\x_mult_f[24][2] ), .B1(n7284), .B2(
        \x_mult_f_int[24][2] ), .ZN(n4694) );
  INV_X1 U5696 ( .A(n4694), .ZN(n9226) );
  OAI21_X1 U5697 ( .B1(n4697), .B2(n4696), .A(n4695), .ZN(n4702) );
  INV_X1 U5698 ( .A(n4698), .ZN(n4700) );
  NAND2_X1 U5699 ( .A1(n4700), .A2(n4699), .ZN(n4701) );
  XNOR2_X1 U5700 ( .A(n4702), .B(n4701), .ZN(n4703) );
  AOI22_X1 U5701 ( .A1(n4713), .A2(\adder_stage3[2][3] ), .B1(n7992), .B2(
        n4703), .ZN(n4704) );
  INV_X1 U5702 ( .A(n4704), .ZN(n9626) );
  AOI22_X1 U5703 ( .A1(n4713), .A2(\x_mult_f[24][1] ), .B1(n7029), .B2(
        \x_mult_f_int[24][1] ), .ZN(n4705) );
  INV_X1 U5704 ( .A(n4705), .ZN(n9340) );
  INV_X1 U5705 ( .A(n4706), .ZN(n4708) );
  NAND2_X1 U5706 ( .A1(n4708), .A2(n4707), .ZN(n4710) );
  XOR2_X1 U5707 ( .A(n4710), .B(n4709), .Z(n4711) );
  AOI22_X1 U5708 ( .A1(n4713), .A2(\adder_stage3[2][1] ), .B1(n8203), .B2(
        n4711), .ZN(n4712) );
  INV_X1 U5709 ( .A(n4712), .ZN(n9628) );
  AOI22_X1 U5710 ( .A1(n4713), .A2(\x_mult_f[25][4] ), .B1(n8363), .B2(
        \x_mult_f_int[25][4] ), .ZN(n4714) );
  INV_X1 U5711 ( .A(n4714), .ZN(n9227) );
  INV_X2 U5712 ( .A(n4715), .ZN(n5678) );
  OR2_X1 U5713 ( .A1(\x_mult_f[26][0] ), .A2(\x_mult_f[27][0] ), .ZN(n4716) );
  AND2_X1 U5714 ( .A1(n4716), .A2(n5166), .ZN(n4717) );
  AOI22_X1 U5715 ( .A1(n5678), .A2(\adder_stage1[13][0] ), .B1(n4596), .B2(
        n4717), .ZN(n4718) );
  INV_X1 U5716 ( .A(n4718), .ZN(n9856) );
  AOI22_X1 U5717 ( .A1(n8202), .A2(\x_mult_f[31][0] ), .B1(n4596), .B2(
        \x_mult_f_int[31][0] ), .ZN(n4719) );
  INV_X1 U5718 ( .A(n4719), .ZN(n9355) );
  AOI21_X1 U5719 ( .B1(n6009), .B2(n4721), .A(n4720), .ZN(n4725) );
  NAND2_X1 U5720 ( .A1(n4723), .A2(n4722), .ZN(n4724) );
  XOR2_X1 U5721 ( .A(n4725), .B(n4724), .Z(n4726) );
  AOI22_X1 U5722 ( .A1(n5294), .A2(\adder_stage1[15][11] ), .B1(n4596), .B2(
        n4726), .ZN(n4727) );
  INV_X1 U5723 ( .A(n4727), .ZN(n9811) );
  AOI22_X1 U5724 ( .A1(n6330), .A2(\x_mult_f[31][2] ), .B1(n4596), .B2(
        \x_mult_f_int[31][2] ), .ZN(n4728) );
  INV_X1 U5725 ( .A(n4728), .ZN(n9291) );
  INV_X1 U5726 ( .A(n4729), .ZN(n4731) );
  NAND2_X1 U5727 ( .A1(n4731), .A2(n4730), .ZN(n4732) );
  XOR2_X1 U5728 ( .A(n4732), .B(n4735), .Z(n4733) );
  AOI22_X1 U5729 ( .A1(n5273), .A2(\adder_stage1[12][1] ), .B1(n4596), .B2(
        n4733), .ZN(n4734) );
  INV_X1 U5730 ( .A(n4734), .ZN(n9872) );
  OR2_X1 U5731 ( .A1(\x_mult_f[24][0] ), .A2(\x_mult_f[25][0] ), .ZN(n4736) );
  AND2_X1 U5732 ( .A1(n4736), .A2(n4735), .ZN(n4737) );
  AOI22_X1 U5733 ( .A1(n5273), .A2(\adder_stage1[12][0] ), .B1(n4596), .B2(
        n4737), .ZN(n4738) );
  INV_X1 U5734 ( .A(n4738), .ZN(n9873) );
  INV_X1 U5735 ( .A(n4739), .ZN(n4741) );
  NAND2_X1 U5736 ( .A1(n4741), .A2(n4740), .ZN(n4742) );
  XOR2_X1 U5737 ( .A(n4743), .B(n4742), .Z(n4744) );
  AOI22_X1 U5738 ( .A1(n4744), .A2(n8150), .B1(n8048), .B2(
        \adder_stage1[0][13] ), .ZN(n4745) );
  INV_X1 U5739 ( .A(n4745), .ZN(n10057) );
  FA_X1 U5740 ( .A(\x_mult_f[0][14] ), .B(\x_mult_f[1][14] ), .CI(n4746), .CO(
        n8148), .S(n4747) );
  AOI22_X1 U5741 ( .A1(n4747), .A2(n8150), .B1(n8048), .B2(
        \adder_stage1[0][14] ), .ZN(n4748) );
  INV_X1 U5742 ( .A(n4748), .ZN(n10056) );
  AOI22_X1 U5743 ( .A1(n5626), .A2(\x_mult_f[28][2] ), .B1(n6643), .B2(
        \x_mult_f_int[28][2] ), .ZN(n4749) );
  INV_X1 U5744 ( .A(n4749), .ZN(n9252) );
  AOI22_X1 U5745 ( .A1(n5626), .A2(\x_mult_f[28][0] ), .B1(n7909), .B2(
        \x_mult_f_int[28][0] ), .ZN(n4750) );
  INV_X1 U5746 ( .A(n4750), .ZN(n9349) );
  INV_X1 U5747 ( .A(n4751), .ZN(n4802) );
  INV_X1 U5748 ( .A(n4752), .ZN(n4800) );
  INV_X1 U5749 ( .A(n4799), .ZN(n4753) );
  AOI21_X1 U5750 ( .B1(n4802), .B2(n4800), .A(n4753), .ZN(n4758) );
  INV_X1 U5751 ( .A(n4754), .ZN(n4756) );
  NAND2_X1 U5752 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  XOR2_X1 U5753 ( .A(n4758), .B(n4757), .Z(n4759) );
  AOI22_X1 U5754 ( .A1(n6337), .A2(\adder_stage2[5][5] ), .B1(n8390), .B2(
        n4759), .ZN(n4760) );
  INV_X1 U5755 ( .A(n4760), .ZN(n9715) );
  AOI22_X1 U5756 ( .A1(n5626), .A2(\x_mult_f[28][4] ), .B1(n5908), .B2(
        \x_mult_f_int[28][4] ), .ZN(n4761) );
  INV_X1 U5757 ( .A(n4761), .ZN(n9250) );
  AOI22_X1 U5758 ( .A1(n5626), .A2(\x_mult_f[28][1] ), .B1(n4596), .B2(
        \x_mult_f_int[28][1] ), .ZN(n4762) );
  INV_X1 U5759 ( .A(n4762), .ZN(n9348) );
  AOI22_X1 U5760 ( .A1(n5626), .A2(\x_mult_f[28][3] ), .B1(n8114), .B2(
        \x_mult_f_int[28][3] ), .ZN(n4763) );
  INV_X1 U5761 ( .A(n4763), .ZN(n9251) );
  AOI21_X1 U5762 ( .B1(n4802), .B2(n4765), .A(n4764), .ZN(n4818) );
  OAI21_X1 U5763 ( .B1(n4818), .B2(n4814), .A(n4815), .ZN(n4770) );
  INV_X1 U5764 ( .A(n4766), .ZN(n4768) );
  NAND2_X1 U5765 ( .A1(n4768), .A2(n4767), .ZN(n4769) );
  XNOR2_X1 U5766 ( .A(n4770), .B(n4769), .ZN(n4771) );
  AOI22_X1 U5767 ( .A1(n6337), .A2(\adder_stage2[5][7] ), .B1(n7909), .B2(
        n4771), .ZN(n4772) );
  INV_X1 U5768 ( .A(n4772), .ZN(n9713) );
  INV_X1 U5769 ( .A(n4773), .ZN(n4775) );
  NAND2_X1 U5770 ( .A1(n4775), .A2(n4774), .ZN(n4776) );
  XOR2_X1 U5771 ( .A(n4777), .B(n4776), .Z(n4778) );
  AOI22_X1 U5772 ( .A1(n6337), .A2(\adder_stage2[5][2] ), .B1(n6643), .B2(
        n4778), .ZN(n4779) );
  INV_X1 U5773 ( .A(n4779), .ZN(n9718) );
  INV_X1 U5774 ( .A(n4780), .ZN(n4824) );
  OAI21_X1 U5775 ( .B1(n4824), .B2(n4781), .A(n4821), .ZN(n4785) );
  NAND2_X1 U5776 ( .A1(n4783), .A2(n4782), .ZN(n4784) );
  XNOR2_X1 U5777 ( .A(n4785), .B(n4784), .ZN(n4786) );
  AOI22_X1 U5778 ( .A1(n6337), .A2(\adder_stage2[5][9] ), .B1(n8318), .B2(
        n4786), .ZN(n4787) );
  INV_X1 U5779 ( .A(n4787), .ZN(n9711) );
  INV_X1 U5780 ( .A(n4788), .ZN(n8322) );
  INV_X1 U5781 ( .A(n8321), .ZN(n4789) );
  NAND2_X1 U5782 ( .A1(n4789), .A2(n8320), .ZN(n4790) );
  XOR2_X1 U5783 ( .A(n8322), .B(n4790), .Z(n4791) );
  AOI22_X1 U5784 ( .A1(n5626), .A2(\adder_stage4[1][2] ), .B1(n6699), .B2(
        n4791), .ZN(n4792) );
  INV_X1 U5785 ( .A(n4792), .ZN(n9565) );
  NAND2_X1 U5786 ( .A1(n3401), .A2(n4794), .ZN(n4795) );
  XOR2_X1 U5787 ( .A(n4796), .B(n4795), .Z(n4797) );
  AOI22_X1 U5788 ( .A1(n6337), .A2(\adder_stage2[5][11] ), .B1(n7909), .B2(
        n4797), .ZN(n4798) );
  INV_X1 U5789 ( .A(n4798), .ZN(n9709) );
  NAND2_X1 U5790 ( .A1(n4800), .A2(n4799), .ZN(n4801) );
  XNOR2_X1 U5791 ( .A(n4802), .B(n4801), .ZN(n4803) );
  AOI22_X1 U5792 ( .A1(n6337), .A2(\adder_stage2[5][4] ), .B1(n5908), .B2(
        n4803), .ZN(n4804) );
  INV_X1 U5793 ( .A(n4804), .ZN(n9716) );
  OAI21_X1 U5794 ( .B1(n4824), .B2(n4806), .A(n4805), .ZN(n4811) );
  INV_X1 U5795 ( .A(n4807), .ZN(n4809) );
  NAND2_X1 U5796 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  XNOR2_X1 U5797 ( .A(n4811), .B(n4810), .ZN(n4812) );
  AOI22_X1 U5798 ( .A1(n6337), .A2(\adder_stage2[5][10] ), .B1(n7117), .B2(
        n4812), .ZN(n4813) );
  INV_X1 U5799 ( .A(n4813), .ZN(n9710) );
  INV_X1 U5800 ( .A(n4814), .ZN(n4816) );
  NAND2_X1 U5801 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  XOR2_X1 U5802 ( .A(n4818), .B(n4817), .Z(n4819) );
  AOI22_X1 U5803 ( .A1(n6337), .A2(\adder_stage2[5][6] ), .B1(n8114), .B2(
        n4819), .ZN(n4820) );
  INV_X1 U5804 ( .A(n4820), .ZN(n9714) );
  NAND2_X1 U5805 ( .A1(n4822), .A2(n4821), .ZN(n4823) );
  XOR2_X1 U5806 ( .A(n4824), .B(n4823), .Z(n4825) );
  AOI22_X1 U5807 ( .A1(n6337), .A2(\adder_stage2[5][8] ), .B1(n7284), .B2(
        n4825), .ZN(n4826) );
  INV_X1 U5808 ( .A(n4826), .ZN(n9712) );
  NAND2_X1 U5809 ( .A1(n4828), .A2(n4827), .ZN(n4829) );
  XNOR2_X1 U5810 ( .A(n4830), .B(n4829), .ZN(n4831) );
  AOI22_X1 U5811 ( .A1(n6337), .A2(\adder_stage2[5][12] ), .B1(n7029), .B2(
        n4831), .ZN(n4832) );
  INV_X1 U5812 ( .A(n4832), .ZN(n9708) );
  BUF_X2 U5813 ( .A(n6699), .Z(n8208) );
  AOI22_X1 U5814 ( .A1(\x_mult_f_int[15][12] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][12] ), .ZN(n4833) );
  INV_X1 U5815 ( .A(n4833), .ZN(n9116) );
  AOI22_X1 U5816 ( .A1(\x_mult_f_int[15][7] ), .A2(n8189), .B1(n8059), .B2(
        \x_mult_f[15][7] ), .ZN(n4834) );
  INV_X1 U5817 ( .A(n4834), .ZN(n9121) );
  AOI22_X1 U5818 ( .A1(\x_mult_f_int[15][6] ), .A2(n8180), .B1(n8059), .B2(
        \x_mult_f[15][6] ), .ZN(n4835) );
  INV_X1 U5819 ( .A(n4835), .ZN(n9122) );
  AOI22_X1 U5820 ( .A1(n8114), .A2(\x_mult_f_int[15][5] ), .B1(n8059), .B2(
        \x_mult_f[15][5] ), .ZN(n4836) );
  INV_X1 U5821 ( .A(n4836), .ZN(n9123) );
  AOI22_X1 U5822 ( .A1(n8208), .A2(\x_mult_f_int[13][5] ), .B1(n8046), .B2(
        \x_mult_f[13][5] ), .ZN(n4837) );
  INV_X1 U5823 ( .A(n4837), .ZN(n9095) );
  BUF_X2 U5824 ( .A(n6699), .Z(n8189) );
  AOI22_X1 U5825 ( .A1(\x_mult_f_int[13][6] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][6] ), .ZN(n4838) );
  INV_X1 U5826 ( .A(n4838), .ZN(n9094) );
  AOI22_X1 U5827 ( .A1(\x_mult_f_int[13][7] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][7] ), .ZN(n4839) );
  INV_X1 U5828 ( .A(n4839), .ZN(n9093) );
  INV_X2 U5829 ( .A(n6736), .ZN(n4891) );
  AOI22_X1 U5830 ( .A1(n4891), .A2(\x_mult_f[22][2] ), .B1(n8216), .B2(
        \x_mult_f_int[22][2] ), .ZN(n4840) );
  INV_X1 U5831 ( .A(n4840), .ZN(n9204) );
  INV_X1 U5832 ( .A(n4841), .ZN(n4889) );
  OAI21_X1 U5833 ( .B1(n4889), .B2(n4885), .A(n4886), .ZN(n4846) );
  INV_X1 U5834 ( .A(n4842), .ZN(n4844) );
  NAND2_X1 U5835 ( .A1(n4844), .A2(n4843), .ZN(n4845) );
  XNOR2_X1 U5836 ( .A(n4846), .B(n4845), .ZN(n4847) );
  AOI22_X1 U5837 ( .A1(n4891), .A2(\adder_stage1[10][3] ), .B1(n8329), .B2(
        n4847), .ZN(n4848) );
  INV_X1 U5838 ( .A(n4848), .ZN(n9902) );
  AOI22_X1 U5839 ( .A1(n4891), .A2(\x_mult_f[22][3] ), .B1(n8363), .B2(
        \x_mult_f_int[22][3] ), .ZN(n4849) );
  INV_X1 U5840 ( .A(n4849), .ZN(n9203) );
  AOI22_X1 U5841 ( .A1(n4891), .A2(\x_mult_f[22][0] ), .B1(n7992), .B2(
        \x_mult_f_int[22][0] ), .ZN(n4850) );
  INV_X1 U5842 ( .A(n4850), .ZN(n9337) );
  INV_X1 U5843 ( .A(n4851), .ZN(n4871) );
  INV_X1 U5844 ( .A(n4852), .ZN(n4869) );
  INV_X1 U5845 ( .A(n4868), .ZN(n4853) );
  AOI21_X1 U5846 ( .B1(n4871), .B2(n4869), .A(n4853), .ZN(n4858) );
  INV_X1 U5847 ( .A(n4854), .ZN(n4856) );
  NAND2_X1 U5848 ( .A1(n4856), .A2(n4855), .ZN(n4857) );
  XOR2_X1 U5849 ( .A(n4858), .B(n4857), .Z(n4859) );
  AOI22_X1 U5850 ( .A1(n4891), .A2(\adder_stage1[10][5] ), .B1(n8318), .B2(
        n4859), .ZN(n4860) );
  INV_X1 U5851 ( .A(n4860), .ZN(n9900) );
  AOI22_X1 U5852 ( .A1(n4891), .A2(\x_mult_f[22][4] ), .B1(n8180), .B2(
        \x_mult_f_int[22][4] ), .ZN(n4861) );
  INV_X1 U5853 ( .A(n4861), .ZN(n9202) );
  AOI21_X1 U5854 ( .B1(n4871), .B2(n4863), .A(n4862), .ZN(n6376) );
  INV_X1 U5855 ( .A(n6375), .ZN(n4864) );
  NAND2_X1 U5856 ( .A1(n4864), .A2(n6374), .ZN(n4865) );
  XOR2_X1 U5857 ( .A(n6376), .B(n4865), .Z(n4866) );
  AOI22_X1 U5858 ( .A1(n4891), .A2(\adder_stage1[10][6] ), .B1(n8387), .B2(
        n4866), .ZN(n4867) );
  INV_X1 U5859 ( .A(n4867), .ZN(n9899) );
  NAND2_X1 U5860 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  XNOR2_X1 U5861 ( .A(n4871), .B(n4870), .ZN(n4872) );
  AOI22_X1 U5862 ( .A1(n4891), .A2(\adder_stage1[10][4] ), .B1(n8329), .B2(
        n4872), .ZN(n4873) );
  INV_X1 U5863 ( .A(n4873), .ZN(n9901) );
  AOI22_X1 U5864 ( .A1(n4891), .A2(\x_mult_f[22][1] ), .B1(n7774), .B2(
        \x_mult_f_int[22][1] ), .ZN(n4874) );
  INV_X1 U5865 ( .A(n4874), .ZN(n9336) );
  INV_X1 U5866 ( .A(n4875), .ZN(n4877) );
  NAND2_X1 U5867 ( .A1(n4877), .A2(n4876), .ZN(n4878) );
  XOR2_X1 U5868 ( .A(n4878), .B(n4881), .Z(n4879) );
  AOI22_X1 U5869 ( .A1(n4891), .A2(\adder_stage1[10][1] ), .B1(n8329), .B2(
        n4879), .ZN(n4880) );
  INV_X1 U5870 ( .A(n4880), .ZN(n9903) );
  OR2_X1 U5871 ( .A1(\x_mult_f[20][0] ), .A2(\x_mult_f[21][0] ), .ZN(n4882) );
  AND2_X1 U5872 ( .A1(n4882), .A2(n4881), .ZN(n4883) );
  AOI22_X1 U5873 ( .A1(n4891), .A2(\adder_stage1[10][0] ), .B1(n8329), .B2(
        n4883), .ZN(n4884) );
  INV_X1 U5874 ( .A(n4884), .ZN(n9904) );
  INV_X1 U5875 ( .A(n4885), .ZN(n4887) );
  NAND2_X1 U5876 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  XOR2_X1 U5877 ( .A(n4889), .B(n4888), .Z(n4890) );
  AOI22_X1 U5878 ( .A1(n4891), .A2(\adder_stage1[10][2] ), .B1(n8329), .B2(
        n4890), .ZN(n8819) );
  INV_X2 U5879 ( .A(n5410), .ZN(n8094) );
  AOI22_X1 U5880 ( .A1(n5908), .A2(\x_mult_f_int[7][5] ), .B1(n8094), .B2(
        \x_mult_f[7][5] ), .ZN(n4893) );
  INV_X1 U5881 ( .A(n4893), .ZN(n9023) );
  AOI22_X1 U5882 ( .A1(\x_mult_f_int[7][7] ), .A2(n7117), .B1(n8094), .B2(
        \x_mult_f[7][7] ), .ZN(n4894) );
  INV_X1 U5883 ( .A(n4894), .ZN(n9021) );
  OAI21_X1 U5884 ( .B1(n4897), .B2(n4896), .A(n4895), .ZN(n4902) );
  INV_X1 U5885 ( .A(n4898), .ZN(n4900) );
  NAND2_X1 U5886 ( .A1(n4900), .A2(n4899), .ZN(n4901) );
  XNOR2_X1 U5887 ( .A(n4902), .B(n4901), .ZN(n4903) );
  AOI22_X1 U5888 ( .A1(n6330), .A2(\adder_stage2[7][3] ), .B1(n6523), .B2(
        n4903), .ZN(n4904) );
  INV_X1 U5889 ( .A(n4904), .ZN(n9683) );
  NOR2_X1 U5890 ( .A1(n4905), .A2(n4909), .ZN(n4912) );
  NAND2_X1 U5891 ( .A1(n4906), .A2(n4912), .ZN(n4914) );
  OAI21_X1 U5892 ( .B1(n4909), .B2(n4908), .A(n4907), .ZN(n4910) );
  AOI21_X1 U5893 ( .B1(n4912), .B2(n4911), .A(n4910), .ZN(n4913) );
  OAI21_X1 U5894 ( .B1(n4915), .B2(n4914), .A(n4913), .ZN(n4924) );
  INV_X1 U5895 ( .A(n4924), .ZN(n4973) );
  NOR2_X1 U5896 ( .A1(\adder_stage2[4][8] ), .A2(\adder_stage2[5][8] ), .ZN(
        n4972) );
  INV_X1 U5897 ( .A(n4972), .ZN(n4916) );
  NAND2_X1 U5898 ( .A1(\adder_stage2[4][8] ), .A2(\adder_stage2[5][8] ), .ZN(
        n4971) );
  NAND2_X1 U5899 ( .A1(n4916), .A2(n4971), .ZN(n4917) );
  XOR2_X1 U5900 ( .A(n4973), .B(n4917), .Z(n4918) );
  AOI22_X1 U5901 ( .A1(n7767), .A2(\adder_stage3[2][8] ), .B1(n5950), .B2(
        n4918), .ZN(n4919) );
  INV_X1 U5902 ( .A(n4919), .ZN(n9621) );
  NOR2_X1 U5903 ( .A1(\adder_stage2[4][9] ), .A2(\adder_stage2[5][9] ), .ZN(
        n4974) );
  NOR2_X1 U5904 ( .A1(n4972), .A2(n4974), .ZN(n4937) );
  NOR2_X1 U5905 ( .A1(\adder_stage2[4][10] ), .A2(\adder_stage2[5][10] ), .ZN(
        n4941) );
  NOR2_X1 U5906 ( .A1(\adder_stage2[4][11] ), .A2(\adder_stage2[5][11] ), .ZN(
        n4943) );
  NOR2_X1 U5907 ( .A1(n4941), .A2(n4943), .ZN(n4921) );
  NAND2_X1 U5908 ( .A1(n4937), .A2(n4921), .ZN(n4963) );
  NOR2_X1 U5909 ( .A1(\adder_stage2[4][12] ), .A2(\adder_stage2[5][12] ), .ZN(
        n4964) );
  NOR2_X1 U5910 ( .A1(n4963), .A2(n4964), .ZN(n4923) );
  NAND2_X1 U5911 ( .A1(\adder_stage2[4][9] ), .A2(\adder_stage2[5][9] ), .ZN(
        n4975) );
  OAI21_X1 U5912 ( .B1(n4974), .B2(n4971), .A(n4975), .ZN(n4938) );
  NAND2_X1 U5913 ( .A1(\adder_stage2[4][10] ), .A2(\adder_stage2[5][10] ), 
        .ZN(n4950) );
  NAND2_X1 U5914 ( .A1(\adder_stage2[4][11] ), .A2(\adder_stage2[5][11] ), 
        .ZN(n4944) );
  OAI21_X1 U5915 ( .B1(n4943), .B2(n4950), .A(n4944), .ZN(n4920) );
  AOI21_X1 U5916 ( .B1(n4921), .B2(n4938), .A(n4920), .ZN(n4962) );
  NAND2_X1 U5917 ( .A1(\adder_stage2[4][12] ), .A2(\adder_stage2[5][12] ), 
        .ZN(n4965) );
  OAI21_X1 U5918 ( .B1(n4962), .B2(n4964), .A(n4965), .ZN(n4922) );
  AOI21_X1 U5919 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4931) );
  NOR2_X1 U5920 ( .A1(\adder_stage2[4][13] ), .A2(\adder_stage2[5][13] ), .ZN(
        n4930) );
  INV_X1 U5921 ( .A(n4930), .ZN(n4925) );
  NAND2_X1 U5922 ( .A1(\adder_stage2[4][13] ), .A2(\adder_stage2[5][13] ), 
        .ZN(n4929) );
  NAND2_X1 U5923 ( .A1(n4925), .A2(n4929), .ZN(n4926) );
  XOR2_X1 U5924 ( .A(n4931), .B(n4926), .Z(n4927) );
  AOI22_X1 U5925 ( .A1(n7910), .A2(\adder_stage3[2][13] ), .B1(n6256), .B2(
        n4927), .ZN(n4928) );
  INV_X1 U5926 ( .A(n4928), .ZN(n9616) );
  OAI21_X1 U5927 ( .B1(n4931), .B2(n4930), .A(n4929), .ZN(n4959) );
  OR2_X1 U5928 ( .A1(\adder_stage2[4][14] ), .A2(\adder_stage2[5][14] ), .ZN(
        n4957) );
  NAND2_X1 U5929 ( .A1(\adder_stage2[4][14] ), .A2(\adder_stage2[5][14] ), 
        .ZN(n4956) );
  INV_X1 U5930 ( .A(n4956), .ZN(n4932) );
  AOI21_X1 U5931 ( .B1(n4959), .B2(n4957), .A(n4932), .ZN(n4986) );
  NOR2_X1 U5932 ( .A1(\adder_stage2[4][15] ), .A2(\adder_stage2[5][15] ), .ZN(
        n4985) );
  INV_X1 U5933 ( .A(n4985), .ZN(n4933) );
  NAND2_X1 U5934 ( .A1(\adder_stage2[4][15] ), .A2(\adder_stage2[5][15] ), 
        .ZN(n4984) );
  NAND2_X1 U5935 ( .A1(n4933), .A2(n4984), .ZN(n4934) );
  XOR2_X1 U5936 ( .A(n4986), .B(n4934), .Z(n4935) );
  AOI22_X1 U5937 ( .A1(n6581), .A2(\adder_stage3[2][15] ), .B1(n7511), .B2(
        n4935), .ZN(n4936) );
  INV_X1 U5938 ( .A(n4936), .ZN(n9614) );
  INV_X1 U5939 ( .A(n4937), .ZN(n4940) );
  INV_X1 U5940 ( .A(n4938), .ZN(n4939) );
  OAI21_X1 U5941 ( .B1(n4973), .B2(n4940), .A(n4939), .ZN(n4953) );
  INV_X1 U5942 ( .A(n4941), .ZN(n4951) );
  INV_X1 U5943 ( .A(n4950), .ZN(n4942) );
  AOI21_X1 U5944 ( .B1(n4953), .B2(n4951), .A(n4942), .ZN(n4947) );
  INV_X1 U5945 ( .A(n4943), .ZN(n4945) );
  NAND2_X1 U5946 ( .A1(n4945), .A2(n4944), .ZN(n4946) );
  XOR2_X1 U5947 ( .A(n4947), .B(n4946), .Z(n4948) );
  AOI22_X1 U5948 ( .A1(n6428), .A2(\adder_stage3[2][11] ), .B1(n6643), .B2(
        n4948), .ZN(n4949) );
  INV_X1 U5949 ( .A(n4949), .ZN(n9618) );
  NAND2_X1 U5950 ( .A1(n4951), .A2(n4950), .ZN(n4952) );
  XNOR2_X1 U5951 ( .A(n4953), .B(n4952), .ZN(n4954) );
  AOI22_X1 U5952 ( .A1(n5909), .A2(\adder_stage3[2][10] ), .B1(n5908), .B2(
        n4954), .ZN(n4955) );
  INV_X1 U5953 ( .A(n4955), .ZN(n9619) );
  NAND2_X1 U5954 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  XNOR2_X1 U5955 ( .A(n4959), .B(n4958), .ZN(n4960) );
  AOI22_X1 U5956 ( .A1(n8048), .A2(\adder_stage3[2][14] ), .B1(n8365), .B2(
        n4960), .ZN(n4961) );
  INV_X1 U5957 ( .A(n4961), .ZN(n9615) );
  OAI21_X1 U5958 ( .B1(n4973), .B2(n4963), .A(n4962), .ZN(n4968) );
  INV_X1 U5959 ( .A(n4964), .ZN(n4966) );
  NAND2_X1 U5960 ( .A1(n4966), .A2(n4965), .ZN(n4967) );
  XNOR2_X1 U5961 ( .A(n4968), .B(n4967), .ZN(n4969) );
  AOI22_X1 U5962 ( .A1(n8157), .A2(\adder_stage3[2][12] ), .B1(n8114), .B2(
        n4969), .ZN(n4970) );
  INV_X1 U5963 ( .A(n4970), .ZN(n9617) );
  OAI21_X1 U5964 ( .B1(n4973), .B2(n4972), .A(n4971), .ZN(n4978) );
  INV_X1 U5965 ( .A(n4974), .ZN(n4976) );
  NAND2_X1 U5966 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  XNOR2_X1 U5967 ( .A(n4978), .B(n4977), .ZN(n4979) );
  AOI22_X1 U5968 ( .A1(n8088), .A2(\adder_stage3[2][9] ), .B1(n8213), .B2(
        n4979), .ZN(n4980) );
  INV_X1 U5969 ( .A(n4980), .ZN(n9620) );
  AOI22_X1 U5970 ( .A1(\x_mult_f_int[11][7] ), .A2(n8186), .B1(n8157), .B2(
        \x_mult_f[11][7] ), .ZN(n4981) );
  INV_X1 U5971 ( .A(n4981), .ZN(n9066) );
  INV_X2 U5972 ( .A(n5378), .ZN(n8212) );
  AOI22_X1 U5973 ( .A1(\x_mult_f_int[6][10] ), .A2(n8114), .B1(n8212), .B2(
        \x_mult_f[6][10] ), .ZN(n4982) );
  INV_X1 U5974 ( .A(n4982), .ZN(n9004) );
  AOI22_X1 U5975 ( .A1(\x_mult_f_int[6][11] ), .A2(n8387), .B1(n8212), .B2(
        \x_mult_f[6][11] ), .ZN(n4983) );
  INV_X1 U5976 ( .A(n4983), .ZN(n9003) );
  OAI21_X1 U5977 ( .B1(n4986), .B2(n4985), .A(n4984), .ZN(n8169) );
  OR2_X1 U5978 ( .A1(\adder_stage2[4][16] ), .A2(\adder_stage2[5][16] ), .ZN(
        n5384) );
  NAND2_X1 U5979 ( .A1(\adder_stage2[4][16] ), .A2(\adder_stage2[5][16] ), 
        .ZN(n4991) );
  INV_X1 U5980 ( .A(n4991), .ZN(n5388) );
  AOI21_X1 U5981 ( .B1(n8169), .B2(n5384), .A(n5388), .ZN(n4988) );
  OR2_X1 U5982 ( .A1(\adder_stage2[4][17] ), .A2(\adder_stage2[5][17] ), .ZN(
        n5387) );
  NAND2_X1 U5983 ( .A1(\adder_stage2[4][17] ), .A2(\adder_stage2[5][17] ), 
        .ZN(n5385) );
  NAND2_X1 U5984 ( .A1(n5387), .A2(n5385), .ZN(n4987) );
  XOR2_X1 U5985 ( .A(n4988), .B(n4987), .Z(n4989) );
  AOI22_X1 U5986 ( .A1(n4989), .A2(n8265), .B1(n8212), .B2(
        \adder_stage3[2][17] ), .ZN(n4990) );
  INV_X1 U5987 ( .A(n4990), .ZN(n9612) );
  NAND2_X1 U5988 ( .A1(n5384), .A2(n4991), .ZN(n4992) );
  XNOR2_X1 U5989 ( .A(n8169), .B(n4992), .ZN(n4993) );
  AOI22_X1 U5990 ( .A1(n6643), .A2(n4993), .B1(n8212), .B2(
        \adder_stage3[2][16] ), .ZN(n4994) );
  INV_X1 U5991 ( .A(n4994), .ZN(n9613) );
  AOI22_X1 U5992 ( .A1(\x_mult_f_int[3][6] ), .A2(n8265), .B1(n8364), .B2(
        \x_mult_f[3][6] ), .ZN(n4995) );
  INV_X1 U5993 ( .A(n4995), .ZN(n8969) );
  AOI22_X1 U5994 ( .A1(n8401), .A2(\x_mult_f_int[3][5] ), .B1(n8364), .B2(
        \x_mult_f[3][5] ), .ZN(n4996) );
  INV_X1 U5995 ( .A(n4996), .ZN(n8970) );
  NAND2_X1 U5996 ( .A1(n3506), .A2(n4998), .ZN(n4999) );
  XOR2_X1 U5997 ( .A(n5000), .B(n4999), .Z(n5001) );
  AOI22_X1 U5998 ( .A1(n5001), .A2(n5950), .B1(n8364), .B2(
        \adder_stage1[14][13] ), .ZN(n5002) );
  INV_X1 U5999 ( .A(n5002), .ZN(n9826) );
  AOI22_X1 U6000 ( .A1(\x_mult_f_int[23][6] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][6] ), .ZN(n5003) );
  INV_X1 U6001 ( .A(n5003), .ZN(n9211) );
  AOI22_X1 U6002 ( .A1(n7992), .A2(\x_mult_f_int[23][5] ), .B1(n8078), .B2(
        \x_mult_f[23][5] ), .ZN(n5004) );
  INV_X1 U6003 ( .A(n5004), .ZN(n9212) );
  AOI22_X1 U6004 ( .A1(\x_mult_f_int[23][7] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][7] ), .ZN(n5005) );
  INV_X1 U6005 ( .A(n5005), .ZN(n9210) );
  AOI22_X1 U6006 ( .A1(n7851), .A2(\x_mult_f[0][4] ), .B1(n8318), .B2(
        \x_mult_f_int[0][4] ), .ZN(n5006) );
  INV_X1 U6007 ( .A(n5006), .ZN(n8934) );
  NAND2_X1 U6008 ( .A1(n5011), .A2(n5010), .ZN(n5012) );
  XNOR2_X1 U6009 ( .A(n5013), .B(n5012), .ZN(n5014) );
  AOI22_X1 U6010 ( .A1(n8046), .A2(\adder_stage1[13][12] ), .B1(n7454), .B2(
        n5014), .ZN(n5015) );
  INV_X1 U6011 ( .A(n5015), .ZN(n9844) );
  NAND2_X1 U6012 ( .A1(n3649), .A2(n5018), .ZN(n5019) );
  XOR2_X1 U6013 ( .A(n5020), .B(n5019), .Z(n5021) );
  AOI22_X1 U6014 ( .A1(n8330), .A2(\adder_stage1[13][11] ), .B1(n6221), .B2(
        n5021), .ZN(n5022) );
  INV_X1 U6015 ( .A(n5022), .ZN(n9845) );
  AOI21_X1 U6016 ( .B1(n5040), .B2(n5024), .A(n5023), .ZN(n5057) );
  INV_X1 U6017 ( .A(n5056), .ZN(n5025) );
  NAND2_X1 U6018 ( .A1(n5025), .A2(n5055), .ZN(n5026) );
  XOR2_X1 U6019 ( .A(n5057), .B(n5026), .Z(n5027) );
  AOI22_X1 U6020 ( .A1(n6337), .A2(\adder_stage1[13][6] ), .B1(n8194), .B2(
        n5027), .ZN(n5028) );
  INV_X1 U6021 ( .A(n5028), .ZN(n9850) );
  INV_X1 U6022 ( .A(n5029), .ZN(n5125) );
  OAI21_X1 U6023 ( .B1(n5125), .B2(n5121), .A(n5122), .ZN(n5034) );
  INV_X1 U6024 ( .A(n5030), .ZN(n5032) );
  NAND2_X1 U6025 ( .A1(n5032), .A2(n5031), .ZN(n5033) );
  XNOR2_X1 U6026 ( .A(n5034), .B(n5033), .ZN(n5035) );
  AOI22_X1 U6027 ( .A1(n8178), .A2(\adder_stage1[13][3] ), .B1(n6915), .B2(
        n5035), .ZN(n5036) );
  INV_X1 U6028 ( .A(n5036), .ZN(n9853) );
  NAND2_X1 U6029 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  XNOR2_X1 U6030 ( .A(n5040), .B(n5039), .ZN(n5041) );
  AOI22_X1 U6031 ( .A1(n6373), .A2(\adder_stage1[13][4] ), .B1(n7356), .B2(
        n5041), .ZN(n5042) );
  INV_X1 U6032 ( .A(n5042), .ZN(n9852) );
  NAND2_X1 U6033 ( .A1(n5044), .A2(n5043), .ZN(n5045) );
  XNOR2_X1 U6034 ( .A(n5046), .B(n5045), .ZN(n5047) );
  AOI22_X1 U6035 ( .A1(n6330), .A2(\adder_stage1[13][10] ), .B1(n8387), .B2(
        n5047), .ZN(n5048) );
  INV_X1 U6036 ( .A(n5048), .ZN(n9846) );
  NAND2_X1 U6037 ( .A1(n5050), .A2(n5049), .ZN(n5051) );
  XNOR2_X1 U6038 ( .A(n5052), .B(n5051), .ZN(n5053) );
  AOI22_X1 U6039 ( .A1(n4689), .A2(\adder_stage1[13][8] ), .B1(n4596), .B2(
        n5053), .ZN(n5054) );
  INV_X1 U6040 ( .A(n5054), .ZN(n9848) );
  OAI21_X1 U6041 ( .B1(n5057), .B2(n5056), .A(n5055), .ZN(n5062) );
  INV_X1 U6042 ( .A(n5058), .ZN(n5060) );
  NAND2_X1 U6043 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  XNOR2_X1 U6044 ( .A(n5062), .B(n5061), .ZN(n5063) );
  AOI22_X1 U6045 ( .A1(n5678), .A2(\adder_stage1[13][7] ), .B1(n8229), .B2(
        n5063), .ZN(n5064) );
  INV_X1 U6046 ( .A(n5064), .ZN(n9849) );
  INV_X1 U6047 ( .A(n5065), .ZN(n5499) );
  INV_X1 U6048 ( .A(n5066), .ZN(n5086) );
  INV_X1 U6049 ( .A(n5085), .ZN(n5067) );
  AOI21_X1 U6050 ( .B1(n5499), .B2(n5086), .A(n5067), .ZN(n5072) );
  INV_X1 U6051 ( .A(n5068), .ZN(n5070) );
  NAND2_X1 U6052 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  XOR2_X1 U6053 ( .A(n5072), .B(n5071), .Z(n5073) );
  AOI22_X1 U6054 ( .A1(n5294), .A2(\adder_stage1[14][5] ), .B1(n4596), .B2(
        n5073), .ZN(n5074) );
  INV_X1 U6055 ( .A(n5074), .ZN(n9834) );
  OAI21_X1 U6056 ( .B1(n5077), .B2(n5076), .A(n5075), .ZN(n5082) );
  INV_X1 U6057 ( .A(n5078), .ZN(n5080) );
  NAND2_X1 U6058 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  XNOR2_X1 U6059 ( .A(n5082), .B(n5081), .ZN(n5083) );
  AOI22_X1 U6060 ( .A1(n5294), .A2(\adder_stage1[14][3] ), .B1(n4596), .B2(
        n5083), .ZN(n5084) );
  INV_X1 U6061 ( .A(n5084), .ZN(n9836) );
  NAND2_X1 U6062 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  XNOR2_X1 U6063 ( .A(n5499), .B(n5087), .ZN(n5088) );
  AOI22_X1 U6064 ( .A1(n5294), .A2(\adder_stage1[14][4] ), .B1(n4596), .B2(
        n5088), .ZN(n5089) );
  INV_X1 U6065 ( .A(n5089), .ZN(n9835) );
  NOR2_X1 U6066 ( .A1(\adder_stage1[12][2] ), .A2(\adder_stage1[13][2] ), .ZN(
        n5618) );
  NOR2_X1 U6067 ( .A1(n5618), .A2(n5620), .ZN(n5094) );
  OAI21_X1 U6068 ( .B1(n5092), .B2(n5091), .A(n5090), .ZN(n5612) );
  NAND2_X1 U6069 ( .A1(\adder_stage1[13][2] ), .A2(\adder_stage1[12][2] ), 
        .ZN(n5617) );
  NAND2_X1 U6070 ( .A1(\adder_stage1[12][3] ), .A2(\adder_stage1[13][3] ), 
        .ZN(n5621) );
  OAI21_X1 U6071 ( .B1(n5620), .B2(n5617), .A(n5621), .ZN(n5093) );
  AOI21_X1 U6072 ( .B1(n5094), .B2(n5612), .A(n5093), .ZN(n5597) );
  NOR2_X1 U6073 ( .A1(\adder_stage1[12][4] ), .A2(\adder_stage1[13][4] ), .ZN(
        n5598) );
  NOR2_X1 U6074 ( .A1(\adder_stage1[12][5] ), .A2(\adder_stage1[13][5] ), .ZN(
        n5605) );
  NOR2_X1 U6075 ( .A1(n5598), .A2(n5605), .ZN(n5663) );
  NOR2_X1 U6076 ( .A1(\adder_stage1[12][6] ), .A2(\adder_stage1[13][6] ), .ZN(
        n5670) );
  NOR2_X1 U6077 ( .A1(\adder_stage1[12][7] ), .A2(\adder_stage1[13][7] ), .ZN(
        n5672) );
  NOR2_X1 U6078 ( .A1(n5670), .A2(n5672), .ZN(n5096) );
  NAND2_X1 U6079 ( .A1(n5663), .A2(n5096), .ZN(n5098) );
  NAND2_X1 U6080 ( .A1(\adder_stage1[12][4] ), .A2(\adder_stage1[13][4] ), 
        .ZN(n5602) );
  NAND2_X1 U6081 ( .A1(\adder_stage1[12][5] ), .A2(\adder_stage1[13][5] ), 
        .ZN(n5606) );
  OAI21_X1 U6082 ( .B1(n5605), .B2(n5602), .A(n5606), .ZN(n5662) );
  NAND2_X1 U6083 ( .A1(\adder_stage1[12][6] ), .A2(\adder_stage1[13][6] ), 
        .ZN(n5669) );
  NAND2_X1 U6084 ( .A1(\adder_stage1[12][7] ), .A2(\adder_stage1[13][7] ), 
        .ZN(n5673) );
  OAI21_X1 U6085 ( .B1(n5672), .B2(n5669), .A(n5673), .ZN(n5095) );
  AOI21_X1 U6086 ( .B1(n5096), .B2(n5662), .A(n5095), .ZN(n5097) );
  OAI21_X1 U6087 ( .B1(n5597), .B2(n5098), .A(n5097), .ZN(n5140) );
  NOR2_X1 U6088 ( .A1(\adder_stage1[12][8] ), .A2(\adder_stage1[13][8] ), .ZN(
        n5155) );
  INV_X1 U6089 ( .A(n5155), .ZN(n5141) );
  OR2_X1 U6090 ( .A1(\adder_stage1[12][9] ), .A2(\adder_stage1[13][9] ), .ZN(
        n5158) );
  NAND2_X1 U6091 ( .A1(n5141), .A2(n5158), .ZN(n5146) );
  NOR2_X1 U6092 ( .A1(\adder_stage1[12][10] ), .A2(\adder_stage1[13][10] ), 
        .ZN(n5147) );
  NOR2_X1 U6093 ( .A1(n5146), .A2(n5147), .ZN(n5102) );
  NAND2_X1 U6094 ( .A1(\adder_stage1[12][8] ), .A2(\adder_stage1[13][8] ), 
        .ZN(n5154) );
  INV_X1 U6095 ( .A(n5154), .ZN(n5100) );
  NAND2_X1 U6096 ( .A1(\adder_stage1[12][9] ), .A2(\adder_stage1[13][9] ), 
        .ZN(n5157) );
  INV_X1 U6097 ( .A(n5157), .ZN(n5099) );
  AOI21_X1 U6098 ( .B1(n5158), .B2(n5100), .A(n5099), .ZN(n5145) );
  NAND2_X1 U6099 ( .A1(\adder_stage1[12][10] ), .A2(\adder_stage1[13][10] ), 
        .ZN(n5148) );
  OAI21_X1 U6100 ( .B1(n5145), .B2(n5147), .A(n5148), .ZN(n5101) );
  OR2_X1 U6101 ( .A1(\adder_stage1[12][12] ), .A2(\adder_stage1[13][12] ), 
        .ZN(n5135) );
  NOR2_X1 U6102 ( .A1(\adder_stage1[12][11] ), .A2(\adder_stage1[13][11] ), 
        .ZN(n5133) );
  INV_X1 U6103 ( .A(n5133), .ZN(n5128) );
  NAND2_X1 U6104 ( .A1(n5135), .A2(n5128), .ZN(n5110) );
  NAND2_X1 U6105 ( .A1(\adder_stage1[12][11] ), .A2(\adder_stage1[13][11] ), 
        .ZN(n5132) );
  INV_X1 U6106 ( .A(n5132), .ZN(n5104) );
  NAND2_X1 U6107 ( .A1(\adder_stage1[12][12] ), .A2(\adder_stage1[13][12] ), 
        .ZN(n5134) );
  INV_X1 U6108 ( .A(n5134), .ZN(n5103) );
  AOI21_X1 U6109 ( .B1(n5135), .B2(n5104), .A(n5103), .ZN(n5115) );
  OAI21_X1 U6110 ( .B1(n5298), .B2(n5110), .A(n5115), .ZN(n5105) );
  INV_X1 U6111 ( .A(n5105), .ZN(n5107) );
  NOR2_X1 U6112 ( .A1(\adder_stage1[12][13] ), .A2(\adder_stage1[13][13] ), 
        .ZN(n5114) );
  INV_X1 U6113 ( .A(n5114), .ZN(n5111) );
  NAND2_X1 U6114 ( .A1(\adder_stage1[12][13] ), .A2(\adder_stage1[13][13] ), 
        .ZN(n5113) );
  NAND2_X1 U6115 ( .A1(n5111), .A2(n5113), .ZN(n5106) );
  XOR2_X1 U6116 ( .A(n5107), .B(n5106), .Z(n5108) );
  AOI22_X1 U6117 ( .A1(n5678), .A2(\adder_stage2[6][13] ), .B1(n4596), .B2(
        n5108), .ZN(n5109) );
  INV_X1 U6118 ( .A(n5109), .ZN(n9690) );
  INV_X1 U6119 ( .A(n5110), .ZN(n5112) );
  NAND2_X1 U6120 ( .A1(n5112), .A2(n5111), .ZN(n5296) );
  OAI21_X1 U6121 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n5116) );
  INV_X1 U6122 ( .A(n5116), .ZN(n5302) );
  OAI21_X1 U6123 ( .B1(n5298), .B2(n5296), .A(n5302), .ZN(n5118) );
  OR2_X1 U6124 ( .A1(\adder_stage1[12][14] ), .A2(\adder_stage1[13][14] ), 
        .ZN(n5299) );
  NAND2_X1 U6125 ( .A1(\adder_stage1[12][14] ), .A2(\adder_stage1[13][14] ), 
        .ZN(n5300) );
  NAND2_X1 U6126 ( .A1(n5299), .A2(n5300), .ZN(n5117) );
  XNOR2_X1 U6127 ( .A(n5118), .B(n5117), .ZN(n5119) );
  AOI22_X1 U6128 ( .A1(n5678), .A2(\adder_stage2[6][14] ), .B1(n7182), .B2(
        n5119), .ZN(n5120) );
  INV_X1 U6129 ( .A(n5120), .ZN(n9689) );
  INV_X1 U6130 ( .A(n5121), .ZN(n5123) );
  NAND2_X1 U6131 ( .A1(n5123), .A2(n5122), .ZN(n5124) );
  XOR2_X1 U6132 ( .A(n5125), .B(n5124), .Z(n5126) );
  AOI22_X1 U6133 ( .A1(n5678), .A2(\adder_stage1[13][2] ), .B1(n8037), .B2(
        n5126), .ZN(n5127) );
  INV_X1 U6134 ( .A(n5127), .ZN(n9854) );
  NAND2_X1 U6135 ( .A1(n5128), .A2(n5132), .ZN(n5129) );
  XOR2_X1 U6136 ( .A(n5298), .B(n5129), .Z(n5130) );
  AOI22_X1 U6137 ( .A1(n5678), .A2(\adder_stage2[6][11] ), .B1(n4596), .B2(
        n5130), .ZN(n5131) );
  INV_X1 U6138 ( .A(n5131), .ZN(n9692) );
  OAI21_X1 U6139 ( .B1(n5298), .B2(n5133), .A(n5132), .ZN(n5137) );
  NAND2_X1 U6140 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  XNOR2_X1 U6141 ( .A(n5137), .B(n5136), .ZN(n5138) );
  AOI22_X1 U6142 ( .A1(n5678), .A2(\adder_stage2[6][12] ), .B1(n7369), .B2(
        n5138), .ZN(n5139) );
  INV_X1 U6143 ( .A(n5139), .ZN(n9691) );
  INV_X1 U6144 ( .A(n5140), .ZN(n5156) );
  NAND2_X1 U6145 ( .A1(n5141), .A2(n5154), .ZN(n5142) );
  XOR2_X1 U6146 ( .A(n5156), .B(n5142), .Z(n5143) );
  AOI22_X1 U6147 ( .A1(n5678), .A2(\adder_stage2[6][8] ), .B1(n7511), .B2(
        n5143), .ZN(n5144) );
  INV_X1 U6148 ( .A(n5144), .ZN(n9695) );
  OAI21_X1 U6149 ( .B1(n5156), .B2(n5146), .A(n5145), .ZN(n5151) );
  INV_X1 U6150 ( .A(n5147), .ZN(n5149) );
  NAND2_X1 U6151 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  XNOR2_X1 U6152 ( .A(n5151), .B(n5150), .ZN(n5152) );
  AOI22_X1 U6153 ( .A1(n5678), .A2(\adder_stage2[6][10] ), .B1(n6256), .B2(
        n5152), .ZN(n5153) );
  INV_X1 U6154 ( .A(n5153), .ZN(n9693) );
  OAI21_X1 U6155 ( .B1(n5156), .B2(n5155), .A(n5154), .ZN(n5160) );
  NAND2_X1 U6156 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  XNOR2_X1 U6157 ( .A(n5160), .B(n5159), .ZN(n5161) );
  AOI22_X1 U6158 ( .A1(n5678), .A2(\adder_stage2[6][9] ), .B1(n8310), .B2(
        n5161), .ZN(n5162) );
  INV_X1 U6159 ( .A(n5162), .ZN(n9694) );
  INV_X1 U6160 ( .A(n5163), .ZN(n5165) );
  NAND2_X1 U6161 ( .A1(n5165), .A2(n5164), .ZN(n5167) );
  XOR2_X1 U6162 ( .A(n5167), .B(n5166), .Z(n5168) );
  AOI22_X1 U6163 ( .A1(n5678), .A2(\adder_stage1[13][1] ), .B1(n8186), .B2(
        n5168), .ZN(n5169) );
  INV_X1 U6164 ( .A(n5169), .ZN(n9855) );
  AOI22_X1 U6165 ( .A1(\x_mult_f_int[19][7] ), .A2(n7454), .B1(n8392), .B2(
        \x_mult_f[19][7] ), .ZN(n5170) );
  INV_X1 U6166 ( .A(n5170), .ZN(n9176) );
  AOI22_X1 U6167 ( .A1(\x_mult_f_int[8][7] ), .A2(n7992), .B1(n8392), .B2(
        \x_mult_f[8][7] ), .ZN(n5171) );
  INV_X1 U6168 ( .A(n5171), .ZN(n9035) );
  AOI22_X1 U6169 ( .A1(\x_mult_f_int[15][13] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][13] ), .ZN(n5172) );
  INV_X1 U6170 ( .A(n5172), .ZN(n9115) );
  AOI22_X1 U6171 ( .A1(\x_mult_f_int[15][8] ), .A2(n8363), .B1(n8059), .B2(
        \x_mult_f[15][8] ), .ZN(n5173) );
  INV_X1 U6172 ( .A(n5173), .ZN(n9120) );
  AOI22_X1 U6173 ( .A1(\x_mult_f_int[15][10] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][10] ), .ZN(n5174) );
  INV_X1 U6174 ( .A(n5174), .ZN(n9118) );
  AOI22_X1 U6175 ( .A1(\x_mult_f_int[15][11] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][11] ), .ZN(n5175) );
  INV_X1 U6176 ( .A(n5175), .ZN(n9117) );
  AOI22_X1 U6177 ( .A1(\x_mult_f_int[15][9] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][9] ), .ZN(n5176) );
  INV_X1 U6178 ( .A(n5176), .ZN(n9119) );
  OR2_X1 U6179 ( .A1(\x_mult_f[4][10] ), .A2(\x_mult_f[5][10] ), .ZN(n7508) );
  OR2_X1 U6180 ( .A1(\x_mult_f[4][11] ), .A2(\x_mult_f[5][11] ), .ZN(n7472) );
  AND2_X1 U6181 ( .A1(n7508), .A2(n7472), .ZN(n7496) );
  OR2_X1 U6182 ( .A1(\x_mult_f[4][12] ), .A2(\x_mult_f[5][12] ), .ZN(n7500) );
  AND2_X1 U6183 ( .A1(n7496), .A2(n7500), .ZN(n8222) );
  OR2_X1 U6184 ( .A1(\x_mult_f[4][13] ), .A2(\x_mult_f[5][13] ), .ZN(n8225) );
  AND2_X1 U6185 ( .A1(n8222), .A2(n8225), .ZN(n5184) );
  NOR2_X1 U6186 ( .A1(\x_mult_f[4][2] ), .A2(\x_mult_f[5][2] ), .ZN(n7363) );
  NOR2_X1 U6187 ( .A1(\x_mult_f[4][3] ), .A2(\x_mult_f[5][3] ), .ZN(n7321) );
  NOR2_X1 U6188 ( .A1(n7363), .A2(n7321), .ZN(n5178) );
  NOR2_X1 U6189 ( .A1(\x_mult_f[4][1] ), .A2(\x_mult_f[5][1] ), .ZN(n6725) );
  NAND2_X1 U6190 ( .A1(\x_mult_f[4][0] ), .A2(\x_mult_f[5][0] ), .ZN(n7298) );
  NAND2_X1 U6191 ( .A1(\x_mult_f[4][1] ), .A2(\x_mult_f[5][1] ), .ZN(n6726) );
  OAI21_X1 U6192 ( .B1(n6725), .B2(n7298), .A(n6726), .ZN(n7320) );
  NAND2_X1 U6193 ( .A1(\x_mult_f[4][2] ), .A2(\x_mult_f[5][2] ), .ZN(n7364) );
  NAND2_X1 U6194 ( .A1(\x_mult_f[4][3] ), .A2(\x_mult_f[5][3] ), .ZN(n7322) );
  OAI21_X1 U6195 ( .B1(n7321), .B2(n7364), .A(n7322), .ZN(n5177) );
  AOI21_X1 U6196 ( .B1(n5178), .B2(n7320), .A(n5177), .ZN(n7304) );
  NOR2_X1 U6197 ( .A1(\x_mult_f[4][5] ), .A2(\x_mult_f[5][5] ), .ZN(n7307) );
  NOR2_X1 U6198 ( .A1(\x_mult_f[4][4] ), .A2(\x_mult_f[5][4] ), .ZN(n7305) );
  NOR2_X1 U6199 ( .A1(n7307), .A2(n7305), .ZN(n7478) );
  NOR2_X1 U6200 ( .A1(\x_mult_f[4][6] ), .A2(\x_mult_f[5][6] ), .ZN(n7486) );
  NOR2_X1 U6201 ( .A1(\x_mult_f[4][7] ), .A2(\x_mult_f[5][7] ), .ZN(n7488) );
  NOR2_X1 U6202 ( .A1(n7486), .A2(n7488), .ZN(n5180) );
  NAND2_X1 U6203 ( .A1(n7478), .A2(n5180), .ZN(n5182) );
  NAND2_X1 U6204 ( .A1(\x_mult_f[4][4] ), .A2(\x_mult_f[5][4] ), .ZN(n7358) );
  NAND2_X1 U6205 ( .A1(\x_mult_f[4][5] ), .A2(\x_mult_f[5][5] ), .ZN(n7308) );
  OAI21_X1 U6206 ( .B1(n7307), .B2(n7358), .A(n7308), .ZN(n7477) );
  NAND2_X1 U6207 ( .A1(\x_mult_f[4][6] ), .A2(\x_mult_f[5][6] ), .ZN(n7485) );
  NAND2_X1 U6208 ( .A1(\x_mult_f[4][7] ), .A2(\x_mult_f[5][7] ), .ZN(n7489) );
  OAI21_X1 U6209 ( .B1(n7488), .B2(n7485), .A(n7489), .ZN(n5179) );
  AOI21_X1 U6210 ( .B1(n7477), .B2(n5180), .A(n5179), .ZN(n5181) );
  OAI21_X1 U6211 ( .B1(n7304), .B2(n5182), .A(n5181), .ZN(n7459) );
  OR2_X1 U6212 ( .A1(\x_mult_f[4][8] ), .A2(\x_mult_f[5][8] ), .ZN(n7457) );
  NAND2_X1 U6213 ( .A1(\x_mult_f[4][8] ), .A2(\x_mult_f[5][8] ), .ZN(n7456) );
  INV_X1 U6214 ( .A(n7456), .ZN(n5183) );
  AOI21_X1 U6215 ( .B1(n7459), .B2(n7457), .A(n5183), .ZN(n7467) );
  NOR2_X1 U6216 ( .A1(\x_mult_f[4][9] ), .A2(\x_mult_f[5][9] ), .ZN(n7463) );
  NAND2_X1 U6217 ( .A1(\x_mult_f[4][9] ), .A2(\x_mult_f[5][9] ), .ZN(n7464) );
  OAI21_X1 U6218 ( .B1(n7467), .B2(n7463), .A(n7464), .ZN(n8223) );
  NAND2_X1 U6219 ( .A1(n5184), .A2(n8223), .ZN(n5189) );
  NAND2_X1 U6220 ( .A1(\x_mult_f[4][10] ), .A2(\x_mult_f[5][10] ), .ZN(n7507)
         );
  INV_X1 U6221 ( .A(n7507), .ZN(n7470) );
  NAND2_X1 U6222 ( .A1(\x_mult_f[4][11] ), .A2(\x_mult_f[5][11] ), .ZN(n7471)
         );
  INV_X1 U6223 ( .A(n7471), .ZN(n5185) );
  AOI21_X1 U6224 ( .B1(n7470), .B2(n7472), .A(n5185), .ZN(n7497) );
  INV_X1 U6225 ( .A(n7500), .ZN(n5186) );
  NAND2_X1 U6226 ( .A1(\x_mult_f[4][12] ), .A2(\x_mult_f[5][12] ), .ZN(n7499)
         );
  OAI21_X1 U6227 ( .B1(n7497), .B2(n5186), .A(n7499), .ZN(n8221) );
  NAND2_X1 U6228 ( .A1(\x_mult_f[4][13] ), .A2(\x_mult_f[5][13] ), .ZN(n8224)
         );
  INV_X1 U6229 ( .A(n8224), .ZN(n5187) );
  AOI21_X1 U6230 ( .B1(n8221), .B2(n8225), .A(n5187), .ZN(n5188) );
  NAND2_X1 U6231 ( .A1(n5189), .A2(n5188), .ZN(n6082) );
  INV_X1 U6232 ( .A(n5190), .ZN(n5191) );
  INV_X2 U6233 ( .A(n4651), .ZN(n8036) );
  AOI22_X1 U6234 ( .A1(n5191), .A2(n8229), .B1(n8036), .B2(
        \adder_stage1[2][20] ), .ZN(n5192) );
  INV_X1 U6235 ( .A(n5192), .ZN(n10021) );
  INV_X2 U6236 ( .A(n5480), .ZN(n8218) );
  AOI22_X1 U6237 ( .A1(n7774), .A2(\x_mult_f_int[31][5] ), .B1(n8218), .B2(
        \x_mult_f[31][5] ), .ZN(n5193) );
  INV_X1 U6238 ( .A(n5193), .ZN(n9288) );
  AOI22_X1 U6239 ( .A1(n8387), .A2(\x_mult_f_int[5][5] ), .B1(n8036), .B2(
        \x_mult_f[5][5] ), .ZN(n5194) );
  INV_X1 U6240 ( .A(n5194), .ZN(n8995) );
  AOI22_X1 U6241 ( .A1(\x_mult_f_int[5][7] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][7] ), .ZN(n5195) );
  INV_X1 U6242 ( .A(n5195), .ZN(n8993) );
  AOI22_X1 U6243 ( .A1(\x_mult_f_int[5][6] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][6] ), .ZN(n5196) );
  INV_X1 U6244 ( .A(n5196), .ZN(n8994) );
  AOI22_X1 U6245 ( .A1(\x_mult_f_int[31][6] ), .A2(n8401), .B1(n8218), .B2(
        \x_mult_f[31][6] ), .ZN(n5197) );
  INV_X1 U6246 ( .A(n5197), .ZN(n9287) );
  INV_X2 U6247 ( .A(n6368), .ZN(n8202) );
  AOI22_X1 U6248 ( .A1(\x_mult_f_int[31][7] ), .A2(n8180), .B1(n8202), .B2(
        \x_mult_f[31][7] ), .ZN(n5198) );
  INV_X1 U6249 ( .A(n5198), .ZN(n9286) );
  INV_X2 U6250 ( .A(n5628), .ZN(n8157) );
  AOI22_X1 U6251 ( .A1(n5908), .A2(\x_mult_f_int[18][5] ), .B1(n8157), .B2(
        \x_mult_f[18][5] ), .ZN(n5199) );
  INV_X1 U6252 ( .A(n5199), .ZN(n9164) );
  INV_X2 U6253 ( .A(n5410), .ZN(n8381) );
  AOI22_X1 U6254 ( .A1(\x_mult_f_int[20][7] ), .A2(n8365), .B1(n8381), .B2(
        \x_mult_f[20][7] ), .ZN(n5200) );
  INV_X1 U6255 ( .A(n5200), .ZN(n9182) );
  AOI22_X1 U6256 ( .A1(n5273), .A2(\x_mult_f[26][1] ), .B1(n5950), .B2(
        \x_mult_f_int[26][1] ), .ZN(n5201) );
  INV_X1 U6257 ( .A(n5201), .ZN(n9344) );
  NAND2_X1 U6258 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  XNOR2_X1 U6259 ( .A(n5208), .B(n5207), .ZN(n5209) );
  AOI22_X1 U6260 ( .A1(n7944), .A2(\adder_stage1[12][12] ), .B1(n7029), .B2(
        n5209), .ZN(n5210) );
  INV_X1 U6261 ( .A(n5210), .ZN(n9861) );
  INV_X1 U6262 ( .A(n5211), .ZN(n5278) );
  INV_X1 U6263 ( .A(n5212), .ZN(n5276) );
  INV_X1 U6264 ( .A(n5275), .ZN(n5213) );
  AOI21_X1 U6265 ( .B1(n5278), .B2(n5276), .A(n5213), .ZN(n5218) );
  INV_X1 U6266 ( .A(n5214), .ZN(n5216) );
  NAND2_X1 U6267 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  XOR2_X1 U6268 ( .A(n5218), .B(n5217), .Z(n5219) );
  AOI22_X1 U6269 ( .A1(n8048), .A2(\adder_stage1[12][5] ), .B1(n8363), .B2(
        n5219), .ZN(n5220) );
  INV_X1 U6270 ( .A(n5220), .ZN(n9868) );
  AOI22_X1 U6271 ( .A1(n5294), .A2(\x_mult_f[30][3] ), .B1(n5950), .B2(
        \x_mult_f_int[30][3] ), .ZN(n5221) );
  INV_X1 U6272 ( .A(n5221), .ZN(n9276) );
  AOI22_X1 U6273 ( .A1(n5294), .A2(\x_mult_f[30][2] ), .B1(n5950), .B2(
        \x_mult_f_int[30][2] ), .ZN(n5222) );
  INV_X1 U6274 ( .A(n5222), .ZN(n9277) );
  AOI22_X1 U6275 ( .A1(n5294), .A2(\x_mult_f[30][1] ), .B1(n5950), .B2(
        \x_mult_f_int[30][1] ), .ZN(n5223) );
  INV_X1 U6276 ( .A(n5223), .ZN(n9352) );
  AOI22_X1 U6277 ( .A1(n5273), .A2(\x_mult_f[26][2] ), .B1(n8229), .B2(
        \x_mult_f_int[26][2] ), .ZN(n5224) );
  INV_X1 U6278 ( .A(n5224), .ZN(n9233) );
  AOI22_X1 U6279 ( .A1(n5273), .A2(\x_mult_f[26][3] ), .B1(n8390), .B2(
        \x_mult_f_int[26][3] ), .ZN(n5225) );
  INV_X1 U6280 ( .A(n5225), .ZN(n9232) );
  AOI22_X1 U6281 ( .A1(n5273), .A2(\x_mult_f[26][0] ), .B1(n5950), .B2(
        \x_mult_f_int[26][0] ), .ZN(n5226) );
  INV_X1 U6282 ( .A(n5226), .ZN(n9345) );
  AOI22_X1 U6283 ( .A1(n5294), .A2(\x_mult_f[30][4] ), .B1(n7774), .B2(
        \x_mult_f_int[30][4] ), .ZN(n5227) );
  INV_X1 U6284 ( .A(n5227), .ZN(n9275) );
  AOI22_X1 U6285 ( .A1(n5273), .A2(\x_mult_f[26][4] ), .B1(n6643), .B2(
        \x_mult_f_int[26][4] ), .ZN(n5228) );
  INV_X1 U6286 ( .A(n5228), .ZN(n9231) );
  AOI22_X1 U6287 ( .A1(n5294), .A2(\x_mult_f[30][0] ), .B1(n5908), .B2(
        \x_mult_f_int[30][0] ), .ZN(n5229) );
  INV_X1 U6288 ( .A(n5229), .ZN(n9353) );
  AOI21_X1 U6289 ( .B1(n5278), .B2(n5231), .A(n5230), .ZN(n5285) );
  OAI21_X1 U6290 ( .B1(n5285), .B2(n5281), .A(n5282), .ZN(n5236) );
  INV_X1 U6291 ( .A(n5232), .ZN(n5234) );
  NAND2_X1 U6292 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  XNOR2_X1 U6293 ( .A(n5236), .B(n5235), .ZN(n5237) );
  AOI22_X1 U6294 ( .A1(n5544), .A2(\adder_stage1[12][7] ), .B1(n7029), .B2(
        n5237), .ZN(n5238) );
  INV_X1 U6295 ( .A(n5238), .ZN(n9866) );
  NAND2_X1 U6296 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  XNOR2_X1 U6297 ( .A(n5242), .B(n5241), .ZN(n5243) );
  AOI22_X1 U6298 ( .A1(n8330), .A2(\adder_stage1[12][8] ), .B1(n7356), .B2(
        n5243), .ZN(n5244) );
  INV_X1 U6299 ( .A(n5244), .ZN(n9865) );
  NAND2_X1 U6300 ( .A1(n3564), .A2(n5247), .ZN(n5248) );
  XOR2_X1 U6301 ( .A(n5249), .B(n5248), .Z(n5250) );
  AOI22_X1 U6302 ( .A1(n8218), .A2(\adder_stage1[12][11] ), .B1(n7110), .B2(
        n5250), .ZN(n5251) );
  INV_X1 U6303 ( .A(n5251), .ZN(n9862) );
  INV_X1 U6304 ( .A(n5252), .ZN(n5271) );
  OAI21_X1 U6305 ( .B1(n5271), .B2(n5267), .A(n5268), .ZN(n5257) );
  INV_X1 U6306 ( .A(n5253), .ZN(n5255) );
  NAND2_X1 U6307 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  XNOR2_X1 U6308 ( .A(n5257), .B(n5256), .ZN(n5258) );
  AOI22_X1 U6309 ( .A1(n5273), .A2(\adder_stage1[12][3] ), .B1(n7454), .B2(
        n5258), .ZN(n5259) );
  INV_X1 U6310 ( .A(n5259), .ZN(n9870) );
  INV_X1 U6311 ( .A(n5260), .ZN(n5262) );
  NAND2_X1 U6312 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  XOR2_X1 U6313 ( .A(n5264), .B(n5263), .Z(n5265) );
  AOI22_X1 U6314 ( .A1(n4689), .A2(\adder_stage1[12][9] ), .B1(n8389), .B2(
        n5265), .ZN(n5266) );
  INV_X1 U6315 ( .A(n5266), .ZN(n9864) );
  INV_X1 U6316 ( .A(n5267), .ZN(n5269) );
  NAND2_X1 U6317 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  XOR2_X1 U6318 ( .A(n5271), .B(n5270), .Z(n5272) );
  AOI22_X1 U6319 ( .A1(n5273), .A2(\adder_stage1[12][2] ), .B1(n8194), .B2(
        n5272), .ZN(n5274) );
  INV_X1 U6320 ( .A(n5274), .ZN(n9871) );
  NAND2_X1 U6321 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  XNOR2_X1 U6322 ( .A(n5278), .B(n5277), .ZN(n5279) );
  AOI22_X1 U6323 ( .A1(n5678), .A2(\adder_stage1[12][4] ), .B1(n6221), .B2(
        n5279), .ZN(n5280) );
  INV_X1 U6324 ( .A(n5280), .ZN(n9869) );
  INV_X1 U6325 ( .A(n5281), .ZN(n5283) );
  NAND2_X1 U6326 ( .A1(n5283), .A2(n5282), .ZN(n5284) );
  XOR2_X1 U6327 ( .A(n5285), .B(n5284), .Z(n5286) );
  AOI22_X1 U6328 ( .A1(n8391), .A2(\adder_stage1[12][6] ), .B1(n6915), .B2(
        n5286), .ZN(n5287) );
  INV_X1 U6329 ( .A(n5287), .ZN(n9867) );
  NAND2_X1 U6330 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  XNOR2_X1 U6331 ( .A(n5291), .B(n5290), .ZN(n5292) );
  AOI22_X1 U6332 ( .A1(n4891), .A2(\adder_stage1[12][10] ), .B1(n8291), .B2(
        n5292), .ZN(n5293) );
  INV_X1 U6333 ( .A(n5293), .ZN(n9863) );
  AOI22_X1 U6334 ( .A1(n5294), .A2(\x_mult_f[31][4] ), .B1(n7992), .B2(
        \x_mult_f_int[31][4] ), .ZN(n5295) );
  INV_X1 U6335 ( .A(n5295), .ZN(n9289) );
  INV_X1 U6336 ( .A(n5296), .ZN(n5297) );
  AND2_X1 U6337 ( .A1(n5297), .A2(n5299), .ZN(n5305) );
  INV_X1 U6338 ( .A(n5298), .ZN(n5304) );
  INV_X1 U6339 ( .A(n5299), .ZN(n5301) );
  OAI21_X1 U6340 ( .B1(n5302), .B2(n5301), .A(n5300), .ZN(n5303) );
  AOI22_X1 U6341 ( .A1(n5306), .A2(n8194), .B1(n8215), .B2(
        \adder_stage2[6][15] ), .ZN(n5307) );
  INV_X1 U6342 ( .A(n5307), .ZN(n9688) );
  NOR2_X1 U6343 ( .A1(\adder_stage1[0][2] ), .A2(\adder_stage1[1][2] ), .ZN(
        n6479) );
  NOR2_X1 U6344 ( .A1(\adder_stage1[0][3] ), .A2(\adder_stage1[1][3] ), .ZN(
        n6451) );
  NOR2_X1 U6345 ( .A1(n6479), .A2(n6451), .ZN(n5309) );
  NOR2_X1 U6346 ( .A1(\adder_stage1[0][1] ), .A2(\adder_stage1[1][1] ), .ZN(
        n6486) );
  NAND2_X1 U6347 ( .A1(\adder_stage1[0][0] ), .A2(\adder_stage1[1][0] ), .ZN(
        n6489) );
  NAND2_X1 U6348 ( .A1(\adder_stage1[0][1] ), .A2(\adder_stage1[1][1] ), .ZN(
        n6487) );
  OAI21_X1 U6349 ( .B1(n6486), .B2(n6489), .A(n6487), .ZN(n6450) );
  NAND2_X1 U6350 ( .A1(\adder_stage1[0][2] ), .A2(\adder_stage1[1][2] ), .ZN(
        n6480) );
  NAND2_X1 U6351 ( .A1(\adder_stage1[0][3] ), .A2(\adder_stage1[1][3] ), .ZN(
        n6452) );
  OAI21_X1 U6352 ( .B1(n6451), .B2(n6480), .A(n6452), .ZN(n5308) );
  AOI21_X1 U6353 ( .B1(n5309), .B2(n6450), .A(n5308), .ZN(n6436) );
  NOR2_X1 U6354 ( .A1(\adder_stage1[0][4] ), .A2(\adder_stage1[1][4] ), .ZN(
        n6437) );
  NOR2_X1 U6355 ( .A1(\adder_stage1[0][5] ), .A2(\adder_stage1[1][5] ), .ZN(
        n6469) );
  NOR2_X1 U6356 ( .A1(n6437), .A2(n6469), .ZN(n6442) );
  NOR2_X1 U6357 ( .A1(\adder_stage1[0][6] ), .A2(\adder_stage1[1][6] ), .ZN(
        n6458) );
  NOR2_X1 U6358 ( .A1(\adder_stage1[0][7] ), .A2(\adder_stage1[1][7] ), .ZN(
        n6443) );
  NOR2_X1 U6359 ( .A1(n6458), .A2(n6443), .ZN(n5311) );
  NAND2_X1 U6360 ( .A1(n6442), .A2(n5311), .ZN(n5313) );
  NAND2_X1 U6361 ( .A1(\adder_stage1[0][4] ), .A2(\adder_stage1[1][4] ), .ZN(
        n6465) );
  NAND2_X1 U6362 ( .A1(\adder_stage1[0][5] ), .A2(\adder_stage1[1][5] ), .ZN(
        n6470) );
  OAI21_X1 U6363 ( .B1(n6465), .B2(n6469), .A(n6470), .ZN(n6441) );
  NAND2_X1 U6364 ( .A1(\adder_stage1[0][6] ), .A2(\adder_stage1[1][6] ), .ZN(
        n6459) );
  NAND2_X1 U6365 ( .A1(\adder_stage1[0][7] ), .A2(\adder_stage1[1][7] ), .ZN(
        n6444) );
  OAI21_X1 U6366 ( .B1(n6443), .B2(n6459), .A(n6444), .ZN(n5310) );
  AOI21_X1 U6367 ( .B1(n5311), .B2(n6441), .A(n5310), .ZN(n5312) );
  OAI21_X1 U6368 ( .B1(n6436), .B2(n5313), .A(n5312), .ZN(n7006) );
  NOR2_X1 U6369 ( .A1(\adder_stage1[0][8] ), .A2(\adder_stage1[1][8] ), .ZN(
        n7007) );
  INV_X1 U6370 ( .A(n7007), .ZN(n7025) );
  OR2_X1 U6371 ( .A1(\adder_stage1[0][9] ), .A2(\adder_stage1[1][9] ), .ZN(
        n7009) );
  NAND2_X1 U6372 ( .A1(n7025), .A2(n7009), .ZN(n7016) );
  NOR2_X1 U6373 ( .A1(\adder_stage1[0][10] ), .A2(\adder_stage1[1][10] ), .ZN(
        n7017) );
  NOR2_X1 U6374 ( .A1(n7016), .A2(n7017), .ZN(n5317) );
  NAND2_X1 U6375 ( .A1(\adder_stage1[0][8] ), .A2(\adder_stage1[1][8] ), .ZN(
        n7024) );
  INV_X1 U6376 ( .A(n7024), .ZN(n5315) );
  NAND2_X1 U6377 ( .A1(\adder_stage1[0][9] ), .A2(\adder_stage1[1][9] ), .ZN(
        n7008) );
  INV_X1 U6378 ( .A(n7008), .ZN(n5314) );
  AOI21_X1 U6379 ( .B1(n7009), .B2(n5315), .A(n5314), .ZN(n7015) );
  NAND2_X1 U6380 ( .A1(\adder_stage1[0][10] ), .A2(\adder_stage1[1][10] ), 
        .ZN(n7018) );
  OAI21_X1 U6381 ( .B1(n7015), .B2(n7017), .A(n7018), .ZN(n5316) );
  AOI21_X1 U6382 ( .B1(n7006), .B2(n5317), .A(n5316), .ZN(n7229) );
  NOR2_X1 U6383 ( .A1(\adder_stage1[0][11] ), .A2(\adder_stage1[1][11] ), .ZN(
        n7225) );
  NAND2_X1 U6384 ( .A1(\adder_stage1[0][11] ), .A2(\adder_stage1[1][11] ), 
        .ZN(n7226) );
  OAI21_X1 U6385 ( .B1(n7229), .B2(n7225), .A(n7226), .ZN(n7242) );
  OR2_X1 U6386 ( .A1(\adder_stage1[0][12] ), .A2(\adder_stage1[1][12] ), .ZN(
        n7240) );
  NAND2_X1 U6387 ( .A1(\adder_stage1[0][12] ), .A2(\adder_stage1[1][12] ), 
        .ZN(n7239) );
  INV_X1 U6388 ( .A(n7239), .ZN(n5318) );
  AOI21_X1 U6389 ( .B1(n7242), .B2(n7240), .A(n5318), .ZN(n7236) );
  NOR2_X1 U6390 ( .A1(\adder_stage1[0][13] ), .A2(\adder_stage1[1][13] ), .ZN(
        n7232) );
  NAND2_X1 U6391 ( .A1(\adder_stage1[0][13] ), .A2(\adder_stage1[1][13] ), 
        .ZN(n7233) );
  OAI21_X1 U6392 ( .B1(n7236), .B2(n7232), .A(n7233), .ZN(n7190) );
  OR2_X1 U6393 ( .A1(\adder_stage1[0][14] ), .A2(\adder_stage1[1][14] ), .ZN(
        n7188) );
  NAND2_X1 U6394 ( .A1(\adder_stage1[0][14] ), .A2(\adder_stage1[1][14] ), 
        .ZN(n7187) );
  INV_X1 U6395 ( .A(n7187), .ZN(n5319) );
  XOR2_X1 U6396 ( .A(\adder_stage1[1][15] ), .B(\adder_stage1[0][15] ), .Z(
        n5320) );
  AOI22_X1 U6397 ( .A1(n5321), .A2(n8213), .B1(n8215), .B2(
        \adder_stage2[0][15] ), .ZN(n5322) );
  INV_X1 U6398 ( .A(n5322), .ZN(n9790) );
  FA_X1 U6399 ( .A(\x_mult_f[26][14] ), .B(\x_mult_f[27][14] ), .CI(n5323), 
        .CO(n7912), .S(n5324) );
  AOI22_X1 U6400 ( .A1(n5324), .A2(n6221), .B1(n8048), .B2(
        \adder_stage1[13][14] ), .ZN(n5325) );
  INV_X1 U6401 ( .A(n5325), .ZN(n9842) );
  AOI22_X1 U6402 ( .A1(n8189), .A2(\x_mult_f_int[12][5] ), .B1(n8046), .B2(
        \x_mult_f[12][5] ), .ZN(n5326) );
  INV_X1 U6403 ( .A(n5326), .ZN(n9082) );
  AOI22_X1 U6404 ( .A1(\x_mult_f_int[13][10] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][10] ), .ZN(n5327) );
  INV_X1 U6405 ( .A(n5327), .ZN(n9090) );
  AOI22_X1 U6406 ( .A1(\x_mult_f_int[13][9] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][9] ), .ZN(n5328) );
  INV_X1 U6407 ( .A(n5328), .ZN(n9091) );
  AOI22_X1 U6408 ( .A1(\x_mult_f_int[12][6] ), .A2(n8114), .B1(n8046), .B2(
        \x_mult_f[12][6] ), .ZN(n5329) );
  INV_X1 U6409 ( .A(n5329), .ZN(n9081) );
  AOI22_X1 U6410 ( .A1(\x_mult_f_int[13][8] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][8] ), .ZN(n5330) );
  INV_X1 U6411 ( .A(n5330), .ZN(n9092) );
  AOI22_X1 U6412 ( .A1(\x_mult_f_int[13][11] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][11] ), .ZN(n5331) );
  INV_X1 U6413 ( .A(n5331), .ZN(n9089) );
  OR2_X1 U6414 ( .A1(\x_mult_f[12][8] ), .A2(\x_mult_f[13][8] ), .ZN(n6979) );
  OR2_X1 U6415 ( .A1(\x_mult_f[12][9] ), .A2(\x_mult_f[13][9] ), .ZN(n6982) );
  AND2_X1 U6416 ( .A1(n6979), .A2(n6982), .ZN(n6964) );
  OR2_X1 U6417 ( .A1(\x_mult_f[12][10] ), .A2(\x_mult_f[13][10] ), .ZN(n6968)
         );
  AND2_X1 U6418 ( .A1(n6964), .A2(n6968), .ZN(n5341) );
  NOR2_X1 U6419 ( .A1(\x_mult_f[12][2] ), .A2(\x_mult_f[13][2] ), .ZN(n7903)
         );
  NOR2_X1 U6420 ( .A1(\x_mult_f[12][3] ), .A2(\x_mult_f[13][3] ), .ZN(n7865)
         );
  NOR2_X1 U6421 ( .A1(n7903), .A2(n7865), .ZN(n5333) );
  NOR2_X1 U6422 ( .A1(\x_mult_f[12][1] ), .A2(\x_mult_f[13][1] ), .ZN(n7858)
         );
  NAND2_X1 U6423 ( .A1(\x_mult_f[12][0] ), .A2(\x_mult_f[13][0] ), .ZN(n7872)
         );
  NAND2_X1 U6424 ( .A1(\x_mult_f[12][1] ), .A2(\x_mult_f[13][1] ), .ZN(n7859)
         );
  OAI21_X1 U6425 ( .B1(n7858), .B2(n7872), .A(n7859), .ZN(n7864) );
  NAND2_X1 U6426 ( .A1(\x_mult_f[12][2] ), .A2(\x_mult_f[13][2] ), .ZN(n7904)
         );
  NAND2_X1 U6427 ( .A1(\x_mult_f[12][3] ), .A2(\x_mult_f[13][3] ), .ZN(n7866)
         );
  OAI21_X1 U6428 ( .B1(n7865), .B2(n7904), .A(n7866), .ZN(n5332) );
  AOI21_X1 U6429 ( .B1(n5333), .B2(n7864), .A(n5332), .ZN(n7853) );
  NOR2_X1 U6430 ( .A1(\x_mult_f[12][4] ), .A2(\x_mult_f[13][4] ), .ZN(n7854)
         );
  NOR2_X1 U6431 ( .A1(\x_mult_f[12][5] ), .A2(\x_mult_f[13][5] ), .ZN(n7879)
         );
  NOR2_X1 U6432 ( .A1(n7854), .A2(n7879), .ZN(n7887) );
  NOR2_X1 U6433 ( .A1(\x_mult_f[12][6] ), .A2(\x_mult_f[13][6] ), .ZN(n7894)
         );
  NOR2_X1 U6434 ( .A1(\x_mult_f[12][7] ), .A2(\x_mult_f[13][7] ), .ZN(n7896)
         );
  NOR2_X1 U6435 ( .A1(n7894), .A2(n7896), .ZN(n5335) );
  NAND2_X1 U6436 ( .A1(n7887), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U6437 ( .A1(\x_mult_f[12][4] ), .A2(\x_mult_f[13][4] ), .ZN(n7876)
         );
  NAND2_X1 U6438 ( .A1(\x_mult_f[12][5] ), .A2(\x_mult_f[13][5] ), .ZN(n7880)
         );
  OAI21_X1 U6439 ( .B1(n7879), .B2(n7876), .A(n7880), .ZN(n7886) );
  NAND2_X1 U6440 ( .A1(\x_mult_f[12][6] ), .A2(\x_mult_f[13][6] ), .ZN(n7893)
         );
  NAND2_X1 U6441 ( .A1(\x_mult_f[12][7] ), .A2(\x_mult_f[13][7] ), .ZN(n7897)
         );
  OAI21_X1 U6442 ( .B1(n7896), .B2(n7893), .A(n7897), .ZN(n5334) );
  AOI21_X1 U6443 ( .B1(n5335), .B2(n7886), .A(n5334), .ZN(n5336) );
  OAI21_X1 U6444 ( .B1(n7853), .B2(n5337), .A(n5336), .ZN(n6975) );
  NAND2_X1 U6445 ( .A1(\x_mult_f[12][8] ), .A2(\x_mult_f[13][8] ), .ZN(n6973)
         );
  INV_X1 U6446 ( .A(n6973), .ZN(n6978) );
  NAND2_X1 U6447 ( .A1(\x_mult_f[12][9] ), .A2(\x_mult_f[13][9] ), .ZN(n6981)
         );
  INV_X1 U6448 ( .A(n6981), .ZN(n5338) );
  AOI21_X1 U6449 ( .B1(n6978), .B2(n6982), .A(n5338), .ZN(n6965) );
  INV_X1 U6450 ( .A(n6968), .ZN(n5339) );
  NAND2_X1 U6451 ( .A1(\x_mult_f[12][10] ), .A2(\x_mult_f[13][10] ), .ZN(n6967) );
  OAI21_X1 U6452 ( .B1(n6965), .B2(n5339), .A(n6967), .ZN(n5340) );
  AOI21_X1 U6453 ( .B1(n5341), .B2(n6975), .A(n5340), .ZN(n6961) );
  NOR2_X1 U6454 ( .A1(\x_mult_f[12][11] ), .A2(\x_mult_f[13][11] ), .ZN(n6957)
         );
  NAND2_X1 U6455 ( .A1(\x_mult_f[12][11] ), .A2(\x_mult_f[13][11] ), .ZN(n6958) );
  OAI21_X1 U6456 ( .B1(n3427), .B2(n6957), .A(n6958), .ZN(n6990) );
  OR2_X1 U6457 ( .A1(\x_mult_f[12][12] ), .A2(\x_mult_f[13][12] ), .ZN(n6988)
         );
  NAND2_X1 U6458 ( .A1(\x_mult_f[12][12] ), .A2(\x_mult_f[13][12] ), .ZN(n6987) );
  INV_X1 U6459 ( .A(n6987), .ZN(n5342) );
  AOI21_X1 U6460 ( .B1(n6990), .B2(n6988), .A(n5342), .ZN(n5354) );
  NOR2_X1 U6461 ( .A1(\x_mult_f[12][13] ), .A2(\x_mult_f[13][13] ), .ZN(n5353)
         );
  INV_X1 U6462 ( .A(n5353), .ZN(n5343) );
  NAND2_X1 U6463 ( .A1(\x_mult_f[12][13] ), .A2(\x_mult_f[13][13] ), .ZN(n5352) );
  NAND2_X1 U6464 ( .A1(n5343), .A2(n5352), .ZN(n5344) );
  XOR2_X1 U6465 ( .A(n5354), .B(n5344), .Z(n5346) );
  INV_X2 U6466 ( .A(n5345), .ZN(n8155) );
  AOI22_X1 U6467 ( .A1(n5346), .A2(n4002), .B1(n8155), .B2(
        \adder_stage1[6][13] ), .ZN(n5347) );
  INV_X1 U6468 ( .A(n5347), .ZN(n9959) );
  AOI22_X1 U6469 ( .A1(\x_mult_f_int[12][10] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][10] ), .ZN(n5348) );
  INV_X1 U6470 ( .A(n5348), .ZN(n9077) );
  AOI22_X1 U6471 ( .A1(\x_mult_f_int[12][7] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][7] ), .ZN(n5349) );
  INV_X1 U6472 ( .A(n5349), .ZN(n9080) );
  AOI22_X1 U6473 ( .A1(\x_mult_f_int[12][8] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][8] ), .ZN(n5350) );
  INV_X1 U6474 ( .A(n5350), .ZN(n9079) );
  AOI22_X1 U6475 ( .A1(\x_mult_f_int[12][9] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][9] ), .ZN(n5351) );
  INV_X1 U6476 ( .A(n5351), .ZN(n9078) );
  OAI21_X1 U6477 ( .B1(n5354), .B2(n5353), .A(n5352), .ZN(n7974) );
  AOI22_X1 U6478 ( .A1(n5355), .A2(n4002), .B1(n8155), .B2(
        \adder_stage1[6][14] ), .ZN(n5356) );
  INV_X1 U6479 ( .A(n5356), .ZN(n9958) );
  AOI22_X1 U6480 ( .A1(n7992), .A2(\x_mult_f_int[29][5] ), .B1(n7944), .B2(
        \x_mult_f[29][5] ), .ZN(n5357) );
  INV_X1 U6481 ( .A(n5357), .ZN(n9260) );
  AOI22_X1 U6482 ( .A1(\x_mult_f_int[29][7] ), .A2(n7774), .B1(n7944), .B2(
        \x_mult_f[29][7] ), .ZN(n5358) );
  INV_X1 U6483 ( .A(n5358), .ZN(n9258) );
  AOI22_X1 U6484 ( .A1(\x_mult_f_int[29][6] ), .A2(n6643), .B1(n7944), .B2(
        \x_mult_f[29][6] ), .ZN(n5359) );
  INV_X1 U6485 ( .A(n5359), .ZN(n9259) );
  AOI22_X1 U6486 ( .A1(\x_mult_f_int[8][9] ), .A2(n8150), .B1(n7285), .B2(
        \x_mult_f[8][9] ), .ZN(n5360) );
  INV_X1 U6487 ( .A(n5360), .ZN(n9033) );
  AOI22_X1 U6488 ( .A1(\x_mult_f_int[8][11] ), .A2(n8150), .B1(n7030), .B2(
        \x_mult_f[8][11] ), .ZN(n5361) );
  INV_X1 U6489 ( .A(n5361), .ZN(n9031) );
  NOR2_X1 U6490 ( .A1(\adder_stage2[0][4] ), .A2(\adder_stage2[1][4] ), .ZN(
        n6817) );
  NOR2_X1 U6491 ( .A1(\adder_stage2[0][5] ), .A2(\adder_stage2[1][5] ), .ZN(
        n6819) );
  NOR2_X1 U6492 ( .A1(n6817), .A2(n6819), .ZN(n6827) );
  NOR2_X1 U6493 ( .A1(\adder_stage2[0][6] ), .A2(\adder_stage2[1][6] ), .ZN(
        n6852) );
  NOR2_X1 U6494 ( .A1(\adder_stage2[0][7] ), .A2(\adder_stage2[1][7] ), .ZN(
        n6828) );
  NOR2_X1 U6495 ( .A1(n6852), .A2(n6828), .ZN(n5366) );
  NAND2_X1 U6496 ( .A1(n6827), .A2(n5366), .ZN(n6784) );
  NOR2_X1 U6497 ( .A1(\adder_stage2[0][13] ), .A2(\adder_stage2[1][13] ), .ZN(
        n6868) );
  OR2_X1 U6498 ( .A1(n6784), .A2(n6868), .ZN(n5367) );
  NOR2_X1 U6499 ( .A1(\adder_stage2[0][2] ), .A2(\adder_stage2[1][2] ), .ZN(
        n6896) );
  NOR2_X1 U6500 ( .A1(\adder_stage2[0][3] ), .A2(\adder_stage2[1][3] ), .ZN(
        n6887) );
  NOR2_X1 U6501 ( .A1(n6896), .A2(n6887), .ZN(n5362) );
  NOR2_X1 U6502 ( .A1(\adder_stage2[0][1] ), .A2(\adder_stage2[1][1] ), .ZN(
        n6909) );
  NAND2_X1 U6503 ( .A1(\adder_stage2[0][0] ), .A2(\adder_stage2[1][0] ), .ZN(
        n6912) );
  NAND2_X1 U6504 ( .A1(\adder_stage2[0][1] ), .A2(\adder_stage2[1][1] ), .ZN(
        n6910) );
  OAI21_X1 U6505 ( .B1(n6909), .B2(n6912), .A(n6910), .ZN(n6886) );
  AND2_X1 U6506 ( .A1(n5362), .A2(n6886), .ZN(n5364) );
  NAND2_X1 U6507 ( .A1(\adder_stage2[1][2] ), .A2(\adder_stage2[0][2] ), .ZN(
        n6897) );
  NAND2_X1 U6508 ( .A1(\adder_stage2[0][3] ), .A2(\adder_stage2[1][3] ), .ZN(
        n6888) );
  OAI21_X1 U6509 ( .B1(n6887), .B2(n6897), .A(n6888), .ZN(n5363) );
  NOR2_X1 U6510 ( .A1(n5364), .A2(n5363), .ZN(n6816) );
  NAND2_X1 U6511 ( .A1(\adder_stage2[0][4] ), .A2(\adder_stage2[1][4] ), .ZN(
        n6903) );
  NAND2_X1 U6512 ( .A1(\adder_stage2[0][5] ), .A2(\adder_stage2[1][5] ), .ZN(
        n6820) );
  OAI21_X1 U6513 ( .B1(n6819), .B2(n6903), .A(n6820), .ZN(n6826) );
  NAND2_X1 U6514 ( .A1(\adder_stage2[0][6] ), .A2(\adder_stage2[1][6] ), .ZN(
        n6853) );
  NAND2_X1 U6515 ( .A1(\adder_stage2[0][7] ), .A2(\adder_stage2[1][7] ), .ZN(
        n6829) );
  OAI21_X1 U6516 ( .B1(n6828), .B2(n6853), .A(n6829), .ZN(n5365) );
  AOI21_X1 U6517 ( .B1(n6826), .B2(n5366), .A(n5365), .ZN(n6783) );
  OAI22_X1 U6518 ( .A1(n5367), .A2(n6816), .B1(n6868), .B2(n6783), .ZN(n5368)
         );
  NOR2_X1 U6519 ( .A1(\adder_stage2[0][8] ), .A2(\adder_stage2[1][8] ), .ZN(
        n6796) );
  NOR2_X1 U6520 ( .A1(\adder_stage2[0][9] ), .A2(\adder_stage2[1][9] ), .ZN(
        n6797) );
  NOR2_X1 U6521 ( .A1(n6796), .A2(n6797), .ZN(n6804) );
  NOR2_X1 U6522 ( .A1(\adder_stage2[0][10] ), .A2(\adder_stage2[1][10] ), .ZN(
        n6807) );
  NOR2_X1 U6523 ( .A1(\adder_stage2[0][11] ), .A2(\adder_stage2[1][11] ), .ZN(
        n6809) );
  NOR2_X1 U6524 ( .A1(n6807), .A2(n6809), .ZN(n6842) );
  NAND2_X1 U6525 ( .A1(n6804), .A2(n6842), .ZN(n6845) );
  NOR2_X1 U6526 ( .A1(\adder_stage2[0][12] ), .A2(\adder_stage2[1][12] ), .ZN(
        n6847) );
  NOR2_X1 U6527 ( .A1(n6845), .A2(n6847), .ZN(n6862) );
  NAND2_X1 U6528 ( .A1(n5368), .A2(n6862), .ZN(n5373) );
  NAND2_X1 U6529 ( .A1(\adder_stage2[0][10] ), .A2(\adder_stage2[1][10] ), 
        .ZN(n6835) );
  NAND2_X1 U6530 ( .A1(\adder_stage2[0][11] ), .A2(\adder_stage2[1][11] ), 
        .ZN(n6810) );
  OAI21_X1 U6531 ( .B1(n6809), .B2(n6835), .A(n6810), .ZN(n6841) );
  OR2_X1 U6532 ( .A1(n6841), .A2(n6842), .ZN(n6860) );
  NOR2_X1 U6533 ( .A1(n6847), .A2(n6868), .ZN(n5369) );
  AND2_X1 U6534 ( .A1(n6860), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6535 ( .A1(\adder_stage2[0][8] ), .A2(\adder_stage2[1][8] ), .ZN(
        n6795) );
  NAND2_X1 U6536 ( .A1(\adder_stage2[0][9] ), .A2(\adder_stage2[1][9] ), .ZN(
        n6798) );
  OAI21_X1 U6537 ( .B1(n6797), .B2(n6795), .A(n6798), .ZN(n6843) );
  OR2_X1 U6538 ( .A1(n6843), .A2(n6841), .ZN(n6861) );
  NAND2_X1 U6539 ( .A1(\adder_stage2[0][12] ), .A2(\adder_stage2[1][12] ), 
        .ZN(n6864) );
  NAND2_X1 U6540 ( .A1(\adder_stage2[0][13] ), .A2(\adder_stage2[1][13] ), 
        .ZN(n6869) );
  OAI21_X1 U6541 ( .B1(n6868), .B2(n6864), .A(n6869), .ZN(n5370) );
  AOI21_X1 U6542 ( .B1(n5371), .B2(n6861), .A(n5370), .ZN(n5372) );
  NAND2_X1 U6543 ( .A1(n5373), .A2(n5372), .ZN(n6792) );
  OR2_X1 U6544 ( .A1(\adder_stage2[0][14] ), .A2(\adder_stage2[1][14] ), .ZN(
        n6790) );
  NAND2_X1 U6545 ( .A1(\adder_stage2[0][14] ), .A2(\adder_stage2[1][14] ), 
        .ZN(n6789) );
  INV_X1 U6546 ( .A(n6789), .ZN(n5374) );
  AOI21_X1 U6547 ( .B1(n6792), .B2(n6790), .A(n5374), .ZN(n8289) );
  NOR2_X1 U6548 ( .A1(\adder_stage2[0][15] ), .A2(\adder_stage2[1][15] ), .ZN(
        n8285) );
  NAND2_X1 U6549 ( .A1(\adder_stage2[0][15] ), .A2(\adder_stage2[1][15] ), 
        .ZN(n8286) );
  OAI21_X1 U6550 ( .B1(n8289), .B2(n8285), .A(n8286), .ZN(n8374) );
  OR2_X1 U6551 ( .A1(\adder_stage2[0][16] ), .A2(\adder_stage2[1][16] ), .ZN(
        n8232) );
  NAND2_X1 U6552 ( .A1(\adder_stage2[0][16] ), .A2(\adder_stage2[1][16] ), 
        .ZN(n5953) );
  NAND2_X1 U6553 ( .A1(n8232), .A2(n5953), .ZN(n5375) );
  XNOR2_X1 U6554 ( .A(n8374), .B(n5375), .ZN(n5376) );
  AOI22_X1 U6555 ( .A1(n7774), .A2(n5376), .B1(n4713), .B2(
        \adder_stage3[0][16] ), .ZN(n5377) );
  INV_X1 U6556 ( .A(n5377), .ZN(n9653) );
  AOI22_X1 U6557 ( .A1(\x_mult_f_int[6][7] ), .A2(n8398), .B1(n8178), .B2(
        \x_mult_f[6][7] ), .ZN(n5379) );
  INV_X1 U6558 ( .A(n5379), .ZN(n9007) );
  AOI22_X1 U6559 ( .A1(\x_mult_f_int[6][8] ), .A2(n8186), .B1(n8178), .B2(
        \x_mult_f[6][8] ), .ZN(n5380) );
  INV_X1 U6560 ( .A(n5380), .ZN(n9006) );
  AOI22_X1 U6561 ( .A1(n8398), .A2(\x_mult_f_int[6][5] ), .B1(n8178), .B2(
        \x_mult_f[6][5] ), .ZN(n5381) );
  INV_X1 U6562 ( .A(n5381), .ZN(n9009) );
  AOI22_X1 U6563 ( .A1(\x_mult_f_int[6][9] ), .A2(n8265), .B1(n8178), .B2(
        \x_mult_f[6][9] ), .ZN(n5382) );
  INV_X1 U6564 ( .A(n5382), .ZN(n9005) );
  AOI22_X1 U6565 ( .A1(\x_mult_f_int[6][6] ), .A2(n8399), .B1(n8178), .B2(
        \x_mult_f[6][6] ), .ZN(n5383) );
  INV_X1 U6566 ( .A(n5383), .ZN(n9008) );
  AND2_X1 U6567 ( .A1(n5384), .A2(n5387), .ZN(n5395) );
  NAND2_X1 U6568 ( .A1(n8169), .A2(n5395), .ZN(n5389) );
  INV_X1 U6569 ( .A(n5385), .ZN(n5386) );
  AOI21_X1 U6570 ( .B1(n5388), .B2(n5387), .A(n5386), .ZN(n5398) );
  NAND2_X1 U6571 ( .A1(n5389), .A2(n5398), .ZN(n5391) );
  NOR2_X1 U6572 ( .A1(\adder_stage2[4][18] ), .A2(\adder_stage2[5][18] ), .ZN(
        n5397) );
  INV_X1 U6573 ( .A(n5397), .ZN(n5394) );
  NAND2_X1 U6574 ( .A1(\adder_stage2[4][18] ), .A2(\adder_stage2[5][18] ), 
        .ZN(n5396) );
  NAND2_X1 U6575 ( .A1(n5394), .A2(n5396), .ZN(n5390) );
  XNOR2_X1 U6576 ( .A(n5391), .B(n5390), .ZN(n5392) );
  BUF_X2 U6577 ( .A(n6699), .Z(n8180) );
  AOI22_X1 U6578 ( .A1(n5392), .A2(n8180), .B1(n8178), .B2(
        \adder_stage3[2][18] ), .ZN(n5393) );
  INV_X1 U6579 ( .A(n5393), .ZN(n9611) );
  AND2_X1 U6580 ( .A1(n5395), .A2(n5394), .ZN(n8167) );
  OAI21_X1 U6581 ( .B1(n5398), .B2(n5397), .A(n5396), .ZN(n8173) );
  AOI21_X1 U6582 ( .B1(n8169), .B2(n8167), .A(n8173), .ZN(n5400) );
  OR2_X1 U6583 ( .A1(\adder_stage2[4][19] ), .A2(\adder_stage2[5][19] ), .ZN(
        n8172) );
  NAND2_X1 U6584 ( .A1(\adder_stage2[4][19] ), .A2(\adder_stage2[5][19] ), 
        .ZN(n8170) );
  NAND2_X1 U6585 ( .A1(n8172), .A2(n8170), .ZN(n5399) );
  XOR2_X1 U6586 ( .A(n5400), .B(n5399), .Z(n5401) );
  AOI22_X1 U6587 ( .A1(n5401), .A2(n8180), .B1(n8178), .B2(
        \adder_stage3[2][19] ), .ZN(n5402) );
  INV_X1 U6588 ( .A(n5402), .ZN(n9610) );
  AOI22_X1 U6589 ( .A1(\x_mult_f_int[7][9] ), .A2(n7029), .B1(n8094), .B2(
        \x_mult_f[7][9] ), .ZN(n5403) );
  INV_X1 U6590 ( .A(n5403), .ZN(n9019) );
  AOI22_X1 U6591 ( .A1(\x_mult_f_int[7][11] ), .A2(n8208), .B1(n8094), .B2(
        \x_mult_f[7][11] ), .ZN(n5404) );
  INV_X1 U6592 ( .A(n5404), .ZN(n9017) );
  AOI22_X1 U6593 ( .A1(\x_mult_f_int[7][8] ), .A2(n8189), .B1(n8094), .B2(
        \x_mult_f[7][8] ), .ZN(n5405) );
  INV_X1 U6594 ( .A(n5405), .ZN(n9020) );
  AOI22_X1 U6595 ( .A1(\x_mult_f_int[7][10] ), .A2(n8114), .B1(n8094), .B2(
        \x_mult_f[7][10] ), .ZN(n5406) );
  INV_X1 U6596 ( .A(n5406), .ZN(n9018) );
  AOI22_X1 U6597 ( .A1(\x_mult_f_int[7][6] ), .A2(n8229), .B1(n8094), .B2(
        \x_mult_f[7][6] ), .ZN(n5407) );
  INV_X1 U6598 ( .A(n5407), .ZN(n9022) );
  AOI22_X1 U6599 ( .A1(\x_mult_f_int[14][6] ), .A2(n8208), .B1(n8381), .B2(
        \x_mult_f[14][6] ), .ZN(n5408) );
  INV_X1 U6600 ( .A(n5408), .ZN(n9108) );
  AOI22_X1 U6601 ( .A1(\x_mult_f_int[14][7] ), .A2(n8208), .B1(n8386), .B2(
        \x_mult_f[14][7] ), .ZN(n5409) );
  INV_X1 U6602 ( .A(n5409), .ZN(n9107) );
  AOI22_X1 U6603 ( .A1(\x_mult_f_int[22][6] ), .A2(n8208), .B1(n7512), .B2(
        \x_mult_f[22][6] ), .ZN(n8820) );
  AOI22_X1 U6604 ( .A1(n8213), .A2(\x_mult_f_int[14][5] ), .B1(n8386), .B2(
        \x_mult_f[14][5] ), .ZN(n5411) );
  INV_X1 U6605 ( .A(n5411), .ZN(n9109) );
  AOI22_X1 U6606 ( .A1(n8229), .A2(\x_mult_f_int[22][5] ), .B1(n8386), .B2(
        \x_mult_f[22][5] ), .ZN(n5412) );
  INV_X1 U6607 ( .A(n5412), .ZN(n9201) );
  BUF_X2 U6608 ( .A(n6699), .Z(n8399) );
  AOI22_X1 U6609 ( .A1(\x_mult_f_int[14][8] ), .A2(n8399), .B1(n8094), .B2(
        \x_mult_f[14][8] ), .ZN(n5413) );
  INV_X1 U6610 ( .A(n5413), .ZN(n9106) );
  AOI22_X1 U6611 ( .A1(\x_mult_f_int[14][10] ), .A2(n8399), .B1(n8386), .B2(
        \x_mult_f[14][10] ), .ZN(n5414) );
  INV_X1 U6612 ( .A(n5414), .ZN(n9104) );
  AOI22_X1 U6613 ( .A1(\x_mult_f_int[14][9] ), .A2(n8399), .B1(n8381), .B2(
        \x_mult_f[14][9] ), .ZN(n5415) );
  INV_X1 U6614 ( .A(n5415), .ZN(n9105) );
  AOI22_X1 U6615 ( .A1(\x_mult_f_int[14][11] ), .A2(n8399), .B1(n8094), .B2(
        \x_mult_f[14][11] ), .ZN(n5416) );
  INV_X1 U6616 ( .A(n5416), .ZN(n9103) );
  OR2_X1 U6617 ( .A1(\x_mult_f[16][8] ), .A2(\x_mult_f[17][8] ), .ZN(n7770) );
  OR2_X1 U6618 ( .A1(\x_mult_f[16][9] ), .A2(\x_mult_f[17][9] ), .ZN(n7702) );
  AND2_X1 U6619 ( .A1(n7770), .A2(n7702), .ZN(n6515) );
  OR2_X1 U6620 ( .A1(\x_mult_f[16][10] ), .A2(\x_mult_f[17][10] ), .ZN(n6519)
         );
  AND2_X1 U6621 ( .A1(n6515), .A2(n6519), .ZN(n5426) );
  NOR2_X1 U6622 ( .A1(\x_mult_f[16][2] ), .A2(\x_mult_f[17][2] ), .ZN(n7755)
         );
  NOR2_X1 U6623 ( .A1(\x_mult_f[16][3] ), .A2(\x_mult_f[17][3] ), .ZN(n7719)
         );
  NOR2_X1 U6624 ( .A1(n7755), .A2(n7719), .ZN(n5418) );
  NOR2_X1 U6625 ( .A1(\x_mult_f[16][1] ), .A2(\x_mult_f[17][1] ), .ZN(n7748)
         );
  NAND2_X1 U6626 ( .A1(\x_mult_f[16][0] ), .A2(\x_mult_f[17][0] ), .ZN(n7751)
         );
  NAND2_X1 U6627 ( .A1(\x_mult_f[16][1] ), .A2(\x_mult_f[17][1] ), .ZN(n7749)
         );
  OAI21_X1 U6628 ( .B1(n7748), .B2(n7751), .A(n7749), .ZN(n7718) );
  NAND2_X1 U6629 ( .A1(\x_mult_f[17][2] ), .A2(\x_mult_f[16][2] ), .ZN(n7756)
         );
  NAND2_X1 U6630 ( .A1(\x_mult_f[16][3] ), .A2(\x_mult_f[17][3] ), .ZN(n7720)
         );
  OAI21_X1 U6631 ( .B1(n7719), .B2(n7756), .A(n7720), .ZN(n5417) );
  AOI21_X1 U6632 ( .B1(n5418), .B2(n7718), .A(n5417), .ZN(n7708) );
  NOR2_X1 U6633 ( .A1(\x_mult_f[16][4] ), .A2(\x_mult_f[17][4] ), .ZN(n7709)
         );
  NOR2_X1 U6634 ( .A1(\x_mult_f[16][5] ), .A2(\x_mult_f[17][5] ), .ZN(n7711)
         );
  NOR2_X1 U6635 ( .A1(n7709), .A2(n7711), .ZN(n7733) );
  NOR2_X1 U6636 ( .A1(\x_mult_f[16][6] ), .A2(\x_mult_f[17][6] ), .ZN(n7741)
         );
  NOR2_X1 U6637 ( .A1(\x_mult_f[16][7] ), .A2(\x_mult_f[17][7] ), .ZN(n7734)
         );
  NOR2_X1 U6638 ( .A1(n7741), .A2(n7734), .ZN(n5420) );
  NAND2_X1 U6639 ( .A1(n7733), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U6640 ( .A1(\x_mult_f[16][4] ), .A2(\x_mult_f[17][4] ), .ZN(n7762)
         );
  NAND2_X1 U6641 ( .A1(\x_mult_f[16][5] ), .A2(\x_mult_f[17][5] ), .ZN(n7712)
         );
  OAI21_X1 U6642 ( .B1(n7711), .B2(n7762), .A(n7712), .ZN(n7732) );
  NAND2_X1 U6643 ( .A1(\x_mult_f[16][6] ), .A2(\x_mult_f[17][6] ), .ZN(n7742)
         );
  NAND2_X1 U6644 ( .A1(\x_mult_f[16][7] ), .A2(\x_mult_f[17][7] ), .ZN(n7735)
         );
  OAI21_X1 U6645 ( .B1(n7734), .B2(n7742), .A(n7735), .ZN(n5419) );
  AOI21_X1 U6646 ( .B1(n5420), .B2(n7732), .A(n5419), .ZN(n5421) );
  OAI21_X1 U6647 ( .B1(n7708), .B2(n5422), .A(n5421), .ZN(n7772) );
  NAND2_X1 U6648 ( .A1(\x_mult_f[16][8] ), .A2(\x_mult_f[17][8] ), .ZN(n7769)
         );
  INV_X1 U6649 ( .A(n7769), .ZN(n7700) );
  NAND2_X1 U6650 ( .A1(\x_mult_f[16][9] ), .A2(\x_mult_f[17][9] ), .ZN(n7701)
         );
  INV_X1 U6651 ( .A(n7701), .ZN(n5423) );
  AOI21_X1 U6652 ( .B1(n7700), .B2(n7702), .A(n5423), .ZN(n6516) );
  INV_X1 U6653 ( .A(n6519), .ZN(n5424) );
  NAND2_X1 U6654 ( .A1(\x_mult_f[16][10] ), .A2(\x_mult_f[17][10] ), .ZN(n6518) );
  OAI21_X1 U6655 ( .B1(n6516), .B2(n5424), .A(n6518), .ZN(n5425) );
  AOI21_X1 U6656 ( .B1(n5426), .B2(n7772), .A(n5425), .ZN(n6502) );
  NOR2_X1 U6657 ( .A1(\x_mult_f[16][11] ), .A2(\x_mult_f[17][11] ), .ZN(n6498)
         );
  NAND2_X1 U6658 ( .A1(\x_mult_f[16][11] ), .A2(\x_mult_f[17][11] ), .ZN(n6499) );
  OAI21_X1 U6659 ( .B1(n3428), .B2(n6498), .A(n6499), .ZN(n6512) );
  OR2_X1 U6660 ( .A1(\x_mult_f[16][12] ), .A2(\x_mult_f[17][12] ), .ZN(n6510)
         );
  NAND2_X1 U6661 ( .A1(\x_mult_f[16][12] ), .A2(\x_mult_f[17][12] ), .ZN(n6509) );
  INV_X1 U6662 ( .A(n6509), .ZN(n5427) );
  AOI21_X1 U6663 ( .B1(n6512), .B2(n6510), .A(n5427), .ZN(n5434) );
  NOR2_X1 U6664 ( .A1(\x_mult_f[16][13] ), .A2(\x_mult_f[17][13] ), .ZN(n5433)
         );
  INV_X1 U6665 ( .A(n5433), .ZN(n5428) );
  NAND2_X1 U6666 ( .A1(\x_mult_f[16][13] ), .A2(\x_mult_f[17][13] ), .ZN(n5432) );
  NAND2_X1 U6667 ( .A1(n5428), .A2(n5432), .ZN(n5429) );
  XOR2_X1 U6668 ( .A(n5434), .B(n5429), .Z(n5430) );
  AOI22_X1 U6669 ( .A1(n5430), .A2(n8387), .B1(n8383), .B2(
        \adder_stage1[8][13] ), .ZN(n5431) );
  INV_X1 U6670 ( .A(n5431), .ZN(n9925) );
  OAI21_X1 U6671 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n7961) );
  AOI22_X1 U6672 ( .A1(n5435), .A2(n8114), .B1(n8386), .B2(
        \adder_stage1[8][14] ), .ZN(n5436) );
  INV_X1 U6673 ( .A(n5436), .ZN(n9924) );
  AOI22_X1 U6674 ( .A1(\x_mult_f_int[17][8] ), .A2(n4596), .B1(n8386), .B2(
        \x_mult_f[17][8] ), .ZN(n5437) );
  INV_X1 U6675 ( .A(n5437), .ZN(n9147) );
  AOI22_X1 U6676 ( .A1(\x_mult_f_int[17][9] ), .A2(n8203), .B1(n8386), .B2(
        \x_mult_f[17][9] ), .ZN(n5438) );
  INV_X1 U6677 ( .A(n5438), .ZN(n9146) );
  FA_X1 U6678 ( .A(\x_mult_f[24][14] ), .B(\x_mult_f[25][14] ), .CI(n5439), 
        .CO(n8144), .S(n5440) );
  AOI22_X1 U6679 ( .A1(n5440), .A2(n7284), .B1(n7944), .B2(
        \adder_stage1[12][14] ), .ZN(n5441) );
  INV_X1 U6680 ( .A(n5441), .ZN(n9859) );
  INV_X1 U6681 ( .A(n5442), .ZN(n5444) );
  NAND2_X1 U6682 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  XOR2_X1 U6683 ( .A(n5446), .B(n5445), .Z(n5448) );
  INV_X2 U6684 ( .A(n5480), .ZN(n8391) );
  AOI22_X1 U6685 ( .A1(n5448), .A2(n8365), .B1(n8391), .B2(
        \adder_stage3[3][17] ), .ZN(n5449) );
  INV_X1 U6686 ( .A(n5449), .ZN(n9592) );
  BUF_X2 U6687 ( .A(n8282), .Z(n8213) );
  AOI22_X1 U6688 ( .A1(\x_mult_f_int[24][10] ), .A2(n8213), .B1(n8391), .B2(
        \x_mult_f[24][10] ), .ZN(n5450) );
  INV_X1 U6689 ( .A(n5450), .ZN(n9220) );
  AOI22_X1 U6690 ( .A1(\x_mult_f_int[24][8] ), .A2(n8213), .B1(n8391), .B2(
        \x_mult_f[24][8] ), .ZN(n5451) );
  INV_X1 U6691 ( .A(n5451), .ZN(n9222) );
  AOI22_X1 U6692 ( .A1(\x_mult_f_int[24][9] ), .A2(n8213), .B1(n8391), .B2(
        \x_mult_f[24][9] ), .ZN(n5452) );
  INV_X1 U6693 ( .A(n5452), .ZN(n9221) );
  AOI22_X1 U6694 ( .A1(\x_mult_f_int[27][9] ), .A2(n8189), .B1(n8391), .B2(
        \x_mult_f[27][9] ), .ZN(n5453) );
  INV_X1 U6695 ( .A(n5453), .ZN(n9240) );
  AOI22_X1 U6696 ( .A1(\x_mult_f_int[0][10] ), .A2(n8189), .B1(n8391), .B2(
        \x_mult_f[0][10] ), .ZN(n5454) );
  INV_X1 U6697 ( .A(n5454), .ZN(n8930) );
  NOR2_X1 U6698 ( .A1(n5455), .A2(n8696), .ZN(n8346) );
  NAND2_X1 U6699 ( .A1(n8346), .A2(n8718), .ZN(n5456) );
  NAND2_X1 U6700 ( .A1(n5457), .A2(n5456), .ZN(n5459) );
  NOR2_X1 U6701 ( .A1(n5459), .A2(n5458), .ZN(n6430) );
  NOR2_X1 U6702 ( .A1(n6430), .A2(reset), .ZN(n6432) );
  NAND2_X1 U6703 ( .A1(n6432), .A2(n5460), .ZN(n6433) );
  INV_X1 U6704 ( .A(n5461), .ZN(n8691) );
  MUX2_X1 U6705 ( .A(n8691), .B(n8714), .S(n6430), .Z(n5462) );
  NAND2_X1 U6706 ( .A1(n6433), .A2(n5462), .ZN(n3387) );
  NAND2_X1 U6707 ( .A1(n3505), .A2(n5464), .ZN(n5465) );
  XOR2_X1 U6708 ( .A(n5466), .B(n5465), .Z(n5467) );
  AOI22_X1 U6709 ( .A1(n5467), .A2(n8363), .B1(n8395), .B2(
        \adder_stage1[10][13] ), .ZN(n8818) );
  INV_X1 U6710 ( .A(n5468), .ZN(n5469) );
  XOR2_X1 U6711 ( .A(\adder_stage1[11][15] ), .B(\adder_stage1[10][15] ), .Z(
        n5472) );
  AOI22_X1 U6712 ( .A1(n5473), .A2(n8216), .B1(n8094), .B2(
        \adder_stage2[5][15] ), .ZN(n5474) );
  INV_X1 U6713 ( .A(n5474), .ZN(n9705) );
  AOI22_X1 U6714 ( .A1(\x_mult_f_int[22][11] ), .A2(n8365), .B1(n8386), .B2(
        \x_mult_f[22][11] ), .ZN(n5475) );
  INV_X1 U6715 ( .A(n5475), .ZN(n9196) );
  AOI22_X1 U6716 ( .A1(\x_mult_f_int[22][9] ), .A2(n8390), .B1(n8381), .B2(
        \x_mult_f[22][9] ), .ZN(n5476) );
  INV_X1 U6717 ( .A(n5476), .ZN(n9198) );
  AOI22_X1 U6718 ( .A1(\x_mult_f_int[22][7] ), .A2(n8186), .B1(n8386), .B2(
        \x_mult_f[22][7] ), .ZN(n5477) );
  INV_X1 U6719 ( .A(n5477), .ZN(n9200) );
  AOI22_X1 U6720 ( .A1(\x_mult_f_int[22][8] ), .A2(n8037), .B1(n8094), .B2(
        \x_mult_f[22][8] ), .ZN(n5478) );
  INV_X1 U6721 ( .A(n5478), .ZN(n9199) );
  AOI22_X1 U6722 ( .A1(\x_mult_f_int[22][10] ), .A2(n8216), .B1(n8381), .B2(
        \x_mult_f[22][10] ), .ZN(n5479) );
  INV_X1 U6723 ( .A(n5479), .ZN(n9197) );
  INV_X2 U6724 ( .A(n5480), .ZN(n8228) );
  AOI22_X1 U6725 ( .A1(\x_mult_f_int[27][11] ), .A2(n4002), .B1(n8228), .B2(
        \x_mult_f[27][11] ), .ZN(n5481) );
  INV_X1 U6726 ( .A(n5481), .ZN(n9238) );
  AOI22_X1 U6727 ( .A1(\x_mult_f_int[0][11] ), .A2(n6523), .B1(n8228), .B2(
        \x_mult_f[0][11] ), .ZN(n5482) );
  INV_X1 U6728 ( .A(n5482), .ZN(n8929) );
  AOI22_X1 U6729 ( .A1(\x_mult_f_int[24][11] ), .A2(n8213), .B1(n8228), .B2(
        \x_mult_f[24][11] ), .ZN(n5483) );
  INV_X1 U6730 ( .A(n5483), .ZN(n9219) );
  AOI22_X1 U6731 ( .A1(\x_mult_f_int[27][10] ), .A2(n8189), .B1(n8228), .B2(
        \x_mult_f[27][10] ), .ZN(n5484) );
  INV_X1 U6732 ( .A(n5484), .ZN(n9239) );
  AOI22_X1 U6733 ( .A1(\x_mult_f_int[26][7] ), .A2(n4002), .B1(n8228), .B2(
        \x_mult_f[26][7] ), .ZN(n5485) );
  INV_X1 U6734 ( .A(n5485), .ZN(n9230) );
  AOI22_X1 U6735 ( .A1(\x_mult_f_int[24][6] ), .A2(n8213), .B1(n8228), .B2(
        \x_mult_f[24][6] ), .ZN(n5486) );
  INV_X1 U6736 ( .A(n5486), .ZN(n9223) );
  AOI22_X1 U6737 ( .A1(\x_mult_f_int[0][7] ), .A2(n7698), .B1(n8228), .B2(
        \x_mult_f[0][7] ), .ZN(n5487) );
  INV_X1 U6738 ( .A(n5487), .ZN(n8932) );
  AOI22_X1 U6739 ( .A1(\x_mult_f_int[0][6] ), .A2(n8180), .B1(n8228), .B2(
        \x_mult_f[0][6] ), .ZN(n5488) );
  INV_X1 U6740 ( .A(n5488), .ZN(n8933) );
  AOI22_X1 U6741 ( .A1(\x_mult_f_int[0][9] ), .A2(n6256), .B1(n8228), .B2(
        \x_mult_f[0][9] ), .ZN(n5489) );
  INV_X1 U6742 ( .A(n5489), .ZN(n8931) );
  AOI22_X1 U6743 ( .A1(\x_mult_f_int[1][7] ), .A2(n8208), .B1(n8228), .B2(
        \x_mult_f[1][7] ), .ZN(n5490) );
  INV_X1 U6744 ( .A(n5490), .ZN(n8942) );
  AOI22_X1 U6745 ( .A1(\x_mult_f_int[0][12] ), .A2(n8399), .B1(n8228), .B2(
        \x_mult_f[0][12] ), .ZN(n5491) );
  INV_X1 U6746 ( .A(n5491), .ZN(n8928) );
  AOI22_X1 U6747 ( .A1(\x_mult_f_int[1][6] ), .A2(n5908), .B1(n8228), .B2(
        \x_mult_f[1][6] ), .ZN(n5492) );
  INV_X1 U6748 ( .A(n5492), .ZN(n8943) );
  NAND2_X1 U6749 ( .A1(n5505), .A2(n5493), .ZN(n5494) );
  XNOR2_X1 U6750 ( .A(n5536), .B(n5494), .ZN(n5495) );
  AOI22_X1 U6751 ( .A1(n5544), .A2(\adder_stage1[14][10] ), .B1(n4002), .B2(
        n5495), .ZN(n5496) );
  INV_X1 U6752 ( .A(n5496), .ZN(n9829) );
  AOI21_X1 U6753 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5521) );
  INV_X1 U6754 ( .A(n5520), .ZN(n5500) );
  NAND2_X1 U6755 ( .A1(n5500), .A2(n5519), .ZN(n5501) );
  XOR2_X1 U6756 ( .A(n5521), .B(n5501), .Z(n5502) );
  AOI22_X1 U6757 ( .A1(n5544), .A2(\adder_stage1[14][6] ), .B1(n8329), .B2(
        n5502), .ZN(n5503) );
  INV_X1 U6758 ( .A(n5503), .ZN(n9833) );
  NAND2_X1 U6759 ( .A1(n3547), .A2(n5507), .ZN(n5508) );
  XOR2_X1 U6760 ( .A(n5509), .B(n5508), .Z(n5510) );
  AOI22_X1 U6761 ( .A1(n5544), .A2(\adder_stage1[14][11] ), .B1(n7909), .B2(
        n5510), .ZN(n5511) );
  INV_X1 U6762 ( .A(n5511), .ZN(n9828) );
  INV_X1 U6763 ( .A(n5512), .ZN(n5514) );
  NAND2_X1 U6764 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  XOR2_X1 U6765 ( .A(n5516), .B(n5515), .Z(n5517) );
  AOI22_X1 U6766 ( .A1(n5544), .A2(\adder_stage1[14][9] ), .B1(n8186), .B2(
        n5517), .ZN(n5518) );
  INV_X1 U6767 ( .A(n5518), .ZN(n9830) );
  OAI21_X1 U6768 ( .B1(n5521), .B2(n5520), .A(n5519), .ZN(n5526) );
  INV_X1 U6769 ( .A(n5522), .ZN(n5524) );
  NAND2_X1 U6770 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  XNOR2_X1 U6771 ( .A(n5526), .B(n5525), .ZN(n5527) );
  AOI22_X1 U6772 ( .A1(n5544), .A2(\adder_stage1[14][7] ), .B1(n5950), .B2(
        n5527), .ZN(n5528) );
  INV_X1 U6773 ( .A(n5528), .ZN(n9832) );
  NAND2_X1 U6774 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  XNOR2_X1 U6775 ( .A(n5532), .B(n5531), .ZN(n5533) );
  AOI22_X1 U6776 ( .A1(n5544), .A2(\adder_stage1[14][8] ), .B1(n8390), .B2(
        n5533), .ZN(n5534) );
  INV_X1 U6777 ( .A(n5534), .ZN(n9831) );
  NAND2_X1 U6778 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  XNOR2_X1 U6779 ( .A(n5542), .B(n5541), .ZN(n5543) );
  AOI22_X1 U6780 ( .A1(n5544), .A2(\adder_stage1[14][12] ), .B1(n7774), .B2(
        n5543), .ZN(n5545) );
  INV_X1 U6781 ( .A(n5545), .ZN(n9827) );
  NOR2_X1 U6782 ( .A1(\adder_stage2[2][2] ), .A2(\adder_stage2[3][2] ), .ZN(
        n6416) );
  NOR2_X1 U6783 ( .A1(\adder_stage2[2][3] ), .A2(\adder_stage2[3][3] ), .ZN(
        n6057) );
  NOR2_X1 U6784 ( .A1(n6416), .A2(n6057), .ZN(n5547) );
  NOR2_X1 U6785 ( .A1(\adder_stage2[2][1] ), .A2(\adder_stage2[3][1] ), .ZN(
        n6049) );
  NAND2_X1 U6786 ( .A1(\adder_stage2[2][0] ), .A2(\adder_stage2[3][0] ), .ZN(
        n6052) );
  NAND2_X1 U6787 ( .A1(\adder_stage2[2][1] ), .A2(\adder_stage2[3][1] ), .ZN(
        n6050) );
  OAI21_X1 U6788 ( .B1(n6049), .B2(n6052), .A(n6050), .ZN(n6056) );
  NAND2_X1 U6789 ( .A1(\adder_stage2[2][2] ), .A2(\adder_stage2[3][2] ), .ZN(
        n6417) );
  NAND2_X1 U6790 ( .A1(\adder_stage2[2][3] ), .A2(\adder_stage2[3][3] ), .ZN(
        n6058) );
  OAI21_X1 U6791 ( .B1(n6057), .B2(n6417), .A(n6058), .ZN(n5546) );
  AOI21_X1 U6792 ( .B1(n5547), .B2(n6056), .A(n5546), .ZN(n6384) );
  NOR2_X1 U6793 ( .A1(\adder_stage2[2][4] ), .A2(\adder_stage2[3][4] ), .ZN(
        n6385) );
  NOR2_X1 U6794 ( .A1(\adder_stage2[2][5] ), .A2(\adder_stage2[3][5] ), .ZN(
        n6387) );
  NOR2_X1 U6795 ( .A1(n6385), .A2(n6387), .ZN(n6395) );
  NOR2_X1 U6796 ( .A1(\adder_stage2[2][7] ), .A2(\adder_stage2[3][7] ), .ZN(
        n6396) );
  NOR2_X1 U6797 ( .A1(\adder_stage2[2][6] ), .A2(\adder_stage2[3][6] ), .ZN(
        n6409) );
  NOR2_X1 U6798 ( .A1(n6396), .A2(n6409), .ZN(n5549) );
  NAND2_X1 U6799 ( .A1(n6395), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U6800 ( .A1(\adder_stage2[2][4] ), .A2(\adder_stage2[3][4] ), .ZN(
        n6403) );
  NAND2_X1 U6801 ( .A1(\adder_stage2[2][5] ), .A2(\adder_stage2[3][5] ), .ZN(
        n6388) );
  OAI21_X1 U6802 ( .B1(n6387), .B2(n6403), .A(n6388), .ZN(n6394) );
  NAND2_X1 U6803 ( .A1(\adder_stage2[2][6] ), .A2(\adder_stage2[3][6] ), .ZN(
        n6410) );
  NAND2_X1 U6804 ( .A1(\adder_stage2[2][7] ), .A2(\adder_stage2[3][7] ), .ZN(
        n6397) );
  OAI21_X1 U6805 ( .B1(n6396), .B2(n6410), .A(n6397), .ZN(n5548) );
  AOI21_X1 U6806 ( .B1(n5549), .B2(n6394), .A(n5548), .ZN(n5550) );
  OAI21_X1 U6807 ( .B1(n6384), .B2(n5551), .A(n5550), .ZN(n5821) );
  NOR2_X1 U6808 ( .A1(\adder_stage2[2][8] ), .A2(\adder_stage2[3][8] ), .ZN(
        n6042) );
  NOR2_X1 U6809 ( .A1(\adder_stage2[2][9] ), .A2(\adder_stage2[3][9] ), .ZN(
        n6035) );
  NOR2_X1 U6810 ( .A1(n6042), .A2(n6035), .ZN(n6022) );
  NOR2_X1 U6811 ( .A1(\adder_stage2[2][10] ), .A2(\adder_stage2[3][10] ), .ZN(
        n6026) );
  NOR2_X1 U6812 ( .A1(\adder_stage2[2][11] ), .A2(\adder_stage2[3][11] ), .ZN(
        n6028) );
  NOR2_X1 U6813 ( .A1(n6026), .A2(n6028), .ZN(n5553) );
  NAND2_X1 U6814 ( .A1(n6022), .A2(n5553), .ZN(n5823) );
  NOR2_X1 U6815 ( .A1(\adder_stage2[2][12] ), .A2(\adder_stage2[3][12] ), .ZN(
        n5824) );
  NOR2_X1 U6816 ( .A1(n5823), .A2(n5824), .ZN(n5555) );
  NAND2_X1 U6817 ( .A1(\adder_stage2[2][8] ), .A2(\adder_stage2[3][8] ), .ZN(
        n6043) );
  NAND2_X1 U6818 ( .A1(\adder_stage2[2][9] ), .A2(\adder_stage2[3][9] ), .ZN(
        n6036) );
  OAI21_X1 U6819 ( .B1(n6035), .B2(n6043), .A(n6036), .ZN(n6023) );
  NAND2_X1 U6820 ( .A1(\adder_stage2[2][10] ), .A2(\adder_stage2[3][10] ), 
        .ZN(n6423) );
  NAND2_X1 U6821 ( .A1(\adder_stage2[2][11] ), .A2(\adder_stage2[3][11] ), 
        .ZN(n6029) );
  OAI21_X1 U6822 ( .B1(n6028), .B2(n6423), .A(n6029), .ZN(n5552) );
  AOI21_X1 U6823 ( .B1(n5553), .B2(n6023), .A(n5552), .ZN(n5822) );
  NAND2_X1 U6824 ( .A1(\adder_stage2[2][12] ), .A2(\adder_stage2[3][12] ), 
        .ZN(n5825) );
  OAI21_X1 U6825 ( .B1(n5822), .B2(n5824), .A(n5825), .ZN(n5554) );
  AOI21_X1 U6826 ( .B1(n5821), .B2(n5555), .A(n5554), .ZN(n5890) );
  OR2_X1 U6827 ( .A1(\adder_stage2[2][14] ), .A2(\adder_stage2[3][14] ), .ZN(
        n5892) );
  NOR2_X1 U6828 ( .A1(\adder_stage2[2][13] ), .A2(\adder_stage2[3][13] ), .ZN(
        n5889) );
  INV_X1 U6829 ( .A(n5889), .ZN(n5807) );
  NAND2_X1 U6830 ( .A1(n5892), .A2(n5807), .ZN(n5813) );
  INV_X1 U6831 ( .A(n5813), .ZN(n5556) );
  NOR2_X1 U6832 ( .A1(\adder_stage2[2][15] ), .A2(\adder_stage2[3][15] ), .ZN(
        n5560) );
  INV_X1 U6833 ( .A(n5560), .ZN(n5816) );
  NAND2_X1 U6834 ( .A1(n5556), .A2(n5816), .ZN(n5575) );
  INV_X1 U6835 ( .A(n5575), .ZN(n5557) );
  OR2_X1 U6836 ( .A1(\adder_stage2[2][16] ), .A2(\adder_stage2[3][16] ), .ZN(
        n5577) );
  NAND2_X1 U6837 ( .A1(n5557), .A2(n5577), .ZN(n5565) );
  NAND2_X1 U6838 ( .A1(\adder_stage2[2][13] ), .A2(\adder_stage2[3][13] ), 
        .ZN(n5888) );
  INV_X1 U6839 ( .A(n5888), .ZN(n5559) );
  NAND2_X1 U6840 ( .A1(\adder_stage2[2][14] ), .A2(\adder_stage2[3][14] ), 
        .ZN(n5891) );
  INV_X1 U6841 ( .A(n5891), .ZN(n5558) );
  AOI21_X1 U6842 ( .B1(n5892), .B2(n5559), .A(n5558), .ZN(n5812) );
  NAND2_X1 U6843 ( .A1(\adder_stage2[2][15] ), .A2(\adder_stage2[3][15] ), 
        .ZN(n5815) );
  OAI21_X1 U6844 ( .B1(n5812), .B2(n5560), .A(n5815), .ZN(n5561) );
  INV_X1 U6845 ( .A(n5561), .ZN(n5574) );
  INV_X1 U6846 ( .A(n5577), .ZN(n5562) );
  NAND2_X1 U6847 ( .A1(\adder_stage2[2][16] ), .A2(\adder_stage2[3][16] ), 
        .ZN(n5576) );
  OAI21_X1 U6848 ( .B1(n5574), .B2(n5562), .A(n5576), .ZN(n5563) );
  INV_X1 U6849 ( .A(n5563), .ZN(n5564) );
  OAI21_X1 U6850 ( .B1(n5890), .B2(n5565), .A(n5564), .ZN(n5566) );
  INV_X1 U6851 ( .A(n5566), .ZN(n5593) );
  NOR2_X1 U6852 ( .A1(\adder_stage2[2][17] ), .A2(\adder_stage2[3][17] ), .ZN(
        n5589) );
  NAND2_X1 U6853 ( .A1(\adder_stage2[2][17] ), .A2(\adder_stage2[3][17] ), 
        .ZN(n5590) );
  OAI21_X1 U6854 ( .B1(n5593), .B2(n5589), .A(n5590), .ZN(n5586) );
  OR2_X1 U6855 ( .A1(\adder_stage2[2][18] ), .A2(\adder_stage2[3][18] ), .ZN(
        n5584) );
  NAND2_X1 U6856 ( .A1(\adder_stage2[2][18] ), .A2(\adder_stage2[3][18] ), 
        .ZN(n5583) );
  INV_X1 U6857 ( .A(n5583), .ZN(n5567) );
  AOI21_X1 U6858 ( .B1(n5586), .B2(n5584), .A(n5567), .ZN(n8001) );
  NOR2_X1 U6859 ( .A1(\adder_stage2[2][19] ), .A2(\adder_stage2[3][19] ), .ZN(
        n8000) );
  INV_X1 U6860 ( .A(n8000), .ZN(n5568) );
  NAND2_X1 U6861 ( .A1(\adder_stage2[2][19] ), .A2(\adder_stage2[3][19] ), 
        .ZN(n7999) );
  NAND2_X1 U6862 ( .A1(n5568), .A2(n7999), .ZN(n5569) );
  XOR2_X1 U6863 ( .A(n8001), .B(n5569), .Z(n5570) );
  AOI22_X1 U6864 ( .A1(n5570), .A2(n8398), .B1(n8212), .B2(
        \adder_stage3[1][19] ), .ZN(n5571) );
  INV_X1 U6865 ( .A(n5571), .ZN(n9631) );
  AOI22_X1 U6866 ( .A1(\x_mult_f_int[11][8] ), .A2(n8186), .B1(n8048), .B2(
        \x_mult_f[11][8] ), .ZN(n5572) );
  INV_X1 U6867 ( .A(n5572), .ZN(n9065) );
  AOI22_X1 U6868 ( .A1(\x_mult_f_int[11][9] ), .A2(n8186), .B1(n8218), .B2(
        \x_mult_f[11][9] ), .ZN(n5573) );
  INV_X1 U6869 ( .A(n5573), .ZN(n9064) );
  OAI21_X1 U6870 ( .B1(n5890), .B2(n5575), .A(n5574), .ZN(n5579) );
  NAND2_X1 U6871 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  XNOR2_X1 U6872 ( .A(n5579), .B(n5578), .ZN(n5580) );
  AOI22_X1 U6873 ( .A1(n8401), .A2(n5580), .B1(n8048), .B2(
        \adder_stage3[1][16] ), .ZN(n5581) );
  INV_X1 U6874 ( .A(n5581), .ZN(n9634) );
  AOI22_X1 U6875 ( .A1(\x_mult_f_int[11][10] ), .A2(n8186), .B1(n8048), .B2(
        \x_mult_f[11][10] ), .ZN(n5582) );
  INV_X1 U6876 ( .A(n5582), .ZN(n9063) );
  NAND2_X1 U6877 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  XNOR2_X1 U6878 ( .A(n5586), .B(n5585), .ZN(n5587) );
  AOI22_X1 U6879 ( .A1(n5587), .A2(n8213), .B1(n8157), .B2(
        \adder_stage3[1][18] ), .ZN(n5588) );
  INV_X1 U6880 ( .A(n5588), .ZN(n9632) );
  INV_X1 U6881 ( .A(n5589), .ZN(n5591) );
  NAND2_X1 U6882 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  XOR2_X1 U6883 ( .A(n5593), .B(n5592), .Z(n5594) );
  AOI22_X1 U6884 ( .A1(n5594), .A2(n8213), .B1(n8212), .B2(
        \adder_stage3[1][17] ), .ZN(n5595) );
  INV_X1 U6885 ( .A(n5595), .ZN(n9633) );
  AOI22_X1 U6886 ( .A1(\x_mult_f_int[11][11] ), .A2(n8186), .B1(n8218), .B2(
        \x_mult_f[11][11] ), .ZN(n5596) );
  INV_X1 U6887 ( .A(n5596), .ZN(n9062) );
  INV_X1 U6888 ( .A(n5597), .ZN(n5664) );
  INV_X1 U6889 ( .A(n5598), .ZN(n5604) );
  NAND2_X1 U6890 ( .A1(n5604), .A2(n5602), .ZN(n5599) );
  XNOR2_X1 U6891 ( .A(n5664), .B(n5599), .ZN(n5600) );
  AOI22_X1 U6892 ( .A1(n5626), .A2(\adder_stage2[6][4] ), .B1(n6643), .B2(
        n5600), .ZN(n5601) );
  INV_X1 U6893 ( .A(n5601), .ZN(n9699) );
  INV_X1 U6894 ( .A(n5602), .ZN(n5603) );
  AOI21_X1 U6895 ( .B1(n5664), .B2(n5604), .A(n5603), .ZN(n5609) );
  INV_X1 U6896 ( .A(n5605), .ZN(n5607) );
  NAND2_X1 U6897 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  XOR2_X1 U6898 ( .A(n5609), .B(n5608), .Z(n5610) );
  AOI22_X1 U6899 ( .A1(n5626), .A2(\adder_stage2[6][5] ), .B1(n5908), .B2(
        n5610), .ZN(n5611) );
  INV_X1 U6900 ( .A(n5611), .ZN(n9698) );
  INV_X1 U6901 ( .A(n5612), .ZN(n5619) );
  INV_X1 U6902 ( .A(n5618), .ZN(n5613) );
  NAND2_X1 U6903 ( .A1(n5613), .A2(n5617), .ZN(n5614) );
  XOR2_X1 U6904 ( .A(n5619), .B(n5614), .Z(n5615) );
  AOI22_X1 U6905 ( .A1(n5626), .A2(\adder_stage2[6][2] ), .B1(n7992), .B2(
        n5615), .ZN(n5616) );
  INV_X1 U6906 ( .A(n5616), .ZN(n9701) );
  OAI21_X1 U6907 ( .B1(n5619), .B2(n5618), .A(n5617), .ZN(n5624) );
  INV_X1 U6908 ( .A(n5620), .ZN(n5622) );
  NAND2_X1 U6909 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  XNOR2_X1 U6910 ( .A(n5624), .B(n5623), .ZN(n5625) );
  AOI22_X1 U6911 ( .A1(n5626), .A2(\adder_stage2[6][3] ), .B1(n4002), .B2(
        n5625), .ZN(n5627) );
  INV_X1 U6912 ( .A(n5627), .ZN(n9700) );
  INV_X2 U6913 ( .A(n5811), .ZN(n6581) );
  BUF_X2 U6914 ( .A(n6955), .Z(n6643) );
  OR2_X1 U6915 ( .A1(\x_mult_f[14][0] ), .A2(\x_mult_f[15][0] ), .ZN(n5629) );
  AND2_X1 U6916 ( .A1(n5629), .A2(n5635), .ZN(n5630) );
  AOI22_X1 U6917 ( .A1(n6581), .A2(\adder_stage1[7][0] ), .B1(n6643), .B2(
        n5630), .ZN(n5631) );
  INV_X1 U6918 ( .A(n5631), .ZN(n9955) );
  INV_X1 U6919 ( .A(n5632), .ZN(n5634) );
  NAND2_X1 U6920 ( .A1(n5634), .A2(n5633), .ZN(n5636) );
  XOR2_X1 U6921 ( .A(n5636), .B(n5635), .Z(n5637) );
  AOI22_X1 U6922 ( .A1(n6581), .A2(\adder_stage1[7][1] ), .B1(n6643), .B2(
        n5637), .ZN(n5638) );
  INV_X1 U6923 ( .A(n5638), .ZN(n9954) );
  INV_X1 U6924 ( .A(n5639), .ZN(n6558) );
  INV_X1 U6925 ( .A(n5640), .ZN(n5658) );
  INV_X1 U6926 ( .A(n5657), .ZN(n5641) );
  AOI21_X1 U6927 ( .B1(n6558), .B2(n5658), .A(n5641), .ZN(n5646) );
  INV_X1 U6928 ( .A(n5642), .ZN(n5644) );
  NAND2_X1 U6929 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  XOR2_X1 U6930 ( .A(n5646), .B(n5645), .Z(n5647) );
  AOI22_X1 U6931 ( .A1(n6581), .A2(\adder_stage1[7][5] ), .B1(n6643), .B2(
        n5647), .ZN(n5648) );
  INV_X1 U6932 ( .A(n5648), .ZN(n9950) );
  INV_X1 U6933 ( .A(n5649), .ZN(n6553) );
  OAI21_X1 U6934 ( .B1(n6553), .B2(n6549), .A(n6550), .ZN(n5654) );
  INV_X1 U6935 ( .A(n5650), .ZN(n5652) );
  NAND2_X1 U6936 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  XNOR2_X1 U6937 ( .A(n5654), .B(n5653), .ZN(n5655) );
  AOI22_X1 U6938 ( .A1(n6581), .A2(\adder_stage1[7][3] ), .B1(n6643), .B2(
        n5655), .ZN(n5656) );
  INV_X1 U6939 ( .A(n5656), .ZN(n9952) );
  NAND2_X1 U6940 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  XNOR2_X1 U6941 ( .A(n6558), .B(n5659), .ZN(n5660) );
  AOI22_X1 U6942 ( .A1(n6581), .A2(\adder_stage1[7][4] ), .B1(n6643), .B2(
        n5660), .ZN(n5661) );
  INV_X1 U6943 ( .A(n5661), .ZN(n9951) );
  AOI21_X1 U6944 ( .B1(n5664), .B2(n5663), .A(n5662), .ZN(n5671) );
  INV_X1 U6945 ( .A(n5670), .ZN(n5665) );
  NAND2_X1 U6946 ( .A1(n5665), .A2(n5669), .ZN(n5666) );
  XOR2_X1 U6947 ( .A(n5671), .B(n5666), .Z(n5667) );
  AOI22_X1 U6948 ( .A1(n5678), .A2(\adder_stage2[6][6] ), .B1(n8318), .B2(
        n5667), .ZN(n5668) );
  INV_X1 U6949 ( .A(n5668), .ZN(n9697) );
  OAI21_X1 U6950 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5676) );
  INV_X1 U6951 ( .A(n5672), .ZN(n5674) );
  NAND2_X1 U6952 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  XNOR2_X1 U6953 ( .A(n5676), .B(n5675), .ZN(n5677) );
  AOI22_X1 U6954 ( .A1(n5678), .A2(\adder_stage2[6][7] ), .B1(n8329), .B2(
        n5677), .ZN(n5679) );
  INV_X1 U6955 ( .A(n5679), .ZN(n9696) );
  AOI22_X1 U6956 ( .A1(\x_mult_f_int[3][10] ), .A2(n8365), .B1(n8364), .B2(
        \x_mult_f[3][10] ), .ZN(n5680) );
  INV_X1 U6957 ( .A(n5680), .ZN(n8966) );
  AND2_X1 U6958 ( .A1(n5681), .A2(n5683), .ZN(n6008) );
  OR2_X1 U6959 ( .A1(\x_mult_f[30][13] ), .A2(\x_mult_f[31][13] ), .ZN(n6011)
         );
  AND2_X1 U6960 ( .A1(n6008), .A2(n6011), .ZN(n5682) );
  NAND2_X1 U6961 ( .A1(n5682), .A2(n6009), .ZN(n5689) );
  INV_X1 U6962 ( .A(n5683), .ZN(n5685) );
  OAI21_X1 U6963 ( .B1(n5686), .B2(n5685), .A(n5684), .ZN(n6007) );
  NAND2_X1 U6964 ( .A1(\x_mult_f[30][13] ), .A2(\x_mult_f[31][13] ), .ZN(n6010) );
  INV_X1 U6965 ( .A(n6010), .ZN(n5687) );
  AOI21_X1 U6966 ( .B1(n6007), .B2(n6011), .A(n5687), .ZN(n5688) );
  NAND2_X1 U6967 ( .A1(n5689), .A2(n5688), .ZN(n7951) );
  AOI22_X1 U6968 ( .A1(n5690), .A2(n8229), .B1(n8364), .B2(
        \adder_stage1[15][14] ), .ZN(n5691) );
  INV_X1 U6969 ( .A(n5691), .ZN(n9808) );
  AOI22_X1 U6970 ( .A1(\x_mult_f_int[3][8] ), .A2(n8365), .B1(n8364), .B2(
        \x_mult_f[3][8] ), .ZN(n5692) );
  INV_X1 U6971 ( .A(n5692), .ZN(n8968) );
  AOI22_X1 U6972 ( .A1(\x_mult_f_int[3][9] ), .A2(n8365), .B1(n8364), .B2(
        \x_mult_f[3][9] ), .ZN(n5693) );
  INV_X1 U6973 ( .A(n5693), .ZN(n8967) );
  INV_X1 U6974 ( .A(n5694), .ZN(n5761) );
  OAI21_X1 U6975 ( .B1(n5761), .B2(n5696), .A(n5695), .ZN(n5701) );
  INV_X1 U6976 ( .A(n5697), .ZN(n5699) );
  NAND2_X1 U6977 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  XNOR2_X1 U6978 ( .A(n5701), .B(n5700), .ZN(n5702) );
  AOI22_X1 U6979 ( .A1(n8088), .A2(\adder_stage4[0][12] ), .B1(n6256), .B2(
        n5702), .ZN(n5703) );
  INV_X1 U6980 ( .A(n5703), .ZN(n9576) );
  INV_X1 U6981 ( .A(n5760), .ZN(n5704) );
  NAND2_X1 U6982 ( .A1(n5704), .A2(n5759), .ZN(n5705) );
  XOR2_X1 U6983 ( .A(n5761), .B(n5705), .Z(n5706) );
  AOI22_X1 U6984 ( .A1(n7244), .A2(\adder_stage4[0][8] ), .B1(n6256), .B2(
        n5706), .ZN(n5707) );
  INV_X1 U6985 ( .A(n5707), .ZN(n9580) );
  INV_X1 U6986 ( .A(n5708), .ZN(n5710) );
  NAND2_X1 U6987 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  XOR2_X1 U6988 ( .A(n5712), .B(n5711), .Z(n5713) );
  AOI22_X1 U6989 ( .A1(n8400), .A2(\adder_stage4[0][13] ), .B1(n6256), .B2(
        n5713), .ZN(n5714) );
  INV_X1 U6990 ( .A(n5714), .ZN(n9575) );
  INV_X1 U6991 ( .A(n5715), .ZN(n5718) );
  INV_X1 U6992 ( .A(n5716), .ZN(n5717) );
  OAI21_X1 U6993 ( .B1(n5761), .B2(n5718), .A(n5717), .ZN(n5731) );
  INV_X1 U6994 ( .A(n5719), .ZN(n5729) );
  INV_X1 U6995 ( .A(n5728), .ZN(n5720) );
  AOI21_X1 U6996 ( .B1(n5731), .B2(n5729), .A(n5720), .ZN(n5725) );
  INV_X1 U6997 ( .A(n5721), .ZN(n5723) );
  NAND2_X1 U6998 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  XOR2_X1 U6999 ( .A(n5725), .B(n5724), .Z(n5726) );
  AOI22_X1 U7000 ( .A1(n7330), .A2(\adder_stage4[0][11] ), .B1(n6256), .B2(
        n5726), .ZN(n5727) );
  INV_X1 U7001 ( .A(n5727), .ZN(n9577) );
  NAND2_X1 U7002 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  XNOR2_X1 U7003 ( .A(n5731), .B(n5730), .ZN(n5732) );
  AOI22_X1 U7004 ( .A1(n6222), .A2(\adder_stage4[0][10] ), .B1(n6256), .B2(
        n5732), .ZN(n5733) );
  INV_X1 U7005 ( .A(n5733), .ZN(n9578) );
  INV_X1 U7006 ( .A(n5734), .ZN(n5772) );
  INV_X1 U7007 ( .A(n5735), .ZN(n5770) );
  INV_X1 U7008 ( .A(n5769), .ZN(n5736) );
  AOI21_X1 U7009 ( .B1(n5772), .B2(n5770), .A(n5736), .ZN(n5741) );
  INV_X1 U7010 ( .A(n5737), .ZN(n5739) );
  NAND2_X1 U7011 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  XOR2_X1 U7012 ( .A(n5741), .B(n5740), .Z(n5742) );
  AOI22_X1 U7013 ( .A1(n8195), .A2(\adder_stage4[0][5] ), .B1(n6256), .B2(
        n5742), .ZN(n5743) );
  INV_X1 U7014 ( .A(n5743), .ZN(n9583) );
  AOI21_X1 U7015 ( .B1(n5772), .B2(n5745), .A(n5744), .ZN(n5779) );
  OAI21_X1 U7016 ( .B1(n5779), .B2(n5775), .A(n5776), .ZN(n5750) );
  INV_X1 U7017 ( .A(n5746), .ZN(n5748) );
  NAND2_X1 U7018 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  XNOR2_X1 U7019 ( .A(n5750), .B(n5749), .ZN(n5751) );
  AOI22_X1 U7020 ( .A1(n7818), .A2(\adder_stage4[0][7] ), .B1(n6256), .B2(
        n5751), .ZN(n5752) );
  INV_X1 U7021 ( .A(n5752), .ZN(n9581) );
  NAND2_X1 U7022 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  XNOR2_X1 U7023 ( .A(n5756), .B(n5755), .ZN(n5757) );
  AOI22_X1 U7024 ( .A1(n8036), .A2(\adder_stage4[0][14] ), .B1(n6256), .B2(
        n5757), .ZN(n5758) );
  INV_X1 U7025 ( .A(n5758), .ZN(n9574) );
  OAI21_X1 U7026 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5766) );
  INV_X1 U7027 ( .A(n5762), .ZN(n5764) );
  NAND2_X1 U7028 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  XNOR2_X1 U7029 ( .A(n5766), .B(n5765), .ZN(n5767) );
  AOI22_X1 U7030 ( .A1(n8048), .A2(\adder_stage4[0][9] ), .B1(n6256), .B2(
        n5767), .ZN(n5768) );
  INV_X1 U7031 ( .A(n5768), .ZN(n9579) );
  NAND2_X1 U7032 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  XNOR2_X1 U7033 ( .A(n5772), .B(n5771), .ZN(n5773) );
  AOI22_X1 U7034 ( .A1(n8195), .A2(\adder_stage4[0][4] ), .B1(n6256), .B2(
        n5773), .ZN(n5774) );
  INV_X1 U7035 ( .A(n5774), .ZN(n9584) );
  INV_X1 U7036 ( .A(n5775), .ZN(n5777) );
  NAND2_X1 U7037 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  XOR2_X1 U7038 ( .A(n5779), .B(n5778), .Z(n5780) );
  AOI22_X1 U7039 ( .A1(n8218), .A2(\adder_stage4[0][6] ), .B1(n6256), .B2(
        n5780), .ZN(n5781) );
  INV_X1 U7040 ( .A(n5781), .ZN(n9582) );
  NOR2_X1 U7041 ( .A1(\x_mult_f[6][2] ), .A2(\x_mult_f[7][2] ), .ZN(n7170) );
  NOR2_X1 U7042 ( .A1(n7170), .A2(n6654), .ZN(n5783) );
  NOR2_X1 U7043 ( .A1(\x_mult_f[6][1] ), .A2(\x_mult_f[7][1] ), .ZN(n6191) );
  NAND2_X1 U7044 ( .A1(\x_mult_f[6][0] ), .A2(\x_mult_f[7][0] ), .ZN(n6194) );
  NAND2_X1 U7045 ( .A1(\x_mult_f[6][1] ), .A2(\x_mult_f[7][1] ), .ZN(n6192) );
  OAI21_X1 U7046 ( .B1(n6191), .B2(n6194), .A(n6192), .ZN(n6653) );
  NAND2_X1 U7047 ( .A1(\x_mult_f[6][2] ), .A2(\x_mult_f[7][2] ), .ZN(n7171) );
  NAND2_X1 U7048 ( .A1(\x_mult_f[6][3] ), .A2(\x_mult_f[7][3] ), .ZN(n6655) );
  OAI21_X1 U7049 ( .B1(n6654), .B2(n7171), .A(n6655), .ZN(n5782) );
  AOI21_X1 U7050 ( .B1(n5783), .B2(n6653), .A(n5782), .ZN(n6646) );
  NOR2_X1 U7051 ( .A1(\x_mult_f[6][4] ), .A2(\x_mult_f[7][4] ), .ZN(n6661) );
  NOR2_X1 U7052 ( .A1(\x_mult_f[6][5] ), .A2(\x_mult_f[7][5] ), .ZN(n6663) );
  NOR2_X1 U7053 ( .A1(n6661), .A2(n6663), .ZN(n6648) );
  NOR2_X1 U7054 ( .A1(\x_mult_f[6][6] ), .A2(\x_mult_f[7][6] ), .ZN(n6676) );
  NOR2_X1 U7055 ( .A1(\x_mult_f[6][7] ), .A2(\x_mult_f[7][7] ), .ZN(n6678) );
  NOR2_X1 U7056 ( .A1(n6676), .A2(n6678), .ZN(n5785) );
  NAND2_X1 U7057 ( .A1(n6648), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U7058 ( .A1(\x_mult_f[6][4] ), .A2(\x_mult_f[7][4] ), .ZN(n7177) );
  NAND2_X1 U7059 ( .A1(\x_mult_f[6][5] ), .A2(\x_mult_f[7][5] ), .ZN(n6664) );
  OAI21_X1 U7060 ( .B1(n6663), .B2(n7177), .A(n6664), .ZN(n6647) );
  NAND2_X1 U7061 ( .A1(\x_mult_f[6][6] ), .A2(\x_mult_f[7][6] ), .ZN(n6675) );
  NAND2_X1 U7062 ( .A1(\x_mult_f[6][7] ), .A2(\x_mult_f[7][7] ), .ZN(n6679) );
  OAI21_X1 U7063 ( .B1(n6678), .B2(n6675), .A(n6679), .ZN(n5784) );
  AOI21_X1 U7064 ( .B1(n5785), .B2(n6647), .A(n5784), .ZN(n5786) );
  OAI21_X1 U7065 ( .B1(n6646), .B2(n5787), .A(n5786), .ZN(n7132) );
  OR2_X1 U7066 ( .A1(\x_mult_f[6][8] ), .A2(\x_mult_f[7][8] ), .ZN(n7130) );
  NAND2_X1 U7067 ( .A1(\x_mult_f[6][8] ), .A2(\x_mult_f[7][8] ), .ZN(n7129) );
  INV_X1 U7068 ( .A(n7129), .ZN(n5788) );
  INV_X1 U7069 ( .A(n7163), .ZN(n5797) );
  OR2_X1 U7070 ( .A1(\x_mult_f[6][10] ), .A2(\x_mult_f[7][10] ), .ZN(n7165) );
  NOR2_X1 U7071 ( .A1(\x_mult_f[6][9] ), .A2(\x_mult_f[7][9] ), .ZN(n7162) );
  INV_X1 U7072 ( .A(n7162), .ZN(n6670) );
  NAND2_X1 U7073 ( .A1(n7165), .A2(n6670), .ZN(n7153) );
  INV_X1 U7074 ( .A(n7153), .ZN(n5789) );
  NOR2_X1 U7075 ( .A1(\x_mult_f[6][11] ), .A2(\x_mult_f[7][11] ), .ZN(n5792)
         );
  INV_X1 U7076 ( .A(n5792), .ZN(n7156) );
  NAND2_X1 U7077 ( .A1(n5789), .A2(n7156), .ZN(n7137) );
  OR2_X1 U7078 ( .A1(\x_mult_f[6][12] ), .A2(\x_mult_f[7][12] ), .ZN(n7139) );
  INV_X1 U7079 ( .A(n7139), .ZN(n5794) );
  NOR2_X1 U7080 ( .A1(n7137), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7081 ( .A1(\x_mult_f[6][9] ), .A2(\x_mult_f[7][9] ), .ZN(n7161) );
  INV_X1 U7082 ( .A(n7161), .ZN(n5791) );
  NAND2_X1 U7083 ( .A1(\x_mult_f[6][10] ), .A2(\x_mult_f[7][10] ), .ZN(n7164)
         );
  INV_X1 U7084 ( .A(n7164), .ZN(n5790) );
  AOI21_X1 U7085 ( .B1(n7165), .B2(n5791), .A(n5790), .ZN(n7152) );
  NAND2_X1 U7086 ( .A1(\x_mult_f[6][11] ), .A2(\x_mult_f[7][11] ), .ZN(n7155)
         );
  OAI21_X1 U7087 ( .B1(n7152), .B2(n5792), .A(n7155), .ZN(n5793) );
  INV_X1 U7088 ( .A(n5793), .ZN(n7136) );
  NAND2_X1 U7089 ( .A1(\x_mult_f[6][12] ), .A2(\x_mult_f[7][12] ), .ZN(n7138)
         );
  OAI21_X1 U7090 ( .B1(n7136), .B2(n5794), .A(n7138), .ZN(n5795) );
  AOI21_X1 U7091 ( .B1(n5797), .B2(n5796), .A(n5795), .ZN(n5804) );
  NOR2_X1 U7092 ( .A1(\x_mult_f[6][13] ), .A2(\x_mult_f[7][13] ), .ZN(n5803)
         );
  INV_X1 U7093 ( .A(n5803), .ZN(n5798) );
  NAND2_X1 U7094 ( .A1(\x_mult_f[6][13] ), .A2(\x_mult_f[7][13] ), .ZN(n5802)
         );
  NAND2_X1 U7095 ( .A1(n5798), .A2(n5802), .ZN(n5799) );
  XOR2_X1 U7096 ( .A(n5804), .B(n5799), .Z(n5800) );
  AOI22_X1 U7097 ( .A1(n5800), .A2(n8150), .B1(n8078), .B2(
        \adder_stage1[3][13] ), .ZN(n5801) );
  INV_X1 U7098 ( .A(n5801), .ZN(n10007) );
  OAI21_X1 U7099 ( .B1(n5804), .B2(n5803), .A(n5802), .ZN(n7979) );
  AOI22_X1 U7100 ( .A1(n5805), .A2(n8186), .B1(n8078), .B2(
        \adder_stage1[3][14] ), .ZN(n5806) );
  INV_X1 U7101 ( .A(n5806), .ZN(n10006) );
  INV_X2 U7102 ( .A(n5811), .ZN(n6428) );
  BUF_X2 U7103 ( .A(n6955), .Z(n5908) );
  NAND2_X1 U7104 ( .A1(n5807), .A2(n5888), .ZN(n5808) );
  XOR2_X1 U7105 ( .A(n5890), .B(n5808), .Z(n5809) );
  AOI22_X1 U7106 ( .A1(n6428), .A2(\adder_stage3[1][13] ), .B1(n5908), .B2(
        n5809), .ZN(n5810) );
  INV_X1 U7107 ( .A(n5810), .ZN(n9637) );
  INV_X2 U7108 ( .A(n5811), .ZN(n5909) );
  OAI21_X1 U7109 ( .B1(n5890), .B2(n5813), .A(n5812), .ZN(n5814) );
  INV_X1 U7110 ( .A(n5814), .ZN(n5818) );
  NAND2_X1 U7111 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  XOR2_X1 U7112 ( .A(n5818), .B(n5817), .Z(n5819) );
  AOI22_X1 U7113 ( .A1(n5909), .A2(\adder_stage3[1][15] ), .B1(n5908), .B2(
        n5819), .ZN(n5820) );
  INV_X1 U7114 ( .A(n5820), .ZN(n9635) );
  INV_X1 U7115 ( .A(n5821), .ZN(n6046) );
  OAI21_X1 U7116 ( .B1(n6046), .B2(n5823), .A(n5822), .ZN(n5828) );
  INV_X1 U7117 ( .A(n5824), .ZN(n5826) );
  NAND2_X1 U7118 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  XNOR2_X1 U7119 ( .A(n5828), .B(n5827), .ZN(n5829) );
  AOI22_X1 U7120 ( .A1(n6428), .A2(\adder_stage3[1][12] ), .B1(n5908), .B2(
        n5829), .ZN(n5830) );
  INV_X1 U7121 ( .A(n5830), .ZN(n9638) );
  INV_X1 U7122 ( .A(n5831), .ZN(n5855) );
  INV_X1 U7123 ( .A(n5832), .ZN(n5854) );
  NAND2_X1 U7124 ( .A1(n5854), .A2(n5852), .ZN(n5833) );
  XNOR2_X1 U7125 ( .A(n5855), .B(n5833), .ZN(n5834) );
  AOI22_X1 U7126 ( .A1(n5909), .A2(\adder_stage2[3][4] ), .B1(n5908), .B2(
        n5834), .ZN(n5835) );
  INV_X1 U7127 ( .A(n5835), .ZN(n9750) );
  AOI21_X1 U7128 ( .B1(n5855), .B2(n5837), .A(n5836), .ZN(n5844) );
  INV_X1 U7129 ( .A(n5843), .ZN(n5838) );
  NAND2_X1 U7130 ( .A1(n5838), .A2(n5842), .ZN(n5839) );
  XOR2_X1 U7131 ( .A(n5844), .B(n5839), .Z(n5840) );
  AOI22_X1 U7132 ( .A1(n5909), .A2(\adder_stage2[3][6] ), .B1(n5908), .B2(
        n5840), .ZN(n5841) );
  INV_X1 U7133 ( .A(n5841), .ZN(n9748) );
  OAI21_X1 U7134 ( .B1(n5844), .B2(n5843), .A(n5842), .ZN(n5849) );
  INV_X1 U7135 ( .A(n5845), .ZN(n5847) );
  NAND2_X1 U7136 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U7137 ( .A(n5849), .B(n5848), .ZN(n5850) );
  AOI22_X1 U7138 ( .A1(n5909), .A2(\adder_stage2[3][7] ), .B1(n5908), .B2(
        n5850), .ZN(n5851) );
  INV_X1 U7139 ( .A(n5851), .ZN(n9747) );
  INV_X1 U7140 ( .A(n5852), .ZN(n5853) );
  AOI21_X1 U7141 ( .B1(n5855), .B2(n5854), .A(n5853), .ZN(n5860) );
  INV_X1 U7142 ( .A(n5856), .ZN(n5858) );
  NAND2_X1 U7143 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  XOR2_X1 U7144 ( .A(n5860), .B(n5859), .Z(n5861) );
  AOI22_X1 U7145 ( .A1(n5909), .A2(\adder_stage2[3][5] ), .B1(n5908), .B2(
        n5861), .ZN(n5862) );
  INV_X1 U7146 ( .A(n5862), .ZN(n9749) );
  INV_X1 U7147 ( .A(n5863), .ZN(n5873) );
  INV_X1 U7148 ( .A(n5872), .ZN(n5864) );
  NAND2_X1 U7149 ( .A1(n5864), .A2(n5871), .ZN(n5865) );
  XOR2_X1 U7150 ( .A(n5873), .B(n5865), .Z(n5866) );
  AOI22_X1 U7151 ( .A1(n5909), .A2(\adder_stage2[3][2] ), .B1(n5908), .B2(
        n5866), .ZN(n5867) );
  INV_X1 U7152 ( .A(n5867), .ZN(n9752) );
  OR2_X1 U7153 ( .A1(\adder_stage1[6][0] ), .A2(\adder_stage1[7][0] ), .ZN(
        n5868) );
  AND2_X1 U7154 ( .A1(n5868), .A2(n5884), .ZN(n5869) );
  AOI22_X1 U7155 ( .A1(n5909), .A2(\adder_stage2[3][0] ), .B1(n5908), .B2(
        n5869), .ZN(n5870) );
  INV_X1 U7156 ( .A(n5870), .ZN(n9754) );
  OAI21_X1 U7157 ( .B1(n5873), .B2(n5872), .A(n5871), .ZN(n5878) );
  INV_X1 U7158 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7159 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  XNOR2_X1 U7160 ( .A(n5878), .B(n5877), .ZN(n5879) );
  AOI22_X1 U7161 ( .A1(n5909), .A2(\adder_stage2[3][3] ), .B1(n5908), .B2(
        n5879), .ZN(n5880) );
  INV_X1 U7162 ( .A(n5880), .ZN(n9751) );
  INV_X1 U7163 ( .A(n5881), .ZN(n5883) );
  NAND2_X1 U7164 ( .A1(n5883), .A2(n5882), .ZN(n5885) );
  XOR2_X1 U7165 ( .A(n5885), .B(n5884), .Z(n5886) );
  AOI22_X1 U7166 ( .A1(n5909), .A2(\adder_stage2[3][1] ), .B1(n5908), .B2(
        n5886), .ZN(n5887) );
  INV_X1 U7167 ( .A(n5887), .ZN(n9753) );
  OAI21_X1 U7168 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(n5894) );
  NAND2_X1 U7169 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  XNOR2_X1 U7170 ( .A(n5894), .B(n5893), .ZN(n5895) );
  AOI22_X1 U7171 ( .A1(n5909), .A2(\adder_stage3[1][14] ), .B1(n5908), .B2(
        n5895), .ZN(n5896) );
  INV_X1 U7172 ( .A(n5896), .ZN(n9636) );
  INV_X1 U7173 ( .A(n6533), .ZN(n6574) );
  NAND2_X1 U7174 ( .A1(n5897), .A2(n5901), .ZN(n5898) );
  XOR2_X1 U7175 ( .A(n6574), .B(n5898), .Z(n5899) );
  AOI22_X1 U7176 ( .A1(n5909), .A2(\adder_stage2[3][8] ), .B1(n5908), .B2(
        n5899), .ZN(n5900) );
  INV_X1 U7177 ( .A(n5900), .ZN(n9746) );
  OAI21_X1 U7178 ( .B1(n6574), .B2(n5902), .A(n5901), .ZN(n5906) );
  NAND2_X1 U7179 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  XNOR2_X1 U7180 ( .A(n5906), .B(n5905), .ZN(n5907) );
  AOI22_X1 U7181 ( .A1(n5909), .A2(\adder_stage2[3][9] ), .B1(n5908), .B2(
        n5907), .ZN(n5910) );
  INV_X1 U7182 ( .A(n5910), .ZN(n9745) );
  FA_X1 U7183 ( .A(\x_mult_f[14][14] ), .B(\x_mult_f[15][14] ), .CI(n5911), 
        .CO(n7938), .S(n5912) );
  AOI22_X1 U7184 ( .A1(n5912), .A2(n7117), .B1(n8088), .B2(
        \adder_stage1[7][14] ), .ZN(n5913) );
  INV_X1 U7185 ( .A(n5913), .ZN(n9941) );
  AOI22_X1 U7186 ( .A1(n8265), .A2(\x_mult_f_int[19][5] ), .B1(n7285), .B2(
        \x_mult_f[19][5] ), .ZN(n5914) );
  INV_X1 U7187 ( .A(n5914), .ZN(n9178) );
  AOI22_X1 U7188 ( .A1(n4002), .A2(\x_mult_f_int[8][5] ), .B1(n7030), .B2(
        \x_mult_f[8][5] ), .ZN(n5915) );
  INV_X1 U7189 ( .A(n5915), .ZN(n9037) );
  AOI22_X1 U7190 ( .A1(\x_mult_f_int[8][6] ), .A2(n8150), .B1(n8195), .B2(
        \x_mult_f[8][6] ), .ZN(n5916) );
  INV_X1 U7191 ( .A(n5916), .ZN(n9036) );
  AOI22_X1 U7192 ( .A1(\x_mult_f_int[31][11] ), .A2(n8189), .B1(n8202), .B2(
        \x_mult_f[31][11] ), .ZN(n5917) );
  INV_X1 U7193 ( .A(n5917), .ZN(n9282) );
  AOI22_X1 U7194 ( .A1(\x_mult_f_int[30][10] ), .A2(n8150), .B1(n8218), .B2(
        \x_mult_f[30][10] ), .ZN(n5918) );
  INV_X1 U7195 ( .A(n5918), .ZN(n9269) );
  AOI22_X1 U7196 ( .A1(\x_mult_f_int[30][8] ), .A2(n8150), .B1(n8218), .B2(
        \x_mult_f[30][8] ), .ZN(n5919) );
  INV_X1 U7197 ( .A(n5919), .ZN(n9271) );
  AOI22_X1 U7198 ( .A1(\x_mult_f_int[30][7] ), .A2(n5921), .B1(n8218), .B2(
        \x_mult_f[30][7] ), .ZN(n5920) );
  INV_X1 U7199 ( .A(n5920), .ZN(n9272) );
  AOI22_X1 U7200 ( .A1(\x_mult_f_int[30][6] ), .A2(n5921), .B1(n8218), .B2(
        \x_mult_f[30][6] ), .ZN(n5922) );
  INV_X1 U7201 ( .A(n5922), .ZN(n9273) );
  AOI22_X1 U7202 ( .A1(n8216), .A2(\x_mult_f_int[30][5] ), .B1(n8202), .B2(
        \x_mult_f[30][5] ), .ZN(n5923) );
  INV_X1 U7203 ( .A(n5923), .ZN(n9274) );
  AOI22_X1 U7204 ( .A1(\x_mult_f_int[31][10] ), .A2(n6643), .B1(n8202), .B2(
        \x_mult_f[31][10] ), .ZN(n5924) );
  INV_X1 U7205 ( .A(n5924), .ZN(n9283) );
  AOI22_X1 U7206 ( .A1(\x_mult_f_int[31][8] ), .A2(n5908), .B1(n8202), .B2(
        \x_mult_f[31][8] ), .ZN(n5925) );
  INV_X1 U7207 ( .A(n5925), .ZN(n9285) );
  AOI22_X1 U7208 ( .A1(\x_mult_f_int[1][11] ), .A2(n7511), .B1(n8036), .B2(
        \x_mult_f[1][11] ), .ZN(n5926) );
  INV_X1 U7209 ( .A(n5926), .ZN(n8939) );
  AOI22_X1 U7210 ( .A1(\x_mult_f_int[30][11] ), .A2(n8150), .B1(n8218), .B2(
        \x_mult_f[30][11] ), .ZN(n5927) );
  INV_X1 U7211 ( .A(n5927), .ZN(n9268) );
  AOI22_X1 U7212 ( .A1(\x_mult_f_int[5][10] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][10] ), .ZN(n5928) );
  INV_X1 U7213 ( .A(n5928), .ZN(n8990) );
  AOI22_X1 U7214 ( .A1(\x_mult_f_int[5][8] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][8] ), .ZN(n5929) );
  INV_X1 U7215 ( .A(n5929), .ZN(n8992) );
  AOI22_X1 U7216 ( .A1(\x_mult_f_int[5][11] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][11] ), .ZN(n5930) );
  INV_X1 U7217 ( .A(n5930), .ZN(n8989) );
  NAND2_X1 U7218 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  XNOR2_X1 U7219 ( .A(n5934), .B(n5933), .ZN(n5935) );
  AOI22_X1 U7220 ( .A1(n8387), .A2(n5935), .B1(n8036), .B2(
        \adder_stage4[1][16] ), .ZN(n5936) );
  INV_X1 U7221 ( .A(n5936), .ZN(n9551) );
  AOI22_X1 U7222 ( .A1(\x_mult_f_int[30][9] ), .A2(n8150), .B1(n8218), .B2(
        \x_mult_f[30][9] ), .ZN(n5937) );
  INV_X1 U7223 ( .A(n5937), .ZN(n9270) );
  AOI22_X1 U7224 ( .A1(\x_mult_f_int[31][9] ), .A2(n7992), .B1(n8202), .B2(
        \x_mult_f[31][9] ), .ZN(n5938) );
  INV_X1 U7225 ( .A(n5938), .ZN(n9284) );
  AOI22_X1 U7226 ( .A1(\x_mult_f_int[5][9] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][9] ), .ZN(n5939) );
  INV_X1 U7227 ( .A(n5939), .ZN(n8991) );
  AOI22_X1 U7228 ( .A1(\x_mult_f_int[3][11] ), .A2(n8365), .B1(n8202), .B2(
        \x_mult_f[3][11] ), .ZN(n5940) );
  INV_X1 U7229 ( .A(n5940), .ZN(n8965) );
  AOI22_X1 U7230 ( .A1(\x_mult_f_int[16][9] ), .A2(n8265), .B1(n8218), .B2(
        \x_mult_f[16][9] ), .ZN(n5941) );
  INV_X1 U7231 ( .A(n5941), .ZN(n9133) );
  AOI22_X1 U7232 ( .A1(\x_mult_f_int[16][10] ), .A2(n8265), .B1(n8046), .B2(
        \x_mult_f[16][10] ), .ZN(n5942) );
  INV_X1 U7233 ( .A(n5942), .ZN(n9132) );
  AOI22_X1 U7234 ( .A1(\x_mult_f_int[16][8] ), .A2(n8180), .B1(n8048), .B2(
        \x_mult_f[16][8] ), .ZN(n5943) );
  INV_X1 U7235 ( .A(n5943), .ZN(n9134) );
  AOI22_X1 U7236 ( .A1(n8265), .A2(\x_mult_f_int[16][5] ), .B1(n8157), .B2(
        \x_mult_f[16][5] ), .ZN(n5944) );
  INV_X1 U7237 ( .A(n5944), .ZN(n9137) );
  AOI22_X1 U7238 ( .A1(\x_mult_f_int[17][10] ), .A2(n8180), .B1(n8157), .B2(
        \x_mult_f[17][10] ), .ZN(n5945) );
  INV_X1 U7239 ( .A(n5945), .ZN(n9145) );
  AOI22_X1 U7240 ( .A1(\x_mult_f_int[16][7] ), .A2(n8180), .B1(n8218), .B2(
        \x_mult_f[16][7] ), .ZN(n5946) );
  INV_X1 U7241 ( .A(n5946), .ZN(n9135) );
  AOI22_X1 U7242 ( .A1(\x_mult_f_int[16][6] ), .A2(n8180), .B1(n8048), .B2(
        \x_mult_f[16][6] ), .ZN(n5947) );
  INV_X1 U7243 ( .A(n5947), .ZN(n9136) );
  AOI22_X1 U7244 ( .A1(\x_mult_f_int[17][11] ), .A2(n8180), .B1(n8157), .B2(
        \x_mult_f[17][11] ), .ZN(n5948) );
  INV_X1 U7245 ( .A(n5948), .ZN(n9144) );
  FA_X1 U7246 ( .A(\x_mult_f[20][14] ), .B(\x_mult_f[21][14] ), .CI(n5949), 
        .CO(n8393), .S(n5951) );
  AOI22_X1 U7247 ( .A1(n5951), .A2(n8389), .B1(n8395), .B2(
        \adder_stage1[10][14] ), .ZN(n5952) );
  INV_X1 U7248 ( .A(n5952), .ZN(n9892) );
  AOI22_X1 U7249 ( .A1(\x_mult_f_int[20][8] ), .A2(n8229), .B1(n8381), .B2(
        \x_mult_f[20][8] ), .ZN(n8810) );
  AOI22_X1 U7250 ( .A1(\x_mult_f_int[20][10] ), .A2(n8399), .B1(n8381), .B2(
        \x_mult_f[20][10] ), .ZN(n8808) );
  INV_X1 U7251 ( .A(n5953), .ZN(n8237) );
  AOI21_X1 U7252 ( .B1(n8374), .B2(n8232), .A(n8237), .ZN(n5955) );
  OR2_X1 U7253 ( .A1(\adder_stage2[0][17] ), .A2(\adder_stage2[1][17] ), .ZN(
        n8236) );
  NAND2_X1 U7254 ( .A1(\adder_stage2[0][17] ), .A2(\adder_stage2[1][17] ), 
        .ZN(n8234) );
  NAND2_X1 U7255 ( .A1(n8236), .A2(n8234), .ZN(n5954) );
  XOR2_X1 U7256 ( .A(n5955), .B(n5954), .Z(n5956) );
  AOI22_X1 U7257 ( .A1(n5956), .A2(n8399), .B1(n8381), .B2(
        \adder_stage3[0][17] ), .ZN(n5957) );
  INV_X1 U7258 ( .A(n5957), .ZN(n9652) );
  AOI22_X1 U7259 ( .A1(\x_mult_f_int[20][11] ), .A2(n8186), .B1(n8381), .B2(
        \x_mult_f[20][11] ), .ZN(n8807) );
  AOI22_X1 U7260 ( .A1(\x_mult_f_int[20][9] ), .A2(n7774), .B1(n8381), .B2(
        \x_mult_f[20][9] ), .ZN(n8809) );
  AOI22_X1 U7261 ( .A1(\x_mult_f_int[23][8] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][8] ), .ZN(n5958) );
  INV_X1 U7262 ( .A(n5958), .ZN(n9209) );
  AOI22_X1 U7263 ( .A1(\x_mult_f_int[23][9] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][9] ), .ZN(n5959) );
  INV_X1 U7264 ( .A(n5959), .ZN(n9208) );
  AOI22_X1 U7265 ( .A1(\x_mult_f_int[23][10] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][10] ), .ZN(n5960) );
  INV_X1 U7266 ( .A(n5960), .ZN(n9207) );
  FA_X1 U7267 ( .A(\x_mult_f[22][14] ), .B(\x_mult_f[23][14] ), .CI(n5961), 
        .CO(n8076), .S(n5962) );
  AOI22_X1 U7268 ( .A1(n5962), .A2(n5950), .B1(n8078), .B2(
        \adder_stage1[11][14] ), .ZN(n5963) );
  INV_X1 U7269 ( .A(n5963), .ZN(n9876) );
  AOI22_X1 U7270 ( .A1(\x_mult_f_int[23][11] ), .A2(n5950), .B1(n8078), .B2(
        \x_mult_f[23][11] ), .ZN(n5964) );
  INV_X1 U7271 ( .A(n5964), .ZN(n9206) );
  AOI22_X1 U7272 ( .A1(\x_mult_f_int[18][7] ), .A2(n8194), .B1(n8157), .B2(
        \x_mult_f[18][7] ), .ZN(n5965) );
  INV_X1 U7273 ( .A(n5965), .ZN(n9162) );
  AOI22_X1 U7274 ( .A1(\x_mult_f_int[18][8] ), .A2(n6221), .B1(n8157), .B2(
        \x_mult_f[18][8] ), .ZN(n5966) );
  INV_X1 U7275 ( .A(n5966), .ZN(n9161) );
  AOI22_X1 U7276 ( .A1(\x_mult_f_int[18][10] ), .A2(n6915), .B1(n8157), .B2(
        \x_mult_f[18][10] ), .ZN(n5967) );
  INV_X1 U7277 ( .A(n5967), .ZN(n9159) );
  AOI22_X1 U7278 ( .A1(\x_mult_f_int[18][9] ), .A2(n7117), .B1(n8157), .B2(
        \x_mult_f[18][9] ), .ZN(n5968) );
  INV_X1 U7279 ( .A(n5968), .ZN(n9160) );
  AOI22_X1 U7280 ( .A1(\x_mult_f_int[18][6] ), .A2(n8213), .B1(n8157), .B2(
        \x_mult_f[18][6] ), .ZN(n5969) );
  INV_X1 U7281 ( .A(n5969), .ZN(n9163) );
  NOR2_X1 U7282 ( .A1(\adder_stage1[8][2] ), .A2(\adder_stage1[9][2] ), .ZN(
        n7343) );
  NOR2_X1 U7283 ( .A1(\adder_stage1[8][3] ), .A2(\adder_stage1[9][3] ), .ZN(
        n7345) );
  NOR2_X1 U7284 ( .A1(n7343), .A2(n7345), .ZN(n5971) );
  NOR2_X1 U7285 ( .A1(\adder_stage1[8][1] ), .A2(\adder_stage1[9][1] ), .ZN(
        n7334) );
  NAND2_X1 U7286 ( .A1(\adder_stage1[8][0] ), .A2(\adder_stage1[9][0] ), .ZN(
        n7337) );
  NAND2_X1 U7287 ( .A1(\adder_stage1[8][1] ), .A2(\adder_stage1[9][1] ), .ZN(
        n7335) );
  OAI21_X1 U7288 ( .B1(n7334), .B2(n7337), .A(n7335), .ZN(n7315) );
  NAND2_X1 U7289 ( .A1(\adder_stage1[8][2] ), .A2(\adder_stage1[9][2] ), .ZN(
        n7342) );
  NAND2_X1 U7290 ( .A1(\adder_stage1[8][3] ), .A2(\adder_stage1[9][3] ), .ZN(
        n7346) );
  OAI21_X1 U7291 ( .B1(n7345), .B2(n7342), .A(n7346), .ZN(n5970) );
  AOI21_X1 U7292 ( .B1(n5971), .B2(n7315), .A(n5970), .ZN(n7287) );
  NOR2_X1 U7293 ( .A1(\adder_stage1[8][4] ), .A2(\adder_stage1[9][4] ), .ZN(
        n7288) );
  NOR2_X1 U7294 ( .A1(\adder_stage1[8][5] ), .A2(\adder_stage1[9][5] ), .ZN(
        n7290) );
  NOR2_X1 U7295 ( .A1(n7288), .A2(n7290), .ZN(n7550) );
  NOR2_X1 U7296 ( .A1(\adder_stage1[8][6] ), .A2(\adder_stage1[9][6] ), .ZN(
        n7607) );
  NOR2_X1 U7297 ( .A1(\adder_stage1[9][7] ), .A2(\adder_stage1[8][7] ), .ZN(
        n7552) );
  NOR2_X1 U7298 ( .A1(n7607), .A2(n7552), .ZN(n5973) );
  NAND2_X1 U7299 ( .A1(n7550), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7300 ( .A1(\adder_stage1[8][4] ), .A2(\adder_stage1[9][4] ), .ZN(
        n7352) );
  NAND2_X1 U7301 ( .A1(\adder_stage1[8][5] ), .A2(\adder_stage1[9][5] ), .ZN(
        n7291) );
  OAI21_X1 U7302 ( .B1(n7290), .B2(n7352), .A(n7291), .ZN(n7549) );
  NAND2_X1 U7303 ( .A1(\adder_stage1[8][6] ), .A2(\adder_stage1[9][6] ), .ZN(
        n7608) );
  NAND2_X1 U7304 ( .A1(\adder_stage1[9][7] ), .A2(\adder_stage1[8][7] ), .ZN(
        n7553) );
  OAI21_X1 U7305 ( .B1(n7552), .B2(n7608), .A(n7553), .ZN(n5972) );
  AOI21_X1 U7306 ( .B1(n5973), .B2(n7549), .A(n5972), .ZN(n5974) );
  OAI21_X1 U7307 ( .B1(n7287), .B2(n5975), .A(n5974), .ZN(n7636) );
  NOR2_X1 U7308 ( .A1(\adder_stage1[8][8] ), .A2(\adder_stage1[9][8] ), .ZN(
        n7646) );
  INV_X1 U7309 ( .A(n7646), .ZN(n7654) );
  OR2_X1 U7310 ( .A1(\adder_stage1[8][9] ), .A2(\adder_stage1[9][9] ), .ZN(
        n7648) );
  NAND2_X1 U7311 ( .A1(n7654), .A2(n7648), .ZN(n7638) );
  NOR2_X1 U7312 ( .A1(\adder_stage1[8][10] ), .A2(\adder_stage1[9][10] ), .ZN(
        n7639) );
  NOR2_X1 U7313 ( .A1(n7638), .A2(n7639), .ZN(n7593) );
  OR2_X1 U7314 ( .A1(\adder_stage1[8][12] ), .A2(\adder_stage1[9][12] ), .ZN(
        n7619) );
  NOR2_X1 U7315 ( .A1(\adder_stage1[8][11] ), .A2(\adder_stage1[9][11] ), .ZN(
        n7616) );
  INV_X1 U7316 ( .A(n7616), .ZN(n7596) );
  NAND2_X1 U7317 ( .A1(n7619), .A2(n7596), .ZN(n5983) );
  INV_X1 U7318 ( .A(n5983), .ZN(n5976) );
  AND2_X1 U7319 ( .A1(n7593), .A2(n5976), .ZN(n5985) );
  NAND2_X1 U7320 ( .A1(\adder_stage1[8][8] ), .A2(\adder_stage1[9][8] ), .ZN(
        n7653) );
  INV_X1 U7321 ( .A(n7653), .ZN(n5978) );
  NAND2_X1 U7322 ( .A1(\adder_stage1[8][9] ), .A2(\adder_stage1[9][9] ), .ZN(
        n7647) );
  INV_X1 U7323 ( .A(n7647), .ZN(n5977) );
  AOI21_X1 U7324 ( .B1(n7648), .B2(n5978), .A(n5977), .ZN(n7637) );
  NAND2_X1 U7325 ( .A1(\adder_stage1[8][10] ), .A2(\adder_stage1[9][10] ), 
        .ZN(n7640) );
  OAI21_X1 U7326 ( .B1(n7637), .B2(n7639), .A(n7640), .ZN(n5979) );
  INV_X1 U7327 ( .A(n5979), .ZN(n7594) );
  NAND2_X1 U7328 ( .A1(\adder_stage1[8][12] ), .A2(\adder_stage1[9][12] ), 
        .ZN(n7618) );
  NAND2_X1 U7329 ( .A1(\adder_stage1[8][11] ), .A2(\adder_stage1[9][11] ), 
        .ZN(n7615) );
  INV_X1 U7330 ( .A(n7615), .ZN(n5980) );
  NAND2_X1 U7331 ( .A1(n7619), .A2(n5980), .ZN(n5981) );
  AND2_X1 U7332 ( .A1(n7618), .A2(n5981), .ZN(n5982) );
  OAI21_X1 U7333 ( .B1(n7594), .B2(n5983), .A(n5982), .ZN(n5984) );
  AOI21_X1 U7334 ( .B1(n7636), .B2(n5985), .A(n5984), .ZN(n7628) );
  NOR2_X1 U7335 ( .A1(\adder_stage1[8][13] ), .A2(\adder_stage1[9][13] ), .ZN(
        n7624) );
  NAND2_X1 U7336 ( .A1(\adder_stage1[8][13] ), .A2(\adder_stage1[9][13] ), 
        .ZN(n7625) );
  OAI21_X1 U7337 ( .B1(n7628), .B2(n7624), .A(n7625), .ZN(n7537) );
  OR2_X1 U7338 ( .A1(\adder_stage1[8][14] ), .A2(\adder_stage1[9][14] ), .ZN(
        n7535) );
  NAND2_X1 U7339 ( .A1(\adder_stage1[8][14] ), .A2(\adder_stage1[9][14] ), 
        .ZN(n7534) );
  INV_X1 U7340 ( .A(n7534), .ZN(n5986) );
  AOI21_X1 U7341 ( .B1(n7537), .B2(n7535), .A(n5986), .ZN(n5987) );
  INV_X1 U7342 ( .A(n5987), .ZN(n8104) );
  AOI22_X1 U7343 ( .A1(n5988), .A2(n5950), .B1(n7285), .B2(
        \adder_stage2[4][15] ), .ZN(n5989) );
  INV_X1 U7344 ( .A(n5989), .ZN(n9722) );
  AOI22_X1 U7345 ( .A1(\x_mult_f_int[18][11] ), .A2(n8229), .B1(n7775), .B2(
        \x_mult_f[18][11] ), .ZN(n5990) );
  INV_X1 U7346 ( .A(n5990), .ZN(n9158) );
  FA_X1 U7347 ( .A(\x_mult_f[28][14] ), .B(\x_mult_f[29][14] ), .CI(n5991), 
        .CO(n7942), .S(n5992) );
  AOI22_X1 U7348 ( .A1(n5992), .A2(n7774), .B1(n7944), .B2(
        \adder_stage1[14][14] ), .ZN(n5993) );
  INV_X1 U7349 ( .A(n5993), .ZN(n9825) );
  AOI22_X1 U7350 ( .A1(\x_mult_f_int[2][6] ), .A2(n8037), .B1(n7944), .B2(
        \x_mult_f[2][6] ), .ZN(n5994) );
  INV_X1 U7351 ( .A(n5994), .ZN(n8956) );
  AOI22_X1 U7352 ( .A1(n5997), .A2(n8387), .B1(n7944), .B2(
        \adder_stage1[1][14] ), .ZN(n5998) );
  INV_X1 U7353 ( .A(n5998), .ZN(n10039) );
  AOI22_X1 U7354 ( .A1(n8365), .A2(\x_mult_f_int[2][5] ), .B1(n7944), .B2(
        \x_mult_f[2][5] ), .ZN(n5999) );
  INV_X1 U7355 ( .A(n5999), .ZN(n8957) );
  INV_X1 U7356 ( .A(n6001), .ZN(n6003) );
  NAND2_X1 U7357 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  XOR2_X1 U7358 ( .A(n6000), .B(n6004), .Z(n6005) );
  AOI22_X1 U7359 ( .A1(n6005), .A2(n8401), .B1(n7944), .B2(
        \adder_stage1[1][13] ), .ZN(n6006) );
  INV_X1 U7360 ( .A(n6006), .ZN(n10040) );
  AOI21_X1 U7361 ( .B1(n6009), .B2(n6008), .A(n6007), .ZN(n6013) );
  NAND2_X1 U7362 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  XOR2_X1 U7363 ( .A(n6013), .B(n6012), .Z(n6014) );
  AOI22_X1 U7364 ( .A1(n6014), .A2(n8229), .B1(n7944), .B2(
        \adder_stage1[15][13] ), .ZN(n6015) );
  INV_X1 U7365 ( .A(n6015), .ZN(n9809) );
  AOI22_X1 U7366 ( .A1(\x_mult_f_int[29][8] ), .A2(n6643), .B1(n7944), .B2(
        \x_mult_f[29][8] ), .ZN(n6016) );
  INV_X1 U7367 ( .A(n6016), .ZN(n9257) );
  BUF_X2 U7368 ( .A(n6955), .Z(n7992) );
  AOI22_X1 U7369 ( .A1(n8048), .A2(\x_mult_f[15][2] ), .B1(n7992), .B2(
        \x_mult_f_int[15][2] ), .ZN(n6017) );
  INV_X1 U7370 ( .A(n6017), .ZN(n9126) );
  AOI22_X1 U7371 ( .A1(n8212), .A2(\x_mult_f[15][4] ), .B1(n7992), .B2(
        \x_mult_f_int[15][4] ), .ZN(n6018) );
  INV_X1 U7372 ( .A(n6018), .ZN(n9124) );
  OR2_X1 U7373 ( .A1(\adder_stage2[2][0] ), .A2(\adder_stage2[3][0] ), .ZN(
        n6019) );
  AND2_X1 U7374 ( .A1(n6019), .A2(n6052), .ZN(n6020) );
  AOI22_X1 U7375 ( .A1(n5294), .A2(\adder_stage3[1][0] ), .B1(n8310), .B2(
        n6020), .ZN(n6021) );
  INV_X1 U7376 ( .A(n6021), .ZN(n9650) );
  INV_X1 U7377 ( .A(n6022), .ZN(n6025) );
  INV_X1 U7378 ( .A(n6023), .ZN(n6024) );
  OAI21_X1 U7379 ( .B1(n6046), .B2(n6025), .A(n6024), .ZN(n6426) );
  INV_X1 U7380 ( .A(n6026), .ZN(n6424) );
  INV_X1 U7381 ( .A(n6423), .ZN(n6027) );
  AOI21_X1 U7382 ( .B1(n6426), .B2(n6424), .A(n6027), .ZN(n6032) );
  INV_X1 U7383 ( .A(n6028), .ZN(n6030) );
  NAND2_X1 U7384 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  XOR2_X1 U7385 ( .A(n6032), .B(n6031), .Z(n6033) );
  AOI22_X1 U7386 ( .A1(n6428), .A2(\adder_stage3[1][11] ), .B1(n8310), .B2(
        n6033), .ZN(n6034) );
  INV_X1 U7387 ( .A(n6034), .ZN(n9639) );
  OAI21_X1 U7388 ( .B1(n6046), .B2(n6042), .A(n6043), .ZN(n6039) );
  INV_X1 U7389 ( .A(n6035), .ZN(n6037) );
  NAND2_X1 U7390 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  XNOR2_X1 U7391 ( .A(n6039), .B(n6038), .ZN(n6040) );
  AOI22_X1 U7392 ( .A1(n6428), .A2(\adder_stage3[1][9] ), .B1(n8310), .B2(
        n6040), .ZN(n6041) );
  INV_X1 U7393 ( .A(n6041), .ZN(n9641) );
  INV_X1 U7394 ( .A(n6042), .ZN(n6044) );
  NAND2_X1 U7395 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  XOR2_X1 U7396 ( .A(n6046), .B(n6045), .Z(n6047) );
  AOI22_X1 U7397 ( .A1(n6428), .A2(\adder_stage3[1][8] ), .B1(n8310), .B2(
        n6047), .ZN(n6048) );
  INV_X1 U7398 ( .A(n6048), .ZN(n9642) );
  INV_X1 U7399 ( .A(n6049), .ZN(n6051) );
  NAND2_X1 U7400 ( .A1(n6051), .A2(n6050), .ZN(n6053) );
  XOR2_X1 U7401 ( .A(n6053), .B(n6052), .Z(n6054) );
  AOI22_X1 U7402 ( .A1(n8157), .A2(\adder_stage3[1][1] ), .B1(n8310), .B2(
        n6054), .ZN(n6055) );
  INV_X1 U7403 ( .A(n6055), .ZN(n9649) );
  INV_X1 U7404 ( .A(n6056), .ZN(n6420) );
  OAI21_X1 U7405 ( .B1(n6420), .B2(n6416), .A(n6417), .ZN(n6061) );
  INV_X1 U7406 ( .A(n6057), .ZN(n6059) );
  NAND2_X1 U7407 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U7408 ( .A(n6061), .B(n6060), .ZN(n6062) );
  AOI22_X1 U7409 ( .A1(n6428), .A2(\adder_stage3[1][3] ), .B1(n8310), .B2(
        n6062), .ZN(n6063) );
  INV_X1 U7410 ( .A(n6063), .ZN(n9647) );
  NOR2_X1 U7411 ( .A1(\adder_stage1[2][2] ), .A2(\adder_stage1[3][2] ), .ZN(
        n6349) );
  NOR2_X1 U7412 ( .A1(\adder_stage1[2][3] ), .A2(\adder_stage1[3][3] ), .ZN(
        n6160) );
  NOR2_X1 U7413 ( .A1(n6349), .A2(n6160), .ZN(n6065) );
  NOR2_X1 U7414 ( .A1(\adder_stage1[2][1] ), .A2(\adder_stage1[3][1] ), .ZN(
        n6343) );
  NAND2_X1 U7415 ( .A1(\adder_stage1[2][0] ), .A2(\adder_stage1[3][0] ), .ZN(
        n6356) );
  NAND2_X1 U7416 ( .A1(\adder_stage1[2][1] ), .A2(\adder_stage1[3][1] ), .ZN(
        n6344) );
  OAI21_X1 U7417 ( .B1(n6343), .B2(n6356), .A(n6344), .ZN(n6159) );
  NAND2_X1 U7418 ( .A1(\adder_stage1[2][2] ), .A2(\adder_stage1[3][2] ), .ZN(
        n6350) );
  NAND2_X1 U7419 ( .A1(\adder_stage1[2][3] ), .A2(\adder_stage1[3][3] ), .ZN(
        n6161) );
  OAI21_X1 U7420 ( .B1(n6160), .B2(n6350), .A(n6161), .ZN(n6064) );
  AOI21_X1 U7421 ( .B1(n6065), .B2(n6159), .A(n6064), .ZN(n6139) );
  NOR2_X1 U7422 ( .A1(\adder_stage1[2][4] ), .A2(\adder_stage1[3][4] ), .ZN(
        n6140) );
  NOR2_X1 U7423 ( .A1(\adder_stage1[2][5] ), .A2(\adder_stage1[3][5] ), .ZN(
        n6142) );
  NOR2_X1 U7424 ( .A1(n6140), .A2(n6142), .ZN(n6168) );
  NAND2_X1 U7425 ( .A1(n3513), .A2(n3475), .ZN(n6170) );
  INV_X1 U7426 ( .A(n6170), .ZN(n6066) );
  NOR2_X1 U7427 ( .A1(\adder_stage1[2][6] ), .A2(\adder_stage1[3][6] ), .ZN(
        n6198) );
  NOR2_X1 U7428 ( .A1(n6066), .A2(n6198), .ZN(n6068) );
  NAND2_X1 U7429 ( .A1(n6168), .A2(n6068), .ZN(n6070) );
  NAND2_X1 U7430 ( .A1(\adder_stage1[2][4] ), .A2(\adder_stage1[3][4] ), .ZN(
        n6205) );
  NAND2_X1 U7431 ( .A1(\adder_stage1[2][5] ), .A2(\adder_stage1[3][5] ), .ZN(
        n6143) );
  OAI21_X1 U7432 ( .B1(n6142), .B2(n6205), .A(n6143), .ZN(n6167) );
  NAND2_X1 U7433 ( .A1(\adder_stage1[2][6] ), .A2(\adder_stage1[3][6] ), .ZN(
        n6199) );
  NAND2_X1 U7434 ( .A1(\adder_stage1[2][7] ), .A2(\adder_stage1[3][7] ), .ZN(
        n6169) );
  OAI21_X1 U7435 ( .B1(n6066), .B2(n6199), .A(n6169), .ZN(n6067) );
  AOI21_X1 U7436 ( .B1(n6068), .B2(n6167), .A(n6067), .ZN(n6069) );
  OAI21_X1 U7437 ( .B1(n6139), .B2(n6070), .A(n6069), .ZN(n6149) );
  NOR2_X1 U7438 ( .A1(\adder_stage1[2][8] ), .A2(\adder_stage1[3][8] ), .ZN(
        n6183) );
  INV_X1 U7439 ( .A(n6183), .ZN(n6175) );
  OR2_X1 U7440 ( .A1(\adder_stage1[2][9] ), .A2(\adder_stage1[3][9] ), .ZN(
        n6186) );
  NAND2_X1 U7441 ( .A1(n6175), .A2(n6186), .ZN(n6151) );
  NOR2_X1 U7442 ( .A1(\adder_stage1[2][10] ), .A2(\adder_stage1[3][10] ), .ZN(
        n6152) );
  NOR2_X1 U7443 ( .A1(n6151), .A2(n6152), .ZN(n6132) );
  OR2_X1 U7444 ( .A1(\adder_stage1[2][11] ), .A2(\adder_stage1[3][11] ), .ZN(
        n6134) );
  OR2_X1 U7445 ( .A1(\adder_stage1[2][12] ), .A2(\adder_stage1[3][12] ), .ZN(
        n6211) );
  OR2_X1 U7446 ( .A1(\adder_stage1[2][13] ), .A2(\adder_stage1[3][13] ), .ZN(
        n6217) );
  NAND2_X1 U7447 ( .A1(n6211), .A2(n6217), .ZN(n6077) );
  NAND2_X1 U7448 ( .A1(\adder_stage1[2][13] ), .A2(\adder_stage1[3][13] ), 
        .ZN(n6216) );
  INV_X1 U7449 ( .A(n6071), .ZN(n6079) );
  NAND2_X1 U7450 ( .A1(\adder_stage1[2][8] ), .A2(\adder_stage1[3][8] ), .ZN(
        n6182) );
  INV_X1 U7451 ( .A(n6182), .ZN(n6073) );
  NAND2_X1 U7452 ( .A1(\adder_stage1[2][9] ), .A2(\adder_stage1[3][9] ), .ZN(
        n6185) );
  INV_X1 U7453 ( .A(n6185), .ZN(n6072) );
  AOI21_X1 U7454 ( .B1(n6186), .B2(n6073), .A(n6072), .ZN(n6150) );
  NAND2_X1 U7455 ( .A1(\adder_stage1[2][10] ), .A2(\adder_stage1[3][10] ), 
        .ZN(n6153) );
  OAI21_X1 U7456 ( .B1(n6150), .B2(n6152), .A(n6153), .ZN(n6131) );
  NAND2_X1 U7457 ( .A1(n6131), .A2(n6134), .ZN(n6124) );
  NAND2_X1 U7458 ( .A1(\adder_stage1[2][11] ), .A2(\adder_stage1[3][11] ), 
        .ZN(n6133) );
  INV_X1 U7459 ( .A(n6133), .ZN(n6075) );
  NAND2_X1 U7460 ( .A1(\adder_stage1[2][12] ), .A2(\adder_stage1[3][12] ), 
        .ZN(n6126) );
  INV_X1 U7461 ( .A(n6126), .ZN(n6074) );
  NOR2_X1 U7462 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  AND2_X1 U7463 ( .A1(n6124), .A2(n6076), .ZN(n6214) );
  OR2_X1 U7464 ( .A1(n6214), .A2(n6077), .ZN(n6078) );
  NAND2_X1 U7465 ( .A1(n6079), .A2(n6078), .ZN(n6116) );
  OR2_X1 U7466 ( .A1(\adder_stage1[2][14] ), .A2(\adder_stage1[3][14] ), .ZN(
        n6118) );
  NAND2_X1 U7467 ( .A1(\adder_stage1[2][14] ), .A2(\adder_stage1[3][14] ), 
        .ZN(n6117) );
  AOI22_X1 U7468 ( .A1(n6080), .A2(n7992), .B1(n8395), .B2(
        \adder_stage2[1][15] ), .ZN(n6081) );
  INV_X1 U7469 ( .A(n6081), .ZN(n9773) );
  INV_X2 U7470 ( .A(n6711), .ZN(n8400) );
  AOI22_X1 U7471 ( .A1(n8363), .A2(\x_mult_f_int[26][5] ), .B1(n8400), .B2(
        \x_mult_f[26][5] ), .ZN(n8835) );
  AOI22_X1 U7472 ( .A1(n8399), .A2(\x_mult_f_int[24][5] ), .B1(n8400), .B2(
        \x_mult_f[24][5] ), .ZN(n8822) );
  AOI22_X1 U7473 ( .A1(\x_mult_f_int[24][7] ), .A2(n8213), .B1(n8400), .B2(
        \x_mult_f[24][7] ), .ZN(n8821) );
  AOI22_X1 U7474 ( .A1(n8180), .A2(\x_mult_f_int[0][5] ), .B1(n8400), .B2(
        \x_mult_f[0][5] ), .ZN(n8785) );
  FA_X1 U7475 ( .A(\x_mult_f[4][14] ), .B(\x_mult_f[5][14] ), .CI(n6082), .CO(
        n7966), .S(n6083) );
  AOI22_X1 U7476 ( .A1(n6083), .A2(n8229), .B1(n8400), .B2(
        \adder_stage1[2][14] ), .ZN(n8792) );
  AOI22_X1 U7477 ( .A1(\x_mult_f_int[27][8] ), .A2(n8114), .B1(n8400), .B2(
        \x_mult_f[27][8] ), .ZN(n8836) );
  NAND2_X1 U7478 ( .A1(n3507), .A2(n6086), .ZN(n6087) );
  XOR2_X1 U7479 ( .A(n6088), .B(n6087), .Z(n6089) );
  AOI22_X1 U7480 ( .A1(n6089), .A2(n5950), .B1(n8094), .B2(
        \adder_stage1[11][13] ), .ZN(n6090) );
  INV_X1 U7481 ( .A(n6090), .ZN(n9877) );
  AOI22_X1 U7482 ( .A1(\x_mult_f_int[19][6] ), .A2(n5950), .B1(n8395), .B2(
        \x_mult_f[19][6] ), .ZN(n6091) );
  INV_X1 U7483 ( .A(n6091), .ZN(n9177) );
  AOI22_X1 U7484 ( .A1(\x_mult_f_int[19][10] ), .A2(n7992), .B1(n8392), .B2(
        \x_mult_f[19][10] ), .ZN(n6092) );
  INV_X1 U7485 ( .A(n6092), .ZN(n9173) );
  AOI22_X1 U7486 ( .A1(\x_mult_f_int[19][8] ), .A2(n7774), .B1(n8392), .B2(
        \x_mult_f[19][8] ), .ZN(n6093) );
  INV_X1 U7487 ( .A(n6093), .ZN(n9175) );
  FA_X1 U7488 ( .A(\x_mult_f[18][14] ), .B(\x_mult_f[19][14] ), .CI(n6094), 
        .CO(n8016), .S(n6095) );
  AOI22_X1 U7489 ( .A1(n6095), .A2(n7284), .B1(n8392), .B2(
        \adder_stage1[9][14] ), .ZN(n6096) );
  INV_X1 U7490 ( .A(n6096), .ZN(n9907) );
  AOI22_X1 U7491 ( .A1(\x_mult_f_int[19][9] ), .A2(n7029), .B1(n8397), .B2(
        \x_mult_f[19][9] ), .ZN(n6097) );
  INV_X1 U7492 ( .A(n6097), .ZN(n9174) );
  AOI22_X1 U7493 ( .A1(\x_mult_f_int[19][11] ), .A2(n8363), .B1(n8157), .B2(
        \x_mult_f[19][11] ), .ZN(n6098) );
  INV_X1 U7494 ( .A(n6098), .ZN(n9172) );
  NAND2_X1 U7495 ( .A1(n3503), .A2(n6100), .ZN(n6101) );
  XOR2_X1 U7496 ( .A(n6102), .B(n6101), .Z(n6103) );
  AOI22_X1 U7497 ( .A1(n6103), .A2(n7992), .B1(n8195), .B2(
        \adder_stage1[9][13] ), .ZN(n6104) );
  INV_X1 U7498 ( .A(n6104), .ZN(n9908) );
  INV_X2 U7499 ( .A(n6105), .ZN(n8154) );
  AOI22_X1 U7500 ( .A1(\x_mult_f_int[2][7] ), .A2(n8037), .B1(n8154), .B2(
        \x_mult_f[2][7] ), .ZN(n6106) );
  INV_X1 U7501 ( .A(n6106), .ZN(n8955) );
  AOI22_X1 U7502 ( .A1(\x_mult_f_int[2][8] ), .A2(n8037), .B1(n8154), .B2(
        \x_mult_f[2][8] ), .ZN(n6107) );
  INV_X1 U7503 ( .A(n6107), .ZN(n8954) );
  AOI22_X1 U7504 ( .A1(\x_mult_f_int[2][10] ), .A2(n8037), .B1(n8154), .B2(
        \x_mult_f[2][10] ), .ZN(n6108) );
  INV_X1 U7505 ( .A(n6108), .ZN(n8952) );
  AOI22_X1 U7506 ( .A1(\x_mult_f_int[2][9] ), .A2(n8037), .B1(n8154), .B2(
        \x_mult_f[2][9] ), .ZN(n6109) );
  INV_X1 U7507 ( .A(n6109), .ZN(n8953) );
  AOI22_X1 U7508 ( .A1(\x_mult_f_int[2][11] ), .A2(n8229), .B1(n8154), .B2(
        \x_mult_f[2][11] ), .ZN(n6110) );
  INV_X1 U7509 ( .A(n6110), .ZN(n8951) );
  AOI22_X1 U7510 ( .A1(\x_mult_f_int[29][11] ), .A2(n8150), .B1(n8154), .B2(
        \x_mult_f[29][11] ), .ZN(n6111) );
  INV_X1 U7511 ( .A(n6111), .ZN(n9254) );
  AOI22_X1 U7512 ( .A1(\x_mult_f_int[29][10] ), .A2(n5908), .B1(n8154), .B2(
        \x_mult_f[29][10] ), .ZN(n6112) );
  INV_X1 U7513 ( .A(n6112), .ZN(n9255) );
  AOI22_X1 U7514 ( .A1(\x_mult_f_int[29][9] ), .A2(n7774), .B1(n8154), .B2(
        \x_mult_f[29][9] ), .ZN(n6113) );
  INV_X1 U7515 ( .A(n6113), .ZN(n9256) );
  AOI22_X1 U7516 ( .A1(\x_mult_f_int[8][8] ), .A2(n8189), .B1(n4713), .B2(
        \x_mult_f[8][8] ), .ZN(n6114) );
  INV_X1 U7517 ( .A(n6114), .ZN(n9034) );
  AOI22_X1 U7518 ( .A1(\x_mult_f_int[8][10] ), .A2(n6643), .B1(n8195), .B2(
        \x_mult_f[8][10] ), .ZN(n6115) );
  INV_X1 U7519 ( .A(n6115), .ZN(n9032) );
  BUF_X1 U7520 ( .A(n3452), .Z(n6122) );
  NAND2_X1 U7521 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  XNOR2_X1 U7522 ( .A(n6116), .B(n6119), .ZN(n6120) );
  AOI22_X1 U7523 ( .A1(n7825), .A2(\adder_stage2[1][14] ), .B1(n6221), .B2(
        n6120), .ZN(n6121) );
  INV_X1 U7524 ( .A(n6121), .ZN(n9774) );
  BUF_X2 U7525 ( .A(n6122), .Z(n6711) );
  INV_X2 U7526 ( .A(n6711), .ZN(n6222) );
  AND2_X1 U7527 ( .A1(n6124), .A2(n6133), .ZN(n6125) );
  NAND2_X1 U7528 ( .A1(n6213), .A2(n6125), .ZN(n6128) );
  NAND2_X1 U7529 ( .A1(n6211), .A2(n6126), .ZN(n6127) );
  XNOR2_X1 U7530 ( .A(n6128), .B(n6127), .ZN(n6129) );
  AOI22_X1 U7531 ( .A1(n6222), .A2(\adder_stage2[1][12] ), .B1(n6221), .B2(
        n6129), .ZN(n6130) );
  INV_X1 U7532 ( .A(n6130), .ZN(n9776) );
  AOI21_X1 U7533 ( .B1(n6149), .B2(n6132), .A(n6131), .ZN(n6136) );
  NAND2_X1 U7534 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  XOR2_X1 U7535 ( .A(n6136), .B(n6135), .Z(n6137) );
  AOI22_X1 U7536 ( .A1(n6222), .A2(\adder_stage2[1][11] ), .B1(n6221), .B2(
        n6137), .ZN(n6138) );
  INV_X1 U7537 ( .A(n6138), .ZN(n9777) );
  INV_X1 U7538 ( .A(n6139), .ZN(n6208) );
  INV_X1 U7539 ( .A(n6140), .ZN(n6206) );
  INV_X1 U7540 ( .A(n6205), .ZN(n6141) );
  AOI21_X1 U7541 ( .B1(n6208), .B2(n6206), .A(n6141), .ZN(n6146) );
  INV_X1 U7542 ( .A(n6142), .ZN(n6144) );
  NAND2_X1 U7543 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  XOR2_X1 U7544 ( .A(n6146), .B(n6145), .Z(n6147) );
  AOI22_X1 U7545 ( .A1(n6222), .A2(\adder_stage2[1][5] ), .B1(n6221), .B2(
        n6147), .ZN(n6148) );
  INV_X1 U7546 ( .A(n6148), .ZN(n9783) );
  INV_X1 U7547 ( .A(n6149), .ZN(n6184) );
  OAI21_X1 U7548 ( .B1(n6184), .B2(n6151), .A(n6150), .ZN(n6156) );
  INV_X1 U7549 ( .A(n6152), .ZN(n6154) );
  NAND2_X1 U7550 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  XNOR2_X1 U7551 ( .A(n6156), .B(n6155), .ZN(n6157) );
  AOI22_X1 U7552 ( .A1(n6222), .A2(\adder_stage2[1][10] ), .B1(n6221), .B2(
        n6157), .ZN(n6158) );
  INV_X1 U7553 ( .A(n6158), .ZN(n9778) );
  INV_X1 U7554 ( .A(n6159), .ZN(n6353) );
  OAI21_X1 U7555 ( .B1(n6353), .B2(n6349), .A(n6350), .ZN(n6164) );
  INV_X1 U7556 ( .A(n6160), .ZN(n6162) );
  NAND2_X1 U7557 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  XNOR2_X1 U7558 ( .A(n6164), .B(n6163), .ZN(n6165) );
  AOI22_X1 U7559 ( .A1(n6222), .A2(\adder_stage2[1][3] ), .B1(n6221), .B2(
        n6165), .ZN(n6166) );
  INV_X1 U7560 ( .A(n6166), .ZN(n9785) );
  AOI21_X1 U7561 ( .B1(n6208), .B2(n6168), .A(n6167), .ZN(n6202) );
  OAI21_X1 U7562 ( .B1(n6202), .B2(n6198), .A(n6199), .ZN(n6172) );
  NAND2_X1 U7563 ( .A1(n6170), .A2(n6169), .ZN(n6171) );
  XNOR2_X1 U7564 ( .A(n6172), .B(n6171), .ZN(n6173) );
  AOI22_X1 U7565 ( .A1(n6222), .A2(\adder_stage2[1][7] ), .B1(n6221), .B2(
        n6173), .ZN(n6174) );
  INV_X1 U7566 ( .A(n6174), .ZN(n9781) );
  NAND2_X1 U7567 ( .A1(n6175), .A2(n6182), .ZN(n6176) );
  XOR2_X1 U7568 ( .A(n6184), .B(n6176), .Z(n6177) );
  AOI22_X1 U7569 ( .A1(n6222), .A2(\adder_stage2[1][8] ), .B1(n6221), .B2(
        n6177), .ZN(n6178) );
  INV_X1 U7570 ( .A(n6178), .ZN(n9780) );
  OR2_X1 U7571 ( .A1(\x_mult_f[6][0] ), .A2(\x_mult_f[7][0] ), .ZN(n6179) );
  AND2_X1 U7572 ( .A1(n6179), .A2(n6194), .ZN(n6180) );
  AOI22_X1 U7573 ( .A1(n6222), .A2(\adder_stage1[3][0] ), .B1(n6221), .B2(
        n6180), .ZN(n6181) );
  INV_X1 U7574 ( .A(n6181), .ZN(n10020) );
  OAI21_X1 U7575 ( .B1(n6184), .B2(n6183), .A(n6182), .ZN(n6188) );
  NAND2_X1 U7576 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  XNOR2_X1 U7577 ( .A(n6188), .B(n6187), .ZN(n6189) );
  AOI22_X1 U7578 ( .A1(n6222), .A2(\adder_stage2[1][9] ), .B1(n6221), .B2(
        n6189), .ZN(n6190) );
  INV_X1 U7579 ( .A(n6190), .ZN(n9779) );
  INV_X1 U7580 ( .A(n6191), .ZN(n6193) );
  NAND2_X1 U7581 ( .A1(n6193), .A2(n6192), .ZN(n6195) );
  XOR2_X1 U7582 ( .A(n6195), .B(n6194), .Z(n6196) );
  AOI22_X1 U7583 ( .A1(n5273), .A2(\adder_stage1[3][1] ), .B1(n6221), .B2(
        n6196), .ZN(n6197) );
  INV_X1 U7584 ( .A(n6197), .ZN(n10019) );
  INV_X1 U7585 ( .A(n6198), .ZN(n6200) );
  NAND2_X1 U7586 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  XOR2_X1 U7587 ( .A(n6202), .B(n6201), .Z(n6203) );
  AOI22_X1 U7588 ( .A1(n6222), .A2(\adder_stage2[1][6] ), .B1(n6221), .B2(
        n6203), .ZN(n6204) );
  INV_X1 U7589 ( .A(n6204), .ZN(n9782) );
  NAND2_X1 U7590 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  XNOR2_X1 U7591 ( .A(n6208), .B(n6207), .ZN(n6209) );
  AOI22_X1 U7592 ( .A1(n6222), .A2(\adder_stage2[1][4] ), .B1(n6221), .B2(
        n6209), .ZN(n6210) );
  INV_X1 U7593 ( .A(n6210), .ZN(n9784) );
  INV_X1 U7594 ( .A(n6211), .ZN(n6212) );
  AOI21_X1 U7595 ( .B1(n6214), .B2(n6213), .A(n6212), .ZN(n6215) );
  INV_X1 U7596 ( .A(n6215), .ZN(n6219) );
  NAND2_X1 U7597 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  XOR2_X1 U7598 ( .A(n6219), .B(n6218), .Z(n6220) );
  AOI22_X1 U7599 ( .A1(n6222), .A2(\adder_stage2[1][13] ), .B1(n6221), .B2(
        n6220), .ZN(n6223) );
  INV_X1 U7600 ( .A(n6223), .ZN(n9775) );
  INV_X1 U7601 ( .A(n6224), .ZN(n6225) );
  XOR2_X1 U7602 ( .A(\adder_stage1[15][15] ), .B(\adder_stage1[14][15] ), .Z(
        n6228) );
  AOI22_X1 U7603 ( .A1(n6229), .A2(n8365), .B1(n8215), .B2(
        \adder_stage2[7][15] ), .ZN(n6230) );
  INV_X1 U7604 ( .A(n6230), .ZN(n9671) );
  AOI22_X1 U7605 ( .A1(n7775), .A2(\x_mult_f[17][1] ), .B1(n6523), .B2(
        \x_mult_f_int[17][1] ), .ZN(n6232) );
  INV_X1 U7606 ( .A(n6232), .ZN(n9326) );
  AOI22_X1 U7607 ( .A1(n8195), .A2(\x_mult_f[17][4] ), .B1(n6523), .B2(
        \x_mult_f_int[17][4] ), .ZN(n6233) );
  INV_X1 U7608 ( .A(n6233), .ZN(n9151) );
  AOI22_X1 U7609 ( .A1(n7775), .A2(\x_mult_f[17][0] ), .B1(n6523), .B2(
        \x_mult_f_int[17][0] ), .ZN(n6234) );
  INV_X1 U7610 ( .A(n6234), .ZN(n9327) );
  AOI22_X1 U7611 ( .A1(n7775), .A2(\x_mult_f[17][3] ), .B1(n6523), .B2(
        \x_mult_f_int[17][3] ), .ZN(n6235) );
  INV_X1 U7612 ( .A(n6235), .ZN(n9152) );
  INV_X1 U7613 ( .A(n6236), .ZN(n6249) );
  INV_X1 U7614 ( .A(n6248), .ZN(n6237) );
  NAND2_X1 U7615 ( .A1(n6237), .A2(n6247), .ZN(n6238) );
  XOR2_X1 U7616 ( .A(n6249), .B(n6238), .Z(n6239) );
  AOI22_X1 U7617 ( .A1(n8195), .A2(\adder_stage4[0][2] ), .B1(n6256), .B2(
        n6239), .ZN(n6240) );
  INV_X1 U7618 ( .A(n6240), .ZN(n9586) );
  INV_X1 U7619 ( .A(n6241), .ZN(n6243) );
  NAND2_X1 U7620 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  XOR2_X1 U7621 ( .A(n6244), .B(n6505), .Z(n6245) );
  AOI22_X1 U7622 ( .A1(n8195), .A2(\adder_stage4[0][1] ), .B1(n6256), .B2(
        n6245), .ZN(n6246) );
  INV_X1 U7623 ( .A(n6246), .ZN(n9587) );
  OAI21_X1 U7624 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6254) );
  INV_X1 U7625 ( .A(n6250), .ZN(n6252) );
  NAND2_X1 U7626 ( .A1(n6252), .A2(n6251), .ZN(n6253) );
  XNOR2_X1 U7627 ( .A(n6254), .B(n6253), .ZN(n6255) );
  AOI22_X1 U7628 ( .A1(n8195), .A2(\adder_stage4[0][3] ), .B1(n6256), .B2(
        n6255), .ZN(n6257) );
  INV_X1 U7629 ( .A(n6257), .ZN(n9585) );
  AOI22_X1 U7630 ( .A1(\x_mult_f_int[1][10] ), .A2(n4002), .B1(n8397), .B2(
        \x_mult_f[1][10] ), .ZN(n6258) );
  INV_X1 U7631 ( .A(n6258), .ZN(n8940) );
  AOI22_X1 U7632 ( .A1(\x_mult_f_int[25][8] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][8] ), .ZN(n8826) );
  AOI22_X1 U7633 ( .A1(\x_mult_f_int[25][10] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][10] ), .ZN(n8824) );
  AOI22_X1 U7634 ( .A1(\x_mult_f_int[26][8] ), .A2(n4002), .B1(n8397), .B2(
        \x_mult_f[26][8] ), .ZN(n8833) );
  AOI22_X1 U7635 ( .A1(\x_mult_f_int[1][9] ), .A2(n7117), .B1(n8397), .B2(
        \x_mult_f[1][9] ), .ZN(n6259) );
  INV_X1 U7636 ( .A(n6259), .ZN(n8941) );
  AOI22_X1 U7637 ( .A1(\x_mult_f_int[25][6] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][6] ), .ZN(n8828) );
  AOI22_X1 U7638 ( .A1(\x_mult_f_int[25][11] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][11] ), .ZN(n8823) );
  AOI22_X1 U7639 ( .A1(\x_mult_f_int[25][9] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][9] ), .ZN(n8825) );
  AOI22_X1 U7640 ( .A1(\x_mult_f_int[1][8] ), .A2(n7029), .B1(n8397), .B2(
        \x_mult_f[1][8] ), .ZN(n8788) );
  INV_X1 U7641 ( .A(n6260), .ZN(n6304) );
  OAI21_X1 U7642 ( .B1(n6304), .B2(n6300), .A(n6301), .ZN(n6265) );
  INV_X1 U7643 ( .A(n6261), .ZN(n6263) );
  NAND2_X1 U7644 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  XNOR2_X1 U7645 ( .A(n6265), .B(n6264), .ZN(n6266) );
  AOI22_X1 U7646 ( .A1(n8383), .A2(\adder_stage1[5][3] ), .B1(n8194), .B2(
        n6266), .ZN(n6267) );
  INV_X1 U7647 ( .A(n6267), .ZN(n9986) );
  INV_X1 U7648 ( .A(n6268), .ZN(n6297) );
  INV_X1 U7649 ( .A(n6269), .ZN(n6295) );
  INV_X1 U7650 ( .A(n6294), .ZN(n6270) );
  AOI21_X1 U7651 ( .B1(n6297), .B2(n6295), .A(n6270), .ZN(n6275) );
  INV_X1 U7652 ( .A(n6271), .ZN(n6273) );
  NAND2_X1 U7653 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  XOR2_X1 U7654 ( .A(n6275), .B(n6274), .Z(n6276) );
  AOI22_X1 U7655 ( .A1(n6222), .A2(\adder_stage1[5][5] ), .B1(n8194), .B2(
        n6276), .ZN(n6277) );
  INV_X1 U7656 ( .A(n6277), .ZN(n9984) );
  AOI21_X1 U7657 ( .B1(n6297), .B2(n6279), .A(n6278), .ZN(n6286) );
  INV_X1 U7658 ( .A(n6285), .ZN(n6280) );
  NAND2_X1 U7659 ( .A1(n6280), .A2(n6284), .ZN(n6281) );
  XOR2_X1 U7660 ( .A(n6286), .B(n6281), .Z(n6282) );
  AOI22_X1 U7661 ( .A1(n7818), .A2(\adder_stage1[5][6] ), .B1(n8194), .B2(
        n6282), .ZN(n6283) );
  INV_X1 U7662 ( .A(n6283), .ZN(n9983) );
  OAI21_X1 U7663 ( .B1(n6286), .B2(n6285), .A(n6284), .ZN(n6291) );
  INV_X1 U7664 ( .A(n6287), .ZN(n6289) );
  NAND2_X1 U7665 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  XNOR2_X1 U7666 ( .A(n6291), .B(n6290), .ZN(n6292) );
  AOI22_X1 U7667 ( .A1(n8400), .A2(\adder_stage1[5][7] ), .B1(n8194), .B2(
        n6292), .ZN(n6293) );
  INV_X1 U7668 ( .A(n6293), .ZN(n9982) );
  NAND2_X1 U7669 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U7670 ( .A(n6297), .B(n6296), .ZN(n6298) );
  AOI22_X1 U7671 ( .A1(n7330), .A2(\adder_stage1[5][4] ), .B1(n8194), .B2(
        n6298), .ZN(n6299) );
  INV_X1 U7672 ( .A(n6299), .ZN(n9985) );
  INV_X1 U7673 ( .A(n6300), .ZN(n6302) );
  NAND2_X1 U7674 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  XOR2_X1 U7675 ( .A(n6304), .B(n6303), .Z(n6305) );
  AOI22_X1 U7676 ( .A1(n6581), .A2(\adder_stage1[5][2] ), .B1(n8194), .B2(
        n6305), .ZN(n6306) );
  INV_X1 U7677 ( .A(n6306), .ZN(n9987) );
  NAND2_X1 U7678 ( .A1(n6592), .A2(n6307), .ZN(n6308) );
  XNOR2_X1 U7679 ( .A(n7120), .B(n6308), .ZN(n6309) );
  AOI22_X1 U7680 ( .A1(n8383), .A2(\adder_stage1[5][8] ), .B1(n8194), .B2(
        n6309), .ZN(n6310) );
  INV_X1 U7681 ( .A(n6310), .ZN(n9981) );
  INV_X1 U7682 ( .A(n6311), .ZN(n6313) );
  NAND2_X1 U7683 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  XOR2_X1 U7684 ( .A(n6314), .B(n6323), .Z(n6315) );
  AOI22_X1 U7685 ( .A1(n6428), .A2(\adder_stage1[5][1] ), .B1(n8194), .B2(
        n6315), .ZN(n6316) );
  INV_X1 U7686 ( .A(n6316), .ZN(n9988) );
  INV_X1 U7687 ( .A(n6317), .ZN(n6319) );
  NAND2_X1 U7688 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  XOR2_X1 U7689 ( .A(n6320), .B(n6327), .Z(n6321) );
  AOI22_X1 U7690 ( .A1(n6330), .A2(\adder_stage2[7][1] ), .B1(n8194), .B2(
        n6321), .ZN(n6322) );
  INV_X1 U7691 ( .A(n6322), .ZN(n9685) );
  OR2_X1 U7692 ( .A1(\x_mult_f[10][0] ), .A2(\x_mult_f[11][0] ), .ZN(n6324) );
  AND2_X1 U7693 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  AOI22_X1 U7694 ( .A1(n5909), .A2(\adder_stage1[5][0] ), .B1(n8194), .B2(
        n6325), .ZN(n6326) );
  INV_X1 U7695 ( .A(n6326), .ZN(n9989) );
  OR2_X1 U7696 ( .A1(\adder_stage1[14][0] ), .A2(\adder_stage1[15][0] ), .ZN(
        n6328) );
  AND2_X1 U7697 ( .A1(n6328), .A2(n6327), .ZN(n6329) );
  AOI22_X1 U7698 ( .A1(n6330), .A2(\adder_stage2[7][0] ), .B1(n8194), .B2(
        n6329), .ZN(n6331) );
  INV_X1 U7699 ( .A(n6331), .ZN(n9686) );
  INV_X1 U7700 ( .A(n6332), .ZN(n6334) );
  NAND2_X1 U7701 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  XOR2_X1 U7702 ( .A(n6339), .B(n6335), .Z(n6336) );
  AOI22_X1 U7703 ( .A1(n6337), .A2(\adder_stage2[5][1] ), .B1(n8194), .B2(
        n6336), .ZN(n6338) );
  INV_X1 U7704 ( .A(n6338), .ZN(n9719) );
  OR2_X1 U7705 ( .A1(\adder_stage1[10][0] ), .A2(\adder_stage1[11][0] ), .ZN(
        n6340) );
  AND2_X1 U7706 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  AOI22_X1 U7707 ( .A1(n8200), .A2(\adder_stage2[5][0] ), .B1(n8194), .B2(
        n6341), .ZN(n6342) );
  INV_X1 U7708 ( .A(n6342), .ZN(n9720) );
  INV_X1 U7709 ( .A(n6343), .ZN(n6345) );
  NAND2_X1 U7710 ( .A1(n6345), .A2(n6344), .ZN(n6346) );
  XOR2_X1 U7711 ( .A(n6346), .B(n6356), .Z(n6347) );
  AOI22_X1 U7712 ( .A1(n8330), .A2(\adder_stage2[1][1] ), .B1(n8291), .B2(
        n6347), .ZN(n6348) );
  INV_X1 U7713 ( .A(n6348), .ZN(n9787) );
  INV_X1 U7714 ( .A(n6349), .ZN(n6351) );
  NAND2_X1 U7715 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  XOR2_X1 U7716 ( .A(n6353), .B(n6352), .Z(n6354) );
  AOI22_X1 U7717 ( .A1(n7443), .A2(\adder_stage2[1][2] ), .B1(n8291), .B2(
        n6354), .ZN(n6355) );
  INV_X1 U7718 ( .A(n6355), .ZN(n9786) );
  OR2_X1 U7719 ( .A1(\adder_stage1[2][0] ), .A2(\adder_stage1[3][0] ), .ZN(
        n6357) );
  AND2_X1 U7720 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  AOI22_X1 U7721 ( .A1(n8330), .A2(\adder_stage2[1][0] ), .B1(n8291), .B2(
        n6358), .ZN(n6359) );
  INV_X1 U7722 ( .A(n6359), .ZN(n9788) );
  INV_X1 U7723 ( .A(n6430), .ZN(n6362) );
  NAND3_X1 U7724 ( .A1(n6432), .A2(\ctrl_inst/state [1]), .A3(n6360), .ZN(
        n6361) );
  OAI211_X1 U7725 ( .C1(n6362), .C2(n8696), .A(n6361), .B(n8347), .ZN(n3386)
         );
  OR2_X1 U7726 ( .A1(\adder_stage2[0][0] ), .A2(\adder_stage2[1][0] ), .ZN(
        n6363) );
  AND2_X1 U7727 ( .A1(n6363), .A2(n6912), .ZN(n6364) );
  AOI22_X1 U7728 ( .A1(n7244), .A2(\adder_stage3[0][0] ), .B1(n6915), .B2(
        n6364), .ZN(n6365) );
  INV_X1 U7729 ( .A(n6365), .ZN(n9669) );
  INV_X2 U7730 ( .A(n6105), .ZN(n7285) );
  AOI22_X1 U7731 ( .A1(n7285), .A2(\x_mult_f[9][2] ), .B1(n6915), .B2(
        \x_mult_f_int[9][2] ), .ZN(n6366) );
  INV_X1 U7732 ( .A(n6366), .ZN(n9045) );
  AOI22_X1 U7733 ( .A1(n7285), .A2(\x_mult_f[9][4] ), .B1(n6915), .B2(
        \x_mult_f_int[9][4] ), .ZN(n6367) );
  INV_X1 U7734 ( .A(n6367), .ZN(n9043) );
  INV_X2 U7735 ( .A(n6368), .ZN(n6373) );
  AOI22_X1 U7736 ( .A1(\x_mult_f_int[28][6] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][6] ), .ZN(n8844) );
  AOI22_X1 U7737 ( .A1(\x_mult_f_int[2][12] ), .A2(n8229), .B1(n6373), .B2(
        \x_mult_f[2][12] ), .ZN(n6369) );
  INV_X1 U7738 ( .A(n6369), .ZN(n8950) );
  AOI22_X1 U7739 ( .A1(\x_mult_f_int[28][10] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][10] ), .ZN(n8840) );
  AOI22_X1 U7740 ( .A1(\x_mult_f_int[28][12] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][12] ), .ZN(n8838) );
  AOI22_X1 U7741 ( .A1(\x_mult_f_int[2][14] ), .A2(n8229), .B1(n6373), .B2(
        \x_mult_f[2][14] ), .ZN(n6370) );
  INV_X1 U7742 ( .A(n6370), .ZN(n8948) );
  AOI22_X1 U7743 ( .A1(\x_mult_f_int[28][7] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][7] ), .ZN(n8843) );
  AOI22_X1 U7744 ( .A1(\x_mult_f_int[28][8] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][8] ), .ZN(n8842) );
  AOI22_X1 U7745 ( .A1(n8180), .A2(\x_mult_f_int[28][5] ), .B1(n6373), .B2(
        \x_mult_f[28][5] ), .ZN(n6371) );
  INV_X1 U7746 ( .A(n6371), .ZN(n9249) );
  AOI22_X1 U7747 ( .A1(\x_mult_f_int[2][13] ), .A2(n8229), .B1(n6373), .B2(
        \x_mult_f[2][13] ), .ZN(n6372) );
  INV_X1 U7748 ( .A(n6372), .ZN(n8949) );
  AOI22_X1 U7749 ( .A1(\x_mult_f_int[28][11] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][11] ), .ZN(n8839) );
  AOI22_X1 U7750 ( .A1(\x_mult_f_int[28][13] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][13] ), .ZN(n8837) );
  AOI22_X1 U7751 ( .A1(\x_mult_f_int[28][9] ), .A2(n8387), .B1(n6373), .B2(
        \x_mult_f[28][9] ), .ZN(n8841) );
  OAI21_X1 U7752 ( .B1(n6376), .B2(n6375), .A(n6374), .ZN(n6381) );
  INV_X1 U7753 ( .A(n6377), .ZN(n6379) );
  NAND2_X1 U7754 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  XNOR2_X1 U7755 ( .A(n6381), .B(n6380), .ZN(n6382) );
  AOI22_X1 U7756 ( .A1(n8059), .A2(\adder_stage1[10][7] ), .B1(n8310), .B2(
        n6382), .ZN(n6383) );
  INV_X1 U7757 ( .A(n6383), .ZN(n9898) );
  INV_X1 U7758 ( .A(n6384), .ZN(n6406) );
  INV_X1 U7759 ( .A(n6385), .ZN(n6404) );
  INV_X1 U7760 ( .A(n6403), .ZN(n6386) );
  AOI21_X1 U7761 ( .B1(n6406), .B2(n6404), .A(n6386), .ZN(n6391) );
  INV_X1 U7762 ( .A(n6387), .ZN(n6389) );
  NAND2_X1 U7763 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  XOR2_X1 U7764 ( .A(n6391), .B(n6390), .Z(n6392) );
  AOI22_X1 U7765 ( .A1(n6428), .A2(\adder_stage3[1][5] ), .B1(n8310), .B2(
        n6392), .ZN(n6393) );
  INV_X1 U7766 ( .A(n6393), .ZN(n9645) );
  AOI21_X1 U7767 ( .B1(n6406), .B2(n6395), .A(n6394), .ZN(n6413) );
  OAI21_X1 U7768 ( .B1(n6413), .B2(n6409), .A(n6410), .ZN(n6400) );
  INV_X1 U7769 ( .A(n6396), .ZN(n6398) );
  NAND2_X1 U7770 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  XNOR2_X1 U7771 ( .A(n6400), .B(n6399), .ZN(n6401) );
  AOI22_X1 U7772 ( .A1(n6428), .A2(\adder_stage3[1][7] ), .B1(n8310), .B2(
        n6401), .ZN(n6402) );
  INV_X1 U7773 ( .A(n6402), .ZN(n9643) );
  NAND2_X1 U7774 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  XNOR2_X1 U7775 ( .A(n6406), .B(n6405), .ZN(n6407) );
  AOI22_X1 U7776 ( .A1(n6428), .A2(\adder_stage3[1][4] ), .B1(n8310), .B2(
        n6407), .ZN(n6408) );
  INV_X1 U7777 ( .A(n6408), .ZN(n9646) );
  INV_X1 U7778 ( .A(n6409), .ZN(n6411) );
  NAND2_X1 U7779 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  XOR2_X1 U7780 ( .A(n6413), .B(n6412), .Z(n6414) );
  AOI22_X1 U7781 ( .A1(n6428), .A2(\adder_stage3[1][6] ), .B1(n8310), .B2(
        n6414), .ZN(n6415) );
  INV_X1 U7782 ( .A(n6415), .ZN(n9644) );
  INV_X1 U7783 ( .A(n6416), .ZN(n6418) );
  NAND2_X1 U7784 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  XOR2_X1 U7785 ( .A(n6420), .B(n6419), .Z(n6421) );
  AOI22_X1 U7786 ( .A1(n6428), .A2(\adder_stage3[1][2] ), .B1(n8310), .B2(
        n6421), .ZN(n6422) );
  INV_X1 U7787 ( .A(n6422), .ZN(n9648) );
  NAND2_X1 U7788 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  XNOR2_X1 U7789 ( .A(n6426), .B(n6425), .ZN(n6427) );
  AOI22_X1 U7790 ( .A1(n6428), .A2(\adder_stage3[1][10] ), .B1(n8310), .B2(
        n6427), .ZN(n6429) );
  INV_X1 U7791 ( .A(n6429), .ZN(n9640) );
  AOI22_X1 U7792 ( .A1(n6432), .A2(n6431), .B1(\ctrl_inst/state [0]), .B2(
        n6430), .ZN(n6434) );
  NAND2_X1 U7793 ( .A1(n6434), .A2(n6433), .ZN(n3388) );
  BUF_X2 U7794 ( .A(n6699), .Z(n7029) );
  INV_X1 U7795 ( .A(n6436), .ZN(n6468) );
  INV_X1 U7796 ( .A(n6437), .ZN(n6467) );
  NAND2_X1 U7797 ( .A1(n6467), .A2(n6465), .ZN(n6438) );
  XNOR2_X1 U7798 ( .A(n6468), .B(n6438), .ZN(n6439) );
  AOI22_X1 U7799 ( .A1(n8330), .A2(\adder_stage2[0][4] ), .B1(n7029), .B2(
        n6439), .ZN(n6440) );
  INV_X1 U7800 ( .A(n6440), .ZN(n9801) );
  INV_X2 U7801 ( .A(n4526), .ZN(n7030) );
  AOI21_X1 U7802 ( .B1(n6468), .B2(n6442), .A(n6441), .ZN(n6462) );
  OAI21_X1 U7803 ( .B1(n6462), .B2(n6458), .A(n6459), .ZN(n6447) );
  INV_X1 U7804 ( .A(n6443), .ZN(n6445) );
  NAND2_X1 U7805 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  XNOR2_X1 U7806 ( .A(n6447), .B(n6446), .ZN(n6448) );
  AOI22_X1 U7807 ( .A1(n7030), .A2(\adder_stage2[0][7] ), .B1(n7029), .B2(
        n6448), .ZN(n6449) );
  INV_X1 U7808 ( .A(n6449), .ZN(n9798) );
  INV_X1 U7809 ( .A(n6450), .ZN(n6483) );
  OAI21_X1 U7810 ( .B1(n6483), .B2(n6479), .A(n6480), .ZN(n6455) );
  INV_X1 U7811 ( .A(n6451), .ZN(n6453) );
  NAND2_X1 U7812 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  XNOR2_X1 U7813 ( .A(n6455), .B(n6454), .ZN(n6456) );
  AOI22_X1 U7814 ( .A1(n7443), .A2(\adder_stage2[0][3] ), .B1(n7029), .B2(
        n6456), .ZN(n6457) );
  INV_X1 U7815 ( .A(n6457), .ZN(n9802) );
  INV_X1 U7816 ( .A(n6458), .ZN(n6460) );
  NAND2_X1 U7817 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  XOR2_X1 U7818 ( .A(n6462), .B(n6461), .Z(n6463) );
  AOI22_X1 U7819 ( .A1(n6222), .A2(\adder_stage2[0][6] ), .B1(n7029), .B2(
        n6463), .ZN(n6464) );
  INV_X1 U7820 ( .A(n6464), .ZN(n9799) );
  INV_X1 U7821 ( .A(n6465), .ZN(n6466) );
  AOI21_X1 U7822 ( .B1(n6468), .B2(n6467), .A(n6466), .ZN(n6473) );
  INV_X1 U7823 ( .A(n6469), .ZN(n6471) );
  NAND2_X1 U7824 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  XOR2_X1 U7825 ( .A(n6473), .B(n6472), .Z(n6474) );
  AOI22_X1 U7826 ( .A1(n7818), .A2(\adder_stage2[0][5] ), .B1(n7029), .B2(
        n6474), .ZN(n6475) );
  INV_X1 U7827 ( .A(n6475), .ZN(n9800) );
  OR2_X1 U7828 ( .A1(\adder_stage1[0][0] ), .A2(\adder_stage1[1][0] ), .ZN(
        n6476) );
  AND2_X1 U7829 ( .A1(n6476), .A2(n6489), .ZN(n6477) );
  AOI22_X1 U7830 ( .A1(n7330), .A2(\adder_stage2[0][0] ), .B1(n7029), .B2(
        n6477), .ZN(n6478) );
  INV_X1 U7831 ( .A(n6478), .ZN(n9805) );
  INV_X1 U7832 ( .A(n6479), .ZN(n6481) );
  NAND2_X1 U7833 ( .A1(n6481), .A2(n6480), .ZN(n6482) );
  XOR2_X1 U7834 ( .A(n6483), .B(n6482), .Z(n6484) );
  AOI22_X1 U7835 ( .A1(n6337), .A2(\adder_stage2[0][2] ), .B1(n7029), .B2(
        n6484), .ZN(n6485) );
  INV_X1 U7836 ( .A(n6485), .ZN(n9803) );
  INV_X1 U7837 ( .A(n6486), .ZN(n6488) );
  NAND2_X1 U7838 ( .A1(n6488), .A2(n6487), .ZN(n6490) );
  XOR2_X1 U7839 ( .A(n6490), .B(n6489), .Z(n6491) );
  AOI22_X1 U7840 ( .A1(n7244), .A2(\adder_stage2[0][1] ), .B1(n7029), .B2(
        n6491), .ZN(n6492) );
  INV_X1 U7841 ( .A(n6492), .ZN(n9804) );
  AOI22_X1 U7842 ( .A1(n8195), .A2(\x_mult_f[16][0] ), .B1(n6523), .B2(
        \x_mult_f_int[16][0] ), .ZN(n6493) );
  INV_X1 U7843 ( .A(n6493), .ZN(n9325) );
  AOI22_X1 U7844 ( .A1(n8195), .A2(\x_mult_f[16][2] ), .B1(n6523), .B2(
        \x_mult_f_int[16][2] ), .ZN(n6494) );
  INV_X1 U7845 ( .A(n6494), .ZN(n9139) );
  AOI22_X1 U7846 ( .A1(n8195), .A2(\x_mult_f[16][3] ), .B1(n6523), .B2(
        \x_mult_f_int[16][3] ), .ZN(n8806) );
  AOI22_X1 U7847 ( .A1(n8195), .A2(\x_mult_f[16][4] ), .B1(n6523), .B2(
        \x_mult_f_int[16][4] ), .ZN(n6495) );
  INV_X1 U7848 ( .A(n6495), .ZN(n9138) );
  AOI22_X1 U7849 ( .A1(n7775), .A2(\x_mult_f[17][2] ), .B1(n6523), .B2(
        \x_mult_f_int[17][2] ), .ZN(n6496) );
  INV_X1 U7850 ( .A(n6496), .ZN(n9153) );
  AOI22_X1 U7851 ( .A1(n8195), .A2(\x_mult_f[16][1] ), .B1(n6523), .B2(
        \x_mult_f_int[16][1] ), .ZN(n6497) );
  INV_X1 U7852 ( .A(n6497), .ZN(n9324) );
  INV_X1 U7853 ( .A(n6498), .ZN(n6500) );
  NAND2_X1 U7854 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  XOR2_X1 U7855 ( .A(n6502), .B(n6501), .Z(n6503) );
  AOI22_X1 U7856 ( .A1(n7775), .A2(\adder_stage1[8][11] ), .B1(n6523), .B2(
        n6503), .ZN(n6504) );
  INV_X1 U7857 ( .A(n6504), .ZN(n9927) );
  OR2_X1 U7858 ( .A1(\adder_stage3[0][0] ), .A2(\adder_stage3[1][0] ), .ZN(
        n6506) );
  AND2_X1 U7859 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  AOI22_X1 U7860 ( .A1(n7443), .A2(\adder_stage4[0][0] ), .B1(n6523), .B2(
        n6507), .ZN(n6508) );
  INV_X1 U7861 ( .A(n6508), .ZN(n9588) );
  NAND2_X1 U7862 ( .A1(n6510), .A2(n6509), .ZN(n6511) );
  XNOR2_X1 U7863 ( .A(n6512), .B(n6511), .ZN(n6513) );
  AOI22_X1 U7864 ( .A1(n7775), .A2(\adder_stage1[8][12] ), .B1(n6523), .B2(
        n6513), .ZN(n6514) );
  INV_X1 U7865 ( .A(n6514), .ZN(n9926) );
  NAND2_X1 U7866 ( .A1(n7772), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U7867 ( .A1(n6517), .A2(n6516), .ZN(n6521) );
  NAND2_X1 U7868 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  XNOR2_X1 U7869 ( .A(n6521), .B(n6520), .ZN(n6522) );
  AOI22_X1 U7870 ( .A1(n7775), .A2(\adder_stage1[8][10] ), .B1(n6523), .B2(
        n6522), .ZN(n6524) );
  INV_X1 U7871 ( .A(n6524), .ZN(n9928) );
  INV_X1 U7872 ( .A(n6537), .ZN(n6525) );
  AOI21_X1 U7873 ( .B1(n6532), .B2(n6538), .A(n6525), .ZN(n6526) );
  NAND2_X1 U7874 ( .A1(n6527), .A2(n6526), .ZN(n6565) );
  NAND2_X1 U7875 ( .A1(n6564), .A2(n6528), .ZN(n6529) );
  XNOR2_X1 U7876 ( .A(n6565), .B(n6529), .ZN(n6530) );
  AOI22_X1 U7877 ( .A1(n6581), .A2(\adder_stage2[3][12] ), .B1(n6643), .B2(
        n6530), .ZN(n6531) );
  INV_X1 U7878 ( .A(n6531), .ZN(n9742) );
  INV_X1 U7879 ( .A(n6532), .ZN(n6536) );
  NAND2_X1 U7880 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  AND2_X1 U7881 ( .A1(n6536), .A2(n6535), .ZN(n6540) );
  NAND2_X1 U7882 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  XOR2_X1 U7883 ( .A(n6540), .B(n6539), .Z(n6541) );
  AOI22_X1 U7884 ( .A1(n6581), .A2(\adder_stage2[3][11] ), .B1(n6643), .B2(
        n6541), .ZN(n6542) );
  INV_X1 U7885 ( .A(n6542), .ZN(n9743) );
  NAND2_X1 U7886 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  XNOR2_X1 U7887 ( .A(n6546), .B(n6545), .ZN(n6547) );
  AOI22_X1 U7888 ( .A1(n6581), .A2(\adder_stage2[3][14] ), .B1(n6643), .B2(
        n6547), .ZN(n6548) );
  INV_X1 U7889 ( .A(n6548), .ZN(n9740) );
  INV_X1 U7890 ( .A(n6549), .ZN(n6551) );
  NAND2_X1 U7891 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  XOR2_X1 U7892 ( .A(n6553), .B(n6552), .Z(n6554) );
  AOI22_X1 U7893 ( .A1(n6581), .A2(\adder_stage1[7][2] ), .B1(n6643), .B2(
        n6554), .ZN(n6555) );
  INV_X1 U7894 ( .A(n6555), .ZN(n9953) );
  AOI21_X1 U7895 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(n6636) );
  INV_X1 U7896 ( .A(n6635), .ZN(n6559) );
  NAND2_X1 U7897 ( .A1(n6559), .A2(n6634), .ZN(n6560) );
  XOR2_X1 U7898 ( .A(n6636), .B(n6560), .Z(n6561) );
  AOI22_X1 U7899 ( .A1(n6581), .A2(\adder_stage1[7][6] ), .B1(n6643), .B2(
        n6561), .ZN(n6562) );
  INV_X1 U7900 ( .A(n6562), .ZN(n9949) );
  AOI21_X1 U7901 ( .B1(n6565), .B2(n6564), .A(n6563), .ZN(n6569) );
  NAND2_X1 U7902 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  XOR2_X1 U7903 ( .A(n6569), .B(n6568), .Z(n6570) );
  AOI22_X1 U7904 ( .A1(n6581), .A2(\adder_stage2[3][13] ), .B1(n6643), .B2(
        n6570), .ZN(n6571) );
  INV_X1 U7905 ( .A(n6571), .ZN(n9741) );
  OAI21_X1 U7906 ( .B1(n6574), .B2(n6573), .A(n6572), .ZN(n6579) );
  INV_X1 U7907 ( .A(n6575), .ZN(n6577) );
  NAND2_X1 U7908 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  XNOR2_X1 U7909 ( .A(n6579), .B(n6578), .ZN(n6580) );
  AOI22_X1 U7910 ( .A1(n6581), .A2(\adder_stage2[3][10] ), .B1(n6643), .B2(
        n6580), .ZN(n6582) );
  INV_X1 U7911 ( .A(n6582), .ZN(n9744) );
  AOI22_X1 U7912 ( .A1(n6222), .A2(\x_mult_f[19][0] ), .B1(n7110), .B2(
        \x_mult_f_int[19][0] ), .ZN(n6583) );
  INV_X1 U7913 ( .A(n6583), .ZN(n9331) );
  AOI22_X1 U7914 ( .A1(n7818), .A2(\x_mult_f[19][1] ), .B1(n7110), .B2(
        \x_mult_f_int[19][1] ), .ZN(n6584) );
  INV_X1 U7915 ( .A(n6584), .ZN(n9330) );
  AOI22_X1 U7916 ( .A1(n7793), .A2(\x_mult_f[11][3] ), .B1(n8389), .B2(
        \x_mult_f_int[11][3] ), .ZN(n6585) );
  INV_X1 U7917 ( .A(n6585), .ZN(n9070) );
  BUF_X2 U7918 ( .A(n6699), .Z(n7117) );
  AOI22_X1 U7919 ( .A1(n7285), .A2(\x_mult_f[3][0] ), .B1(n7117), .B2(
        \x_mult_f_int[3][0] ), .ZN(n6586) );
  INV_X1 U7920 ( .A(n6586), .ZN(n9299) );
  AOI22_X1 U7921 ( .A1(n7793), .A2(\x_mult_f[11][1] ), .B1(n8389), .B2(
        \x_mult_f_int[11][1] ), .ZN(n6587) );
  INV_X1 U7922 ( .A(n6587), .ZN(n9314) );
  AOI22_X1 U7923 ( .A1(n8330), .A2(\x_mult_f[3][2] ), .B1(n7117), .B2(
        \x_mult_f_int[3][2] ), .ZN(n6589) );
  INV_X1 U7924 ( .A(n6589), .ZN(n8973) );
  AOI21_X1 U7925 ( .B1(n7120), .B2(n6592), .A(n6591), .ZN(n6596) );
  NAND2_X1 U7926 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  XOR2_X1 U7927 ( .A(n6596), .B(n6595), .Z(n6597) );
  AOI22_X1 U7928 ( .A1(n7512), .A2(\adder_stage1[5][9] ), .B1(n8389), .B2(
        n6597), .ZN(n6598) );
  INV_X1 U7929 ( .A(n6598), .ZN(n9980) );
  AOI22_X1 U7930 ( .A1(n7793), .A2(\x_mult_f[11][0] ), .B1(n8389), .B2(
        \x_mult_f_int[11][0] ), .ZN(n6599) );
  INV_X1 U7931 ( .A(n6599), .ZN(n9315) );
  INV_X1 U7932 ( .A(n6600), .ZN(n7682) );
  AOI21_X1 U7933 ( .B1(n7682), .B2(n6602), .A(n6601), .ZN(n7061) );
  INV_X1 U7934 ( .A(n7060), .ZN(n6603) );
  NAND2_X1 U7935 ( .A1(n6603), .A2(n7059), .ZN(n6604) );
  XOR2_X1 U7936 ( .A(n7061), .B(n6604), .Z(n6605) );
  AOI22_X1 U7937 ( .A1(n7825), .A2(\adder_stage1[9][6] ), .B1(n7110), .B2(
        n6605), .ZN(n6606) );
  INV_X1 U7938 ( .A(n6606), .ZN(n9915) );
  INV_X1 U7939 ( .A(n6607), .ZN(n6609) );
  NAND2_X1 U7940 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  XOR2_X1 U7941 ( .A(n6611), .B(n6610), .Z(n6612) );
  AOI22_X1 U7942 ( .A1(n5273), .A2(\adder_stage1[9][9] ), .B1(n7110), .B2(
        n6612), .ZN(n6613) );
  INV_X1 U7943 ( .A(n6613), .ZN(n9912) );
  AOI22_X1 U7944 ( .A1(n8391), .A2(\x_mult_f[2][2] ), .B1(n7117), .B2(
        \x_mult_f_int[2][2] ), .ZN(n6614) );
  INV_X1 U7945 ( .A(n6614), .ZN(n8960) );
  AOI22_X1 U7946 ( .A1(n8391), .A2(\x_mult_f[2][3] ), .B1(n7117), .B2(
        \x_mult_f_int[2][3] ), .ZN(n6615) );
  INV_X1 U7947 ( .A(n6615), .ZN(n8959) );
  NAND2_X1 U7948 ( .A1(n6617), .A2(n6616), .ZN(n6618) );
  XNOR2_X1 U7949 ( .A(n6619), .B(n6618), .ZN(n6620) );
  AOI22_X1 U7950 ( .A1(n6337), .A2(\adder_stage1[9][8] ), .B1(n7110), .B2(
        n6620), .ZN(n6621) );
  INV_X1 U7951 ( .A(n6621), .ZN(n9913) );
  AOI22_X1 U7952 ( .A1(n7767), .A2(\x_mult_f[19][4] ), .B1(n7110), .B2(
        \x_mult_f_int[19][4] ), .ZN(n6622) );
  INV_X1 U7953 ( .A(n6622), .ZN(n9179) );
  AOI22_X1 U7954 ( .A1(n7030), .A2(\x_mult_f[19][3] ), .B1(n7110), .B2(
        \x_mult_f_int[19][3] ), .ZN(n6623) );
  INV_X1 U7955 ( .A(n6623), .ZN(n9180) );
  AOI22_X1 U7956 ( .A1(n7793), .A2(\x_mult_f[11][2] ), .B1(n8389), .B2(
        \x_mult_f_int[11][2] ), .ZN(n6624) );
  INV_X1 U7957 ( .A(n6624), .ZN(n9071) );
  AOI22_X1 U7958 ( .A1(n8178), .A2(\x_mult_f[3][4] ), .B1(n7117), .B2(
        \x_mult_f_int[3][4] ), .ZN(n6625) );
  INV_X1 U7959 ( .A(n6625), .ZN(n8971) );
  AOI22_X1 U7960 ( .A1(n6337), .A2(\x_mult_f[3][3] ), .B1(n7117), .B2(
        \x_mult_f_int[3][3] ), .ZN(n6626) );
  INV_X1 U7961 ( .A(n6626), .ZN(n8972) );
  AOI22_X1 U7962 ( .A1(n7285), .A2(\x_mult_f[3][1] ), .B1(n7117), .B2(
        \x_mult_f_int[3][1] ), .ZN(n6627) );
  INV_X1 U7963 ( .A(n6627), .ZN(n9298) );
  NAND2_X1 U7964 ( .A1(n6629), .A2(n6628), .ZN(n6630) );
  XNOR2_X1 U7965 ( .A(n6631), .B(n6630), .ZN(n6632) );
  AOI22_X1 U7966 ( .A1(n7512), .A2(\adder_stage1[7][8] ), .B1(n6643), .B2(
        n6632), .ZN(n6633) );
  INV_X1 U7967 ( .A(n6633), .ZN(n9947) );
  OAI21_X1 U7968 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6641) );
  INV_X1 U7969 ( .A(n6637), .ZN(n6639) );
  NAND2_X1 U7970 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  XNOR2_X1 U7971 ( .A(n6641), .B(n6640), .ZN(n6642) );
  AOI22_X1 U7972 ( .A1(n8036), .A2(\adder_stage1[7][7] ), .B1(n6643), .B2(
        n6642), .ZN(n6644) );
  INV_X1 U7973 ( .A(n6644), .ZN(n9948) );
  INV_X1 U7974 ( .A(n6646), .ZN(n7180) );
  AOI21_X1 U7975 ( .B1(n7180), .B2(n6648), .A(n6647), .ZN(n6677) );
  INV_X1 U7976 ( .A(n6676), .ZN(n6649) );
  NAND2_X1 U7977 ( .A1(n6649), .A2(n6675), .ZN(n6650) );
  XOR2_X1 U7978 ( .A(n6677), .B(n6650), .Z(n6651) );
  AOI22_X1 U7979 ( .A1(n4689), .A2(\adder_stage1[3][6] ), .B1(n7182), .B2(
        n6651), .ZN(n6652) );
  INV_X1 U7980 ( .A(n6652), .ZN(n10014) );
  INV_X1 U7981 ( .A(n6653), .ZN(n7174) );
  OAI21_X1 U7982 ( .B1(n7174), .B2(n7170), .A(n7171), .ZN(n6658) );
  INV_X1 U7983 ( .A(n6654), .ZN(n6656) );
  NAND2_X1 U7984 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  XNOR2_X1 U7985 ( .A(n6658), .B(n6657), .ZN(n6659) );
  AOI22_X1 U7986 ( .A1(n5678), .A2(\adder_stage1[3][3] ), .B1(n7182), .B2(
        n6659), .ZN(n6660) );
  INV_X1 U7987 ( .A(n6660), .ZN(n10017) );
  INV_X1 U7988 ( .A(n6661), .ZN(n7178) );
  INV_X1 U7989 ( .A(n7177), .ZN(n6662) );
  AOI21_X1 U7990 ( .B1(n7180), .B2(n7178), .A(n6662), .ZN(n6667) );
  INV_X1 U7991 ( .A(n6663), .ZN(n6665) );
  NAND2_X1 U7992 ( .A1(n6665), .A2(n6664), .ZN(n6666) );
  XOR2_X1 U7993 ( .A(n6667), .B(n6666), .Z(n6668) );
  AOI22_X1 U7994 ( .A1(n5273), .A2(\adder_stage1[3][5] ), .B1(n7182), .B2(
        n6668), .ZN(n6669) );
  INV_X1 U7995 ( .A(n6669), .ZN(n10015) );
  INV_X2 U7996 ( .A(n6711), .ZN(n7330) );
  NAND2_X1 U7997 ( .A1(n6670), .A2(n7161), .ZN(n6671) );
  XOR2_X1 U7998 ( .A(n7163), .B(n6671), .Z(n6672) );
  AOI22_X1 U7999 ( .A1(n7330), .A2(\adder_stage1[3][9] ), .B1(n7182), .B2(
        n6672), .ZN(n6673) );
  INV_X1 U8000 ( .A(n6673), .ZN(n10011) );
  AOI22_X1 U8001 ( .A1(n7330), .A2(\x_mult_f[7][0] ), .B1(n7182), .B2(
        \x_mult_f_int[7][0] ), .ZN(n6674) );
  INV_X1 U8002 ( .A(n6674), .ZN(n9307) );
  OAI21_X1 U8003 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6682) );
  INV_X1 U8004 ( .A(n6678), .ZN(n6680) );
  NAND2_X1 U8005 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  XNOR2_X1 U8006 ( .A(n6682), .B(n6681), .ZN(n6683) );
  AOI22_X1 U8007 ( .A1(n4689), .A2(\adder_stage1[3][7] ), .B1(n7182), .B2(
        n6683), .ZN(n6684) );
  INV_X1 U8008 ( .A(n6684), .ZN(n10013) );
  BUF_X2 U8009 ( .A(n6699), .Z(n7284) );
  INV_X1 U8010 ( .A(n6685), .ZN(n7249) );
  AOI21_X1 U8011 ( .B1(n7249), .B2(n6687), .A(n6686), .ZN(n6716) );
  INV_X1 U8012 ( .A(n6715), .ZN(n6688) );
  NAND2_X1 U8013 ( .A1(n6688), .A2(n6714), .ZN(n6689) );
  XOR2_X1 U8014 ( .A(n6716), .B(n6689), .Z(n6690) );
  AOI22_X1 U8015 ( .A1(n4891), .A2(\adder_stage1[1][6] ), .B1(n7284), .B2(
        n6690), .ZN(n6691) );
  INV_X1 U8016 ( .A(n6691), .ZN(n10047) );
  INV_X1 U8017 ( .A(n6692), .ZN(n7276) );
  OAI21_X1 U8018 ( .B1(n7276), .B2(n7272), .A(n7273), .ZN(n6696) );
  NAND2_X1 U8019 ( .A1(n3435), .A2(n6694), .ZN(n6695) );
  XNOR2_X1 U8020 ( .A(n6696), .B(n6695), .ZN(n6697) );
  AOI22_X1 U8021 ( .A1(n4891), .A2(\adder_stage1[1][3] ), .B1(n7284), .B2(
        n6697), .ZN(n6698) );
  INV_X1 U8022 ( .A(n6698), .ZN(n10050) );
  BUF_X2 U8023 ( .A(n6699), .Z(n8363) );
  AOI22_X1 U8024 ( .A1(n8212), .A2(\x_mult_f[21][0] ), .B1(n8363), .B2(
        \x_mult_f_int[21][0] ), .ZN(n6700) );
  INV_X1 U8025 ( .A(n6700), .ZN(n9335) );
  INV_X1 U8026 ( .A(n6701), .ZN(n6703) );
  NAND2_X1 U8027 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  XOR2_X1 U8028 ( .A(n6705), .B(n6704), .Z(n6706) );
  AOI22_X1 U8029 ( .A1(n7285), .A2(\adder_stage1[1][9] ), .B1(n7284), .B2(
        n6706), .ZN(n6707) );
  INV_X1 U8030 ( .A(n6707), .ZN(n10044) );
  OR2_X1 U8031 ( .A1(\x_mult_f[2][0] ), .A2(\x_mult_f[3][0] ), .ZN(n6708) );
  AND2_X1 U8032 ( .A1(n6708), .A2(n7268), .ZN(n6709) );
  AOI22_X1 U8033 ( .A1(n7244), .A2(\adder_stage1[1][0] ), .B1(n7284), .B2(
        n6709), .ZN(n6710) );
  INV_X1 U8034 ( .A(n6710), .ZN(n10053) );
  INV_X2 U8035 ( .A(n6711), .ZN(n7818) );
  AOI22_X1 U8036 ( .A1(n7818), .A2(\x_mult_f[1][2] ), .B1(n8363), .B2(
        \x_mult_f_int[1][2] ), .ZN(n6712) );
  INV_X1 U8037 ( .A(n6712), .ZN(n8946) );
  AOI22_X1 U8038 ( .A1(n7818), .A2(\x_mult_f[1][3] ), .B1(n8363), .B2(
        \x_mult_f_int[1][3] ), .ZN(n6713) );
  INV_X1 U8039 ( .A(n6713), .ZN(n8945) );
  OAI21_X1 U8040 ( .B1(n6716), .B2(n6715), .A(n6714), .ZN(n6721) );
  INV_X1 U8041 ( .A(n6717), .ZN(n6719) );
  NAND2_X1 U8042 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  XNOR2_X1 U8043 ( .A(n6721), .B(n6720), .ZN(n6722) );
  AOI22_X1 U8044 ( .A1(n5678), .A2(\adder_stage1[1][7] ), .B1(n7284), .B2(
        n6722), .ZN(n6723) );
  INV_X1 U8045 ( .A(n6723), .ZN(n10046) );
  AOI22_X1 U8046 ( .A1(n8036), .A2(\x_mult_f[21][2] ), .B1(n7356), .B2(
        \x_mult_f_int[21][2] ), .ZN(n6724) );
  INV_X1 U8047 ( .A(n6724), .ZN(n9195) );
  INV_X1 U8048 ( .A(n6725), .ZN(n6727) );
  NAND2_X1 U8049 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  XOR2_X1 U8050 ( .A(n6728), .B(n7298), .Z(n6729) );
  AOI22_X1 U8051 ( .A1(n7825), .A2(\adder_stage1[2][1] ), .B1(n7369), .B2(
        n6729), .ZN(n6730) );
  INV_X1 U8052 ( .A(n6730), .ZN(n10035) );
  AOI22_X1 U8053 ( .A1(n8088), .A2(\x_mult_f[21][4] ), .B1(n7356), .B2(
        \x_mult_f_int[21][4] ), .ZN(n6731) );
  INV_X1 U8054 ( .A(n6731), .ZN(n9193) );
  AOI22_X1 U8055 ( .A1(n4891), .A2(\x_mult_f[21][3] ), .B1(n7356), .B2(
        \x_mult_f_int[21][3] ), .ZN(n6732) );
  INV_X1 U8056 ( .A(n6732), .ZN(n9194) );
  AOI22_X1 U8057 ( .A1(n7330), .A2(\x_mult_f[7][2] ), .B1(n7369), .B2(
        \x_mult_f_int[7][2] ), .ZN(n6733) );
  INV_X1 U8058 ( .A(n6733), .ZN(n9026) );
  AOI22_X1 U8059 ( .A1(n7330), .A2(\x_mult_f[7][3] ), .B1(n7369), .B2(
        \x_mult_f_int[7][3] ), .ZN(n6734) );
  INV_X1 U8060 ( .A(n6734), .ZN(n9025) );
  INV_X2 U8061 ( .A(n6711), .ZN(n7512) );
  AOI22_X1 U8062 ( .A1(n7512), .A2(\x_mult_f[6][0] ), .B1(n7369), .B2(
        \x_mult_f_int[6][0] ), .ZN(n6735) );
  INV_X1 U8063 ( .A(n6735), .ZN(n9305) );
  OR2_X1 U8064 ( .A1(\adder_stage1[8][0] ), .A2(\adder_stage1[9][0] ), .ZN(
        n6737) );
  AND2_X1 U8065 ( .A1(n6737), .A2(n7337), .ZN(n6738) );
  AOI22_X1 U8066 ( .A1(n7613), .A2(\adder_stage2[4][0] ), .B1(n7356), .B2(
        n6738), .ZN(n6739) );
  INV_X1 U8067 ( .A(n6739), .ZN(n9737) );
  NAND2_X1 U8068 ( .A1(n6746), .A2(n6740), .ZN(n6741) );
  XNOR2_X1 U8069 ( .A(n6763), .B(n6741), .ZN(n6742) );
  AOI22_X1 U8070 ( .A1(n5294), .A2(\adder_stage1[7][10] ), .B1(n7992), .B2(
        n6742), .ZN(n6743) );
  INV_X1 U8071 ( .A(n6743), .ZN(n9945) );
  AOI22_X1 U8072 ( .A1(n7818), .A2(\x_mult_f[14][0] ), .B1(n7992), .B2(
        \x_mult_f_int[14][0] ), .ZN(n6744) );
  INV_X1 U8073 ( .A(n6744), .ZN(n9321) );
  NAND2_X1 U8074 ( .A1(n3598), .A2(n6748), .ZN(n6749) );
  XOR2_X1 U8075 ( .A(n6750), .B(n6749), .Z(n6751) );
  AOI22_X1 U8076 ( .A1(n6222), .A2(\adder_stage1[7][11] ), .B1(n7992), .B2(
        n6751), .ZN(n6752) );
  INV_X1 U8077 ( .A(n6752), .ZN(n9944) );
  AOI22_X1 U8078 ( .A1(n8088), .A2(\x_mult_f[15][1] ), .B1(n7992), .B2(
        \x_mult_f_int[15][1] ), .ZN(n6753) );
  INV_X1 U8079 ( .A(n6753), .ZN(n9322) );
  INV_X1 U8080 ( .A(n6754), .ZN(n6756) );
  NAND2_X1 U8081 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  XOR2_X1 U8082 ( .A(n6758), .B(n6757), .Z(n6759) );
  AOI22_X1 U8083 ( .A1(n8157), .A2(\adder_stage1[7][9] ), .B1(n7992), .B2(
        n6759), .ZN(n6760) );
  INV_X1 U8084 ( .A(n6760), .ZN(n9946) );
  AOI22_X1 U8085 ( .A1(n7793), .A2(\x_mult_f[15][0] ), .B1(n7992), .B2(
        \x_mult_f_int[15][0] ), .ZN(n6761) );
  INV_X1 U8086 ( .A(n6761), .ZN(n9323) );
  NAND2_X1 U8087 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  XNOR2_X1 U8088 ( .A(n6769), .B(n6768), .ZN(n6770) );
  AOI22_X1 U8089 ( .A1(n8078), .A2(\adder_stage1[7][12] ), .B1(n7992), .B2(
        n6770), .ZN(n6771) );
  INV_X1 U8090 ( .A(n6771), .ZN(n9943) );
  AOI22_X1 U8091 ( .A1(n7285), .A2(\x_mult_f[9][0] ), .B1(n7454), .B2(
        \x_mult_f_int[9][0] ), .ZN(n6772) );
  INV_X1 U8092 ( .A(n6772), .ZN(n9311) );
  OR2_X1 U8093 ( .A1(\x_mult_f[8][0] ), .A2(\x_mult_f[9][0] ), .ZN(n6773) );
  AND2_X1 U8094 ( .A1(n6773), .A2(n7390), .ZN(n6774) );
  AOI22_X1 U8095 ( .A1(n8036), .A2(\adder_stage1[4][0] ), .B1(n7454), .B2(
        n6774), .ZN(n6775) );
  INV_X1 U8096 ( .A(n6775), .ZN(n10003) );
  INV_X1 U8097 ( .A(n6776), .ZN(n7426) );
  AOI21_X1 U8098 ( .B1(n7426), .B2(n6778), .A(n6777), .ZN(n7396) );
  INV_X1 U8099 ( .A(n7395), .ZN(n6779) );
  NAND2_X1 U8100 ( .A1(n6779), .A2(n7394), .ZN(n6780) );
  XOR2_X1 U8101 ( .A(n7396), .B(n6780), .Z(n6781) );
  AOI22_X1 U8102 ( .A1(n7244), .A2(\adder_stage1[4][6] ), .B1(n7454), .B2(
        n6781), .ZN(n6782) );
  INV_X1 U8103 ( .A(n6782), .ZN(n9997) );
  OAI21_X1 U8104 ( .B1(n6816), .B2(n6784), .A(n6783), .ZN(n6863) );
  INV_X1 U8105 ( .A(n6863), .ZN(n6846) );
  INV_X1 U8106 ( .A(n6796), .ZN(n6785) );
  NAND2_X1 U8107 ( .A1(n6785), .A2(n6795), .ZN(n6786) );
  XOR2_X1 U8108 ( .A(n6846), .B(n6786), .Z(n6787) );
  AOI22_X1 U8109 ( .A1(n7030), .A2(\adder_stage3[0][8] ), .B1(n8291), .B2(
        n6787), .ZN(n6788) );
  INV_X1 U8110 ( .A(n6788), .ZN(n9661) );
  NAND2_X1 U8111 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  XNOR2_X1 U8112 ( .A(n6792), .B(n6791), .ZN(n6793) );
  AOI22_X1 U8113 ( .A1(n7030), .A2(\adder_stage3[0][14] ), .B1(n8291), .B2(
        n6793), .ZN(n6794) );
  INV_X1 U8114 ( .A(n6794), .ZN(n9655) );
  OAI21_X1 U8115 ( .B1(n6846), .B2(n6796), .A(n6795), .ZN(n6801) );
  INV_X1 U8116 ( .A(n6797), .ZN(n6799) );
  NAND2_X1 U8117 ( .A1(n6799), .A2(n6798), .ZN(n6800) );
  XNOR2_X1 U8118 ( .A(n6801), .B(n6800), .ZN(n6802) );
  AOI22_X1 U8119 ( .A1(n7030), .A2(\adder_stage3[0][9] ), .B1(n8291), .B2(
        n6802), .ZN(n6803) );
  INV_X1 U8120 ( .A(n6803), .ZN(n9660) );
  INV_X1 U8121 ( .A(n6804), .ZN(n6806) );
  INV_X1 U8122 ( .A(n6843), .ZN(n6805) );
  OAI21_X1 U8123 ( .B1(n6846), .B2(n6806), .A(n6805), .ZN(n6838) );
  INV_X1 U8124 ( .A(n6807), .ZN(n6836) );
  INV_X1 U8125 ( .A(n6835), .ZN(n6808) );
  AOI21_X1 U8126 ( .B1(n6838), .B2(n6836), .A(n6808), .ZN(n6813) );
  INV_X1 U8127 ( .A(n6809), .ZN(n6811) );
  NAND2_X1 U8128 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  XOR2_X1 U8129 ( .A(n6813), .B(n6812), .Z(n6814) );
  AOI22_X1 U8130 ( .A1(n7030), .A2(\adder_stage3[0][11] ), .B1(n8291), .B2(
        n6814), .ZN(n6815) );
  INV_X1 U8131 ( .A(n6815), .ZN(n9658) );
  INV_X1 U8132 ( .A(n6816), .ZN(n6906) );
  INV_X1 U8133 ( .A(n6817), .ZN(n6904) );
  INV_X1 U8134 ( .A(n6903), .ZN(n6818) );
  AOI21_X1 U8135 ( .B1(n6906), .B2(n6904), .A(n6818), .ZN(n6823) );
  INV_X1 U8136 ( .A(n6819), .ZN(n6821) );
  NAND2_X1 U8137 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  XOR2_X1 U8138 ( .A(n6823), .B(n6822), .Z(n6824) );
  AOI22_X1 U8139 ( .A1(n7030), .A2(\adder_stage3[0][5] ), .B1(n8291), .B2(
        n6824), .ZN(n6825) );
  INV_X1 U8140 ( .A(n6825), .ZN(n9664) );
  AOI21_X1 U8141 ( .B1(n6906), .B2(n6827), .A(n6826), .ZN(n6856) );
  OAI21_X1 U8142 ( .B1(n6856), .B2(n6852), .A(n6853), .ZN(n6832) );
  INV_X1 U8143 ( .A(n6828), .ZN(n6830) );
  NAND2_X1 U8144 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  XNOR2_X1 U8145 ( .A(n6832), .B(n6831), .ZN(n6833) );
  AOI22_X1 U8146 ( .A1(n7030), .A2(\adder_stage3[0][7] ), .B1(n8291), .B2(
        n6833), .ZN(n6834) );
  INV_X1 U8147 ( .A(n6834), .ZN(n9662) );
  NAND2_X1 U8148 ( .A1(n6836), .A2(n6835), .ZN(n6837) );
  XNOR2_X1 U8149 ( .A(n6838), .B(n6837), .ZN(n6839) );
  AOI22_X1 U8150 ( .A1(n7030), .A2(\adder_stage3[0][10] ), .B1(n8291), .B2(
        n6839), .ZN(n6840) );
  INV_X1 U8151 ( .A(n6840), .ZN(n9659) );
  AOI21_X1 U8152 ( .B1(n6843), .B2(n6842), .A(n6841), .ZN(n6844) );
  OAI21_X1 U8153 ( .B1(n6846), .B2(n6845), .A(n6844), .ZN(n6849) );
  INV_X1 U8154 ( .A(n6847), .ZN(n6859) );
  NAND2_X1 U8155 ( .A1(n6859), .A2(n6864), .ZN(n6848) );
  XNOR2_X1 U8156 ( .A(n6849), .B(n6848), .ZN(n6850) );
  AOI22_X1 U8157 ( .A1(n7030), .A2(\adder_stage3[0][12] ), .B1(n8291), .B2(
        n6850), .ZN(n6851) );
  INV_X1 U8158 ( .A(n6851), .ZN(n9657) );
  INV_X1 U8159 ( .A(n6852), .ZN(n6854) );
  NAND2_X1 U8160 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  XOR2_X1 U8161 ( .A(n6856), .B(n6855), .Z(n6857) );
  AOI22_X1 U8162 ( .A1(n7030), .A2(\adder_stage3[0][6] ), .B1(n8291), .B2(
        n6857), .ZN(n6858) );
  INV_X1 U8163 ( .A(n6858), .ZN(n9663) );
  AND3_X1 U8164 ( .A1(n6861), .A2(n6860), .A3(n6859), .ZN(n6867) );
  NAND2_X1 U8165 ( .A1(n6863), .A2(n6862), .ZN(n6865) );
  NAND2_X1 U8166 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  NOR2_X1 U8167 ( .A1(n6867), .A2(n6866), .ZN(n6872) );
  INV_X1 U8168 ( .A(n6868), .ZN(n6870) );
  NAND2_X1 U8169 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  XOR2_X1 U8170 ( .A(n6872), .B(n6871), .Z(n6873) );
  AOI22_X1 U8171 ( .A1(n7030), .A2(\adder_stage3[0][13] ), .B1(n8291), .B2(
        n6873), .ZN(n6874) );
  INV_X1 U8172 ( .A(n6874), .ZN(n9656) );
  AOI22_X1 U8173 ( .A1(n7910), .A2(\x_mult_f[14][3] ), .B1(n7992), .B2(
        \x_mult_f_int[14][3] ), .ZN(n6875) );
  INV_X1 U8174 ( .A(n6875), .ZN(n9111) );
  AOI22_X1 U8175 ( .A1(n7910), .A2(\x_mult_f[14][1] ), .B1(n7992), .B2(
        \x_mult_f_int[14][1] ), .ZN(n6876) );
  INV_X1 U8176 ( .A(n6876), .ZN(n9320) );
  AOI22_X1 U8177 ( .A1(n7910), .A2(\x_mult_f[14][4] ), .B1(n7992), .B2(
        \x_mult_f_int[14][4] ), .ZN(n6877) );
  INV_X1 U8178 ( .A(n6877), .ZN(n9110) );
  AOI22_X1 U8179 ( .A1(n7910), .A2(\x_mult_f[14][2] ), .B1(n7992), .B2(
        \x_mult_f_int[14][2] ), .ZN(n6878) );
  INV_X1 U8180 ( .A(n6878), .ZN(n9112) );
  AOI22_X1 U8181 ( .A1(n7330), .A2(\x_mult_f[5][4] ), .B1(n7511), .B2(
        \x_mult_f_int[5][4] ), .ZN(n6879) );
  INV_X1 U8182 ( .A(n6879), .ZN(n8996) );
  AOI22_X1 U8183 ( .A1(n7330), .A2(\x_mult_f[5][3] ), .B1(n7511), .B2(
        \x_mult_f_int[5][3] ), .ZN(n6880) );
  INV_X1 U8184 ( .A(n6880), .ZN(n8997) );
  AOI22_X1 U8185 ( .A1(n7285), .A2(\x_mult_f[9][3] ), .B1(n6915), .B2(
        \x_mult_f_int[9][3] ), .ZN(n6881) );
  INV_X1 U8186 ( .A(n6881), .ZN(n9044) );
  AOI22_X1 U8187 ( .A1(n8195), .A2(\x_mult_f[8][1] ), .B1(n6915), .B2(
        \x_mult_f_int[8][1] ), .ZN(n6882) );
  INV_X1 U8188 ( .A(n6882), .ZN(n9308) );
  AOI22_X1 U8189 ( .A1(n7285), .A2(\x_mult_f[9][1] ), .B1(n6915), .B2(
        \x_mult_f_int[9][1] ), .ZN(n6883) );
  INV_X1 U8190 ( .A(n6883), .ZN(n9310) );
  AOI22_X1 U8191 ( .A1(n7330), .A2(\x_mult_f[8][3] ), .B1(n6915), .B2(
        \x_mult_f_int[8][3] ), .ZN(n6884) );
  INV_X1 U8192 ( .A(n6884), .ZN(n9039) );
  AOI22_X1 U8193 ( .A1(n8195), .A2(\x_mult_f[8][4] ), .B1(n6915), .B2(
        \x_mult_f_int[8][4] ), .ZN(n6885) );
  INV_X1 U8194 ( .A(n6885), .ZN(n9038) );
  INV_X1 U8195 ( .A(n6886), .ZN(n6900) );
  OAI21_X1 U8196 ( .B1(n6900), .B2(n6896), .A(n6897), .ZN(n6891) );
  INV_X1 U8197 ( .A(n6887), .ZN(n6889) );
  NAND2_X1 U8198 ( .A1(n6889), .A2(n6888), .ZN(n6890) );
  XNOR2_X1 U8199 ( .A(n6891), .B(n6890), .ZN(n6892) );
  AOI22_X1 U8200 ( .A1(n7244), .A2(\adder_stage3[0][3] ), .B1(n6915), .B2(
        n6892), .ZN(n6893) );
  INV_X1 U8201 ( .A(n6893), .ZN(n9666) );
  AOI22_X1 U8202 ( .A1(n6330), .A2(\x_mult_f[8][2] ), .B1(n6915), .B2(
        \x_mult_f_int[8][2] ), .ZN(n6894) );
  INV_X1 U8203 ( .A(n6894), .ZN(n9040) );
  AOI22_X1 U8204 ( .A1(n7443), .A2(\x_mult_f[8][0] ), .B1(n6915), .B2(
        \x_mult_f_int[8][0] ), .ZN(n6895) );
  INV_X1 U8205 ( .A(n6895), .ZN(n9309) );
  INV_X1 U8206 ( .A(n6896), .ZN(n6898) );
  NAND2_X1 U8207 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  XOR2_X1 U8208 ( .A(n6900), .B(n6899), .Z(n6901) );
  AOI22_X1 U8209 ( .A1(n7244), .A2(\adder_stage3[0][2] ), .B1(n6915), .B2(
        n6901), .ZN(n6902) );
  INV_X1 U8210 ( .A(n6902), .ZN(n9667) );
  NAND2_X1 U8211 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  XNOR2_X1 U8212 ( .A(n6906), .B(n6905), .ZN(n6907) );
  AOI22_X1 U8213 ( .A1(n7244), .A2(\adder_stage3[0][4] ), .B1(n6915), .B2(
        n6907), .ZN(n6908) );
  INV_X1 U8214 ( .A(n6908), .ZN(n9665) );
  INV_X1 U8215 ( .A(n6909), .ZN(n6911) );
  NAND2_X1 U8216 ( .A1(n6911), .A2(n6910), .ZN(n6913) );
  XOR2_X1 U8217 ( .A(n6913), .B(n6912), .Z(n6914) );
  AOI22_X1 U8218 ( .A1(n7244), .A2(\adder_stage3[0][1] ), .B1(n6915), .B2(
        n6914), .ZN(n6916) );
  INV_X1 U8219 ( .A(n6916), .ZN(n9668) );
  INV_X2 U8220 ( .A(n6917), .ZN(n8330) );
  BUF_X2 U8221 ( .A(n6955), .Z(n8390) );
  AOI22_X1 U8222 ( .A1(n8330), .A2(\x_mult_f[12][0] ), .B1(n8390), .B2(
        \x_mult_f_int[12][0] ), .ZN(n6918) );
  INV_X1 U8223 ( .A(n6918), .ZN(n9317) );
  AOI22_X1 U8224 ( .A1(n8330), .A2(\x_mult_f[13][3] ), .B1(n8390), .B2(
        \x_mult_f_int[13][3] ), .ZN(n6919) );
  INV_X1 U8225 ( .A(n6919), .ZN(n9097) );
  AOI22_X1 U8226 ( .A1(n8330), .A2(\x_mult_f[13][1] ), .B1(n8390), .B2(
        \x_mult_f_int[13][1] ), .ZN(n6920) );
  INV_X1 U8227 ( .A(n6920), .ZN(n9318) );
  AOI22_X1 U8228 ( .A1(n8330), .A2(\x_mult_f[13][4] ), .B1(n8390), .B2(
        \x_mult_f_int[13][4] ), .ZN(n6921) );
  INV_X1 U8229 ( .A(n6921), .ZN(n9096) );
  AOI22_X1 U8230 ( .A1(n8330), .A2(\x_mult_f[13][2] ), .B1(n8390), .B2(
        \x_mult_f_int[13][2] ), .ZN(n6922) );
  INV_X1 U8231 ( .A(n6922), .ZN(n9098) );
  OR2_X1 U8232 ( .A1(\adder_stage1[4][0] ), .A2(\adder_stage1[5][0] ), .ZN(
        n6923) );
  AND2_X1 U8233 ( .A1(n6923), .A2(n7790), .ZN(n6924) );
  AOI22_X1 U8234 ( .A1(n7793), .A2(\adder_stage2[2][0] ), .B1(n8390), .B2(
        n6924), .ZN(n6925) );
  INV_X1 U8235 ( .A(n6925), .ZN(n9771) );
  INV_X1 U8236 ( .A(n6926), .ZN(n7779) );
  INV_X1 U8237 ( .A(n7778), .ZN(n6927) );
  NAND2_X1 U8238 ( .A1(n6927), .A2(n7777), .ZN(n6928) );
  XOR2_X1 U8239 ( .A(n7779), .B(n6928), .Z(n6929) );
  AOI22_X1 U8240 ( .A1(n7793), .A2(\adder_stage2[2][2] ), .B1(n8390), .B2(
        n6929), .ZN(n6930) );
  INV_X1 U8241 ( .A(n6930), .ZN(n9769) );
  INV_X1 U8242 ( .A(n6931), .ZN(n6996) );
  INV_X1 U8243 ( .A(n6932), .ZN(n6995) );
  NAND2_X1 U8244 ( .A1(n6995), .A2(n6993), .ZN(n6933) );
  XNOR2_X1 U8245 ( .A(n6996), .B(n6933), .ZN(n6934) );
  AOI22_X1 U8246 ( .A1(n7818), .A2(\adder_stage2[2][4] ), .B1(n8390), .B2(
        n6934), .ZN(n6935) );
  INV_X1 U8247 ( .A(n6935), .ZN(n9767) );
  AOI21_X1 U8248 ( .B1(n6996), .B2(n6937), .A(n6936), .ZN(n7807) );
  OAI21_X1 U8249 ( .B1(n7807), .B2(n7803), .A(n7804), .ZN(n6942) );
  INV_X1 U8250 ( .A(n6938), .ZN(n6940) );
  NAND2_X1 U8251 ( .A1(n6940), .A2(n6939), .ZN(n6941) );
  XNOR2_X1 U8252 ( .A(n6942), .B(n6941), .ZN(n6943) );
  AOI22_X1 U8253 ( .A1(n7825), .A2(\adder_stage2[2][7] ), .B1(n8390), .B2(
        n6943), .ZN(n6944) );
  INV_X1 U8254 ( .A(n6944), .ZN(n9764) );
  AOI22_X1 U8255 ( .A1(n7818), .A2(\x_mult_f[1][0] ), .B1(n8208), .B2(
        \x_mult_f_int[1][0] ), .ZN(n6945) );
  INV_X1 U8256 ( .A(n6945), .ZN(n9295) );
  AOI22_X1 U8257 ( .A1(n8391), .A2(\x_mult_f[12][3] ), .B1(n8390), .B2(
        \x_mult_f_int[12][3] ), .ZN(n6946) );
  INV_X1 U8258 ( .A(n6946), .ZN(n9083) );
  BUF_X2 U8259 ( .A(n6645), .Z(n7698) );
  INV_X1 U8260 ( .A(n6947), .ZN(n7696) );
  OAI21_X1 U8261 ( .B1(n7696), .B2(n7692), .A(n7693), .ZN(n6952) );
  INV_X1 U8262 ( .A(n6948), .ZN(n6950) );
  NAND2_X1 U8263 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  XNOR2_X1 U8264 ( .A(n6952), .B(n6951), .ZN(n6953) );
  AOI22_X1 U8265 ( .A1(n7443), .A2(\adder_stage1[9][3] ), .B1(n7698), .B2(
        n6953), .ZN(n6954) );
  INV_X1 U8266 ( .A(n6954), .ZN(n9918) );
  BUF_X2 U8267 ( .A(n6955), .Z(n7909) );
  AOI22_X1 U8268 ( .A1(n8330), .A2(\x_mult_f[13][0] ), .B1(n7909), .B2(
        \x_mult_f_int[13][0] ), .ZN(n6956) );
  INV_X1 U8269 ( .A(n6956), .ZN(n9319) );
  INV_X1 U8270 ( .A(n6957), .ZN(n6959) );
  NAND2_X1 U8271 ( .A1(n6959), .A2(n6958), .ZN(n6960) );
  XOR2_X1 U8272 ( .A(n6961), .B(n6960), .Z(n6962) );
  AOI22_X1 U8273 ( .A1(n8330), .A2(\adder_stage1[6][11] ), .B1(n7909), .B2(
        n6962), .ZN(n6963) );
  INV_X1 U8274 ( .A(n6963), .ZN(n9961) );
  NAND2_X1 U8275 ( .A1(n6980), .A2(n6964), .ZN(n6966) );
  NAND2_X1 U8276 ( .A1(n6966), .A2(n6965), .ZN(n6970) );
  NAND2_X1 U8277 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  XNOR2_X1 U8278 ( .A(n6970), .B(n6969), .ZN(n6971) );
  AOI22_X1 U8279 ( .A1(n8330), .A2(\adder_stage1[6][10] ), .B1(n7909), .B2(
        n6971), .ZN(n6972) );
  INV_X1 U8280 ( .A(n6972), .ZN(n9962) );
  NAND2_X1 U8281 ( .A1(n6979), .A2(n6973), .ZN(n6974) );
  XNOR2_X1 U8282 ( .A(n6980), .B(n6974), .ZN(n6976) );
  AOI22_X1 U8283 ( .A1(n8330), .A2(\adder_stage1[6][8] ), .B1(n7909), .B2(
        n6976), .ZN(n6977) );
  INV_X1 U8284 ( .A(n6977), .ZN(n9964) );
  AOI21_X1 U8285 ( .B1(n6980), .B2(n6979), .A(n6978), .ZN(n6984) );
  NAND2_X1 U8286 ( .A1(n6982), .A2(n6981), .ZN(n6983) );
  XOR2_X1 U8287 ( .A(n6984), .B(n6983), .Z(n6985) );
  AOI22_X1 U8288 ( .A1(n8330), .A2(\adder_stage1[6][9] ), .B1(n7909), .B2(
        n6985), .ZN(n6986) );
  INV_X1 U8289 ( .A(n6986), .ZN(n9963) );
  NAND2_X1 U8290 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  XNOR2_X1 U8291 ( .A(n6990), .B(n6989), .ZN(n6991) );
  AOI22_X1 U8292 ( .A1(n8330), .A2(\adder_stage1[6][12] ), .B1(n7909), .B2(
        n6991), .ZN(n6992) );
  INV_X1 U8293 ( .A(n6992), .ZN(n9960) );
  INV_X1 U8294 ( .A(n6993), .ZN(n6994) );
  AOI21_X1 U8295 ( .B1(n6996), .B2(n6995), .A(n6994), .ZN(n7001) );
  INV_X1 U8296 ( .A(n6997), .ZN(n6999) );
  NAND2_X1 U8297 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  XOR2_X1 U8298 ( .A(n7001), .B(n7000), .Z(n7002) );
  AOI22_X1 U8299 ( .A1(n7818), .A2(\adder_stage2[2][5] ), .B1(n7909), .B2(
        n7002), .ZN(n7003) );
  INV_X1 U8300 ( .A(n7003), .ZN(n9766) );
  AOI22_X1 U8301 ( .A1(n5678), .A2(\x_mult_f[4][3] ), .B1(n7029), .B2(
        \x_mult_f_int[4][3] ), .ZN(n7004) );
  INV_X1 U8302 ( .A(n7004), .ZN(n8986) );
  AOI22_X1 U8303 ( .A1(n7285), .A2(\x_mult_f[4][4] ), .B1(n7029), .B2(
        \x_mult_f_int[4][4] ), .ZN(n7005) );
  INV_X1 U8304 ( .A(n7005), .ZN(n8985) );
  INV_X1 U8305 ( .A(n7006), .ZN(n7027) );
  OAI21_X1 U8306 ( .B1(n7027), .B2(n7007), .A(n7024), .ZN(n7011) );
  NAND2_X1 U8307 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  XNOR2_X1 U8308 ( .A(n7011), .B(n7010), .ZN(n7012) );
  AOI22_X1 U8309 ( .A1(n7244), .A2(\adder_stage2[0][9] ), .B1(n7029), .B2(
        n7012), .ZN(n7013) );
  INV_X1 U8310 ( .A(n7013), .ZN(n9796) );
  AOI22_X1 U8311 ( .A1(n8400), .A2(\x_mult_f[4][2] ), .B1(n7029), .B2(
        \x_mult_f_int[4][2] ), .ZN(n7014) );
  INV_X1 U8312 ( .A(n7014), .ZN(n8987) );
  OAI21_X1 U8313 ( .B1(n7027), .B2(n7016), .A(n7015), .ZN(n7021) );
  INV_X1 U8314 ( .A(n7017), .ZN(n7019) );
  NAND2_X1 U8315 ( .A1(n7019), .A2(n7018), .ZN(n7020) );
  XNOR2_X1 U8316 ( .A(n7021), .B(n7020), .ZN(n7022) );
  AOI22_X1 U8317 ( .A1(n7244), .A2(\adder_stage2[0][10] ), .B1(n7029), .B2(
        n7022), .ZN(n7023) );
  INV_X1 U8318 ( .A(n7023), .ZN(n9795) );
  NAND2_X1 U8319 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  XOR2_X1 U8320 ( .A(n7027), .B(n7026), .Z(n7028) );
  AOI22_X1 U8321 ( .A1(n7030), .A2(\adder_stage2[0][8] ), .B1(n7029), .B2(
        n7028), .ZN(n7031) );
  INV_X1 U8322 ( .A(n7031), .ZN(n9797) );
  AOI22_X1 U8323 ( .A1(n7851), .A2(\x_mult_f[2][0] ), .B1(n7117), .B2(
        \x_mult_f_int[2][0] ), .ZN(n7032) );
  INV_X1 U8324 ( .A(n7032), .ZN(n9297) );
  AOI22_X1 U8325 ( .A1(n7851), .A2(\x_mult_f[2][4] ), .B1(n7117), .B2(
        \x_mult_f_int[2][4] ), .ZN(n7033) );
  INV_X1 U8326 ( .A(n7033), .ZN(n8958) );
  AOI22_X1 U8327 ( .A1(n7851), .A2(\x_mult_f[2][1] ), .B1(n7117), .B2(
        \x_mult_f_int[2][1] ), .ZN(n7034) );
  INV_X1 U8328 ( .A(n7034), .ZN(n9296) );
  AOI22_X1 U8329 ( .A1(n7767), .A2(\x_mult_f[18][0] ), .B1(n7110), .B2(
        \x_mult_f_int[18][0] ), .ZN(n7035) );
  INV_X1 U8330 ( .A(n7035), .ZN(n9329) );
  INV_X1 U8331 ( .A(n7036), .ZN(n7038) );
  NAND2_X1 U8332 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  XOR2_X1 U8333 ( .A(n7040), .B(n7039), .Z(n7041) );
  AOI22_X1 U8334 ( .A1(n6222), .A2(\adder_stage1[5][11] ), .B1(n8389), .B2(
        n7041), .ZN(n7042) );
  INV_X1 U8335 ( .A(n7042), .ZN(n9978) );
  NAND2_X1 U8336 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  XNOR2_X1 U8337 ( .A(n7046), .B(n7045), .ZN(n7047) );
  AOI22_X1 U8338 ( .A1(n7285), .A2(\adder_stage1[1][12] ), .B1(n7117), .B2(
        n7047), .ZN(n7048) );
  INV_X1 U8339 ( .A(n7048), .ZN(n10041) );
  NAND2_X1 U8340 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  XNOR2_X1 U8341 ( .A(n7052), .B(n7051), .ZN(n7053) );
  AOI22_X1 U8342 ( .A1(n7818), .A2(\adder_stage1[5][12] ), .B1(n8389), .B2(
        n7053), .ZN(n7054) );
  INV_X1 U8343 ( .A(n7054), .ZN(n9977) );
  OR2_X1 U8344 ( .A1(\x_mult_f[0][0] ), .A2(\x_mult_f[1][0] ), .ZN(n7055) );
  AND2_X1 U8345 ( .A1(n7055), .A2(n7675), .ZN(n7056) );
  AOI22_X1 U8346 ( .A1(n7793), .A2(\adder_stage1[0][0] ), .B1(n7117), .B2(
        n7056), .ZN(n7057) );
  INV_X1 U8347 ( .A(n7057), .ZN(n10069) );
  AOI22_X1 U8348 ( .A1(n7851), .A2(\x_mult_f[10][0] ), .B1(n8389), .B2(
        \x_mult_f_int[10][0] ), .ZN(n7058) );
  INV_X1 U8349 ( .A(n7058), .ZN(n9313) );
  OAI21_X1 U8350 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(n7066) );
  INV_X1 U8351 ( .A(n7062), .ZN(n7064) );
  NAND2_X1 U8352 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  XNOR2_X1 U8353 ( .A(n7066), .B(n7065), .ZN(n7067) );
  AOI22_X1 U8354 ( .A1(n7512), .A2(\adder_stage1[9][7] ), .B1(n7110), .B2(
        n7067), .ZN(n7068) );
  INV_X1 U8355 ( .A(n7068), .ZN(n9914) );
  INV_X1 U8356 ( .A(n7069), .ZN(n7680) );
  INV_X1 U8357 ( .A(n7679), .ZN(n7070) );
  AOI21_X1 U8358 ( .B1(n7682), .B2(n7680), .A(n7070), .ZN(n7075) );
  INV_X1 U8359 ( .A(n7071), .ZN(n7073) );
  NAND2_X1 U8360 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  XOR2_X1 U8361 ( .A(n7075), .B(n7074), .Z(n7076) );
  AOI22_X1 U8362 ( .A1(n6428), .A2(\adder_stage1[9][5] ), .B1(n7110), .B2(
        n7076), .ZN(n7077) );
  INV_X1 U8363 ( .A(n7077), .ZN(n9916) );
  NAND2_X1 U8364 ( .A1(n3632), .A2(n7080), .ZN(n7081) );
  XOR2_X1 U8365 ( .A(n7082), .B(n7081), .Z(n7083) );
  AOI22_X1 U8366 ( .A1(n5544), .A2(\adder_stage1[9][11] ), .B1(n7110), .B2(
        n7083), .ZN(n7084) );
  INV_X1 U8367 ( .A(n7084), .ZN(n9910) );
  AOI22_X1 U8368 ( .A1(n7793), .A2(\x_mult_f[11][4] ), .B1(n8389), .B2(
        \x_mult_f_int[11][4] ), .ZN(n7085) );
  INV_X1 U8369 ( .A(n7085), .ZN(n9069) );
  AOI22_X1 U8370 ( .A1(n7775), .A2(\x_mult_f[19][2] ), .B1(n7110), .B2(
        \x_mult_f_int[19][2] ), .ZN(n7086) );
  INV_X1 U8371 ( .A(n7086), .ZN(n9181) );
  NAND2_X1 U8372 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  XNOR2_X1 U8373 ( .A(n7093), .B(n7092), .ZN(n7094) );
  AOI22_X1 U8374 ( .A1(n7767), .A2(\adder_stage1[9][12] ), .B1(n7110), .B2(
        n7094), .ZN(n7095) );
  INV_X1 U8375 ( .A(n7095), .ZN(n9909) );
  AOI22_X1 U8376 ( .A1(n7851), .A2(\x_mult_f[10][3] ), .B1(n8389), .B2(
        \x_mult_f_int[10][3] ), .ZN(n7096) );
  INV_X1 U8377 ( .A(n7096), .ZN(n9057) );
  AOI22_X1 U8378 ( .A1(n7851), .A2(\x_mult_f[10][1] ), .B1(n8389), .B2(
        \x_mult_f_int[10][1] ), .ZN(n7097) );
  INV_X1 U8379 ( .A(n7097), .ZN(n9312) );
  INV_X1 U8380 ( .A(n7098), .ZN(n7100) );
  NAND2_X1 U8381 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  XOR2_X1 U8382 ( .A(n7102), .B(n7101), .Z(n7103) );
  AOI22_X1 U8383 ( .A1(n7285), .A2(\adder_stage1[1][11] ), .B1(n7117), .B2(
        n7103), .ZN(n7104) );
  INV_X1 U8384 ( .A(n7104), .ZN(n10042) );
  NAND2_X1 U8385 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  XNOR2_X1 U8386 ( .A(n7108), .B(n7107), .ZN(n7109) );
  AOI22_X1 U8387 ( .A1(n4891), .A2(\adder_stage1[9][10] ), .B1(n7110), .B2(
        n7109), .ZN(n7111) );
  INV_X1 U8388 ( .A(n7111), .ZN(n9911) );
  NAND2_X1 U8389 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  XNOR2_X1 U8390 ( .A(n7115), .B(n7114), .ZN(n7116) );
  AOI22_X1 U8391 ( .A1(n7285), .A2(\adder_stage1[1][10] ), .B1(n7117), .B2(
        n7116), .ZN(n7118) );
  INV_X1 U8392 ( .A(n7118), .ZN(n10043) );
  NAND2_X1 U8393 ( .A1(n7120), .A2(n7119), .ZN(n7122) );
  NAND2_X1 U8394 ( .A1(n7122), .A2(n7121), .ZN(n7126) );
  NAND2_X1 U8395 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  XNOR2_X1 U8396 ( .A(n7126), .B(n7125), .ZN(n7127) );
  AOI22_X1 U8397 ( .A1(n8155), .A2(\adder_stage1[5][10] ), .B1(n8389), .B2(
        n7127), .ZN(n7128) );
  INV_X1 U8398 ( .A(n7128), .ZN(n9979) );
  NAND2_X1 U8399 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  XNOR2_X1 U8400 ( .A(n7132), .B(n7131), .ZN(n7133) );
  AOI22_X1 U8401 ( .A1(n7330), .A2(\adder_stage1[3][8] ), .B1(n7182), .B2(
        n7133), .ZN(n7134) );
  INV_X1 U8402 ( .A(n7134), .ZN(n10012) );
  AOI22_X1 U8403 ( .A1(n7330), .A2(\x_mult_f[7][1] ), .B1(n7182), .B2(
        \x_mult_f_int[7][1] ), .ZN(n7135) );
  INV_X1 U8404 ( .A(n7135), .ZN(n9306) );
  OAI21_X1 U8405 ( .B1(n7163), .B2(n7137), .A(n7136), .ZN(n7141) );
  NAND2_X1 U8406 ( .A1(n7139), .A2(n7138), .ZN(n7140) );
  XNOR2_X1 U8407 ( .A(n7141), .B(n7140), .ZN(n7142) );
  AOI22_X1 U8408 ( .A1(n7330), .A2(\adder_stage1[3][12] ), .B1(n7182), .B2(
        n7142), .ZN(n7143) );
  INV_X1 U8409 ( .A(n7143), .ZN(n10008) );
  OAI21_X1 U8410 ( .B1(n7843), .B2(n7145), .A(n7144), .ZN(n7149) );
  NAND2_X1 U8411 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  XNOR2_X1 U8412 ( .A(n7149), .B(n7148), .ZN(n7150) );
  AOI22_X1 U8413 ( .A1(n7851), .A2(\adder_stage2[2][14] ), .B1(n7182), .B2(
        n7150), .ZN(n7151) );
  INV_X1 U8414 ( .A(n7151), .ZN(n9757) );
  OAI21_X1 U8415 ( .B1(n7163), .B2(n7153), .A(n7152), .ZN(n7154) );
  INV_X1 U8416 ( .A(n7154), .ZN(n7158) );
  NAND2_X1 U8417 ( .A1(n7156), .A2(n7155), .ZN(n7157) );
  XOR2_X1 U8418 ( .A(n7158), .B(n7157), .Z(n7159) );
  AOI22_X1 U8419 ( .A1(n7330), .A2(\adder_stage1[3][11] ), .B1(n7182), .B2(
        n7159), .ZN(n7160) );
  INV_X1 U8420 ( .A(n7160), .ZN(n10009) );
  OAI21_X1 U8421 ( .B1(n7163), .B2(n7162), .A(n7161), .ZN(n7167) );
  NAND2_X1 U8422 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  XNOR2_X1 U8423 ( .A(n7167), .B(n7166), .ZN(n7168) );
  AOI22_X1 U8424 ( .A1(n7330), .A2(\adder_stage1[3][10] ), .B1(n7182), .B2(
        n7168), .ZN(n7169) );
  INV_X1 U8425 ( .A(n7169), .ZN(n10010) );
  INV_X1 U8426 ( .A(n7170), .ZN(n7172) );
  NAND2_X1 U8427 ( .A1(n7172), .A2(n7171), .ZN(n7173) );
  XOR2_X1 U8428 ( .A(n7174), .B(n7173), .Z(n7175) );
  AOI22_X1 U8429 ( .A1(n8381), .A2(\adder_stage1[3][2] ), .B1(n7182), .B2(
        n7175), .ZN(n7176) );
  INV_X1 U8430 ( .A(n7176), .ZN(n10018) );
  NAND2_X1 U8431 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  XNOR2_X1 U8432 ( .A(n7180), .B(n7179), .ZN(n7181) );
  AOI22_X1 U8433 ( .A1(n8400), .A2(\adder_stage1[3][4] ), .B1(n7182), .B2(
        n7181), .ZN(n7183) );
  INV_X1 U8434 ( .A(n7183), .ZN(n10016) );
  AOI22_X1 U8435 ( .A1(n8078), .A2(\x_mult_f[21][1] ), .B1(n8363), .B2(
        \x_mult_f_int[21][1] ), .ZN(n7184) );
  INV_X1 U8436 ( .A(n7184), .ZN(n9334) );
  AOI22_X1 U8437 ( .A1(n7851), .A2(\x_mult_f[0][0] ), .B1(n8363), .B2(
        \x_mult_f_int[0][0] ), .ZN(n7185) );
  INV_X1 U8438 ( .A(n7185), .ZN(n9293) );
  AOI22_X1 U8439 ( .A1(n7818), .A2(\x_mult_f[1][4] ), .B1(n8363), .B2(
        \x_mult_f_int[1][4] ), .ZN(n7186) );
  INV_X1 U8440 ( .A(n7186), .ZN(n8944) );
  NAND2_X1 U8441 ( .A1(n7188), .A2(n7187), .ZN(n7189) );
  XNOR2_X1 U8442 ( .A(n7190), .B(n7189), .ZN(n7191) );
  AOI22_X1 U8443 ( .A1(n7244), .A2(\adder_stage2[0][14] ), .B1(n7284), .B2(
        n7191), .ZN(n7192) );
  INV_X1 U8444 ( .A(n7192), .ZN(n9791) );
  NAND2_X1 U8445 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  XNOR2_X1 U8446 ( .A(n7199), .B(n7198), .ZN(n7200) );
  AOI22_X1 U8447 ( .A1(n8228), .A2(\adder_stage1[10][12] ), .B1(n8363), .B2(
        n7200), .ZN(n7201) );
  INV_X1 U8448 ( .A(n7201), .ZN(n9893) );
  NAND2_X1 U8449 ( .A1(n7203), .A2(n7202), .ZN(n7204) );
  XNOR2_X1 U8450 ( .A(n7205), .B(n7204), .ZN(n7206) );
  AOI22_X1 U8451 ( .A1(n8154), .A2(\adder_stage1[10][8] ), .B1(n8363), .B2(
        n7206), .ZN(n7207) );
  INV_X1 U8452 ( .A(n7207), .ZN(n9897) );
  INV_X1 U8453 ( .A(n7208), .ZN(n7247) );
  INV_X1 U8454 ( .A(n7246), .ZN(n7209) );
  AOI21_X1 U8455 ( .B1(n7249), .B2(n7247), .A(n7209), .ZN(n7214) );
  INV_X1 U8456 ( .A(n7210), .ZN(n7212) );
  NAND2_X1 U8457 ( .A1(n7212), .A2(n7211), .ZN(n7213) );
  XOR2_X1 U8458 ( .A(n7214), .B(n7213), .Z(n7215) );
  AOI22_X1 U8459 ( .A1(n8154), .A2(\adder_stage1[1][5] ), .B1(n7284), .B2(
        n7215), .ZN(n7216) );
  INV_X1 U8460 ( .A(n7216), .ZN(n10048) );
  INV_X1 U8461 ( .A(n7217), .ZN(n7219) );
  NAND2_X1 U8462 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  XOR2_X1 U8463 ( .A(n7221), .B(n7220), .Z(n7222) );
  AOI22_X1 U8464 ( .A1(n6373), .A2(\adder_stage1[10][9] ), .B1(n8363), .B2(
        n7222), .ZN(n7223) );
  INV_X1 U8465 ( .A(n7223), .ZN(n9896) );
  AOI22_X1 U8466 ( .A1(n7851), .A2(\x_mult_f[0][1] ), .B1(n8363), .B2(
        \x_mult_f_int[0][1] ), .ZN(n7224) );
  INV_X1 U8467 ( .A(n7224), .ZN(n9292) );
  INV_X1 U8468 ( .A(n7225), .ZN(n7227) );
  NAND2_X1 U8469 ( .A1(n7227), .A2(n7226), .ZN(n7228) );
  XOR2_X1 U8470 ( .A(n7229), .B(n7228), .Z(n7230) );
  AOI22_X1 U8471 ( .A1(n7244), .A2(\adder_stage2[0][11] ), .B1(n7284), .B2(
        n7230), .ZN(n7231) );
  INV_X1 U8472 ( .A(n7231), .ZN(n9794) );
  INV_X1 U8473 ( .A(n7232), .ZN(n7234) );
  NAND2_X1 U8474 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  XOR2_X1 U8475 ( .A(n7236), .B(n7235), .Z(n7237) );
  AOI22_X1 U8476 ( .A1(n7244), .A2(\adder_stage2[0][13] ), .B1(n7284), .B2(
        n7237), .ZN(n7238) );
  INV_X1 U8477 ( .A(n7238), .ZN(n9792) );
  NAND2_X1 U8478 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  XNOR2_X1 U8479 ( .A(n7242), .B(n7241), .ZN(n7243) );
  AOI22_X1 U8480 ( .A1(n7244), .A2(\adder_stage2[0][12] ), .B1(n7284), .B2(
        n7243), .ZN(n7245) );
  INV_X1 U8481 ( .A(n7245), .ZN(n9793) );
  NAND2_X1 U8482 ( .A1(n7247), .A2(n7246), .ZN(n7248) );
  XNOR2_X1 U8483 ( .A(n7249), .B(n7248), .ZN(n7250) );
  AOI22_X1 U8484 ( .A1(n7613), .A2(\adder_stage1[1][4] ), .B1(n7284), .B2(
        n7250), .ZN(n7251) );
  INV_X1 U8485 ( .A(n7251), .ZN(n10049) );
  NAND2_X1 U8486 ( .A1(n7257), .A2(n7252), .ZN(n7253) );
  XNOR2_X1 U8487 ( .A(n7258), .B(n7253), .ZN(n7254) );
  AOI22_X1 U8488 ( .A1(n8154), .A2(\adder_stage1[10][10] ), .B1(n8363), .B2(
        n7254), .ZN(n7255) );
  INV_X1 U8489 ( .A(n7255), .ZN(n9895) );
  NAND2_X1 U8490 ( .A1(n3581), .A2(n7260), .ZN(n7261) );
  XOR2_X1 U8491 ( .A(n7262), .B(n7261), .Z(n7263) );
  AOI22_X1 U8492 ( .A1(n8202), .A2(\adder_stage1[10][11] ), .B1(n8363), .B2(
        n7263), .ZN(n7264) );
  INV_X1 U8493 ( .A(n7264), .ZN(n9894) );
  INV_X1 U8494 ( .A(n7265), .ZN(n7267) );
  NAND2_X1 U8495 ( .A1(n7267), .A2(n7266), .ZN(n7269) );
  XOR2_X1 U8496 ( .A(n7268), .B(n7269), .Z(n7270) );
  AOI22_X1 U8497 ( .A1(n4891), .A2(\adder_stage1[1][1] ), .B1(n7284), .B2(
        n7270), .ZN(n7271) );
  INV_X1 U8498 ( .A(n7271), .ZN(n10052) );
  INV_X1 U8499 ( .A(n7272), .ZN(n7274) );
  NAND2_X1 U8500 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  XOR2_X1 U8501 ( .A(n7276), .B(n7275), .Z(n7277) );
  AOI22_X1 U8502 ( .A1(n6337), .A2(\adder_stage1[1][2] ), .B1(n7284), .B2(
        n7277), .ZN(n7278) );
  INV_X1 U8503 ( .A(n7278), .ZN(n10051) );
  NAND2_X1 U8504 ( .A1(n7280), .A2(n7279), .ZN(n7281) );
  XNOR2_X1 U8505 ( .A(n7282), .B(n7281), .ZN(n7283) );
  AOI22_X1 U8506 ( .A1(n7285), .A2(\adder_stage1[1][8] ), .B1(n7284), .B2(
        n7283), .ZN(n7286) );
  INV_X1 U8507 ( .A(n7286), .ZN(n10045) );
  INV_X1 U8508 ( .A(n7287), .ZN(n7551) );
  INV_X1 U8509 ( .A(n7288), .ZN(n7353) );
  INV_X1 U8510 ( .A(n7352), .ZN(n7289) );
  AOI21_X1 U8511 ( .B1(n7551), .B2(n7353), .A(n7289), .ZN(n7294) );
  INV_X1 U8512 ( .A(n7290), .ZN(n7292) );
  NAND2_X1 U8513 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  XOR2_X1 U8514 ( .A(n7294), .B(n7293), .Z(n7295) );
  AOI22_X1 U8515 ( .A1(n7613), .A2(\adder_stage2[4][5] ), .B1(n7356), .B2(
        n7295), .ZN(n7296) );
  INV_X1 U8516 ( .A(n7296), .ZN(n9732) );
  AOI22_X1 U8517 ( .A1(n7512), .A2(\x_mult_f[6][4] ), .B1(n7369), .B2(
        \x_mult_f_int[6][4] ), .ZN(n7297) );
  INV_X1 U8518 ( .A(n7297), .ZN(n9010) );
  OR2_X1 U8519 ( .A1(\x_mult_f[4][0] ), .A2(\x_mult_f[5][0] ), .ZN(n7299) );
  AND2_X1 U8520 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  AOI22_X1 U8521 ( .A1(n7512), .A2(\adder_stage1[2][0] ), .B1(n7369), .B2(
        n7300), .ZN(n7301) );
  INV_X1 U8522 ( .A(n7301), .ZN(n10036) );
  AOI22_X1 U8523 ( .A1(n7613), .A2(\x_mult_f[20][4] ), .B1(n7356), .B2(
        \x_mult_f_int[20][4] ), .ZN(n7302) );
  INV_X1 U8524 ( .A(n7302), .ZN(n9185) );
  AOI22_X1 U8525 ( .A1(n7613), .A2(\x_mult_f[20][2] ), .B1(n7356), .B2(
        \x_mult_f_int[20][2] ), .ZN(n7303) );
  INV_X1 U8526 ( .A(n7303), .ZN(n9187) );
  INV_X1 U8527 ( .A(n7304), .ZN(n7479) );
  INV_X1 U8528 ( .A(n7305), .ZN(n7359) );
  INV_X1 U8529 ( .A(n7358), .ZN(n7306) );
  AOI21_X1 U8530 ( .B1(n7479), .B2(n7359), .A(n7306), .ZN(n7311) );
  INV_X1 U8531 ( .A(n7307), .ZN(n7309) );
  NAND2_X1 U8532 ( .A1(n7309), .A2(n7308), .ZN(n7310) );
  XOR2_X1 U8533 ( .A(n7311), .B(n7310), .Z(n7312) );
  AOI22_X1 U8534 ( .A1(n7825), .A2(\adder_stage1[2][5] ), .B1(n7369), .B2(
        n7312), .ZN(n7313) );
  INV_X1 U8535 ( .A(n7313), .ZN(n10031) );
  AOI22_X1 U8536 ( .A1(n7944), .A2(\x_mult_f[20][0] ), .B1(n7356), .B2(
        \x_mult_f_int[20][0] ), .ZN(n7314) );
  INV_X1 U8537 ( .A(n7314), .ZN(n9333) );
  INV_X1 U8538 ( .A(n7315), .ZN(n7344) );
  INV_X1 U8539 ( .A(n7343), .ZN(n7316) );
  NAND2_X1 U8540 ( .A1(n7316), .A2(n7342), .ZN(n7317) );
  XOR2_X1 U8541 ( .A(n7344), .B(n7317), .Z(n7318) );
  AOI22_X1 U8542 ( .A1(n7613), .A2(\adder_stage2[4][2] ), .B1(n7356), .B2(
        n7318), .ZN(n7319) );
  INV_X1 U8543 ( .A(n7319), .ZN(n9735) );
  INV_X1 U8544 ( .A(n7320), .ZN(n7367) );
  OAI21_X1 U8545 ( .B1(n7367), .B2(n7363), .A(n7364), .ZN(n7325) );
  INV_X1 U8546 ( .A(n7321), .ZN(n7323) );
  NAND2_X1 U8547 ( .A1(n7323), .A2(n7322), .ZN(n7324) );
  XNOR2_X1 U8548 ( .A(n7325), .B(n7324), .ZN(n7326) );
  AOI22_X1 U8549 ( .A1(n7825), .A2(\adder_stage1[2][3] ), .B1(n7369), .B2(
        n7326), .ZN(n7327) );
  INV_X1 U8550 ( .A(n7327), .ZN(n10033) );
  AOI22_X1 U8551 ( .A1(n7613), .A2(\x_mult_f[20][1] ), .B1(n7356), .B2(
        \x_mult_f_int[20][1] ), .ZN(n7328) );
  INV_X1 U8552 ( .A(n7328), .ZN(n9332) );
  AOI22_X1 U8553 ( .A1(n7512), .A2(\x_mult_f[6][2] ), .B1(n7369), .B2(
        \x_mult_f_int[6][2] ), .ZN(n7329) );
  INV_X1 U8554 ( .A(n7329), .ZN(n9012) );
  AOI22_X1 U8555 ( .A1(n7330), .A2(\x_mult_f[7][4] ), .B1(n7369), .B2(
        \x_mult_f_int[7][4] ), .ZN(n7331) );
  INV_X1 U8556 ( .A(n7331), .ZN(n9024) );
  AOI22_X1 U8557 ( .A1(n7512), .A2(\x_mult_f[6][3] ), .B1(n7369), .B2(
        \x_mult_f_int[6][3] ), .ZN(n7332) );
  INV_X1 U8558 ( .A(n7332), .ZN(n9011) );
  AOI22_X1 U8559 ( .A1(n7613), .A2(\x_mult_f[20][3] ), .B1(n7356), .B2(
        \x_mult_f_int[20][3] ), .ZN(n7333) );
  INV_X1 U8560 ( .A(n7333), .ZN(n9186) );
  INV_X1 U8561 ( .A(n7334), .ZN(n7336) );
  NAND2_X1 U8562 ( .A1(n7336), .A2(n7335), .ZN(n7338) );
  XOR2_X1 U8563 ( .A(n7338), .B(n7337), .Z(n7339) );
  AOI22_X1 U8564 ( .A1(n7613), .A2(\adder_stage2[4][1] ), .B1(n7356), .B2(
        n7339), .ZN(n7340) );
  INV_X1 U8565 ( .A(n7340), .ZN(n9736) );
  AOI22_X1 U8566 ( .A1(n7512), .A2(\x_mult_f[6][1] ), .B1(n7369), .B2(
        \x_mult_f_int[6][1] ), .ZN(n7341) );
  INV_X1 U8567 ( .A(n7341), .ZN(n9304) );
  OAI21_X1 U8568 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n7349) );
  INV_X1 U8569 ( .A(n7345), .ZN(n7347) );
  NAND2_X1 U8570 ( .A1(n7347), .A2(n7346), .ZN(n7348) );
  XNOR2_X1 U8571 ( .A(n7349), .B(n7348), .ZN(n7350) );
  AOI22_X1 U8572 ( .A1(n7613), .A2(\adder_stage2[4][3] ), .B1(n7356), .B2(
        n7350), .ZN(n7351) );
  INV_X1 U8573 ( .A(n7351), .ZN(n9734) );
  NAND2_X1 U8574 ( .A1(n7353), .A2(n7352), .ZN(n7354) );
  XNOR2_X1 U8575 ( .A(n7551), .B(n7354), .ZN(n7355) );
  AOI22_X1 U8576 ( .A1(n7613), .A2(\adder_stage2[4][4] ), .B1(n7356), .B2(
        n7355), .ZN(n7357) );
  INV_X1 U8577 ( .A(n7357), .ZN(n9733) );
  NAND2_X1 U8578 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  XNOR2_X1 U8579 ( .A(n7479), .B(n7360), .ZN(n7361) );
  AOI22_X1 U8580 ( .A1(n7825), .A2(\adder_stage1[2][4] ), .B1(n7369), .B2(
        n7361), .ZN(n7362) );
  INV_X1 U8581 ( .A(n7362), .ZN(n10032) );
  INV_X1 U8582 ( .A(n7363), .ZN(n7365) );
  NAND2_X1 U8583 ( .A1(n7365), .A2(n7364), .ZN(n7366) );
  XOR2_X1 U8584 ( .A(n7367), .B(n7366), .Z(n7368) );
  AOI22_X1 U8585 ( .A1(n7825), .A2(\adder_stage1[2][2] ), .B1(n7369), .B2(
        n7368), .ZN(n7370) );
  INV_X1 U8586 ( .A(n7370), .ZN(n10034) );
  INV_X1 U8587 ( .A(n7371), .ZN(n7424) );
  INV_X1 U8588 ( .A(n7423), .ZN(n7372) );
  AOI21_X1 U8589 ( .B1(n7426), .B2(n7424), .A(n7372), .ZN(n7377) );
  INV_X1 U8590 ( .A(n7373), .ZN(n7375) );
  NAND2_X1 U8591 ( .A1(n7375), .A2(n7374), .ZN(n7376) );
  XOR2_X1 U8592 ( .A(n7377), .B(n7376), .Z(n7378) );
  AOI22_X1 U8593 ( .A1(n7443), .A2(\adder_stage1[4][5] ), .B1(n7454), .B2(
        n7378), .ZN(n7379) );
  INV_X1 U8594 ( .A(n7379), .ZN(n9998) );
  INV_X1 U8595 ( .A(n7380), .ZN(n7382) );
  NAND2_X1 U8596 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  XOR2_X1 U8597 ( .A(n7384), .B(n7383), .Z(n7385) );
  AOI22_X1 U8598 ( .A1(n8330), .A2(\adder_stage1[4][11] ), .B1(n7454), .B2(
        n7385), .ZN(n7386) );
  INV_X1 U8599 ( .A(n7386), .ZN(n9992) );
  INV_X1 U8600 ( .A(n7387), .ZN(n7389) );
  NAND2_X1 U8601 ( .A1(n7389), .A2(n7388), .ZN(n7391) );
  XOR2_X1 U8602 ( .A(n7391), .B(n7390), .Z(n7392) );
  AOI22_X1 U8603 ( .A1(n7443), .A2(\adder_stage1[4][1] ), .B1(n7454), .B2(
        n7392), .ZN(n7393) );
  INV_X1 U8604 ( .A(n7393), .ZN(n10002) );
  OAI21_X1 U8605 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7401) );
  INV_X1 U8606 ( .A(n7397), .ZN(n7399) );
  NAND2_X1 U8607 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  XNOR2_X1 U8608 ( .A(n7401), .B(n7400), .ZN(n7402) );
  AOI22_X1 U8609 ( .A1(n8178), .A2(\adder_stage1[4][7] ), .B1(n7454), .B2(
        n7402), .ZN(n7403) );
  INV_X1 U8610 ( .A(n7403), .ZN(n9996) );
  AOI21_X1 U8611 ( .B1(n7446), .B2(n7418), .A(n7404), .ZN(n7408) );
  NAND2_X1 U8612 ( .A1(n7406), .A2(n7405), .ZN(n7407) );
  XOR2_X1 U8613 ( .A(n7408), .B(n7407), .Z(n7409) );
  AOI22_X1 U8614 ( .A1(n6581), .A2(\adder_stage1[4][9] ), .B1(n7454), .B2(
        n7409), .ZN(n7410) );
  INV_X1 U8615 ( .A(n7410), .ZN(n9994) );
  NAND2_X1 U8616 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  XNOR2_X1 U8617 ( .A(n7414), .B(n7413), .ZN(n7415) );
  AOI22_X1 U8618 ( .A1(n8154), .A2(\adder_stage1[4][12] ), .B1(n7454), .B2(
        n7415), .ZN(n7416) );
  INV_X1 U8619 ( .A(n7416), .ZN(n9991) );
  NAND2_X1 U8620 ( .A1(n7418), .A2(n7417), .ZN(n7419) );
  XNOR2_X1 U8621 ( .A(n7446), .B(n7419), .ZN(n7421) );
  AOI22_X1 U8622 ( .A1(n8381), .A2(\adder_stage1[4][8] ), .B1(n7454), .B2(
        n7421), .ZN(n7422) );
  INV_X1 U8623 ( .A(n7422), .ZN(n9995) );
  NAND2_X1 U8624 ( .A1(n7424), .A2(n7423), .ZN(n7425) );
  XNOR2_X1 U8625 ( .A(n7426), .B(n7425), .ZN(n7427) );
  AOI22_X1 U8626 ( .A1(n6222), .A2(\adder_stage1[4][4] ), .B1(n7454), .B2(
        n7427), .ZN(n7428) );
  INV_X1 U8627 ( .A(n7428), .ZN(n9999) );
  INV_X1 U8628 ( .A(n7429), .ZN(n7441) );
  OAI21_X1 U8629 ( .B1(n7441), .B2(n7437), .A(n7438), .ZN(n7434) );
  INV_X1 U8630 ( .A(n7430), .ZN(n7432) );
  NAND2_X1 U8631 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  XNOR2_X1 U8632 ( .A(n7434), .B(n7433), .ZN(n7435) );
  AOI22_X1 U8633 ( .A1(n7443), .A2(\adder_stage1[4][3] ), .B1(n7454), .B2(
        n7435), .ZN(n7436) );
  INV_X1 U8634 ( .A(n7436), .ZN(n10000) );
  INV_X1 U8635 ( .A(n7437), .ZN(n7439) );
  NAND2_X1 U8636 ( .A1(n7439), .A2(n7438), .ZN(n7440) );
  XOR2_X1 U8637 ( .A(n7441), .B(n7440), .Z(n7442) );
  AOI22_X1 U8638 ( .A1(n7443), .A2(\adder_stage1[4][2] ), .B1(n7454), .B2(
        n7442), .ZN(n7444) );
  INV_X1 U8639 ( .A(n7444), .ZN(n10001) );
  NAND2_X1 U8640 ( .A1(n7446), .A2(n7445), .ZN(n7448) );
  NAND2_X1 U8641 ( .A1(n7448), .A2(n7447), .ZN(n7452) );
  NAND2_X1 U8642 ( .A1(n7450), .A2(n7449), .ZN(n7451) );
  XNOR2_X1 U8643 ( .A(n7452), .B(n7451), .ZN(n7453) );
  AOI22_X1 U8644 ( .A1(n7818), .A2(\adder_stage1[4][10] ), .B1(n7454), .B2(
        n7453), .ZN(n7455) );
  INV_X1 U8645 ( .A(n7455), .ZN(n9993) );
  NAND2_X1 U8646 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  XNOR2_X1 U8647 ( .A(n7459), .B(n7458), .ZN(n7460) );
  AOI22_X1 U8648 ( .A1(n7825), .A2(\adder_stage1[2][8] ), .B1(n7511), .B2(
        n7460), .ZN(n7461) );
  INV_X1 U8649 ( .A(n7461), .ZN(n10028) );
  AOI22_X1 U8650 ( .A1(n7512), .A2(\x_mult_f[5][2] ), .B1(n7511), .B2(
        \x_mult_f_int[5][2] ), .ZN(n7462) );
  INV_X1 U8651 ( .A(n7462), .ZN(n8998) );
  INV_X1 U8652 ( .A(n7463), .ZN(n7465) );
  NAND2_X1 U8653 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  XOR2_X1 U8654 ( .A(n7467), .B(n7466), .Z(n7468) );
  AOI22_X1 U8655 ( .A1(n7825), .A2(\adder_stage1[2][9] ), .B1(n7511), .B2(
        n7468), .ZN(n7469) );
  INV_X1 U8656 ( .A(n7469), .ZN(n10027) );
  AOI21_X1 U8657 ( .B1(n8223), .B2(n7508), .A(n7470), .ZN(n7474) );
  NAND2_X1 U8658 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  XOR2_X1 U8659 ( .A(n7474), .B(n7473), .Z(n7475) );
  AOI22_X1 U8660 ( .A1(n7512), .A2(\adder_stage1[2][11] ), .B1(n7511), .B2(
        n7475), .ZN(n7476) );
  INV_X1 U8661 ( .A(n7476), .ZN(n10025) );
  AOI21_X1 U8662 ( .B1(n7479), .B2(n7478), .A(n7477), .ZN(n7487) );
  INV_X1 U8663 ( .A(n7486), .ZN(n7480) );
  NAND2_X1 U8664 ( .A1(n7480), .A2(n7485), .ZN(n7481) );
  XOR2_X1 U8665 ( .A(n7487), .B(n7481), .Z(n7482) );
  AOI22_X1 U8666 ( .A1(n7825), .A2(\adder_stage1[2][6] ), .B1(n7511), .B2(
        n7482), .ZN(n7483) );
  INV_X1 U8667 ( .A(n7483), .ZN(n10030) );
  AOI22_X1 U8668 ( .A1(n7512), .A2(\x_mult_f[5][0] ), .B1(n7511), .B2(
        \x_mult_f_int[5][0] ), .ZN(n7484) );
  INV_X1 U8669 ( .A(n7484), .ZN(n9303) );
  OAI21_X1 U8670 ( .B1(n7487), .B2(n7486), .A(n7485), .ZN(n7492) );
  INV_X1 U8671 ( .A(n7488), .ZN(n7490) );
  NAND2_X1 U8672 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  XNOR2_X1 U8673 ( .A(n7492), .B(n7491), .ZN(n7493) );
  AOI22_X1 U8674 ( .A1(n7825), .A2(\adder_stage1[2][7] ), .B1(n7511), .B2(
        n7493), .ZN(n7494) );
  INV_X1 U8675 ( .A(n7494), .ZN(n10029) );
  AOI22_X1 U8676 ( .A1(n8330), .A2(\x_mult_f[4][0] ), .B1(n7511), .B2(
        \x_mult_f_int[4][0] ), .ZN(n7495) );
  INV_X1 U8677 ( .A(n7495), .ZN(n9301) );
  NAND2_X1 U8678 ( .A1(n8223), .A2(n7496), .ZN(n7498) );
  NAND2_X1 U8679 ( .A1(n7498), .A2(n7497), .ZN(n7502) );
  NAND2_X1 U8680 ( .A1(n7500), .A2(n7499), .ZN(n7501) );
  XNOR2_X1 U8681 ( .A(n7502), .B(n7501), .ZN(n7503) );
  AOI22_X1 U8682 ( .A1(n7512), .A2(\adder_stage1[2][12] ), .B1(n7511), .B2(
        n7503), .ZN(n7504) );
  INV_X1 U8683 ( .A(n7504), .ZN(n10024) );
  AOI22_X1 U8684 ( .A1(n7512), .A2(\x_mult_f[5][1] ), .B1(n7511), .B2(
        \x_mult_f_int[5][1] ), .ZN(n7505) );
  INV_X1 U8685 ( .A(n7505), .ZN(n9302) );
  AOI22_X1 U8686 ( .A1(n4713), .A2(\x_mult_f[4][1] ), .B1(n7511), .B2(
        \x_mult_f_int[4][1] ), .ZN(n7506) );
  INV_X1 U8687 ( .A(n7506), .ZN(n9300) );
  NAND2_X1 U8688 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  XNOR2_X1 U8689 ( .A(n8223), .B(n7509), .ZN(n7510) );
  AOI22_X1 U8690 ( .A1(n7512), .A2(\adder_stage1[2][10] ), .B1(n7511), .B2(
        n7510), .ZN(n7513) );
  INV_X1 U8691 ( .A(n7513), .ZN(n10026) );
  INV_X1 U8692 ( .A(n7514), .ZN(n7562) );
  INV_X1 U8693 ( .A(n7515), .ZN(n7560) );
  INV_X1 U8694 ( .A(n7559), .ZN(n7516) );
  AOI21_X1 U8695 ( .B1(n7562), .B2(n7560), .A(n7516), .ZN(n7521) );
  INV_X1 U8696 ( .A(n7517), .ZN(n7519) );
  NAND2_X1 U8697 ( .A1(n7519), .A2(n7518), .ZN(n7520) );
  XOR2_X1 U8698 ( .A(n7521), .B(n7520), .Z(n7522) );
  AOI22_X1 U8699 ( .A1(n5544), .A2(\adder_stage1[0][5] ), .B1(n8399), .B2(
        n7522), .ZN(n7523) );
  INV_X1 U8700 ( .A(n7523), .ZN(n10065) );
  OR2_X1 U8701 ( .A1(\x_mult_f[18][0] ), .A2(\x_mult_f[19][0] ), .ZN(n7524) );
  AND2_X1 U8702 ( .A1(n7524), .A2(n7688), .ZN(n7525) );
  AOI22_X1 U8703 ( .A1(n7910), .A2(\adder_stage1[9][0] ), .B1(n7698), .B2(
        n7525), .ZN(n7526) );
  INV_X1 U8704 ( .A(n7526), .ZN(n9921) );
  AOI21_X1 U8705 ( .B1(n7664), .B2(n7632), .A(n7527), .ZN(n7531) );
  NAND2_X1 U8706 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  XOR2_X1 U8707 ( .A(n7531), .B(n7530), .Z(n7532) );
  AOI22_X1 U8708 ( .A1(n6581), .A2(\adder_stage1[0][9] ), .B1(n6699), .B2(
        n7532), .ZN(n7533) );
  INV_X1 U8709 ( .A(n7533), .ZN(n10061) );
  NAND2_X1 U8710 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  XNOR2_X1 U8711 ( .A(n7537), .B(n7536), .ZN(n7538) );
  AOI22_X1 U8712 ( .A1(n6581), .A2(\adder_stage2[4][14] ), .B1(n7698), .B2(
        n7538), .ZN(n7539) );
  INV_X1 U8713 ( .A(n7539), .ZN(n9723) );
  AOI21_X1 U8714 ( .B1(n7562), .B2(n7541), .A(n7540), .ZN(n7583) );
  OAI21_X1 U8715 ( .B1(n7583), .B2(n7579), .A(n7580), .ZN(n7546) );
  INV_X1 U8716 ( .A(n7542), .ZN(n7544) );
  NAND2_X1 U8717 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  XNOR2_X1 U8718 ( .A(n7546), .B(n7545), .ZN(n7547) );
  AOI22_X1 U8719 ( .A1(n6428), .A2(\adder_stage1[0][7] ), .B1(n7698), .B2(
        n7547), .ZN(n7548) );
  INV_X1 U8720 ( .A(n7548), .ZN(n10063) );
  AOI21_X1 U8721 ( .B1(n7551), .B2(n7550), .A(n7549), .ZN(n7611) );
  OAI21_X1 U8722 ( .B1(n7611), .B2(n7607), .A(n7608), .ZN(n7556) );
  INV_X1 U8723 ( .A(n7552), .ZN(n7554) );
  NAND2_X1 U8724 ( .A1(n7554), .A2(n7553), .ZN(n7555) );
  XNOR2_X1 U8725 ( .A(n7556), .B(n7555), .ZN(n7557) );
  AOI22_X1 U8726 ( .A1(n7613), .A2(\adder_stage2[4][7] ), .B1(n7698), .B2(
        n7557), .ZN(n7558) );
  INV_X1 U8727 ( .A(n7558), .ZN(n9730) );
  NAND2_X1 U8728 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  XNOR2_X1 U8729 ( .A(n7562), .B(n7561), .ZN(n7563) );
  AOI22_X1 U8730 ( .A1(n8094), .A2(\adder_stage1[0][4] ), .B1(n8390), .B2(
        n7563), .ZN(n7564) );
  INV_X1 U8731 ( .A(n7564), .ZN(n10066) );
  INV_X1 U8732 ( .A(n7565), .ZN(n7591) );
  OAI21_X1 U8733 ( .B1(n7591), .B2(n7587), .A(n7588), .ZN(n7570) );
  INV_X1 U8734 ( .A(n7566), .ZN(n7568) );
  NAND2_X1 U8735 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  XNOR2_X1 U8736 ( .A(n7570), .B(n7569), .ZN(n7571) );
  AOI22_X1 U8737 ( .A1(n8059), .A2(\adder_stage1[0][3] ), .B1(n8114), .B2(
        n7571), .ZN(n7572) );
  INV_X1 U8738 ( .A(n7572), .ZN(n10067) );
  NAND2_X1 U8739 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  XNOR2_X1 U8740 ( .A(n7576), .B(n7575), .ZN(n7577) );
  AOI22_X1 U8741 ( .A1(n7818), .A2(\adder_stage1[0][12] ), .B1(n6523), .B2(
        n7577), .ZN(n7578) );
  INV_X1 U8742 ( .A(n7578), .ZN(n10058) );
  INV_X1 U8743 ( .A(n7579), .ZN(n7581) );
  NAND2_X1 U8744 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  XOR2_X1 U8745 ( .A(n7583), .B(n7582), .Z(n7584) );
  AOI22_X1 U8746 ( .A1(n5909), .A2(\adder_stage1[0][6] ), .B1(n8318), .B2(
        n7584), .ZN(n7585) );
  INV_X1 U8747 ( .A(n7585), .ZN(n10064) );
  AOI22_X1 U8748 ( .A1(n7818), .A2(\x_mult_f[1][1] ), .B1(n7909), .B2(
        \x_mult_f_int[1][1] ), .ZN(n7586) );
  INV_X1 U8749 ( .A(n7586), .ZN(n9294) );
  INV_X1 U8750 ( .A(n7587), .ZN(n7589) );
  NAND2_X1 U8751 ( .A1(n7589), .A2(n7588), .ZN(n7590) );
  XOR2_X1 U8752 ( .A(n7591), .B(n7590), .Z(n7592) );
  AOI22_X1 U8753 ( .A1(n7793), .A2(\adder_stage1[0][2] ), .B1(n6256), .B2(
        n7592), .ZN(n8790) );
  NAND2_X1 U8754 ( .A1(n7636), .A2(n7593), .ZN(n7595) );
  AND2_X1 U8755 ( .A1(n7595), .A2(n7594), .ZN(n7617) );
  NAND2_X1 U8756 ( .A1(n7596), .A2(n7615), .ZN(n7597) );
  XOR2_X1 U8757 ( .A(n7617), .B(n7597), .Z(n7598) );
  AOI22_X1 U8758 ( .A1(n6428), .A2(\adder_stage2[4][11] ), .B1(n7698), .B2(
        n7598), .ZN(n7599) );
  INV_X1 U8759 ( .A(n7599), .ZN(n9726) );
  NAND2_X1 U8760 ( .A1(n7664), .A2(n7600), .ZN(n7601) );
  NAND2_X1 U8761 ( .A1(n7601), .A2(n7662), .ZN(n7604) );
  NAND2_X1 U8762 ( .A1(n7602), .A2(n7660), .ZN(n7603) );
  XNOR2_X1 U8763 ( .A(n7604), .B(n7603), .ZN(n7605) );
  AOI22_X1 U8764 ( .A1(n7910), .A2(\adder_stage1[0][10] ), .B1(n7774), .B2(
        n7605), .ZN(n7606) );
  INV_X1 U8765 ( .A(n7606), .ZN(n10060) );
  INV_X1 U8766 ( .A(n7607), .ZN(n7609) );
  NAND2_X1 U8767 ( .A1(n7609), .A2(n7608), .ZN(n7610) );
  XOR2_X1 U8768 ( .A(n7611), .B(n7610), .Z(n7612) );
  AOI22_X1 U8769 ( .A1(n7613), .A2(\adder_stage2[4][6] ), .B1(n7698), .B2(
        n7612), .ZN(n7614) );
  INV_X1 U8770 ( .A(n7614), .ZN(n9731) );
  OAI21_X1 U8771 ( .B1(n7617), .B2(n7616), .A(n7615), .ZN(n7621) );
  NAND2_X1 U8772 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  XNOR2_X1 U8773 ( .A(n7621), .B(n7620), .ZN(n7622) );
  AOI22_X1 U8774 ( .A1(n5909), .A2(\adder_stage2[4][12] ), .B1(n7698), .B2(
        n7622), .ZN(n7623) );
  INV_X1 U8775 ( .A(n7623), .ZN(n9725) );
  INV_X1 U8776 ( .A(n7624), .ZN(n7626) );
  NAND2_X1 U8777 ( .A1(n7626), .A2(n7625), .ZN(n7627) );
  XOR2_X1 U8778 ( .A(n7628), .B(n7627), .Z(n7629) );
  AOI22_X1 U8779 ( .A1(n5273), .A2(\adder_stage2[4][13] ), .B1(n7698), .B2(
        n7629), .ZN(n7630) );
  INV_X1 U8780 ( .A(n7630), .ZN(n9724) );
  NAND2_X1 U8781 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  XNOR2_X1 U8782 ( .A(n7664), .B(n7633), .ZN(n7634) );
  AOI22_X1 U8783 ( .A1(n5909), .A2(\adder_stage1[0][8] ), .B1(n7284), .B2(
        n7634), .ZN(n7635) );
  INV_X1 U8784 ( .A(n7635), .ZN(n10062) );
  INV_X1 U8785 ( .A(n7636), .ZN(n7656) );
  OAI21_X1 U8786 ( .B1(n7656), .B2(n7638), .A(n7637), .ZN(n7643) );
  INV_X1 U8787 ( .A(n7639), .ZN(n7641) );
  NAND2_X1 U8788 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  XNOR2_X1 U8789 ( .A(n7643), .B(n7642), .ZN(n7644) );
  AOI22_X1 U8790 ( .A1(n8383), .A2(\adder_stage2[4][10] ), .B1(n7698), .B2(
        n7644), .ZN(n7645) );
  INV_X1 U8791 ( .A(n7645), .ZN(n9727) );
  OAI21_X1 U8792 ( .B1(n7656), .B2(n7646), .A(n7653), .ZN(n7650) );
  NAND2_X1 U8793 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  XNOR2_X1 U8794 ( .A(n7650), .B(n7649), .ZN(n7651) );
  AOI22_X1 U8795 ( .A1(n8048), .A2(\adder_stage2[4][9] ), .B1(n7698), .B2(
        n7651), .ZN(n7652) );
  INV_X1 U8796 ( .A(n7652), .ZN(n9728) );
  NAND2_X1 U8797 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  XOR2_X1 U8798 ( .A(n7656), .B(n7655), .Z(n7657) );
  AOI22_X1 U8799 ( .A1(n8154), .A2(\adder_stage2[4][8] ), .B1(n7698), .B2(
        n7657), .ZN(n7658) );
  INV_X1 U8800 ( .A(n7658), .ZN(n9729) );
  INV_X1 U8801 ( .A(n7659), .ZN(n7665) );
  OAI21_X1 U8802 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7663) );
  AOI21_X1 U8803 ( .B1(n7665), .B2(n7664), .A(n7663), .ZN(n7669) );
  NAND2_X1 U8804 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  XOR2_X1 U8805 ( .A(n7669), .B(n7668), .Z(n7670) );
  AOI22_X1 U8806 ( .A1(n7818), .A2(\adder_stage1[0][11] ), .B1(n6643), .B2(
        n7670), .ZN(n7671) );
  INV_X1 U8807 ( .A(n7671), .ZN(n10059) );
  INV_X1 U8808 ( .A(n7672), .ZN(n7674) );
  NAND2_X1 U8809 ( .A1(n7674), .A2(n7673), .ZN(n7676) );
  XOR2_X1 U8810 ( .A(n7676), .B(n7675), .Z(n7677) );
  AOI22_X1 U8811 ( .A1(n7793), .A2(\adder_stage1[0][1] ), .B1(n5908), .B2(
        n7677), .ZN(n7678) );
  INV_X1 U8812 ( .A(n7678), .ZN(n10068) );
  NAND2_X1 U8813 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  XNOR2_X1 U8814 ( .A(n7682), .B(n7681), .ZN(n7683) );
  AOI22_X1 U8815 ( .A1(n8364), .A2(\adder_stage1[9][4] ), .B1(n7698), .B2(
        n7683), .ZN(n7684) );
  INV_X1 U8816 ( .A(n7684), .ZN(n9917) );
  INV_X1 U8817 ( .A(n7685), .ZN(n7687) );
  NAND2_X1 U8818 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  XOR2_X1 U8819 ( .A(n7689), .B(n7688), .Z(n7690) );
  AOI22_X1 U8820 ( .A1(n8215), .A2(\adder_stage1[9][1] ), .B1(n7698), .B2(
        n7690), .ZN(n7691) );
  INV_X1 U8821 ( .A(n7691), .ZN(n9920) );
  INV_X1 U8822 ( .A(n7692), .ZN(n7694) );
  NAND2_X1 U8823 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  XOR2_X1 U8824 ( .A(n7696), .B(n7695), .Z(n7697) );
  AOI22_X1 U8825 ( .A1(n8155), .A2(\adder_stage1[9][2] ), .B1(n7698), .B2(
        n7697), .ZN(n7699) );
  INV_X1 U8826 ( .A(n7699), .ZN(n9919) );
  BUF_X2 U8827 ( .A(n6955), .Z(n7774) );
  AOI21_X1 U8828 ( .B1(n3429), .B2(n7770), .A(n7700), .ZN(n7704) );
  NAND2_X1 U8829 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  XOR2_X1 U8830 ( .A(n7704), .B(n7703), .Z(n7705) );
  AOI22_X1 U8831 ( .A1(n7775), .A2(\adder_stage1[8][9] ), .B1(n7774), .B2(
        n7705), .ZN(n7706) );
  INV_X1 U8832 ( .A(n7706), .ZN(n9929) );
  AOI22_X1 U8833 ( .A1(n7767), .A2(\x_mult_f[18][4] ), .B1(n7774), .B2(
        \x_mult_f_int[18][4] ), .ZN(n7707) );
  INV_X1 U8834 ( .A(n7707), .ZN(n9165) );
  INV_X1 U8835 ( .A(n7708), .ZN(n7765) );
  INV_X1 U8836 ( .A(n7709), .ZN(n7763) );
  INV_X1 U8837 ( .A(n7762), .ZN(n7710) );
  AOI21_X1 U8838 ( .B1(n7765), .B2(n7763), .A(n7710), .ZN(n7715) );
  INV_X1 U8839 ( .A(n7711), .ZN(n7713) );
  NAND2_X1 U8840 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  XOR2_X1 U8841 ( .A(n7715), .B(n7714), .Z(n7716) );
  AOI22_X1 U8842 ( .A1(n7767), .A2(\adder_stage1[8][5] ), .B1(n7774), .B2(
        n7716), .ZN(n7717) );
  INV_X1 U8843 ( .A(n7717), .ZN(n9933) );
  INV_X1 U8844 ( .A(n7718), .ZN(n7759) );
  OAI21_X1 U8845 ( .B1(n7759), .B2(n7755), .A(n7756), .ZN(n7723) );
  INV_X1 U8846 ( .A(n7719), .ZN(n7721) );
  NAND2_X1 U8847 ( .A1(n7721), .A2(n7720), .ZN(n7722) );
  XNOR2_X1 U8848 ( .A(n7723), .B(n7722), .ZN(n7724) );
  AOI22_X1 U8849 ( .A1(n7767), .A2(\adder_stage1[8][3] ), .B1(n7774), .B2(
        n7724), .ZN(n7725) );
  INV_X1 U8850 ( .A(n7725), .ZN(n9935) );
  AOI22_X1 U8851 ( .A1(n7767), .A2(\x_mult_f[18][3] ), .B1(n7774), .B2(
        \x_mult_f_int[18][3] ), .ZN(n7726) );
  INV_X1 U8852 ( .A(n7726), .ZN(n9166) );
  AOI22_X1 U8853 ( .A1(n7767), .A2(\x_mult_f[18][1] ), .B1(n7774), .B2(
        \x_mult_f_int[18][1] ), .ZN(n7727) );
  INV_X1 U8854 ( .A(n7727), .ZN(n9328) );
  OR2_X1 U8855 ( .A1(\x_mult_f[16][0] ), .A2(\x_mult_f[17][0] ), .ZN(n7728) );
  AND2_X1 U8856 ( .A1(n7728), .A2(n7751), .ZN(n7729) );
  AOI22_X1 U8857 ( .A1(n7767), .A2(\adder_stage1[8][0] ), .B1(n7774), .B2(
        n7729), .ZN(n7730) );
  INV_X1 U8858 ( .A(n7730), .ZN(n9938) );
  AOI22_X1 U8859 ( .A1(n7767), .A2(\x_mult_f[18][2] ), .B1(n7774), .B2(
        \x_mult_f_int[18][2] ), .ZN(n7731) );
  INV_X1 U8860 ( .A(n7731), .ZN(n9167) );
  AOI21_X1 U8861 ( .B1(n7765), .B2(n7733), .A(n7732), .ZN(n7745) );
  OAI21_X1 U8862 ( .B1(n7745), .B2(n7741), .A(n7742), .ZN(n7738) );
  INV_X1 U8863 ( .A(n7734), .ZN(n7736) );
  NAND2_X1 U8864 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  XNOR2_X1 U8865 ( .A(n7738), .B(n7737), .ZN(n7739) );
  AOI22_X1 U8866 ( .A1(n7775), .A2(\adder_stage1[8][7] ), .B1(n7774), .B2(
        n7739), .ZN(n7740) );
  INV_X1 U8867 ( .A(n7740), .ZN(n9931) );
  INV_X1 U8868 ( .A(n7741), .ZN(n7743) );
  NAND2_X1 U8869 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  XOR2_X1 U8870 ( .A(n7745), .B(n7744), .Z(n7746) );
  AOI22_X1 U8871 ( .A1(n7775), .A2(\adder_stage1[8][6] ), .B1(n7774), .B2(
        n7746), .ZN(n7747) );
  INV_X1 U8872 ( .A(n7747), .ZN(n9932) );
  INV_X1 U8873 ( .A(n7748), .ZN(n7750) );
  NAND2_X1 U8874 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  XOR2_X1 U8875 ( .A(n7752), .B(n7751), .Z(n7753) );
  AOI22_X1 U8876 ( .A1(n7767), .A2(\adder_stage1[8][1] ), .B1(n7774), .B2(
        n7753), .ZN(n7754) );
  INV_X1 U8877 ( .A(n7754), .ZN(n9937) );
  INV_X1 U8878 ( .A(n7755), .ZN(n7757) );
  NAND2_X1 U8879 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  XOR2_X1 U8880 ( .A(n7759), .B(n7758), .Z(n7760) );
  AOI22_X1 U8881 ( .A1(n7767), .A2(\adder_stage1[8][2] ), .B1(n7774), .B2(
        n7760), .ZN(n7761) );
  INV_X1 U8882 ( .A(n7761), .ZN(n9936) );
  NAND2_X1 U8883 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  XNOR2_X1 U8884 ( .A(n7765), .B(n7764), .ZN(n7766) );
  AOI22_X1 U8885 ( .A1(n7767), .A2(\adder_stage1[8][4] ), .B1(n7774), .B2(
        n7766), .ZN(n7768) );
  INV_X1 U8886 ( .A(n7768), .ZN(n9934) );
  NAND2_X1 U8887 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  XNOR2_X1 U8888 ( .A(n3429), .B(n7771), .ZN(n7773) );
  AOI22_X1 U8889 ( .A1(n7775), .A2(\adder_stage1[8][8] ), .B1(n7774), .B2(
        n7773), .ZN(n7776) );
  INV_X1 U8890 ( .A(n7776), .ZN(n9930) );
  OAI21_X1 U8891 ( .B1(n7779), .B2(n7778), .A(n7777), .ZN(n7784) );
  INV_X1 U8892 ( .A(n7780), .ZN(n7782) );
  NAND2_X1 U8893 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  XNOR2_X1 U8894 ( .A(n7784), .B(n7783), .ZN(n7785) );
  AOI22_X1 U8895 ( .A1(n7793), .A2(\adder_stage2[2][3] ), .B1(n8390), .B2(
        n7785), .ZN(n7786) );
  INV_X1 U8896 ( .A(n7786), .ZN(n9768) );
  INV_X1 U8897 ( .A(n7787), .ZN(n7789) );
  NAND2_X1 U8898 ( .A1(n7789), .A2(n7788), .ZN(n7791) );
  XOR2_X1 U8899 ( .A(n7791), .B(n7790), .Z(n7792) );
  AOI22_X1 U8900 ( .A1(n7793), .A2(\adder_stage2[2][1] ), .B1(n8390), .B2(
        n7792), .ZN(n7794) );
  INV_X1 U8901 ( .A(n7794), .ZN(n9770) );
  INV_X1 U8902 ( .A(n7795), .ZN(n7823) );
  OAI21_X1 U8903 ( .B1(n7823), .B2(n7796), .A(n7820), .ZN(n7800) );
  NAND2_X1 U8904 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  XNOR2_X1 U8905 ( .A(n7800), .B(n7799), .ZN(n7801) );
  AOI22_X1 U8906 ( .A1(n7818), .A2(\adder_stage2[2][9] ), .B1(n8390), .B2(
        n7801), .ZN(n7802) );
  INV_X1 U8907 ( .A(n7802), .ZN(n9762) );
  INV_X1 U8908 ( .A(n7803), .ZN(n7805) );
  NAND2_X1 U8909 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  XOR2_X1 U8910 ( .A(n7807), .B(n7806), .Z(n7808) );
  AOI22_X1 U8911 ( .A1(n7818), .A2(\adder_stage2[2][6] ), .B1(n7909), .B2(
        n7808), .ZN(n7809) );
  INV_X1 U8912 ( .A(n7809), .ZN(n9765) );
  OAI21_X1 U8913 ( .B1(n7823), .B2(n7811), .A(n7810), .ZN(n7816) );
  INV_X1 U8914 ( .A(n7812), .ZN(n7814) );
  NAND2_X1 U8915 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  XNOR2_X1 U8916 ( .A(n7816), .B(n7815), .ZN(n7817) );
  AOI22_X1 U8917 ( .A1(n7818), .A2(\adder_stage2[2][10] ), .B1(n7909), .B2(
        n7817), .ZN(n7819) );
  INV_X1 U8918 ( .A(n7819), .ZN(n9761) );
  NAND2_X1 U8919 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  XOR2_X1 U8920 ( .A(n7823), .B(n7822), .Z(n7824) );
  AOI22_X1 U8921 ( .A1(n7825), .A2(\adder_stage2[2][8] ), .B1(n8390), .B2(
        n7824), .ZN(n7826) );
  INV_X1 U8922 ( .A(n7826), .ZN(n9763) );
  NAND2_X1 U8923 ( .A1(n7827), .A2(n7841), .ZN(n7828) );
  XOR2_X1 U8924 ( .A(n7843), .B(n7828), .Z(n7829) );
  AOI22_X1 U8925 ( .A1(n6581), .A2(\adder_stage2[2][11] ), .B1(n8390), .B2(
        n7829), .ZN(n7830) );
  INV_X1 U8926 ( .A(n7830), .ZN(n9760) );
  NOR2_X1 U8927 ( .A1(n7843), .A2(n7831), .ZN(n7834) );
  INV_X1 U8928 ( .A(n7832), .ZN(n7833) );
  NOR2_X1 U8929 ( .A1(n7834), .A2(n7833), .ZN(n7838) );
  NAND2_X1 U8930 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  XOR2_X1 U8931 ( .A(n7838), .B(n7837), .Z(n7839) );
  AOI22_X1 U8932 ( .A1(n7512), .A2(\adder_stage2[2][13] ), .B1(n8390), .B2(
        n7839), .ZN(n7840) );
  INV_X1 U8933 ( .A(n7840), .ZN(n9758) );
  OAI21_X1 U8934 ( .B1(n7843), .B2(n7842), .A(n7841), .ZN(n7847) );
  NAND2_X1 U8935 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  XNOR2_X1 U8936 ( .A(n7847), .B(n7846), .ZN(n7848) );
  AOI22_X1 U8937 ( .A1(n7825), .A2(\adder_stage2[2][12] ), .B1(n7909), .B2(
        n7848), .ZN(n7849) );
  INV_X1 U8938 ( .A(n7849), .ZN(n9759) );
  AOI22_X1 U8939 ( .A1(n7851), .A2(\x_mult_f[12][1] ), .B1(n8390), .B2(
        \x_mult_f_int[12][1] ), .ZN(n7850) );
  INV_X1 U8940 ( .A(n7850), .ZN(n9316) );
  AOI22_X1 U8941 ( .A1(n7851), .A2(\x_mult_f[12][2] ), .B1(n8390), .B2(
        \x_mult_f_int[12][2] ), .ZN(n7852) );
  INV_X1 U8942 ( .A(n7852), .ZN(n9084) );
  INV_X1 U8943 ( .A(n7853), .ZN(n7888) );
  INV_X1 U8944 ( .A(n7854), .ZN(n7878) );
  NAND2_X1 U8945 ( .A1(n7878), .A2(n7876), .ZN(n7855) );
  XNOR2_X1 U8946 ( .A(n7888), .B(n7855), .ZN(n7856) );
  AOI22_X1 U8947 ( .A1(n7910), .A2(\adder_stage1[6][4] ), .B1(n7909), .B2(
        n7856), .ZN(n7857) );
  INV_X1 U8948 ( .A(n7857), .ZN(n9968) );
  INV_X1 U8949 ( .A(n7858), .ZN(n7860) );
  NAND2_X1 U8950 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  XOR2_X1 U8951 ( .A(n7861), .B(n7872), .Z(n7862) );
  AOI22_X1 U8952 ( .A1(n7910), .A2(\adder_stage1[6][1] ), .B1(n7909), .B2(
        n7862), .ZN(n7863) );
  INV_X1 U8953 ( .A(n7863), .ZN(n9971) );
  INV_X1 U8954 ( .A(n7864), .ZN(n7907) );
  OAI21_X1 U8955 ( .B1(n7907), .B2(n7903), .A(n7904), .ZN(n7869) );
  INV_X1 U8956 ( .A(n7865), .ZN(n7867) );
  NAND2_X1 U8957 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  XNOR2_X1 U8958 ( .A(n7869), .B(n7868), .ZN(n7870) );
  AOI22_X1 U8959 ( .A1(n7910), .A2(\adder_stage1[6][3] ), .B1(n7909), .B2(
        n7870), .ZN(n7871) );
  INV_X1 U8960 ( .A(n7871), .ZN(n9969) );
  OR2_X1 U8961 ( .A1(\x_mult_f[12][0] ), .A2(\x_mult_f[13][0] ), .ZN(n7873) );
  AND2_X1 U8962 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  AOI22_X1 U8963 ( .A1(n7910), .A2(\adder_stage1[6][0] ), .B1(n7909), .B2(
        n7874), .ZN(n7875) );
  INV_X1 U8964 ( .A(n7875), .ZN(n9972) );
  INV_X1 U8965 ( .A(n7876), .ZN(n7877) );
  AOI21_X1 U8966 ( .B1(n7888), .B2(n7878), .A(n7877), .ZN(n7883) );
  INV_X1 U8967 ( .A(n7879), .ZN(n7881) );
  NAND2_X1 U8968 ( .A1(n7881), .A2(n7880), .ZN(n7882) );
  XOR2_X1 U8969 ( .A(n7883), .B(n7882), .Z(n7884) );
  AOI22_X1 U8970 ( .A1(n7910), .A2(\adder_stage1[6][5] ), .B1(n7909), .B2(
        n7884), .ZN(n7885) );
  INV_X1 U8971 ( .A(n7885), .ZN(n9967) );
  AOI21_X1 U8972 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7895) );
  INV_X1 U8973 ( .A(n7894), .ZN(n7889) );
  NAND2_X1 U8974 ( .A1(n7889), .A2(n7893), .ZN(n7890) );
  XOR2_X1 U8975 ( .A(n7895), .B(n7890), .Z(n7891) );
  AOI22_X1 U8976 ( .A1(n7910), .A2(\adder_stage1[6][6] ), .B1(n7909), .B2(
        n7891), .ZN(n7892) );
  INV_X1 U8977 ( .A(n7892), .ZN(n9966) );
  OAI21_X1 U8978 ( .B1(n7895), .B2(n7894), .A(n7893), .ZN(n7900) );
  INV_X1 U8979 ( .A(n7896), .ZN(n7898) );
  NAND2_X1 U8980 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  XNOR2_X1 U8981 ( .A(n7900), .B(n7899), .ZN(n7901) );
  AOI22_X1 U8982 ( .A1(n7910), .A2(\adder_stage1[6][7] ), .B1(n7909), .B2(
        n7901), .ZN(n7902) );
  INV_X1 U8983 ( .A(n7902), .ZN(n9965) );
  INV_X1 U8984 ( .A(n7903), .ZN(n7905) );
  NAND2_X1 U8985 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  XOR2_X1 U8986 ( .A(n7907), .B(n7906), .Z(n7908) );
  AOI22_X1 U8987 ( .A1(n7910), .A2(\adder_stage1[6][2] ), .B1(n7909), .B2(
        n7908), .ZN(n7911) );
  INV_X1 U8988 ( .A(n7911), .ZN(n9970) );
  FA_X1 U8989 ( .A(n8704), .B(n3482), .CI(n7912), .CO(n7913), .S(n3654) );
  INV_X1 U8990 ( .A(n7913), .ZN(n7914) );
  AOI22_X1 U8991 ( .A1(n7914), .A2(n7454), .B1(n8048), .B2(
        \adder_stage1[13][20] ), .ZN(n7915) );
  INV_X1 U8992 ( .A(n7915), .ZN(n9840) );
  NAND2_X1 U8993 ( .A1(\x_mult_f[3][15] ), .A2(\x_mult_f[2][15] ), .ZN(n7916)
         );
  NAND2_X1 U8994 ( .A1(n7917), .A2(n7916), .ZN(n7919) );
  NAND2_X1 U8995 ( .A1(n3476), .A2(n3451), .ZN(n7918) );
  INV_X1 U8996 ( .A(n7920), .ZN(n10037) );
  INV_X1 U8997 ( .A(n7921), .ZN(n8159) );
  AOI21_X1 U8998 ( .B1(n3431), .B2(n8160), .A(n8159), .ZN(n7924) );
  NOR2_X1 U8999 ( .A1(\adder_stage2[6][19] ), .A2(\adder_stage2[7][19] ), .ZN(
        n8163) );
  INV_X1 U9000 ( .A(n8163), .ZN(n7922) );
  NAND2_X1 U9001 ( .A1(\adder_stage2[6][19] ), .A2(\adder_stage2[7][19] ), 
        .ZN(n8162) );
  NAND2_X1 U9002 ( .A1(n7922), .A2(n8162), .ZN(n7923) );
  XOR2_X1 U9003 ( .A(n7924), .B(n7923), .Z(n7925) );
  AOI22_X1 U9004 ( .A1(n7925), .A2(n8213), .B1(n8200), .B2(
        \adder_stage3[3][19] ), .ZN(n7926) );
  INV_X1 U9005 ( .A(n7926), .ZN(n9590) );
  INV_X1 U9006 ( .A(n8278), .ZN(n7927) );
  NAND2_X1 U9007 ( .A1(n7927), .A2(n7931), .ZN(n8268) );
  INV_X1 U9008 ( .A(n8279), .ZN(n7930) );
  INV_X1 U9009 ( .A(n7928), .ZN(n7929) );
  AOI21_X1 U9010 ( .B1(n7931), .B2(n7930), .A(n7929), .ZN(n8271) );
  NOR2_X1 U9011 ( .A1(\adder_stage3[2][19] ), .A2(\adder_stage3[3][19] ), .ZN(
        n8270) );
  INV_X1 U9012 ( .A(n8270), .ZN(n7933) );
  NAND2_X1 U9013 ( .A1(\adder_stage3[2][19] ), .A2(\adder_stage3[3][19] ), 
        .ZN(n8269) );
  NAND2_X1 U9014 ( .A1(n7933), .A2(n8269), .ZN(n7934) );
  XOR2_X1 U9015 ( .A(n7935), .B(n7934), .Z(n7936) );
  AOI22_X1 U9016 ( .A1(n7936), .A2(n8037), .B1(n8381), .B2(
        \adder_stage4[1][19] ), .ZN(n7937) );
  INV_X1 U9017 ( .A(n7937), .ZN(n9548) );
  FA_X1 U9018 ( .A(n3453), .B(n3483), .CI(n7938), .CO(n7939), .S(n3603) );
  INV_X1 U9019 ( .A(n7939), .ZN(n7940) );
  AOI22_X1 U9020 ( .A1(n7940), .A2(n7029), .B1(n8059), .B2(
        \adder_stage1[7][20] ), .ZN(n7941) );
  INV_X1 U9021 ( .A(n7941), .ZN(n9939) );
  FA_X1 U9022 ( .A(n3477), .B(n8705), .CI(n7942), .CO(n7943), .S(n3552) );
  INV_X1 U9023 ( .A(n7943), .ZN(n7945) );
  AOI22_X1 U9024 ( .A1(n7945), .A2(n8390), .B1(n7944), .B2(
        \adder_stage1[14][20] ), .ZN(n7946) );
  INV_X1 U9025 ( .A(n7946), .ZN(n9823) );
  FA_X1 U9026 ( .A(\x_mult_f[8][14] ), .B(\x_mult_f[9][14] ), .CI(n7947), .CO(
        n8384), .S(n3909) );
  NAND2_X1 U9027 ( .A1(n7948), .A2(n8387), .ZN(n7950) );
  NAND2_X1 U9028 ( .A1(n8386), .A2(\adder_stage1[4][15] ), .ZN(n7949) );
  NAND2_X1 U9029 ( .A1(n7950), .A2(n7949), .ZN(n9990) );
  FA_X1 U9030 ( .A(\x_mult_f[30][14] ), .B(\x_mult_f[31][14] ), .CI(n7951), 
        .CO(n8068), .S(n5690) );
  NAND2_X1 U9031 ( .A1(n7952), .A2(n8229), .ZN(n7954) );
  NAND2_X1 U9032 ( .A1(n8364), .A2(\adder_stage1[15][15] ), .ZN(n7953) );
  NAND2_X1 U9033 ( .A1(n7954), .A2(n7953), .ZN(n9807) );
  NAND2_X1 U9034 ( .A1(n7958), .A2(n8213), .ZN(n7960) );
  NAND2_X1 U9035 ( .A1(n8215), .A2(\adder_stage2[0][16] ), .ZN(n7959) );
  NAND2_X1 U9036 ( .A1(n7960), .A2(n7959), .ZN(n9789) );
  FA_X1 U9037 ( .A(\x_mult_f[16][14] ), .B(\x_mult_f[17][14] ), .CI(n7961), 
        .CO(n8110), .S(n5435) );
  INV_X1 U9038 ( .A(n7962), .ZN(n7963) );
  NAND2_X1 U9039 ( .A1(n7963), .A2(n8401), .ZN(n7965) );
  NAND2_X1 U9040 ( .A1(n8386), .A2(\adder_stage1[8][20] ), .ZN(n7964) );
  NAND2_X1 U9041 ( .A1(n7965), .A2(n7964), .ZN(n9922) );
  FA_X1 U9042 ( .A(n3478), .B(n8698), .CI(n7966), .CO(n5190), .S(n7967) );
  NAND2_X1 U9043 ( .A1(n7967), .A2(n8229), .ZN(n7969) );
  NAND2_X1 U9044 ( .A1(n8400), .A2(\adder_stage1[2][15] ), .ZN(n7968) );
  NAND2_X1 U9045 ( .A1(n7969), .A2(n7968), .ZN(n10022) );
  FA_X1 U9046 ( .A(\adder_stage1[12][15] ), .B(\adder_stage1[13][15] ), .CI(
        n7970), .CO(n8142), .S(n5306) );
  NAND2_X1 U9047 ( .A1(n7971), .A2(n8216), .ZN(n7973) );
  NAND2_X1 U9048 ( .A1(n8215), .A2(\adder_stage2[6][16] ), .ZN(n7972) );
  NAND2_X1 U9049 ( .A1(n7973), .A2(n7972), .ZN(n9687) );
  FA_X1 U9050 ( .A(\x_mult_f[12][14] ), .B(\x_mult_f[13][14] ), .CI(n7974), 
        .CO(n8062), .S(n5355) );
  INV_X1 U9051 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U9052 ( .A1(n7976), .A2(n4002), .ZN(n7978) );
  NAND2_X1 U9053 ( .A1(n8046), .A2(\adder_stage1[6][20] ), .ZN(n7977) );
  NAND2_X1 U9054 ( .A1(n7978), .A2(n7977), .ZN(n9956) );
  FA_X1 U9055 ( .A(\x_mult_f[6][14] ), .B(\x_mult_f[7][14] ), .CI(n7979), .CO(
        n8072), .S(n5805) );
  NAND2_X1 U9056 ( .A1(n7980), .A2(n7356), .ZN(n7982) );
  NAND2_X1 U9057 ( .A1(n8094), .A2(\adder_stage1[3][15] ), .ZN(n7981) );
  NAND2_X1 U9058 ( .A1(n7982), .A2(n7981), .ZN(n10005) );
  FA_X1 U9059 ( .A(\adder_stage1[4][15] ), .B(\adder_stage1[5][15] ), .CI(
        n7983), .CO(n8116), .S(n4180) );
  NAND2_X1 U9060 ( .A1(n7984), .A2(n8203), .ZN(n7986) );
  NAND2_X1 U9061 ( .A1(n8088), .A2(\adder_stage2[2][16] ), .ZN(n7985) );
  NAND2_X1 U9062 ( .A1(n7986), .A2(n7985), .ZN(n9755) );
  FA_X1 U9063 ( .A(n3454), .B(n3484), .CI(n7987), .CO(n3894), .S(n7988) );
  NAND2_X1 U9064 ( .A1(n7988), .A2(n8186), .ZN(n7990) );
  NAND2_X1 U9065 ( .A1(n8088), .A2(\adder_stage1[5][15] ), .ZN(n7989) );
  NAND2_X1 U9066 ( .A1(n7990), .A2(n7989), .ZN(n9974) );
  AOI22_X1 U9067 ( .A1(n6330), .A2(\x_mult_f[25][2] ), .B1(n7117), .B2(
        \x_mult_f_int[25][2] ), .ZN(n7991) );
  INV_X1 U9068 ( .A(n7991), .ZN(n9229) );
  AOI22_X1 U9069 ( .A1(n5294), .A2(\x_mult_f[15][3] ), .B1(n7992), .B2(
        \x_mult_f_int[15][3] ), .ZN(n7993) );
  INV_X1 U9070 ( .A(n7993), .ZN(n9125) );
  AOI22_X1 U9071 ( .A1(n7997), .A2(n8365), .B1(n8215), .B2(
        \adder_stage2[7][16] ), .ZN(n7998) );
  INV_X1 U9072 ( .A(n7998), .ZN(n9670) );
  OAI21_X1 U9073 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(n8003) );
  XOR2_X1 U9074 ( .A(\adder_stage2[3][20] ), .B(\adder_stage2[2][20] ), .Z(
        n8002) );
  XOR2_X1 U9075 ( .A(n8003), .B(n8002), .Z(n8005) );
  AND2_X1 U9076 ( .A1(n8178), .A2(\adder_stage3[1][20] ), .ZN(n8004) );
  AOI21_X1 U9077 ( .B1(n8005), .B2(n8398), .A(n8004), .ZN(n8006) );
  INV_X1 U9078 ( .A(n8006), .ZN(n9630) );
  FA_X1 U9079 ( .A(n3455), .B(n3485), .CI(n8007), .CO(n8008), .S(n7997) );
  INV_X1 U9080 ( .A(n8008), .ZN(n8009) );
  NAND2_X1 U9081 ( .A1(n8009), .A2(n3950), .ZN(n8010) );
  OAI21_X1 U9082 ( .B1(n8141), .B2(n8720), .A(n8010), .ZN(n1912) );
  OAI21_X1 U9083 ( .B1(n8141), .B2(n8721), .A(n8010), .ZN(n1911) );
  OAI21_X1 U9084 ( .B1(n8141), .B2(n8722), .A(n8010), .ZN(n1910) );
  OAI21_X1 U9085 ( .B1(n8136), .B2(n8751), .A(n8010), .ZN(n1909) );
  AOI22_X1 U9086 ( .A1(\x_mult_f_int[27][13] ), .A2(n4002), .B1(n8228), .B2(
        \x_mult_f[27][13] ), .ZN(n8011) );
  INV_X1 U9087 ( .A(n8011), .ZN(n9236) );
  AOI22_X1 U9088 ( .A1(\x_mult_f_int[27][12] ), .A2(n4002), .B1(n8391), .B2(
        \x_mult_f[27][12] ), .ZN(n8012) );
  INV_X1 U9089 ( .A(n8012), .ZN(n9237) );
  AOI22_X1 U9090 ( .A1(\x_mult_f_int[17][15] ), .A2(n8180), .B1(n8048), .B2(
        \x_mult_f[17][15] ), .ZN(n8013) );
  INV_X1 U9091 ( .A(n8013), .ZN(n9140) );
  AOI22_X1 U9092 ( .A1(\x_mult_f_int[8][13] ), .A2(n5908), .B1(n7775), .B2(
        \x_mult_f[8][13] ), .ZN(n8014) );
  INV_X1 U9093 ( .A(n8014), .ZN(n9029) );
  AOI22_X1 U9094 ( .A1(\x_mult_f_int[13][13] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][13] ), .ZN(n8015) );
  INV_X1 U9095 ( .A(n8015), .ZN(n9087) );
  FA_X1 U9096 ( .A(n3456), .B(n3486), .CI(n8016), .CO(n8017), .S(n3637) );
  INV_X1 U9097 ( .A(n8017), .ZN(n8018) );
  AOI22_X1 U9098 ( .A1(n8018), .A2(n7356), .B1(n4713), .B2(
        \adder_stage1[9][20] ), .ZN(n8019) );
  INV_X1 U9099 ( .A(n8019), .ZN(n9905) );
  AOI22_X1 U9100 ( .A1(\x_mult_f_int[22][12] ), .A2(n8401), .B1(n7825), .B2(
        \x_mult_f[22][12] ), .ZN(n8755) );
  AOI22_X1 U9101 ( .A1(\x_mult_f_int[7][13] ), .A2(n7774), .B1(n8178), .B2(
        \x_mult_f[7][13] ), .ZN(n8020) );
  INV_X1 U9102 ( .A(n8020), .ZN(n9015) );
  AOI22_X1 U9103 ( .A1(\x_mult_f_int[7][12] ), .A2(n8180), .B1(n8178), .B2(
        \x_mult_f[7][12] ), .ZN(n8021) );
  INV_X1 U9104 ( .A(n8021), .ZN(n9016) );
  AOI22_X1 U9105 ( .A1(\x_mult_f_int[7][15] ), .A2(n8399), .B1(n8178), .B2(
        \x_mult_f[7][15] ), .ZN(n8022) );
  INV_X1 U9106 ( .A(n8022), .ZN(n9013) );
  AOI22_X1 U9107 ( .A1(\x_mult_f_int[17][14] ), .A2(n8180), .B1(n8218), .B2(
        \x_mult_f[17][14] ), .ZN(n8023) );
  INV_X1 U9108 ( .A(n8023), .ZN(n9141) );
  AOI22_X1 U9109 ( .A1(\x_mult_f_int[17][12] ), .A2(n8180), .B1(n8157), .B2(
        \x_mult_f[17][12] ), .ZN(n8024) );
  INV_X1 U9110 ( .A(n8024), .ZN(n9143) );
  AOI22_X1 U9111 ( .A1(\x_mult_f_int[6][13] ), .A2(n8365), .B1(n8212), .B2(
        \x_mult_f[6][13] ), .ZN(n8025) );
  INV_X1 U9112 ( .A(n8025), .ZN(n9001) );
  AOI22_X1 U9113 ( .A1(\x_mult_f_int[6][12] ), .A2(n8203), .B1(n8212), .B2(
        \x_mult_f[6][12] ), .ZN(n8026) );
  INV_X1 U9114 ( .A(n8026), .ZN(n9002) );
  AOI22_X1 U9115 ( .A1(\x_mult_f_int[18][13] ), .A2(n5950), .B1(n8200), .B2(
        \x_mult_f[18][13] ), .ZN(n8027) );
  INV_X1 U9116 ( .A(n8027), .ZN(n9156) );
  AOI22_X1 U9117 ( .A1(\x_mult_f_int[18][12] ), .A2(n8399), .B1(n8212), .B2(
        \x_mult_f[18][12] ), .ZN(n8028) );
  INV_X1 U9118 ( .A(n8028), .ZN(n9157) );
  AOI22_X1 U9119 ( .A1(\x_mult_f_int[3][14] ), .A2(n8203), .B1(n8202), .B2(
        \x_mult_f[3][14] ), .ZN(n8029) );
  INV_X1 U9120 ( .A(n8029), .ZN(n8962) );
  AOI22_X1 U9121 ( .A1(\x_mult_f_int[4][13] ), .A2(n8365), .B1(n8215), .B2(
        \x_mult_f[4][13] ), .ZN(n8030) );
  INV_X1 U9122 ( .A(n8030), .ZN(n8976) );
  AOI22_X1 U9123 ( .A1(\x_mult_f_int[14][13] ), .A2(n8399), .B1(n8094), .B2(
        \x_mult_f[14][13] ), .ZN(n8031) );
  INV_X1 U9124 ( .A(n8031), .ZN(n9101) );
  AOI22_X1 U9125 ( .A1(\x_mult_f_int[30][13] ), .A2(n7992), .B1(n8218), .B2(
        \x_mult_f[30][13] ), .ZN(n8032) );
  INV_X1 U9126 ( .A(n8032), .ZN(n9266) );
  AOI22_X1 U9127 ( .A1(\x_mult_f_int[10][13] ), .A2(n8216), .B1(n8395), .B2(
        \x_mult_f[10][13] ), .ZN(n8033) );
  INV_X1 U9128 ( .A(n8033), .ZN(n9048) );
  AOI22_X1 U9129 ( .A1(\x_mult_f_int[10][12] ), .A2(n8216), .B1(n8392), .B2(
        \x_mult_f[10][12] ), .ZN(n8034) );
  INV_X1 U9130 ( .A(n8034), .ZN(n9049) );
  AOI22_X1 U9131 ( .A1(\x_mult_f_int[1][12] ), .A2(n7774), .B1(n8036), .B2(
        \x_mult_f[1][12] ), .ZN(n8035) );
  INV_X1 U9132 ( .A(n8035), .ZN(n8938) );
  AOI22_X1 U9133 ( .A1(\x_mult_f_int[5][12] ), .A2(n8037), .B1(n8036), .B2(
        \x_mult_f[5][12] ), .ZN(n8038) );
  INV_X1 U9134 ( .A(n8038), .ZN(n8988) );
  AOI22_X1 U9135 ( .A1(\x_mult_f_int[23][14] ), .A2(n6523), .B1(n8154), .B2(
        \x_mult_f[23][14] ), .ZN(n8756) );
  AOI22_X1 U9136 ( .A1(\x_mult_f_int[23][13] ), .A2(n6256), .B1(n8094), .B2(
        \x_mult_f[23][13] ), .ZN(n8757) );
  AOI22_X1 U9137 ( .A1(\x_mult_f_int[24][12] ), .A2(n8213), .B1(n8395), .B2(
        \x_mult_f[24][12] ), .ZN(n8758) );
  AOI22_X1 U9138 ( .A1(\x_mult_f_int[23][12] ), .A2(n5950), .B1(n8094), .B2(
        \x_mult_f[23][12] ), .ZN(n8039) );
  INV_X1 U9139 ( .A(n8039), .ZN(n9205) );
  AOI22_X1 U9140 ( .A1(\x_mult_f_int[24][13] ), .A2(n8213), .B1(n8212), .B2(
        \x_mult_f[24][13] ), .ZN(n8040) );
  INV_X1 U9141 ( .A(n8040), .ZN(n9218) );
  AOI22_X1 U9142 ( .A1(\x_mult_f_int[10][14] ), .A2(n8216), .B1(n8200), .B2(
        \x_mult_f[10][14] ), .ZN(n8041) );
  INV_X1 U9143 ( .A(n8041), .ZN(n9047) );
  AOI22_X1 U9144 ( .A1(\x_mult_f_int[3][13] ), .A2(n8203), .B1(n8202), .B2(
        \x_mult_f[3][13] ), .ZN(n8042) );
  INV_X1 U9145 ( .A(n8042), .ZN(n8963) );
  AOI22_X1 U9146 ( .A1(\x_mult_f_int[25][12] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][12] ), .ZN(n8759) );
  AOI22_X1 U9147 ( .A1(\x_mult_f_int[25][13] ), .A2(n8398), .B1(n8400), .B2(
        \x_mult_f[25][13] ), .ZN(n8760) );
  AOI22_X1 U9148 ( .A1(\x_mult_f_int[22][13] ), .A2(n8401), .B1(n8395), .B2(
        \x_mult_f[22][13] ), .ZN(n8761) );
  AOI22_X1 U9149 ( .A1(\x_mult_f_int[5][14] ), .A2(n8203), .B1(n8391), .B2(
        \x_mult_f[5][14] ), .ZN(n8762) );
  AOI22_X1 U9150 ( .A1(\x_mult_f_int[13][14] ), .A2(n8189), .B1(n8212), .B2(
        \x_mult_f[13][14] ), .ZN(n8043) );
  INV_X1 U9151 ( .A(n8043), .ZN(n9086) );
  AOI22_X1 U9152 ( .A1(\x_mult_f_int[17][13] ), .A2(n8180), .B1(n8048), .B2(
        \x_mult_f[17][13] ), .ZN(n8044) );
  INV_X1 U9153 ( .A(n8044), .ZN(n9142) );
  AOI22_X1 U9154 ( .A1(\x_mult_f_int[8][12] ), .A2(n8150), .B1(n7285), .B2(
        \x_mult_f[8][12] ), .ZN(n8045) );
  INV_X1 U9155 ( .A(n8045), .ZN(n9030) );
  AOI22_X1 U9156 ( .A1(\x_mult_f_int[13][12] ), .A2(n8189), .B1(n8046), .B2(
        \x_mult_f[13][12] ), .ZN(n8047) );
  INV_X1 U9157 ( .A(n8047), .ZN(n9088) );
  AOI22_X1 U9158 ( .A1(\x_mult_f_int[4][12] ), .A2(n8365), .B1(n8048), .B2(
        \x_mult_f[4][12] ), .ZN(n8049) );
  INV_X1 U9159 ( .A(n8049), .ZN(n8977) );
  AOI22_X1 U9160 ( .A1(\x_mult_f_int[14][12] ), .A2(n8399), .B1(n8386), .B2(
        \x_mult_f[14][12] ), .ZN(n8050) );
  INV_X1 U9161 ( .A(n8050), .ZN(n9102) );
  AOI22_X1 U9162 ( .A1(\x_mult_f_int[30][12] ), .A2(n8150), .B1(n8218), .B2(
        \x_mult_f[30][12] ), .ZN(n8051) );
  INV_X1 U9163 ( .A(n8051), .ZN(n9267) );
  AOI22_X1 U9164 ( .A1(\x_mult_f_int[3][12] ), .A2(n8203), .B1(n8202), .B2(
        \x_mult_f[3][12] ), .ZN(n8052) );
  INV_X1 U9165 ( .A(n8052), .ZN(n8964) );
  AOI22_X1 U9166 ( .A1(\x_mult_f_int[1][13] ), .A2(n7284), .B1(n6373), .B2(
        \x_mult_f[1][13] ), .ZN(n8053) );
  INV_X1 U9167 ( .A(n8053), .ZN(n8937) );
  AOI22_X1 U9168 ( .A1(\x_mult_f_int[5][13] ), .A2(n8203), .B1(n8048), .B2(
        \x_mult_f[5][13] ), .ZN(n8763) );
  AOI22_X1 U9169 ( .A1(\x_mult_f_int[6][14] ), .A2(n8365), .B1(n8212), .B2(
        \x_mult_f[6][14] ), .ZN(n8054) );
  INV_X1 U9170 ( .A(n8054), .ZN(n9000) );
  AOI22_X1 U9171 ( .A1(\x_mult_f_int[31][12] ), .A2(n6915), .B1(n8202), .B2(
        \x_mult_f[31][12] ), .ZN(n8055) );
  INV_X1 U9172 ( .A(n8055), .ZN(n9281) );
  AOI22_X1 U9173 ( .A1(\x_mult_f_int[31][13] ), .A2(n8194), .B1(n7944), .B2(
        \x_mult_f[31][13] ), .ZN(n8056) );
  INV_X1 U9174 ( .A(n8056), .ZN(n9280) );
  AOI22_X1 U9175 ( .A1(\x_mult_f_int[20][12] ), .A2(n7511), .B1(n8381), .B2(
        \x_mult_f[20][12] ), .ZN(n8764) );
  AOI22_X1 U9176 ( .A1(\x_mult_f_int[26][13] ), .A2(n8208), .B1(n7613), .B2(
        \x_mult_f[26][13] ), .ZN(n8765) );
  AOI22_X1 U9177 ( .A1(\x_mult_f_int[12][11] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][11] ), .ZN(n8057) );
  INV_X1 U9178 ( .A(n8057), .ZN(n9076) );
  AOI22_X1 U9179 ( .A1(\x_mult_f_int[24][14] ), .A2(n8213), .B1(n8212), .B2(
        \x_mult_f[24][14] ), .ZN(n8058) );
  INV_X1 U9180 ( .A(n8058), .ZN(n9217) );
  AOI22_X1 U9181 ( .A1(\x_mult_f_int[15][14] ), .A2(n8208), .B1(n8059), .B2(
        \x_mult_f[15][14] ), .ZN(n8060) );
  INV_X1 U9182 ( .A(n8060), .ZN(n9114) );
  AOI22_X1 U9183 ( .A1(\x_mult_f_int[31][14] ), .A2(n6221), .B1(n8154), .B2(
        \x_mult_f[31][14] ), .ZN(n8061) );
  INV_X1 U9184 ( .A(n8061), .ZN(n9279) );
  FA_X1 U9185 ( .A(n3457), .B(n3487), .CI(n8062), .CO(n7975), .S(n8063) );
  AOI22_X1 U9186 ( .A1(n8063), .A2(n4002), .B1(n8155), .B2(
        \adder_stage1[6][15] ), .ZN(n8064) );
  INV_X1 U9187 ( .A(n8064), .ZN(n9957) );
  AOI22_X1 U9188 ( .A1(\x_mult_f_int[21][14] ), .A2(n8189), .B1(n8392), .B2(
        \x_mult_f[21][14] ), .ZN(n8065) );
  INV_X1 U9189 ( .A(n8065), .ZN(n9189) );
  AOI22_X1 U9190 ( .A1(\x_mult_f_int[11][12] ), .A2(n8186), .B1(n8048), .B2(
        \x_mult_f[11][12] ), .ZN(n8066) );
  INV_X1 U9191 ( .A(n8066), .ZN(n9061) );
  AOI22_X1 U9192 ( .A1(\x_mult_f_int[21][13] ), .A2(n6643), .B1(n8392), .B2(
        \x_mult_f[21][13] ), .ZN(n8067) );
  INV_X1 U9193 ( .A(n8067), .ZN(n9190) );
  AOI22_X1 U9194 ( .A1(\x_mult_f_int[20][13] ), .A2(n8180), .B1(n8381), .B2(
        \x_mult_f[20][13] ), .ZN(n8766) );
  FA_X1 U9195 ( .A(n3458), .B(n3488), .CI(n8068), .CO(n8069), .S(n7952) );
  INV_X1 U9196 ( .A(n8069), .ZN(n8070) );
  AOI22_X1 U9197 ( .A1(n8070), .A2(n8229), .B1(n8364), .B2(
        \adder_stage1[15][20] ), .ZN(n8071) );
  INV_X1 U9198 ( .A(n8071), .ZN(n9806) );
  FA_X1 U9199 ( .A(n3459), .B(n3489), .CI(n8072), .CO(n8073), .S(n7980) );
  INV_X1 U9200 ( .A(n8073), .ZN(n8074) );
  AOI22_X1 U9201 ( .A1(n8074), .A2(n7454), .B1(n8094), .B2(
        \adder_stage1[3][20] ), .ZN(n8075) );
  INV_X1 U9202 ( .A(n8075), .ZN(n10004) );
  FA_X1 U9203 ( .A(n8701), .B(n8702), .CI(n8076), .CO(n8077), .S(n3620) );
  INV_X1 U9204 ( .A(n8077), .ZN(n8079) );
  AOI22_X1 U9205 ( .A1(n8079), .A2(n5950), .B1(n8078), .B2(
        \adder_stage1[11][20] ), .ZN(n8080) );
  INV_X1 U9206 ( .A(n8080), .ZN(n9874) );
  AOI22_X1 U9207 ( .A1(\x_mult_f_int[28][14] ), .A2(n8216), .B1(n8215), .B2(
        \x_mult_f[28][14] ), .ZN(n8081) );
  INV_X1 U9208 ( .A(n8081), .ZN(n9248) );
  AOI22_X1 U9209 ( .A1(\x_mult_f_int[0][14] ), .A2(n7909), .B1(n8391), .B2(
        \x_mult_f[0][14] ), .ZN(n8082) );
  INV_X1 U9210 ( .A(n8082), .ZN(n8926) );
  AOI22_X1 U9211 ( .A1(\x_mult_f_int[16][14] ), .A2(n8265), .B1(n4713), .B2(
        \x_mult_f[16][14] ), .ZN(n8083) );
  INV_X1 U9212 ( .A(n8083), .ZN(n9128) );
  AOI22_X1 U9213 ( .A1(\x_mult_f_int[7][14] ), .A2(n8208), .B1(n8178), .B2(
        \x_mult_f[7][14] ), .ZN(n8084) );
  INV_X1 U9214 ( .A(n8084), .ZN(n9014) );
  AOI22_X1 U9215 ( .A1(\x_mult_f_int[0][13] ), .A2(n7117), .B1(n8228), .B2(
        \x_mult_f[0][13] ), .ZN(n8085) );
  INV_X1 U9216 ( .A(n8085), .ZN(n8927) );
  AOI22_X1 U9217 ( .A1(\x_mult_f_int[26][12] ), .A2(n8399), .B1(n7030), .B2(
        \x_mult_f[26][12] ), .ZN(n8767) );
  AOI22_X1 U9218 ( .A1(\x_mult_f_int[14][14] ), .A2(n8399), .B1(n8381), .B2(
        \x_mult_f[14][14] ), .ZN(n8086) );
  INV_X1 U9219 ( .A(n8086), .ZN(n9100) );
  FA_X1 U9220 ( .A(\adder_stage1[6][15] ), .B(\adder_stage1[7][15] ), .CI(
        n8087), .CO(n8128), .S(n4214) );
  AOI22_X1 U9221 ( .A1(n8089), .A2(n8114), .B1(n8088), .B2(
        \adder_stage2[3][16] ), .ZN(n8090) );
  INV_X1 U9222 ( .A(n8090), .ZN(n9738) );
  AOI22_X1 U9223 ( .A1(\x_mult_f_int[23][15] ), .A2(n8318), .B1(n8400), .B2(
        \x_mult_f[23][15] ), .ZN(n8768) );
  AOI22_X1 U9224 ( .A1(\x_mult_f_int[18][14] ), .A2(n8398), .B1(n8383), .B2(
        \x_mult_f[18][14] ), .ZN(n8096) );
  INV_X1 U9225 ( .A(n8096), .ZN(n9155) );
  AOI22_X1 U9226 ( .A1(\x_mult_f_int[4][14] ), .A2(n8365), .B1(n8215), .B2(
        \x_mult_f[4][14] ), .ZN(n8097) );
  INV_X1 U9227 ( .A(n8097), .ZN(n8975) );
  AOI22_X1 U9228 ( .A1(\x_mult_f_int[9][14] ), .A2(n8213), .B1(n8157), .B2(
        \x_mult_f[9][14] ), .ZN(n8769) );
  AOI22_X1 U9229 ( .A1(\x_mult_f_int[29][14] ), .A2(n8365), .B1(n8154), .B2(
        \x_mult_f[29][14] ), .ZN(n8770) );
  AOI22_X1 U9230 ( .A1(\x_mult_f_int[19][13] ), .A2(n7909), .B1(n8157), .B2(
        \x_mult_f[19][13] ), .ZN(n8098) );
  INV_X1 U9231 ( .A(n8098), .ZN(n9170) );
  AOI22_X1 U9232 ( .A1(\x_mult_f_int[30][14] ), .A2(n7698), .B1(n8218), .B2(
        \x_mult_f[30][14] ), .ZN(n8099) );
  INV_X1 U9233 ( .A(n8099), .ZN(n9265) );
  AOI22_X1 U9234 ( .A1(\x_mult_f_int[8][14] ), .A2(n8150), .B1(n7775), .B2(
        \x_mult_f[8][14] ), .ZN(n8100) );
  INV_X1 U9235 ( .A(n8100), .ZN(n9028) );
  AOI22_X1 U9236 ( .A1(\x_mult_f_int[19][12] ), .A2(n7110), .B1(n8157), .B2(
        \x_mult_f[19][12] ), .ZN(n8101) );
  INV_X1 U9237 ( .A(n8101), .ZN(n9171) );
  AOI22_X1 U9238 ( .A1(\x_mult_f_int[19][14] ), .A2(n8180), .B1(n8157), .B2(
        \x_mult_f[19][14] ), .ZN(n8102) );
  INV_X1 U9239 ( .A(n8102), .ZN(n9169) );
  AOI22_X1 U9240 ( .A1(\x_mult_f_int[29][12] ), .A2(n8282), .B1(n8154), .B2(
        \x_mult_f[29][12] ), .ZN(n8103) );
  INV_X1 U9241 ( .A(n8103), .ZN(n9253) );
  AOI22_X1 U9242 ( .A1(\x_mult_f_int[9][12] ), .A2(n8265), .B1(n8383), .B2(
        \x_mult_f[9][12] ), .ZN(n8771) );
  AOI22_X1 U9243 ( .A1(\x_mult_f_int[9][13] ), .A2(n8387), .B1(n8383), .B2(
        \x_mult_f[9][13] ), .ZN(n8772) );
  FA_X1 U9244 ( .A(\adder_stage1[8][15] ), .B(\adder_stage1[9][15] ), .CI(
        n8104), .CO(n8132), .S(n5988) );
  AOI22_X1 U9245 ( .A1(n8105), .A2(n5950), .B1(n7030), .B2(
        \adder_stage2[4][16] ), .ZN(n8106) );
  INV_X1 U9246 ( .A(n8106), .ZN(n9721) );
  FA_X1 U9247 ( .A(\adder_stage1[2][15] ), .B(\adder_stage1[3][15] ), .CI(
        n8107), .CO(n8124), .S(n6080) );
  AOI22_X1 U9248 ( .A1(n8108), .A2(n7698), .B1(n8395), .B2(
        \adder_stage2[1][16] ), .ZN(n8109) );
  INV_X1 U9249 ( .A(n8109), .ZN(n9772) );
  FA_X1 U9250 ( .A(n3460), .B(n3490), .CI(n8110), .CO(n7962), .S(n8111) );
  AOI22_X1 U9251 ( .A1(n8111), .A2(n8037), .B1(n8386), .B2(
        \adder_stage1[8][15] ), .ZN(n8112) );
  INV_X1 U9252 ( .A(n8112), .ZN(n9923) );
  AOI22_X1 U9253 ( .A1(\x_mult_f_int[12][12] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][12] ), .ZN(n8113) );
  INV_X1 U9254 ( .A(n8113), .ZN(n9075) );
  AOI22_X1 U9255 ( .A1(\x_mult_f_int[12][13] ), .A2(n8114), .B1(n8155), .B2(
        \x_mult_f[12][13] ), .ZN(n8115) );
  INV_X1 U9256 ( .A(n8115), .ZN(n9074) );
  FA_X1 U9257 ( .A(n8707), .B(n3491), .CI(n8116), .CO(n8117), .S(n7984) );
  INV_X1 U9258 ( .A(n8117), .ZN(n8118) );
  NAND2_X1 U9259 ( .A1(n8118), .A2(n6645), .ZN(n8119) );
  OAI21_X1 U9260 ( .B1(n8141), .B2(n8732), .A(n8119), .ZN(n2017) );
  OAI21_X1 U9261 ( .B1(n8136), .B2(n8733), .A(n8119), .ZN(n2016) );
  OAI21_X1 U9262 ( .B1(n8141), .B2(n8734), .A(n8119), .ZN(n2015) );
  OAI21_X1 U9263 ( .B1(n8136), .B2(n8747), .A(n8119), .ZN(n2014) );
  AOI22_X1 U9264 ( .A1(\x_mult_f_int[26][14] ), .A2(n8208), .B1(n8212), .B2(
        \x_mult_f[26][14] ), .ZN(n8773) );
  FA_X1 U9265 ( .A(n3479), .B(n8706), .CI(n8120), .CO(n8121), .S(n7958) );
  INV_X1 U9266 ( .A(n8121), .ZN(n8122) );
  NAND2_X1 U9267 ( .A1(n8122), .A2(n7511), .ZN(n8123) );
  OAI21_X1 U9268 ( .B1(n8136), .B2(n8735), .A(n8123), .ZN(n2059) );
  OAI21_X1 U9269 ( .B1(n8141), .B2(n8736), .A(n8123), .ZN(n2058) );
  OAI21_X1 U9270 ( .B1(n8136), .B2(n8737), .A(n3432), .ZN(n2057) );
  OAI21_X1 U9271 ( .B1(n8136), .B2(n8748), .A(n3432), .ZN(n2056) );
  FA_X1 U9272 ( .A(n3461), .B(n3492), .CI(n8124), .CO(n8125), .S(n8108) );
  INV_X1 U9273 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U9274 ( .A1(n8126), .A2(n6699), .ZN(n8127) );
  OAI21_X1 U9275 ( .B1(n8141), .B2(n8752), .A(n8127), .ZN(n2035) );
  OAI21_X1 U9276 ( .B1(n8136), .B2(n8723), .A(n8127), .ZN(n2038) );
  OAI21_X1 U9277 ( .B1(n8141), .B2(n8724), .A(n8127), .ZN(n2037) );
  OAI21_X1 U9278 ( .B1(n8136), .B2(n8725), .A(n8127), .ZN(n2036) );
  FA_X1 U9279 ( .A(n3464), .B(n3493), .CI(n8128), .CO(n8129), .S(n8089) );
  INV_X1 U9280 ( .A(n8129), .ZN(n8130) );
  NAND2_X1 U9281 ( .A1(n8130), .A2(n3950), .ZN(n8131) );
  OAI21_X1 U9282 ( .B1(n8136), .B2(n8726), .A(n8131), .ZN(n1996) );
  OAI21_X1 U9283 ( .B1(n8136), .B2(n8727), .A(n8131), .ZN(n1995) );
  OAI21_X1 U9284 ( .B1(n8136), .B2(n8728), .A(n8131), .ZN(n1994) );
  OAI21_X1 U9285 ( .B1(n8136), .B2(n8753), .A(n8131), .ZN(n1993) );
  FA_X1 U9286 ( .A(n3465), .B(n3494), .CI(n8132), .CO(n8133), .S(n8105) );
  INV_X1 U9287 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9288 ( .A1(n8134), .A2(n6955), .ZN(n8135) );
  OAI21_X1 U9289 ( .B1(n8136), .B2(n8749), .A(n8135), .ZN(n1972) );
  OAI21_X1 U9290 ( .B1(n8141), .B2(n8738), .A(n8135), .ZN(n1975) );
  OAI21_X1 U9291 ( .B1(n8141), .B2(n8739), .A(n8135), .ZN(n1974) );
  OAI21_X1 U9292 ( .B1(n8136), .B2(n8740), .A(n8135), .ZN(n1973) );
  FA_X1 U9293 ( .A(n8708), .B(n3495), .CI(n8137), .CO(n8138), .S(n8095) );
  INV_X1 U9294 ( .A(n8138), .ZN(n8139) );
  NAND2_X1 U9295 ( .A1(n8139), .A2(n3950), .ZN(n8140) );
  OAI21_X1 U9296 ( .B1(n8141), .B2(n8729), .A(n8140), .ZN(n1954) );
  OAI21_X1 U9297 ( .B1(n8141), .B2(n8730), .A(n8140), .ZN(n1953) );
  OAI21_X1 U9298 ( .B1(n8141), .B2(n8731), .A(n8140), .ZN(n1952) );
  OAI21_X1 U9299 ( .B1(n8141), .B2(n8754), .A(n8140), .ZN(n1951) );
  NAND2_X1 U9300 ( .A1(n3413), .A2(n3950), .ZN(n8143) );
  OAI21_X1 U9301 ( .B1(n8136), .B2(n8750), .A(n8143), .ZN(n1930) );
  OAI21_X1 U9302 ( .B1(n8141), .B2(n8741), .A(n8143), .ZN(n1933) );
  OAI21_X1 U9303 ( .B1(n8136), .B2(n8742), .A(n8143), .ZN(n1932) );
  OAI21_X1 U9304 ( .B1(n8141), .B2(n8743), .A(n8143), .ZN(n1931) );
  FA_X1 U9305 ( .A(n3480), .B(n8703), .CI(n8144), .CO(n8145), .S(n3569) );
  INV_X1 U9306 ( .A(n8145), .ZN(n8146) );
  AOI22_X1 U9307 ( .A1(n8146), .A2(n8208), .B1(n8202), .B2(
        \adder_stage1[12][20] ), .ZN(n8147) );
  INV_X1 U9308 ( .A(n8147), .ZN(n9857) );
  AOI22_X1 U9309 ( .A1(\x_mult_f_int[20][14] ), .A2(n7774), .B1(n8381), .B2(
        \x_mult_f[20][14] ), .ZN(n8774) );
  FA_X1 U9310 ( .A(n3463), .B(n3497), .CI(n8148), .CO(n4584), .S(n8151) );
  AND2_X1 U9311 ( .A1(n8200), .A2(\adder_stage1[0][15] ), .ZN(n8149) );
  AOI21_X1 U9312 ( .B1(n8151), .B2(n8150), .A(n8149), .ZN(n8152) );
  INV_X1 U9313 ( .A(n8152), .ZN(n10055) );
  AOI22_X1 U9314 ( .A1(\x_mult_f_int[25][14] ), .A2(n8398), .B1(n8400), .B2(
        \x_mult_f[25][14] ), .ZN(n8775) );
  AOI22_X1 U9315 ( .A1(\x_mult_f_int[20][15] ), .A2(n7698), .B1(n8381), .B2(
        \x_mult_f[20][15] ), .ZN(n8776) );
  AOI22_X1 U9316 ( .A1(\x_mult_f_int[25][15] ), .A2(n8398), .B1(n8400), .B2(
        \x_mult_f[25][15] ), .ZN(n8777) );
  AOI22_X1 U9317 ( .A1(\x_mult_f_int[12][14] ), .A2(n8389), .B1(n8155), .B2(
        \x_mult_f[12][14] ), .ZN(n8153) );
  INV_X1 U9318 ( .A(n8153), .ZN(n9073) );
  AOI22_X1 U9319 ( .A1(\x_mult_f_int[22][14] ), .A2(n8401), .B1(n8395), .B2(
        \x_mult_f[22][14] ), .ZN(n8778) );
  AOI22_X1 U9320 ( .A1(\x_mult_f_int[9][15] ), .A2(n8401), .B1(n8157), .B2(
        \x_mult_f[9][15] ), .ZN(n8779) );
  AOI22_X1 U9321 ( .A1(\x_mult_f_int[29][15] ), .A2(n8213), .B1(n8154), .B2(
        \x_mult_f[29][15] ), .ZN(n8780) );
  AOI22_X1 U9322 ( .A1(\x_mult_f_int[12][15] ), .A2(n7110), .B1(n8155), .B2(
        \x_mult_f[12][15] ), .ZN(n8156) );
  INV_X1 U9323 ( .A(n8156), .ZN(n9072) );
  AOI22_X1 U9324 ( .A1(\x_mult_f_int[19][15] ), .A2(n8208), .B1(n8157), .B2(
        \x_mult_f[19][15] ), .ZN(n8158) );
  INV_X1 U9325 ( .A(n8158), .ZN(n9168) );
  AOI21_X1 U9326 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n8164) );
  OAI21_X1 U9327 ( .B1(n8164), .B2(n8163), .A(n8162), .ZN(n8165) );
  XNOR2_X1 U9328 ( .A(n8165), .B(n3500), .ZN(n8166) );
  AND2_X1 U9329 ( .A1(n8167), .A2(n8172), .ZN(n8168) );
  NAND2_X1 U9330 ( .A1(n8169), .A2(n8168), .ZN(n8175) );
  INV_X1 U9331 ( .A(n8170), .ZN(n8171) );
  AOI21_X1 U9332 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8174) );
  NAND2_X1 U9333 ( .A1(n8175), .A2(n8174), .ZN(n8177) );
  XOR2_X1 U9334 ( .A(\adder_stage2[5][20] ), .B(\adder_stage2[4][20] ), .Z(
        n8176) );
  XOR2_X1 U9335 ( .A(n8177), .B(n8176), .Z(n8181) );
  AND2_X1 U9336 ( .A1(n8178), .A2(\adder_stage3[2][20] ), .ZN(n8179) );
  AOI22_X1 U9337 ( .A1(\x_mult_f_int[11][14] ), .A2(n8186), .B1(n8397), .B2(
        \x_mult_f[11][14] ), .ZN(n8183) );
  INV_X1 U9338 ( .A(n8183), .ZN(n9059) );
  AOI22_X1 U9339 ( .A1(\x_mult_f_int[27][14] ), .A2(n4002), .B1(n8228), .B2(
        \x_mult_f[27][14] ), .ZN(n8184) );
  INV_X1 U9340 ( .A(n8184), .ZN(n9235) );
  AOI22_X1 U9341 ( .A1(\x_mult_f_int[1][15] ), .A2(n7992), .B1(n8202), .B2(
        \x_mult_f[1][15] ), .ZN(n8185) );
  INV_X1 U9342 ( .A(n8185), .ZN(n8935) );
  AOI22_X1 U9343 ( .A1(\x_mult_f_int[5][15] ), .A2(n8203), .B1(n8202), .B2(
        \x_mult_f[5][15] ), .ZN(n8781) );
  AOI22_X1 U9344 ( .A1(\x_mult_f_int[11][15] ), .A2(n8186), .B1(n8395), .B2(
        \x_mult_f[11][15] ), .ZN(n8187) );
  INV_X1 U9345 ( .A(n8187), .ZN(n9058) );
  AOI22_X1 U9346 ( .A1(\x_mult_f_int[21][15] ), .A2(n5908), .B1(n8392), .B2(
        \x_mult_f[21][15] ), .ZN(n8188) );
  INV_X1 U9347 ( .A(n8188), .ZN(n9188) );
  AOI22_X1 U9348 ( .A1(\x_mult_f_int[26][15] ), .A2(n8208), .B1(n8078), .B2(
        \x_mult_f[26][15] ), .ZN(n8782) );
  AOI22_X1 U9349 ( .A1(\x_mult_f_int[13][15] ), .A2(n8189), .B1(n8228), .B2(
        \x_mult_f[13][15] ), .ZN(n8190) );
  INV_X1 U9350 ( .A(n8190), .ZN(n9085) );
  AOI22_X1 U9351 ( .A1(\x_mult_f_int[27][15] ), .A2(n4002), .B1(n8228), .B2(
        \x_mult_f[27][15] ), .ZN(n8191) );
  INV_X1 U9352 ( .A(n8191), .ZN(n9234) );
  OR2_X1 U9353 ( .A1(\adder_stage3[2][0] ), .A2(\adder_stage3[3][0] ), .ZN(
        n8192) );
  AND2_X1 U9354 ( .A1(n8192), .A2(n8315), .ZN(n8193) );
  AOI22_X1 U9355 ( .A1(n8195), .A2(\adder_stage4[1][0] ), .B1(n8194), .B2(
        n8193), .ZN(n8196) );
  INV_X1 U9356 ( .A(n8196), .ZN(n9567) );
  AOI22_X1 U9357 ( .A1(\x_mult_f_int[2][15] ), .A2(n8186), .B1(n8215), .B2(
        \x_mult_f[2][15] ), .ZN(n8197) );
  INV_X1 U9358 ( .A(n8197), .ZN(n8947) );
  AOI22_X1 U9359 ( .A1(\x_mult_f_int[4][15] ), .A2(n8365), .B1(n8215), .B2(
        \x_mult_f[4][15] ), .ZN(n8198) );
  INV_X1 U9360 ( .A(n8198), .ZN(n8974) );
  AOI22_X1 U9361 ( .A1(\x_mult_f_int[10][15] ), .A2(n8216), .B1(n7285), .B2(
        \x_mult_f[10][15] ), .ZN(n8199) );
  INV_X1 U9362 ( .A(n8199), .ZN(n9046) );
  AOI22_X1 U9363 ( .A1(\x_mult_f_int[0][15] ), .A2(n8282), .B1(n8200), .B2(
        \x_mult_f[0][15] ), .ZN(n8201) );
  INV_X1 U9364 ( .A(n8201), .ZN(n8925) );
  AOI22_X1 U9365 ( .A1(\x_mult_f_int[3][15] ), .A2(n8203), .B1(n8202), .B2(
        \x_mult_f[3][15] ), .ZN(n8204) );
  INV_X1 U9366 ( .A(n8204), .ZN(n8961) );
  AOI22_X1 U9367 ( .A1(\x_mult_f_int[6][15] ), .A2(n8037), .B1(n8212), .B2(
        \x_mult_f[6][15] ), .ZN(n8205) );
  INV_X1 U9368 ( .A(n8205), .ZN(n8999) );
  AOI22_X1 U9369 ( .A1(\x_mult_f_int[8][15] ), .A2(n8363), .B1(n8195), .B2(
        \x_mult_f[8][15] ), .ZN(n8206) );
  INV_X1 U9370 ( .A(n8206), .ZN(n9027) );
  AOI22_X1 U9371 ( .A1(\x_mult_f_int[14][15] ), .A2(n8399), .B1(n8381), .B2(
        \x_mult_f[14][15] ), .ZN(n8207) );
  INV_X1 U9372 ( .A(n8207), .ZN(n9099) );
  AOI22_X1 U9373 ( .A1(\x_mult_f_int[15][15] ), .A2(n8208), .B1(n8094), .B2(
        \x_mult_f[15][15] ), .ZN(n8209) );
  INV_X1 U9374 ( .A(n8209), .ZN(n9113) );
  AOI22_X1 U9375 ( .A1(\x_mult_f_int[16][15] ), .A2(n8265), .B1(n4891), .B2(
        \x_mult_f[16][15] ), .ZN(n8210) );
  INV_X1 U9376 ( .A(n8210), .ZN(n9127) );
  AOI22_X1 U9377 ( .A1(\x_mult_f_int[18][15] ), .A2(n8387), .B1(n8383), .B2(
        \x_mult_f[18][15] ), .ZN(n8211) );
  INV_X1 U9378 ( .A(n8211), .ZN(n9154) );
  AOI22_X1 U9379 ( .A1(\x_mult_f_int[24][15] ), .A2(n8213), .B1(n8212), .B2(
        \x_mult_f[24][15] ), .ZN(n8214) );
  INV_X1 U9380 ( .A(n8214), .ZN(n9216) );
  AOI22_X1 U9381 ( .A1(\x_mult_f_int[28][15] ), .A2(n8216), .B1(n8215), .B2(
        \x_mult_f[28][15] ), .ZN(n8217) );
  INV_X1 U9382 ( .A(n8217), .ZN(n9247) );
  AOI22_X1 U9383 ( .A1(\x_mult_f_int[30][15] ), .A2(n8213), .B1(n8218), .B2(
        \x_mult_f[30][15] ), .ZN(n8219) );
  INV_X1 U9384 ( .A(n8219), .ZN(n9264) );
  AOI22_X1 U9385 ( .A1(\x_mult_f_int[31][15] ), .A2(n8389), .B1(n8397), .B2(
        \x_mult_f[31][15] ), .ZN(n8220) );
  INV_X1 U9386 ( .A(n8220), .ZN(n9278) );
  AOI22_X1 U9387 ( .A1(\x_mult_f_int[22][15] ), .A2(n8401), .B1(n8395), .B2(
        \x_mult_f[22][15] ), .ZN(n8783) );
  AOI21_X1 U9388 ( .B1(n8223), .B2(n8222), .A(n8221), .ZN(n8227) );
  NAND2_X1 U9389 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  XOR2_X1 U9390 ( .A(n8227), .B(n8226), .Z(n8230) );
  AOI22_X1 U9391 ( .A1(n8230), .A2(n8229), .B1(n8228), .B2(
        \adder_stage1[2][13] ), .ZN(n8231) );
  INV_X1 U9392 ( .A(n8231), .ZN(n10023) );
  AND2_X1 U9393 ( .A1(n8232), .A2(n8236), .ZN(n8373) );
  NOR2_X1 U9394 ( .A1(\adder_stage2[0][18] ), .A2(\adder_stage2[1][18] ), .ZN(
        n8238) );
  INV_X1 U9395 ( .A(n8238), .ZN(n8378) );
  AND2_X1 U9396 ( .A1(n8373), .A2(n8378), .ZN(n8367) );
  OR2_X1 U9397 ( .A1(\adder_stage2[0][19] ), .A2(\adder_stage2[1][19] ), .ZN(
        n8369) );
  AND2_X1 U9398 ( .A1(n8367), .A2(n8369), .ZN(n8233) );
  NAND2_X1 U9399 ( .A1(n8374), .A2(n8233), .ZN(n8241) );
  INV_X1 U9400 ( .A(n8234), .ZN(n8235) );
  AOI21_X1 U9401 ( .B1(n8237), .B2(n8236), .A(n8235), .ZN(n8375) );
  NAND2_X1 U9402 ( .A1(\adder_stage2[0][18] ), .A2(\adder_stage2[1][18] ), 
        .ZN(n8377) );
  OAI21_X1 U9403 ( .B1(n8375), .B2(n8238), .A(n8377), .ZN(n8366) );
  NAND2_X1 U9404 ( .A1(\adder_stage2[0][19] ), .A2(\adder_stage2[1][19] ), 
        .ZN(n8368) );
  INV_X1 U9405 ( .A(n8368), .ZN(n8239) );
  AOI21_X1 U9406 ( .B1(n8366), .B2(n8369), .A(n8239), .ZN(n8240) );
  NAND2_X1 U9407 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  XOR2_X1 U9408 ( .A(\adder_stage2[1][20] ), .B(\adder_stage2[0][20] ), .Z(
        n8242) );
  XOR2_X1 U9409 ( .A(n8243), .B(n8242), .Z(n8245) );
  AND2_X1 U9410 ( .A1(n8392), .A2(\adder_stage3[0][20] ), .ZN(n8244) );
  AOI21_X1 U9411 ( .B1(n8245), .B2(n5950), .A(n8244), .ZN(n8246) );
  INV_X1 U9412 ( .A(n8246), .ZN(n9651) );
  NAND2_X1 U9413 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  XNOR2_X1 U9414 ( .A(n3447), .B(n8249), .ZN(n8251) );
  AOI22_X1 U9415 ( .A1(n7909), .A2(n8251), .B1(n8391), .B2(
        \adder_stage3[3][16] ), .ZN(n8252) );
  INV_X1 U9416 ( .A(n8252), .ZN(n9593) );
  AND2_X1 U9417 ( .A1(n8253), .A2(n8258), .ZN(n8254) );
  NAND2_X1 U9418 ( .A1(n8255), .A2(n8254), .ZN(n8261) );
  INV_X1 U9419 ( .A(n8256), .ZN(n8257) );
  AOI21_X1 U9420 ( .B1(n8259), .B2(n8258), .A(n8257), .ZN(n8260) );
  NAND2_X1 U9421 ( .A1(n8261), .A2(n8260), .ZN(n8263) );
  XOR2_X1 U9422 ( .A(\adder_stage3[1][20] ), .B(\adder_stage3[0][20] ), .Z(
        n8262) );
  XOR2_X1 U9423 ( .A(n8263), .B(n8262), .Z(n8266) );
  AND2_X1 U9424 ( .A1(n8200), .A2(\adder_stage4[0][20] ), .ZN(n8264) );
  AOI21_X1 U9425 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8267) );
  INV_X1 U9426 ( .A(n8267), .ZN(n9568) );
  XNOR2_X1 U9427 ( .A(n8275), .B(n3499), .ZN(n8276) );
  AOI22_X1 U9428 ( .A1(n8276), .A2(n8216), .B1(n7944), .B2(
        \adder_stage4[1][20] ), .ZN(n8277) );
  INV_X1 U9429 ( .A(n8277), .ZN(n9547) );
  NAND2_X1 U9430 ( .A1(n7927), .A2(n8279), .ZN(n8280) );
  XOR2_X1 U9431 ( .A(n8281), .B(n8280), .Z(n8283) );
  AOI22_X1 U9432 ( .A1(n8283), .A2(n8282), .B1(n8391), .B2(
        \adder_stage4[1][17] ), .ZN(n8284) );
  INV_X1 U9433 ( .A(n8284), .ZN(n9550) );
  INV_X1 U9434 ( .A(n8285), .ZN(n8287) );
  NAND2_X1 U9435 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  XOR2_X1 U9436 ( .A(n8289), .B(n8288), .Z(n8290) );
  AOI22_X1 U9437 ( .A1(n7030), .A2(\adder_stage3[0][15] ), .B1(n8291), .B2(
        n8290), .ZN(n8292) );
  INV_X1 U9438 ( .A(n8292), .ZN(n9654) );
  INV_X1 U9439 ( .A(n8293), .ZN(n8294) );
  AOI21_X1 U9440 ( .B1(n8296), .B2(n8295), .A(n8294), .ZN(n8301) );
  INV_X1 U9441 ( .A(n8297), .ZN(n8299) );
  NAND2_X1 U9442 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  XOR2_X1 U9443 ( .A(n8301), .B(n8300), .Z(n8302) );
  AOI22_X1 U9444 ( .A1(n5544), .A2(\adder_stage3[3][11] ), .B1(n7698), .B2(
        n8302), .ZN(n8303) );
  INV_X1 U9445 ( .A(n8303), .ZN(n9598) );
  INV_X1 U9446 ( .A(n8304), .ZN(n8306) );
  NAND2_X1 U9447 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  XOR2_X1 U9448 ( .A(n8308), .B(n8307), .Z(n8309) );
  AOI22_X1 U9449 ( .A1(n7330), .A2(\adder_stage4[0][15] ), .B1(n8310), .B2(
        n8309), .ZN(n8311) );
  INV_X1 U9450 ( .A(n8311), .ZN(n9573) );
  INV_X1 U9451 ( .A(n8312), .ZN(n8314) );
  NAND2_X1 U9452 ( .A1(n8314), .A2(n8313), .ZN(n8316) );
  XOR2_X1 U9453 ( .A(n8316), .B(n8315), .Z(n8317) );
  AOI22_X1 U9454 ( .A1(n7330), .A2(\adder_stage4[1][1] ), .B1(n8318), .B2(
        n8317), .ZN(n8319) );
  INV_X1 U9455 ( .A(n8319), .ZN(n9566) );
  OAI21_X1 U9456 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8327) );
  INV_X1 U9457 ( .A(n8323), .ZN(n8325) );
  NAND2_X1 U9458 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  XNOR2_X1 U9459 ( .A(n8327), .B(n8326), .ZN(n8328) );
  AOI22_X1 U9460 ( .A1(n8330), .A2(\adder_stage4[1][3] ), .B1(n8329), .B2(
        n8328), .ZN(n8331) );
  INV_X1 U9461 ( .A(n8331), .ZN(n9564) );
  NAND2_X1 U9462 ( .A1(n8332), .A2(\ctrl_inst/xmem_tracker [0]), .ZN(n8333) );
  OAI21_X1 U9463 ( .B1(\ctrl_inst/xmem_tracker [0]), .B2(n8667), .A(n8333), 
        .ZN(n3383) );
  AND2_X1 U9464 ( .A1(n8342), .A2(\ctrl_inst/pline_cntr [2]), .ZN(n8334) );
  OR2_X1 U9465 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  NOR2_X1 U9466 ( .A1(n8337), .A2(n8336), .ZN(n8341) );
  INV_X1 U9467 ( .A(n8338), .ZN(n8339) );
  NAND4_X1 U9468 ( .A1(n8344), .A2(\ctrl_inst/pline_cntr [2]), .A3(n8717), 
        .A4(n8339), .ZN(n8340) );
  OAI21_X1 U9469 ( .B1(n8341), .B2(n8717), .A(n8340), .ZN(n3118) );
  NAND3_X1 U9470 ( .A1(n8342), .A2(n8713), .A3(n8349), .ZN(n8690) );
  NAND2_X1 U9471 ( .A1(n8690), .A2(n8343), .ZN(n8345) );
  MUX2_X1 U9472 ( .A(\ctrl_inst/pline_cntr [0]), .B(n8345), .S(n8344), .Z(
        n3121) );
  OAI33_X1 U9473 ( .A1(n8349), .A2(n8348), .A3(n8347), .B1(n8718), .B2(n8346), 
        .B3(reset), .ZN(n3390) );
  MUX2_X1 U9474 ( .A(s_data_in_x[0]), .B(\xmem_data[31][0] ), .S(n8355), .Z(
        n3370) );
  MUX2_X1 U9475 ( .A(\xmem_data[31][0] ), .B(\xmem_data[30][0] ), .S(n8356), 
        .Z(n10310) );
  MUX2_X1 U9476 ( .A(\xmem_data[30][0] ), .B(\xmem_data[29][0] ), .S(n8353), 
        .Z(n10302) );
  MUX2_X1 U9477 ( .A(\xmem_data[29][0] ), .B(\xmem_data[28][0] ), .S(n8354), 
        .Z(n10294) );
  MUX2_X1 U9478 ( .A(\xmem_data[28][0] ), .B(\xmem_data[27][0] ), .S(n8352), 
        .Z(n10286) );
  BUF_X2 U9479 ( .A(n3835), .Z(n8351) );
  MUX2_X1 U9480 ( .A(\xmem_data[27][0] ), .B(\xmem_data[26][0] ), .S(n8351), 
        .Z(n10278) );
  BUF_X2 U9481 ( .A(n3835), .Z(n8352) );
  MUX2_X1 U9482 ( .A(\xmem_data[26][0] ), .B(\xmem_data[25][0] ), .S(n8352), 
        .Z(n10145) );
  MUX2_X1 U9483 ( .A(\xmem_data[25][0] ), .B(\xmem_data[24][0] ), .S(n8351), 
        .Z(n10144) );
  BUF_X2 U9484 ( .A(n3835), .Z(n8354) );
  MUX2_X1 U9485 ( .A(\xmem_data[24][0] ), .B(\xmem_data[23][0] ), .S(n8354), 
        .Z(n10143) );
  MUX2_X1 U9486 ( .A(\xmem_data[23][0] ), .B(\xmem_data[22][0] ), .S(n8355), 
        .Z(n10142) );
  MUX2_X1 U9487 ( .A(\xmem_data[22][0] ), .B(\xmem_data[21][0] ), .S(n8353), 
        .Z(n10141) );
  MUX2_X1 U9488 ( .A(\xmem_data[21][0] ), .B(\xmem_data[20][0] ), .S(n8351), 
        .Z(n10140) );
  MUX2_X1 U9489 ( .A(\xmem_data[20][0] ), .B(\xmem_data[19][0] ), .S(n8355), 
        .Z(n10139) );
  MUX2_X1 U9490 ( .A(\xmem_data[19][0] ), .B(\xmem_data[18][0] ), .S(n8354), 
        .Z(n10138) );
  MUX2_X1 U9491 ( .A(\xmem_data[18][0] ), .B(\xmem_data[17][0] ), .S(n8353), 
        .Z(n10137) );
  MUX2_X1 U9492 ( .A(\xmem_data[17][0] ), .B(\xmem_data[16][0] ), .S(n8356), 
        .Z(n10136) );
  MUX2_X1 U9493 ( .A(\xmem_data[16][0] ), .B(\xmem_data[15][0] ), .S(n8351), 
        .Z(n10135) );
  BUF_X2 U9494 ( .A(n3835), .Z(n8353) );
  MUX2_X1 U9495 ( .A(\xmem_data[15][0] ), .B(\xmem_data[14][0] ), .S(n8353), 
        .Z(n10134) );
  MUX2_X1 U9496 ( .A(\xmem_data[14][0] ), .B(\xmem_data[13][0] ), .S(n8351), 
        .Z(n10133) );
  MUX2_X1 U9497 ( .A(\xmem_data[13][0] ), .B(\xmem_data[12][0] ), .S(n8352), 
        .Z(n10132) );
  MUX2_X1 U9498 ( .A(\xmem_data[12][0] ), .B(\xmem_data[11][0] ), .S(n8354), 
        .Z(n10131) );
  MUX2_X1 U9499 ( .A(\xmem_data[11][0] ), .B(\xmem_data[10][0] ), .S(n8353), 
        .Z(n10130) );
  MUX2_X1 U9500 ( .A(\xmem_data[10][0] ), .B(\xmem_data[9][0] ), .S(n8354), 
        .Z(n10129) );
  MUX2_X1 U9501 ( .A(\xmem_data[9][0] ), .B(\xmem_data[8][0] ), .S(n8356), .Z(
        n10128) );
  MUX2_X1 U9502 ( .A(\xmem_data[8][0] ), .B(\xmem_data[7][0] ), .S(n8354), .Z(
        n10127) );
  MUX2_X1 U9503 ( .A(\xmem_data[7][0] ), .B(\xmem_data[6][0] ), .S(n8353), .Z(
        n10126) );
  MUX2_X1 U9504 ( .A(\xmem_data[6][0] ), .B(\xmem_data[5][0] ), .S(n8352), .Z(
        n10125) );
  MUX2_X1 U9505 ( .A(\xmem_data[5][0] ), .B(\xmem_data[4][0] ), .S(n8351), .Z(
        n10124) );
  MUX2_X1 U9506 ( .A(\xmem_data[4][0] ), .B(\xmem_data[3][0] ), .S(n8352), .Z(
        n10123) );
  MUX2_X1 U9507 ( .A(\xmem_data[3][0] ), .B(\xmem_data[2][0] ), .S(n8355), .Z(
        n10122) );
  MUX2_X1 U9508 ( .A(\xmem_data[2][0] ), .B(\xmem_data[1][0] ), .S(n8352), .Z(
        n10121) );
  MUX2_X1 U9509 ( .A(\xmem_data[1][0] ), .B(\xmem_data[0][0] ), .S(n8353), .Z(
        n10120) );
  MUX2_X1 U9510 ( .A(s_data_in_x[1]), .B(\xmem_data[31][1] ), .S(n8352), .Z(
        n3371) );
  MUX2_X1 U9511 ( .A(\xmem_data[31][1] ), .B(\xmem_data[30][1] ), .S(n8354), 
        .Z(n10311) );
  MUX2_X1 U9512 ( .A(\xmem_data[30][1] ), .B(\xmem_data[29][1] ), .S(n8354), 
        .Z(n10303) );
  MUX2_X1 U9513 ( .A(\xmem_data[29][1] ), .B(\xmem_data[28][1] ), .S(n8356), 
        .Z(n10295) );
  MUX2_X1 U9514 ( .A(\xmem_data[28][1] ), .B(\xmem_data[27][1] ), .S(n8353), 
        .Z(n10287) );
  MUX2_X1 U9515 ( .A(\xmem_data[27][1] ), .B(\xmem_data[26][1] ), .S(n8356), 
        .Z(n10279) );
  MUX2_X1 U9516 ( .A(\xmem_data[26][1] ), .B(\xmem_data[25][1] ), .S(n8352), 
        .Z(n10171) );
  MUX2_X1 U9517 ( .A(\xmem_data[25][1] ), .B(\xmem_data[24][1] ), .S(n8355), 
        .Z(n10170) );
  BUF_X4 U9518 ( .A(n3835), .Z(n8356) );
  MUX2_X1 U9519 ( .A(\xmem_data[24][1] ), .B(\xmem_data[23][1] ), .S(n8356), 
        .Z(n10169) );
  MUX2_X1 U9520 ( .A(\xmem_data[23][1] ), .B(\xmem_data[22][1] ), .S(n8356), 
        .Z(n10168) );
  MUX2_X1 U9521 ( .A(\xmem_data[22][1] ), .B(\xmem_data[21][1] ), .S(n8351), 
        .Z(n10167) );
  MUX2_X1 U9522 ( .A(\xmem_data[21][1] ), .B(\xmem_data[20][1] ), .S(n8355), 
        .Z(n10166) );
  MUX2_X1 U9523 ( .A(\xmem_data[20][1] ), .B(\xmem_data[19][1] ), .S(n8353), 
        .Z(n10165) );
  MUX2_X1 U9524 ( .A(\xmem_data[19][1] ), .B(\xmem_data[18][1] ), .S(n8355), 
        .Z(n10164) );
  MUX2_X1 U9525 ( .A(\xmem_data[18][1] ), .B(\xmem_data[17][1] ), .S(n8355), 
        .Z(n10163) );
  MUX2_X1 U9526 ( .A(\xmem_data[17][1] ), .B(\xmem_data[16][1] ), .S(n8355), 
        .Z(n10162) );
  MUX2_X1 U9527 ( .A(\xmem_data[16][1] ), .B(\xmem_data[15][1] ), .S(n8352), 
        .Z(n10161) );
  MUX2_X1 U9528 ( .A(\xmem_data[15][1] ), .B(\xmem_data[14][1] ), .S(n8351), 
        .Z(n10160) );
  MUX2_X1 U9529 ( .A(\xmem_data[14][1] ), .B(\xmem_data[13][1] ), .S(n8352), 
        .Z(n10159) );
  MUX2_X1 U9530 ( .A(\xmem_data[13][1] ), .B(\xmem_data[12][1] ), .S(n8354), 
        .Z(n10158) );
  MUX2_X1 U9531 ( .A(\xmem_data[12][1] ), .B(\xmem_data[11][1] ), .S(n8355), 
        .Z(n10157) );
  MUX2_X1 U9532 ( .A(\xmem_data[11][1] ), .B(\xmem_data[10][1] ), .S(n8352), 
        .Z(n10156) );
  MUX2_X1 U9533 ( .A(\xmem_data[10][1] ), .B(\xmem_data[9][1] ), .S(n8355), 
        .Z(n10155) );
  MUX2_X1 U9534 ( .A(\xmem_data[9][1] ), .B(\xmem_data[8][1] ), .S(n8356), .Z(
        n10154) );
  MUX2_X1 U9535 ( .A(\xmem_data[8][1] ), .B(\xmem_data[7][1] ), .S(n8355), .Z(
        n10153) );
  MUX2_X1 U9536 ( .A(\xmem_data[7][1] ), .B(\xmem_data[6][1] ), .S(n8354), .Z(
        n10152) );
  MUX2_X1 U9537 ( .A(\xmem_data[6][1] ), .B(\xmem_data[5][1] ), .S(n8354), .Z(
        n10151) );
  MUX2_X1 U9538 ( .A(\xmem_data[5][1] ), .B(\xmem_data[4][1] ), .S(n8352), .Z(
        n10150) );
  MUX2_X1 U9539 ( .A(\xmem_data[4][1] ), .B(\xmem_data[3][1] ), .S(n8353), .Z(
        n10149) );
  MUX2_X1 U9540 ( .A(\xmem_data[3][1] ), .B(\xmem_data[2][1] ), .S(n8353), .Z(
        n10148) );
  MUX2_X1 U9541 ( .A(\xmem_data[2][1] ), .B(\xmem_data[1][1] ), .S(n8356), .Z(
        n10147) );
  MUX2_X1 U9542 ( .A(\xmem_data[1][1] ), .B(\xmem_data[0][1] ), .S(n8356), .Z(
        n10146) );
  MUX2_X1 U9543 ( .A(s_data_in_x[2]), .B(\xmem_data[31][2] ), .S(n8356), .Z(
        n3372) );
  MUX2_X1 U9544 ( .A(\xmem_data[31][2] ), .B(\xmem_data[30][2] ), .S(n8354), 
        .Z(n10312) );
  MUX2_X1 U9545 ( .A(\xmem_data[30][2] ), .B(\xmem_data[29][2] ), .S(n8352), 
        .Z(n10304) );
  MUX2_X1 U9546 ( .A(\xmem_data[29][2] ), .B(\xmem_data[28][2] ), .S(n8352), 
        .Z(n10296) );
  MUX2_X1 U9547 ( .A(\xmem_data[28][2] ), .B(\xmem_data[27][2] ), .S(n8356), 
        .Z(n10288) );
  MUX2_X1 U9548 ( .A(\xmem_data[27][2] ), .B(\xmem_data[26][2] ), .S(n8356), 
        .Z(n10280) );
  MUX2_X1 U9549 ( .A(\xmem_data[26][2] ), .B(\xmem_data[25][2] ), .S(n8356), 
        .Z(n10197) );
  MUX2_X1 U9550 ( .A(\xmem_data[25][2] ), .B(\xmem_data[24][2] ), .S(n8351), 
        .Z(n10196) );
  MUX2_X1 U9551 ( .A(\xmem_data[24][2] ), .B(\xmem_data[23][2] ), .S(n8356), 
        .Z(n10195) );
  MUX2_X1 U9552 ( .A(\xmem_data[23][2] ), .B(\xmem_data[22][2] ), .S(n8355), 
        .Z(n10194) );
  MUX2_X1 U9553 ( .A(\xmem_data[22][2] ), .B(\xmem_data[21][2] ), .S(n8355), 
        .Z(n10193) );
  MUX2_X1 U9554 ( .A(\xmem_data[21][2] ), .B(\xmem_data[20][2] ), .S(n8351), 
        .Z(n10192) );
  MUX2_X1 U9555 ( .A(\xmem_data[20][2] ), .B(\xmem_data[19][2] ), .S(n8355), 
        .Z(n10191) );
  MUX2_X1 U9556 ( .A(\xmem_data[19][2] ), .B(\xmem_data[18][2] ), .S(n8356), 
        .Z(n10190) );
  MUX2_X1 U9557 ( .A(\xmem_data[18][2] ), .B(\xmem_data[17][2] ), .S(n8353), 
        .Z(n10189) );
  MUX2_X1 U9558 ( .A(\xmem_data[17][2] ), .B(\xmem_data[16][2] ), .S(n8352), 
        .Z(n10188) );
  MUX2_X1 U9559 ( .A(\xmem_data[16][2] ), .B(\xmem_data[15][2] ), .S(n8352), 
        .Z(n10187) );
  MUX2_X1 U9560 ( .A(\xmem_data[15][2] ), .B(\xmem_data[14][2] ), .S(n8353), 
        .Z(n10186) );
  MUX2_X1 U9561 ( .A(\xmem_data[14][2] ), .B(\xmem_data[13][2] ), .S(n8356), 
        .Z(n10185) );
  MUX2_X1 U9562 ( .A(\xmem_data[13][2] ), .B(\xmem_data[12][2] ), .S(n8353), 
        .Z(n10184) );
  MUX2_X1 U9563 ( .A(\xmem_data[12][2] ), .B(\xmem_data[11][2] ), .S(n8352), 
        .Z(n10183) );
  MUX2_X1 U9564 ( .A(\xmem_data[11][2] ), .B(\xmem_data[10][2] ), .S(n8354), 
        .Z(n10182) );
  MUX2_X1 U9565 ( .A(\xmem_data[10][2] ), .B(\xmem_data[9][2] ), .S(n8356), 
        .Z(n10181) );
  MUX2_X1 U9566 ( .A(\xmem_data[9][2] ), .B(\xmem_data[8][2] ), .S(n8353), .Z(
        n10180) );
  MUX2_X1 U9567 ( .A(\xmem_data[8][2] ), .B(\xmem_data[7][2] ), .S(n8356), .Z(
        n10179) );
  MUX2_X1 U9568 ( .A(\xmem_data[7][2] ), .B(\xmem_data[6][2] ), .S(n8352), .Z(
        n10178) );
  MUX2_X1 U9569 ( .A(\xmem_data[6][2] ), .B(\xmem_data[5][2] ), .S(n8356), .Z(
        n10177) );
  MUX2_X1 U9570 ( .A(\xmem_data[5][2] ), .B(\xmem_data[4][2] ), .S(n8356), .Z(
        n10176) );
  MUX2_X1 U9571 ( .A(\xmem_data[4][2] ), .B(\xmem_data[3][2] ), .S(n8356), .Z(
        n10175) );
  MUX2_X1 U9572 ( .A(\xmem_data[3][2] ), .B(\xmem_data[2][2] ), .S(n8354), .Z(
        n10174) );
  MUX2_X1 U9573 ( .A(\xmem_data[2][2] ), .B(\xmem_data[1][2] ), .S(n8353), .Z(
        n10173) );
  MUX2_X1 U9574 ( .A(\xmem_data[1][2] ), .B(\xmem_data[0][2] ), .S(n8352), .Z(
        n10172) );
  MUX2_X1 U9575 ( .A(s_data_in_x[3]), .B(\xmem_data[31][3] ), .S(n8353), .Z(
        n3373) );
  MUX2_X1 U9576 ( .A(\xmem_data[31][3] ), .B(\xmem_data[30][3] ), .S(n8355), 
        .Z(n10313) );
  MUX2_X1 U9577 ( .A(\xmem_data[30][3] ), .B(\xmem_data[29][3] ), .S(n8351), 
        .Z(n10305) );
  MUX2_X1 U9578 ( .A(\xmem_data[29][3] ), .B(\xmem_data[28][3] ), .S(n8352), 
        .Z(n10297) );
  MUX2_X1 U9579 ( .A(\xmem_data[28][3] ), .B(\xmem_data[27][3] ), .S(n8351), 
        .Z(n10289) );
  MUX2_X1 U9580 ( .A(\xmem_data[27][3] ), .B(\xmem_data[26][3] ), .S(n8354), 
        .Z(n10281) );
  MUX2_X1 U9581 ( .A(\xmem_data[26][3] ), .B(\xmem_data[25][3] ), .S(n8355), 
        .Z(n10223) );
  MUX2_X1 U9582 ( .A(\xmem_data[25][3] ), .B(\xmem_data[24][3] ), .S(n8354), 
        .Z(n10222) );
  MUX2_X1 U9583 ( .A(\xmem_data[24][3] ), .B(\xmem_data[23][3] ), .S(n8355), 
        .Z(n10221) );
  MUX2_X1 U9584 ( .A(\xmem_data[23][3] ), .B(\xmem_data[22][3] ), .S(n8354), 
        .Z(n10220) );
  MUX2_X1 U9585 ( .A(\xmem_data[22][3] ), .B(\xmem_data[21][3] ), .S(n8356), 
        .Z(n10219) );
  MUX2_X1 U9586 ( .A(\xmem_data[21][3] ), .B(\xmem_data[20][3] ), .S(n8352), 
        .Z(n10218) );
  MUX2_X1 U9587 ( .A(\xmem_data[20][3] ), .B(\xmem_data[19][3] ), .S(n8355), 
        .Z(n10217) );
  MUX2_X1 U9588 ( .A(\xmem_data[19][3] ), .B(\xmem_data[18][3] ), .S(n8356), 
        .Z(n10216) );
  MUX2_X1 U9589 ( .A(\xmem_data[18][3] ), .B(\xmem_data[17][3] ), .S(n8351), 
        .Z(n10215) );
  MUX2_X1 U9590 ( .A(\xmem_data[17][3] ), .B(\xmem_data[16][3] ), .S(n8355), 
        .Z(n10214) );
  MUX2_X1 U9591 ( .A(\xmem_data[16][3] ), .B(\xmem_data[15][3] ), .S(n8354), 
        .Z(n10213) );
  MUX2_X1 U9592 ( .A(\xmem_data[15][3] ), .B(\xmem_data[14][3] ), .S(n8351), 
        .Z(n10212) );
  MUX2_X1 U9593 ( .A(\xmem_data[14][3] ), .B(\xmem_data[13][3] ), .S(n8351), 
        .Z(n10211) );
  MUX2_X1 U9594 ( .A(\xmem_data[13][3] ), .B(\xmem_data[12][3] ), .S(n8351), 
        .Z(n10210) );
  MUX2_X1 U9595 ( .A(\xmem_data[12][3] ), .B(\xmem_data[11][3] ), .S(n8352), 
        .Z(n10209) );
  MUX2_X1 U9596 ( .A(\xmem_data[11][3] ), .B(\xmem_data[10][3] ), .S(n8351), 
        .Z(n10208) );
  MUX2_X1 U9597 ( .A(\xmem_data[10][3] ), .B(\xmem_data[9][3] ), .S(n8352), 
        .Z(n10207) );
  MUX2_X1 U9598 ( .A(\xmem_data[9][3] ), .B(\xmem_data[8][3] ), .S(n8353), .Z(
        n10206) );
  MUX2_X1 U9599 ( .A(\xmem_data[8][3] ), .B(\xmem_data[7][3] ), .S(n8355), .Z(
        n10205) );
  MUX2_X1 U9600 ( .A(\xmem_data[7][3] ), .B(\xmem_data[6][3] ), .S(n8355), .Z(
        n10204) );
  MUX2_X1 U9601 ( .A(\xmem_data[6][3] ), .B(\xmem_data[5][3] ), .S(n8351), .Z(
        n10203) );
  MUX2_X1 U9602 ( .A(\xmem_data[5][3] ), .B(\xmem_data[4][3] ), .S(n8354), .Z(
        n10202) );
  MUX2_X1 U9603 ( .A(\xmem_data[4][3] ), .B(\xmem_data[3][3] ), .S(n8353), .Z(
        n10201) );
  MUX2_X1 U9604 ( .A(\xmem_data[3][3] ), .B(\xmem_data[2][3] ), .S(n8356), .Z(
        n10200) );
  MUX2_X1 U9605 ( .A(\xmem_data[2][3] ), .B(\xmem_data[1][3] ), .S(n8351), .Z(
        n10199) );
  MUX2_X1 U9606 ( .A(\xmem_data[1][3] ), .B(\xmem_data[0][3] ), .S(n8355), .Z(
        n10198) );
  MUX2_X1 U9607 ( .A(s_data_in_x[4]), .B(\xmem_data[31][4] ), .S(n8354), .Z(
        n3374) );
  MUX2_X1 U9608 ( .A(\xmem_data[31][4] ), .B(\xmem_data[30][4] ), .S(n8355), 
        .Z(n10314) );
  MUX2_X1 U9609 ( .A(\xmem_data[30][4] ), .B(\xmem_data[29][4] ), .S(n8356), 
        .Z(n10306) );
  MUX2_X1 U9610 ( .A(\xmem_data[29][4] ), .B(\xmem_data[28][4] ), .S(n8353), 
        .Z(n10298) );
  MUX2_X1 U9611 ( .A(\xmem_data[28][4] ), .B(\xmem_data[27][4] ), .S(n8354), 
        .Z(n10290) );
  MUX2_X1 U9612 ( .A(\xmem_data[27][4] ), .B(\xmem_data[26][4] ), .S(n8352), 
        .Z(n10282) );
  MUX2_X1 U9613 ( .A(\xmem_data[26][4] ), .B(\xmem_data[25][4] ), .S(n8351), 
        .Z(n10249) );
  MUX2_X1 U9614 ( .A(\xmem_data[25][4] ), .B(\xmem_data[24][4] ), .S(n3835), 
        .Z(n10248) );
  MUX2_X1 U9615 ( .A(\xmem_data[24][4] ), .B(\xmem_data[23][4] ), .S(n8352), 
        .Z(n10247) );
  MUX2_X1 U9616 ( .A(\xmem_data[23][4] ), .B(\xmem_data[22][4] ), .S(n8354), 
        .Z(n10246) );
  MUX2_X1 U9617 ( .A(\xmem_data[22][4] ), .B(\xmem_data[21][4] ), .S(n8353), 
        .Z(n10245) );
  MUX2_X1 U9618 ( .A(\xmem_data[21][4] ), .B(\xmem_data[20][4] ), .S(n8353), 
        .Z(n10244) );
  MUX2_X1 U9619 ( .A(\xmem_data[20][4] ), .B(\xmem_data[19][4] ), .S(n8356), 
        .Z(n10243) );
  MUX2_X1 U9620 ( .A(\xmem_data[19][4] ), .B(\xmem_data[18][4] ), .S(n8353), 
        .Z(n10242) );
  MUX2_X1 U9621 ( .A(\xmem_data[18][4] ), .B(\xmem_data[17][4] ), .S(n8356), 
        .Z(n10241) );
  MUX2_X1 U9622 ( .A(\xmem_data[17][4] ), .B(\xmem_data[16][4] ), .S(n8351), 
        .Z(n10240) );
  MUX2_X1 U9623 ( .A(\xmem_data[16][4] ), .B(\xmem_data[15][4] ), .S(n8353), 
        .Z(n10239) );
  MUX2_X1 U9624 ( .A(\xmem_data[15][4] ), .B(\xmem_data[14][4] ), .S(n8355), 
        .Z(n10238) );
  MUX2_X1 U9625 ( .A(\xmem_data[14][4] ), .B(\xmem_data[13][4] ), .S(n8353), 
        .Z(n10237) );
  MUX2_X1 U9626 ( .A(\xmem_data[13][4] ), .B(\xmem_data[12][4] ), .S(n8356), 
        .Z(n10236) );
  MUX2_X1 U9627 ( .A(\xmem_data[12][4] ), .B(\xmem_data[11][4] ), .S(n8356), 
        .Z(n10235) );
  MUX2_X1 U9628 ( .A(\xmem_data[11][4] ), .B(\xmem_data[10][4] ), .S(n8353), 
        .Z(n10234) );
  MUX2_X1 U9629 ( .A(\xmem_data[10][4] ), .B(\xmem_data[9][4] ), .S(n3835), 
        .Z(n10233) );
  MUX2_X1 U9630 ( .A(\xmem_data[9][4] ), .B(\xmem_data[8][4] ), .S(n8355), .Z(
        n10232) );
  MUX2_X1 U9631 ( .A(\xmem_data[8][4] ), .B(\xmem_data[7][4] ), .S(n8353), .Z(
        n10231) );
  MUX2_X1 U9632 ( .A(\xmem_data[7][4] ), .B(\xmem_data[6][4] ), .S(n8353), .Z(
        n10230) );
  MUX2_X1 U9633 ( .A(\xmem_data[6][4] ), .B(\xmem_data[5][4] ), .S(n8353), .Z(
        n10229) );
  MUX2_X1 U9634 ( .A(\xmem_data[5][4] ), .B(\xmem_data[4][4] ), .S(n8354), .Z(
        n10228) );
  MUX2_X1 U9635 ( .A(\xmem_data[4][4] ), .B(\xmem_data[3][4] ), .S(n8354), .Z(
        n10227) );
  MUX2_X1 U9636 ( .A(\xmem_data[3][4] ), .B(\xmem_data[2][4] ), .S(n3835), .Z(
        n10226) );
  MUX2_X1 U9637 ( .A(\xmem_data[2][4] ), .B(\xmem_data[1][4] ), .S(n8353), .Z(
        n10225) );
  MUX2_X1 U9638 ( .A(\xmem_data[1][4] ), .B(\xmem_data[0][4] ), .S(n8353), .Z(
        n10224) );
  MUX2_X1 U9639 ( .A(s_data_in_x[5]), .B(\xmem_data[31][5] ), .S(n8352), .Z(
        n3375) );
  MUX2_X1 U9640 ( .A(\xmem_data[31][5] ), .B(\xmem_data[30][5] ), .S(n8351), 
        .Z(n10315) );
  MUX2_X1 U9641 ( .A(\xmem_data[30][5] ), .B(\xmem_data[29][5] ), .S(n8352), 
        .Z(n10307) );
  MUX2_X1 U9642 ( .A(\xmem_data[29][5] ), .B(\xmem_data[28][5] ), .S(n8356), 
        .Z(n10299) );
  MUX2_X1 U9643 ( .A(\xmem_data[28][5] ), .B(\xmem_data[27][5] ), .S(n8354), 
        .Z(n10291) );
  MUX2_X1 U9644 ( .A(\xmem_data[27][5] ), .B(\xmem_data[26][5] ), .S(n8355), 
        .Z(n10283) );
  MUX2_X1 U9645 ( .A(\xmem_data[26][5] ), .B(\xmem_data[25][5] ), .S(n8354), 
        .Z(n10275) );
  MUX2_X1 U9646 ( .A(\xmem_data[25][5] ), .B(\xmem_data[24][5] ), .S(n8355), 
        .Z(n10274) );
  MUX2_X1 U9647 ( .A(\xmem_data[24][5] ), .B(\xmem_data[23][5] ), .S(n8354), 
        .Z(n10273) );
  MUX2_X1 U9648 ( .A(\xmem_data[23][5] ), .B(\xmem_data[22][5] ), .S(n8354), 
        .Z(n10272) );
  MUX2_X1 U9649 ( .A(\xmem_data[22][5] ), .B(\xmem_data[21][5] ), .S(n8351), 
        .Z(n10271) );
  MUX2_X1 U9650 ( .A(\xmem_data[21][5] ), .B(\xmem_data[20][5] ), .S(n8352), 
        .Z(n10270) );
  MUX2_X1 U9651 ( .A(\xmem_data[20][5] ), .B(\xmem_data[19][5] ), .S(n8351), 
        .Z(n10269) );
  MUX2_X1 U9652 ( .A(\xmem_data[19][5] ), .B(\xmem_data[18][5] ), .S(n3835), 
        .Z(n10268) );
  MUX2_X1 U9653 ( .A(\xmem_data[18][5] ), .B(\xmem_data[17][5] ), .S(n8356), 
        .Z(n10267) );
  MUX2_X1 U9654 ( .A(\xmem_data[17][5] ), .B(\xmem_data[16][5] ), .S(n8356), 
        .Z(n10266) );
  MUX2_X1 U9655 ( .A(\xmem_data[16][5] ), .B(\xmem_data[15][5] ), .S(n8352), 
        .Z(n10265) );
  MUX2_X1 U9656 ( .A(\xmem_data[15][5] ), .B(\xmem_data[14][5] ), .S(n8355), 
        .Z(n10264) );
  MUX2_X1 U9657 ( .A(\xmem_data[14][5] ), .B(\xmem_data[13][5] ), .S(n8356), 
        .Z(n10263) );
  MUX2_X1 U9658 ( .A(\xmem_data[13][5] ), .B(\xmem_data[12][5] ), .S(n8354), 
        .Z(n10262) );
  MUX2_X1 U9659 ( .A(\xmem_data[12][5] ), .B(\xmem_data[11][5] ), .S(n3835), 
        .Z(n10261) );
  MUX2_X1 U9660 ( .A(\xmem_data[11][5] ), .B(\xmem_data[10][5] ), .S(n8352), 
        .Z(n10260) );
  MUX2_X1 U9661 ( .A(\xmem_data[10][5] ), .B(\xmem_data[9][5] ), .S(n8355), 
        .Z(n10259) );
  MUX2_X1 U9662 ( .A(\xmem_data[9][5] ), .B(\xmem_data[8][5] ), .S(n3835), .Z(
        n10258) );
  MUX2_X1 U9663 ( .A(\xmem_data[8][5] ), .B(\xmem_data[7][5] ), .S(n8353), .Z(
        n10257) );
  MUX2_X1 U9664 ( .A(\xmem_data[7][5] ), .B(\xmem_data[6][5] ), .S(n8351), .Z(
        n10256) );
  MUX2_X1 U9665 ( .A(\xmem_data[6][5] ), .B(\xmem_data[5][5] ), .S(n8352), .Z(
        n10255) );
  MUX2_X1 U9666 ( .A(\xmem_data[5][5] ), .B(\xmem_data[4][5] ), .S(n8354), .Z(
        n10254) );
  MUX2_X1 U9667 ( .A(\xmem_data[4][5] ), .B(\xmem_data[3][5] ), .S(n8355), .Z(
        n10253) );
  MUX2_X1 U9668 ( .A(\xmem_data[3][5] ), .B(\xmem_data[2][5] ), .S(n8355), .Z(
        n10252) );
  MUX2_X1 U9669 ( .A(\xmem_data[2][5] ), .B(\xmem_data[1][5] ), .S(n3835), .Z(
        n10251) );
  MUX2_X1 U9670 ( .A(\xmem_data[1][5] ), .B(\xmem_data[0][5] ), .S(n8356), .Z(
        n10250) );
  MUX2_X1 U9671 ( .A(s_data_in_x[6]), .B(\xmem_data[31][6] ), .S(n8355), .Z(
        n3376) );
  MUX2_X1 U9672 ( .A(\xmem_data[31][6] ), .B(\xmem_data[30][6] ), .S(n8353), 
        .Z(n10316) );
  MUX2_X1 U9673 ( .A(\xmem_data[30][6] ), .B(\xmem_data[29][6] ), .S(n8353), 
        .Z(n10308) );
  MUX2_X1 U9674 ( .A(\xmem_data[29][6] ), .B(\xmem_data[28][6] ), .S(n8353), 
        .Z(n10300) );
  MUX2_X1 U9675 ( .A(\xmem_data[28][6] ), .B(\xmem_data[27][6] ), .S(n8354), 
        .Z(n10292) );
  MUX2_X1 U9676 ( .A(\xmem_data[27][6] ), .B(\xmem_data[26][6] ), .S(n3835), 
        .Z(n10284) );
  MUX2_X1 U9677 ( .A(\xmem_data[26][6] ), .B(\xmem_data[25][6] ), .S(n8356), 
        .Z(n10276) );
  MUX2_X1 U9678 ( .A(\xmem_data[25][6] ), .B(\xmem_data[24][6] ), .S(n8356), 
        .Z(n10094) );
  MUX2_X1 U9679 ( .A(\xmem_data[24][6] ), .B(\xmem_data[23][6] ), .S(n8351), 
        .Z(n10093) );
  MUX2_X1 U9680 ( .A(\xmem_data[23][6] ), .B(\xmem_data[22][6] ), .S(n8351), 
        .Z(n10092) );
  MUX2_X1 U9681 ( .A(\xmem_data[22][6] ), .B(\xmem_data[21][6] ), .S(n8351), 
        .Z(n10091) );
  MUX2_X1 U9682 ( .A(\xmem_data[21][6] ), .B(\xmem_data[20][6] ), .S(n8354), 
        .Z(n10090) );
  MUX2_X1 U9683 ( .A(\xmem_data[20][6] ), .B(\xmem_data[19][6] ), .S(n8355), 
        .Z(n10089) );
  MUX2_X1 U9684 ( .A(\xmem_data[19][6] ), .B(\xmem_data[18][6] ), .S(n8351), 
        .Z(n10088) );
  MUX2_X1 U9685 ( .A(\xmem_data[18][6] ), .B(\xmem_data[17][6] ), .S(n8356), 
        .Z(n10087) );
  MUX2_X1 U9686 ( .A(\xmem_data[17][6] ), .B(\xmem_data[16][6] ), .S(n8353), 
        .Z(n10086) );
  MUX2_X1 U9687 ( .A(\xmem_data[16][6] ), .B(\xmem_data[15][6] ), .S(n8356), 
        .Z(n10085) );
  MUX2_X1 U9688 ( .A(\xmem_data[15][6] ), .B(\xmem_data[14][6] ), .S(n8352), 
        .Z(n10084) );
  MUX2_X1 U9689 ( .A(\xmem_data[14][6] ), .B(\xmem_data[13][6] ), .S(n8351), 
        .Z(n10083) );
  MUX2_X1 U9690 ( .A(\xmem_data[13][6] ), .B(\xmem_data[12][6] ), .S(n8351), 
        .Z(n10082) );
  MUX2_X1 U9691 ( .A(\xmem_data[12][6] ), .B(\xmem_data[11][6] ), .S(n8352), 
        .Z(n10081) );
  MUX2_X1 U9692 ( .A(\xmem_data[11][6] ), .B(\xmem_data[10][6] ), .S(n8356), 
        .Z(n10080) );
  MUX2_X1 U9693 ( .A(\xmem_data[10][6] ), .B(\xmem_data[9][6] ), .S(n8353), 
        .Z(n10079) );
  MUX2_X1 U9694 ( .A(\xmem_data[9][6] ), .B(\xmem_data[8][6] ), .S(n8352), .Z(
        n10078) );
  MUX2_X1 U9695 ( .A(\xmem_data[8][6] ), .B(\xmem_data[7][6] ), .S(n8351), .Z(
        n10077) );
  MUX2_X1 U9696 ( .A(\xmem_data[7][6] ), .B(\xmem_data[6][6] ), .S(n8352), .Z(
        n10076) );
  MUX2_X1 U9697 ( .A(\xmem_data[6][6] ), .B(\xmem_data[5][6] ), .S(n8351), .Z(
        n10075) );
  MUX2_X1 U9698 ( .A(\xmem_data[5][6] ), .B(\xmem_data[4][6] ), .S(n8356), .Z(
        n10074) );
  MUX2_X1 U9699 ( .A(\xmem_data[4][6] ), .B(\xmem_data[3][6] ), .S(n8354), .Z(
        n10073) );
  MUX2_X1 U9700 ( .A(\xmem_data[3][6] ), .B(\xmem_data[2][6] ), .S(n8353), .Z(
        n10072) );
  MUX2_X1 U9701 ( .A(\xmem_data[2][6] ), .B(\xmem_data[1][6] ), .S(n8356), .Z(
        n10071) );
  MUX2_X1 U9702 ( .A(\xmem_data[1][6] ), .B(\xmem_data[0][6] ), .S(n3835), .Z(
        n10070) );
  MUX2_X1 U9703 ( .A(s_data_in_x[7]), .B(\xmem_data[31][7] ), .S(n8354), .Z(
        n3377) );
  MUX2_X1 U9704 ( .A(\xmem_data[31][7] ), .B(\xmem_data[30][7] ), .S(n8356), 
        .Z(n10317) );
  MUX2_X1 U9705 ( .A(\xmem_data[30][7] ), .B(\xmem_data[29][7] ), .S(n3835), 
        .Z(n10309) );
  MUX2_X1 U9706 ( .A(\xmem_data[29][7] ), .B(\xmem_data[28][7] ), .S(n8351), 
        .Z(n10301) );
  MUX2_X1 U9707 ( .A(\xmem_data[28][7] ), .B(\xmem_data[27][7] ), .S(n8355), 
        .Z(n10293) );
  MUX2_X1 U9708 ( .A(\xmem_data[27][7] ), .B(\xmem_data[26][7] ), .S(n8356), 
        .Z(n10285) );
  MUX2_X1 U9709 ( .A(\xmem_data[26][7] ), .B(\xmem_data[25][7] ), .S(n3835), 
        .Z(n10277) );
  MUX2_X1 U9710 ( .A(\xmem_data[25][7] ), .B(\xmem_data[24][7] ), .S(n8352), 
        .Z(n10119) );
  MUX2_X1 U9711 ( .A(\xmem_data[24][7] ), .B(\xmem_data[23][7] ), .S(n8351), 
        .Z(n10118) );
  MUX2_X1 U9712 ( .A(\xmem_data[23][7] ), .B(\xmem_data[22][7] ), .S(n8354), 
        .Z(n10117) );
  MUX2_X1 U9713 ( .A(\xmem_data[22][7] ), .B(\xmem_data[21][7] ), .S(n8355), 
        .Z(n10116) );
  MUX2_X1 U9714 ( .A(\xmem_data[21][7] ), .B(\xmem_data[20][7] ), .S(n8354), 
        .Z(n10115) );
  MUX2_X1 U9715 ( .A(\xmem_data[20][7] ), .B(\xmem_data[19][7] ), .S(n8355), 
        .Z(n10114) );
  MUX2_X1 U9716 ( .A(\xmem_data[19][7] ), .B(\xmem_data[18][7] ), .S(n8355), 
        .Z(n10113) );
  MUX2_X1 U9717 ( .A(\xmem_data[18][7] ), .B(\xmem_data[17][7] ), .S(n8356), 
        .Z(n10112) );
  MUX2_X1 U9718 ( .A(\xmem_data[17][7] ), .B(\xmem_data[16][7] ), .S(n8354), 
        .Z(n10111) );
  MUX2_X1 U9719 ( .A(\xmem_data[16][7] ), .B(\xmem_data[15][7] ), .S(n8356), 
        .Z(n10110) );
  MUX2_X1 U9720 ( .A(\xmem_data[15][7] ), .B(\xmem_data[14][7] ), .S(n8356), 
        .Z(n10109) );
  MUX2_X1 U9721 ( .A(\xmem_data[14][7] ), .B(\xmem_data[13][7] ), .S(n8356), 
        .Z(n10108) );
  MUX2_X1 U9722 ( .A(\xmem_data[13][7] ), .B(\xmem_data[12][7] ), .S(n8352), 
        .Z(n10107) );
  MUX2_X1 U9723 ( .A(\xmem_data[12][7] ), .B(\xmem_data[11][7] ), .S(n8354), 
        .Z(n10106) );
  MUX2_X1 U9724 ( .A(\xmem_data[11][7] ), .B(\xmem_data[10][7] ), .S(n8351), 
        .Z(n10105) );
  MUX2_X1 U9725 ( .A(\xmem_data[10][7] ), .B(\xmem_data[9][7] ), .S(n3835), 
        .Z(n10104) );
  MUX2_X1 U9726 ( .A(\xmem_data[9][7] ), .B(\xmem_data[8][7] ), .S(n8353), .Z(
        n10103) );
  MUX2_X1 U9727 ( .A(\xmem_data[8][7] ), .B(\xmem_data[7][7] ), .S(n8351), .Z(
        n10102) );
  MUX2_X1 U9728 ( .A(\xmem_data[7][7] ), .B(\xmem_data[6][7] ), .S(n3835), .Z(
        n10101) );
  MUX2_X1 U9729 ( .A(\xmem_data[6][7] ), .B(\xmem_data[5][7] ), .S(n8351), .Z(
        n10100) );
  MUX2_X1 U9730 ( .A(\xmem_data[5][7] ), .B(\xmem_data[4][7] ), .S(n3835), .Z(
        n10099) );
  MUX2_X1 U9731 ( .A(\xmem_data[4][7] ), .B(\xmem_data[3][7] ), .S(n8352), .Z(
        n10098) );
  MUX2_X1 U9732 ( .A(\xmem_data[3][7] ), .B(\xmem_data[2][7] ), .S(n8354), .Z(
        n10097) );
  MUX2_X1 U9733 ( .A(\xmem_data[2][7] ), .B(\xmem_data[1][7] ), .S(n8356), .Z(
        n10096) );
  MUX2_X1 U9734 ( .A(\xmem_data[1][7] ), .B(\xmem_data[0][7] ), .S(n8351), .Z(
        n10095) );
  NOR2_X1 U9735 ( .A1(n8357), .A2(reset), .ZN(n8362) );
  NAND3_X1 U9736 ( .A1(n8360), .A2(n8359), .A3(n8358), .ZN(n8361) );
  MUX2_X1 U9737 ( .A(xmem_full), .B(n8362), .S(n8361), .Z(n3391) );
  AOI22_X1 U9738 ( .A1(\x_mult_f_int[0][8] ), .A2(n8401), .B1(n8400), .B2(
        \x_mult_f[0][8] ), .ZN(n8784) );
  AOI22_X1 U9739 ( .A1(n8391), .A2(\x_mult_f[0][3] ), .B1(n8363), .B2(
        \x_mult_f_int[0][3] ), .ZN(n8786) );
  AOI22_X1 U9740 ( .A1(n8391), .A2(\x_mult_f[0][2] ), .B1(n8363), .B2(
        \x_mult_f_int[0][2] ), .ZN(n8787) );
  AOI22_X1 U9741 ( .A1(n8208), .A2(\x_mult_f_int[1][5] ), .B1(n8400), .B2(
        \x_mult_f[1][5] ), .ZN(n8789) );
  AOI22_X1 U9742 ( .A1(\x_mult_f_int[3][7] ), .A2(n8365), .B1(n8364), .B2(
        \x_mult_f[3][7] ), .ZN(n8791) );
  AOI21_X1 U9743 ( .B1(n8374), .B2(n8367), .A(n8366), .ZN(n8371) );
  NAND2_X1 U9744 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  XOR2_X1 U9745 ( .A(n8371), .B(n8370), .Z(n8372) );
  AOI22_X1 U9746 ( .A1(n8372), .A2(n8213), .B1(n8381), .B2(
        \adder_stage3[0][19] ), .ZN(n8793) );
  NAND2_X1 U9747 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  NAND2_X1 U9748 ( .A1(n8376), .A2(n8375), .ZN(n8380) );
  NAND2_X1 U9749 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  XNOR2_X1 U9750 ( .A(n8380), .B(n8379), .ZN(n8382) );
  AOI22_X1 U9751 ( .A1(n8382), .A2(n8114), .B1(n8381), .B2(
        \adder_stage3[0][18] ), .ZN(n8794) );
  AOI22_X1 U9752 ( .A1(\x_mult_f_int[9][6] ), .A2(n8365), .B1(n8383), .B2(
        \x_mult_f[9][6] ), .ZN(n8799) );
  FA_X1 U9753 ( .A(n3481), .B(n8699), .CI(n8384), .CO(n8385), .S(n7948) );
  INV_X1 U9754 ( .A(n8385), .ZN(n8388) );
  AOI22_X1 U9755 ( .A1(n8388), .A2(n8387), .B1(n8386), .B2(
        \adder_stage1[4][20] ), .ZN(n8800) );
  AOI22_X1 U9756 ( .A1(n8391), .A2(\x_mult_f[10][4] ), .B1(n8389), .B2(
        \x_mult_f_int[10][4] ), .ZN(n8803) );
  AOI22_X1 U9757 ( .A1(n8391), .A2(\x_mult_f[10][2] ), .B1(n8389), .B2(
        \x_mult_f_int[10][2] ), .ZN(n8804) );
  AOI22_X1 U9758 ( .A1(n8391), .A2(\x_mult_f[12][4] ), .B1(n8390), .B2(
        \x_mult_f_int[12][4] ), .ZN(n8805) );
  AOI22_X1 U9759 ( .A1(\x_mult_f_int[21][10] ), .A2(n8401), .B1(n8392), .B2(
        \x_mult_f[21][10] ), .ZN(n8811) );
  AOI22_X1 U9760 ( .A1(\x_mult_f_int[21][9] ), .A2(n8401), .B1(n8392), .B2(
        \x_mult_f[21][9] ), .ZN(n8812) );
  AOI22_X1 U9761 ( .A1(\x_mult_f_int[21][8] ), .A2(n8401), .B1(n8392), .B2(
        \x_mult_f[21][8] ), .ZN(n8813) );
  AOI22_X1 U9762 ( .A1(\x_mult_f_int[21][7] ), .A2(n8401), .B1(n8392), .B2(
        \x_mult_f[21][7] ), .ZN(n8814) );
  AOI22_X1 U9763 ( .A1(\x_mult_f_int[21][6] ), .A2(n8401), .B1(n8395), .B2(
        \x_mult_f[21][6] ), .ZN(n8815) );
  AOI22_X1 U9764 ( .A1(n8186), .A2(\x_mult_f_int[21][5] ), .B1(n8395), .B2(
        \x_mult_f[21][5] ), .ZN(n8816) );
  FA_X1 U9765 ( .A(n8700), .B(n3498), .CI(n8393), .CO(n8394), .S(n3586) );
  INV_X1 U9766 ( .A(n8394), .ZN(n8396) );
  AOI22_X1 U9767 ( .A1(n8396), .A2(n8401), .B1(n8395), .B2(
        \adder_stage1[10][20] ), .ZN(n8817) );
  AOI22_X1 U9768 ( .A1(\x_mult_f_int[25][7] ), .A2(n8398), .B1(n8397), .B2(
        \x_mult_f[25][7] ), .ZN(n8827) );
  AOI22_X1 U9769 ( .A1(n8037), .A2(\x_mult_f_int[25][5] ), .B1(n5294), .B2(
        \x_mult_f[25][5] ), .ZN(n8829) );
  AOI22_X1 U9770 ( .A1(\x_mult_f_int[26][11] ), .A2(n8399), .B1(n8400), .B2(
        \x_mult_f[26][11] ), .ZN(n8830) );
  AOI22_X1 U9771 ( .A1(\x_mult_f_int[26][10] ), .A2(n8399), .B1(n8157), .B2(
        \x_mult_f[26][10] ), .ZN(n8831) );
  AOI22_X1 U9772 ( .A1(\x_mult_f_int[26][9] ), .A2(n8399), .B1(n6330), .B2(
        \x_mult_f[26][9] ), .ZN(n8832) );
  AOI22_X1 U9773 ( .A1(\x_mult_f_int[26][6] ), .A2(n4002), .B1(n8400), .B2(
        \x_mult_f[26][6] ), .ZN(n8834) );
  AOI22_X1 U9774 ( .A1(\x_mult_f_int[29][13] ), .A2(n8401), .B1(n7512), .B2(
        \x_mult_f[29][13] ), .ZN(n8845) );
  NAND3_X1 U9775 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .A3(fmem_addr[2]), 
        .ZN(n8676) );
  NAND2_X1 U9776 ( .A1(n8681), .A2(fmem_addr[4]), .ZN(n8481) );
  OAI22_X1 U9777 ( .A1(n8675), .A2(s_data_in_f[7]), .B1(\fmem_data[31][7] ), 
        .B2(n8689), .ZN(n8402) );
  INV_X1 U9778 ( .A(n8402), .ZN(n9356) );
  OAI22_X1 U9779 ( .A1(n8675), .A2(s_data_in_f[6]), .B1(\fmem_data[31][6] ), 
        .B2(n8689), .ZN(n8403) );
  INV_X1 U9780 ( .A(n8403), .ZN(n9357) );
  OAI22_X1 U9781 ( .A1(n8675), .A2(s_data_in_f[5]), .B1(\fmem_data[31][5] ), 
        .B2(n8689), .ZN(n8404) );
  INV_X1 U9782 ( .A(n8404), .ZN(n9358) );
  OAI22_X1 U9783 ( .A1(n8675), .A2(s_data_in_f[4]), .B1(\fmem_data[31][4] ), 
        .B2(n8689), .ZN(n8405) );
  INV_X1 U9784 ( .A(n8405), .ZN(n9359) );
  OAI22_X1 U9785 ( .A1(n8675), .A2(s_data_in_f[3]), .B1(\fmem_data[31][3] ), 
        .B2(n8689), .ZN(n8406) );
  INV_X1 U9786 ( .A(n8406), .ZN(n9360) );
  OAI22_X1 U9787 ( .A1(n8675), .A2(s_data_in_f[2]), .B1(\fmem_data[31][2] ), 
        .B2(n8689), .ZN(n8407) );
  INV_X1 U9788 ( .A(n8407), .ZN(n9361) );
  OAI22_X1 U9789 ( .A1(n8675), .A2(s_data_in_f[1]), .B1(\fmem_data[31][1] ), 
        .B2(n8689), .ZN(n8408) );
  INV_X1 U9790 ( .A(n8408), .ZN(n9362) );
  OAI22_X1 U9791 ( .A1(n8675), .A2(s_data_in_f[0]), .B1(\fmem_data[31][0] ), 
        .B2(n8689), .ZN(n8409) );
  INV_X1 U9792 ( .A(n8409), .ZN(n9363) );
  NAND3_X1 U9793 ( .A1(fmem_addr[1]), .A2(fmem_addr[2]), .A3(n8710), .ZN(n8590) );
  OAI22_X1 U9794 ( .A1(n8418), .A2(s_data_in_f[7]), .B1(\fmem_data[30][7] ), 
        .B2(n8417), .ZN(n8410) );
  INV_X1 U9795 ( .A(n8410), .ZN(n9364) );
  OAI22_X1 U9796 ( .A1(n8418), .A2(s_data_in_f[6]), .B1(\fmem_data[30][6] ), 
        .B2(n8417), .ZN(n8411) );
  INV_X1 U9797 ( .A(n8411), .ZN(n9365) );
  OAI22_X1 U9798 ( .A1(n8418), .A2(s_data_in_f[5]), .B1(\fmem_data[30][5] ), 
        .B2(n8417), .ZN(n8412) );
  INV_X1 U9799 ( .A(n8412), .ZN(n9366) );
  OAI22_X1 U9800 ( .A1(n8418), .A2(s_data_in_f[4]), .B1(\fmem_data[30][4] ), 
        .B2(n8417), .ZN(n8413) );
  INV_X1 U9801 ( .A(n8413), .ZN(n9367) );
  OAI22_X1 U9802 ( .A1(n8418), .A2(s_data_in_f[3]), .B1(\fmem_data[30][3] ), 
        .B2(n8417), .ZN(n8414) );
  INV_X1 U9803 ( .A(n8414), .ZN(n9368) );
  OAI22_X1 U9804 ( .A1(n8418), .A2(s_data_in_f[2]), .B1(\fmem_data[30][2] ), 
        .B2(n8417), .ZN(n8415) );
  INV_X1 U9805 ( .A(n8415), .ZN(n9369) );
  OAI22_X1 U9806 ( .A1(n8418), .A2(s_data_in_f[1]), .B1(\fmem_data[30][1] ), 
        .B2(n8417), .ZN(n8416) );
  INV_X1 U9807 ( .A(n8416), .ZN(n9370) );
  OAI22_X1 U9808 ( .A1(n8418), .A2(s_data_in_f[0]), .B1(\fmem_data[30][0] ), 
        .B2(n8417), .ZN(n8419) );
  INV_X1 U9809 ( .A(n8419), .ZN(n9371) );
  NAND3_X1 U9810 ( .A1(fmem_addr[0]), .A2(fmem_addr[2]), .A3(n8711), .ZN(n8601) );
  OAI22_X1 U9811 ( .A1(n8428), .A2(s_data_in_f[7]), .B1(\fmem_data[29][7] ), 
        .B2(n8427), .ZN(n8420) );
  INV_X1 U9812 ( .A(n8420), .ZN(n9372) );
  OAI22_X1 U9813 ( .A1(n8428), .A2(s_data_in_f[6]), .B1(\fmem_data[29][6] ), 
        .B2(n8427), .ZN(n8421) );
  INV_X1 U9814 ( .A(n8421), .ZN(n9373) );
  OAI22_X1 U9815 ( .A1(n8428), .A2(s_data_in_f[5]), .B1(\fmem_data[29][5] ), 
        .B2(n8427), .ZN(n8422) );
  INV_X1 U9816 ( .A(n8422), .ZN(n9374) );
  OAI22_X1 U9817 ( .A1(n8428), .A2(s_data_in_f[4]), .B1(\fmem_data[29][4] ), 
        .B2(n8427), .ZN(n8423) );
  INV_X1 U9818 ( .A(n8423), .ZN(n9375) );
  OAI22_X1 U9819 ( .A1(n8428), .A2(s_data_in_f[3]), .B1(\fmem_data[29][3] ), 
        .B2(n8427), .ZN(n8424) );
  INV_X1 U9820 ( .A(n8424), .ZN(n9376) );
  OAI22_X1 U9821 ( .A1(n8428), .A2(s_data_in_f[2]), .B1(\fmem_data[29][2] ), 
        .B2(n8427), .ZN(n8425) );
  INV_X1 U9822 ( .A(n8425), .ZN(n9377) );
  OAI22_X1 U9823 ( .A1(n8428), .A2(s_data_in_f[1]), .B1(\fmem_data[29][1] ), 
        .B2(n8427), .ZN(n8426) );
  INV_X1 U9824 ( .A(n8426), .ZN(n9378) );
  OAI22_X1 U9825 ( .A1(n8428), .A2(s_data_in_f[0]), .B1(\fmem_data[29][0] ), 
        .B2(n8427), .ZN(n8429) );
  INV_X1 U9826 ( .A(n8429), .ZN(n9379) );
  NAND3_X1 U9827 ( .A1(fmem_addr[2]), .A2(n8710), .A3(n8711), .ZN(n8612) );
  OAI22_X1 U9828 ( .A1(n8438), .A2(s_data_in_f[7]), .B1(\fmem_data[28][7] ), 
        .B2(n8437), .ZN(n8430) );
  INV_X1 U9829 ( .A(n8430), .ZN(n9380) );
  OAI22_X1 U9830 ( .A1(n8438), .A2(s_data_in_f[6]), .B1(\fmem_data[28][6] ), 
        .B2(n8437), .ZN(n8431) );
  INV_X1 U9831 ( .A(n8431), .ZN(n9381) );
  OAI22_X1 U9832 ( .A1(n8438), .A2(s_data_in_f[5]), .B1(\fmem_data[28][5] ), 
        .B2(n8437), .ZN(n8432) );
  INV_X1 U9833 ( .A(n8432), .ZN(n9382) );
  OAI22_X1 U9834 ( .A1(n8438), .A2(s_data_in_f[4]), .B1(\fmem_data[28][4] ), 
        .B2(n8437), .ZN(n8433) );
  INV_X1 U9835 ( .A(n8433), .ZN(n9383) );
  OAI22_X1 U9836 ( .A1(n8438), .A2(s_data_in_f[3]), .B1(\fmem_data[28][3] ), 
        .B2(n8437), .ZN(n8434) );
  INV_X1 U9837 ( .A(n8434), .ZN(n9384) );
  OAI22_X1 U9838 ( .A1(n8438), .A2(s_data_in_f[2]), .B1(\fmem_data[28][2] ), 
        .B2(n8437), .ZN(n8435) );
  INV_X1 U9839 ( .A(n8435), .ZN(n9385) );
  OAI22_X1 U9840 ( .A1(n8438), .A2(s_data_in_f[1]), .B1(\fmem_data[28][1] ), 
        .B2(n8437), .ZN(n8436) );
  INV_X1 U9841 ( .A(n8436), .ZN(n9386) );
  OAI22_X1 U9842 ( .A1(n8438), .A2(s_data_in_f[0]), .B1(\fmem_data[28][0] ), 
        .B2(n8437), .ZN(n8439) );
  INV_X1 U9843 ( .A(n8439), .ZN(n9387) );
  NAND3_X1 U9844 ( .A1(fmem_addr[1]), .A2(fmem_addr[0]), .A3(n8709), .ZN(n8685) );
  OAI22_X1 U9845 ( .A1(n8448), .A2(s_data_in_f[7]), .B1(\fmem_data[27][7] ), 
        .B2(n8447), .ZN(n8440) );
  INV_X1 U9846 ( .A(n8440), .ZN(n9388) );
  OAI22_X1 U9847 ( .A1(n8448), .A2(s_data_in_f[6]), .B1(\fmem_data[27][6] ), 
        .B2(n8447), .ZN(n8441) );
  INV_X1 U9848 ( .A(n8441), .ZN(n9389) );
  OAI22_X1 U9849 ( .A1(n8448), .A2(s_data_in_f[5]), .B1(\fmem_data[27][5] ), 
        .B2(n8447), .ZN(n8442) );
  INV_X1 U9850 ( .A(n8442), .ZN(n9390) );
  OAI22_X1 U9851 ( .A1(n8448), .A2(s_data_in_f[4]), .B1(\fmem_data[27][4] ), 
        .B2(n8447), .ZN(n8443) );
  INV_X1 U9852 ( .A(n8443), .ZN(n9391) );
  OAI22_X1 U9853 ( .A1(n8448), .A2(s_data_in_f[3]), .B1(\fmem_data[27][3] ), 
        .B2(n8447), .ZN(n8444) );
  INV_X1 U9854 ( .A(n8444), .ZN(n9392) );
  OAI22_X1 U9855 ( .A1(n8448), .A2(s_data_in_f[2]), .B1(\fmem_data[27][2] ), 
        .B2(n8447), .ZN(n8445) );
  INV_X1 U9856 ( .A(n8445), .ZN(n9393) );
  OAI22_X1 U9857 ( .A1(n8448), .A2(s_data_in_f[1]), .B1(\fmem_data[27][1] ), 
        .B2(n8447), .ZN(n8446) );
  INV_X1 U9858 ( .A(n8446), .ZN(n9394) );
  OAI22_X1 U9859 ( .A1(n8448), .A2(s_data_in_f[0]), .B1(\fmem_data[27][0] ), 
        .B2(n8447), .ZN(n8449) );
  INV_X1 U9860 ( .A(n8449), .ZN(n9395) );
  NAND3_X1 U9861 ( .A1(fmem_addr[1]), .A2(n8710), .A3(n8709), .ZN(n8632) );
  OAI22_X1 U9862 ( .A1(n8458), .A2(s_data_in_f[7]), .B1(\fmem_data[26][7] ), 
        .B2(n8457), .ZN(n8450) );
  INV_X1 U9863 ( .A(n8450), .ZN(n9396) );
  OAI22_X1 U9864 ( .A1(n8458), .A2(s_data_in_f[6]), .B1(\fmem_data[26][6] ), 
        .B2(n8457), .ZN(n8451) );
  INV_X1 U9865 ( .A(n8451), .ZN(n9397) );
  OAI22_X1 U9866 ( .A1(n8458), .A2(s_data_in_f[5]), .B1(\fmem_data[26][5] ), 
        .B2(n8457), .ZN(n8452) );
  INV_X1 U9867 ( .A(n8452), .ZN(n9398) );
  OAI22_X1 U9868 ( .A1(n8458), .A2(s_data_in_f[4]), .B1(\fmem_data[26][4] ), 
        .B2(n8457), .ZN(n8453) );
  INV_X1 U9869 ( .A(n8453), .ZN(n9399) );
  OAI22_X1 U9870 ( .A1(n8458), .A2(s_data_in_f[3]), .B1(\fmem_data[26][3] ), 
        .B2(n8457), .ZN(n8454) );
  INV_X1 U9871 ( .A(n8454), .ZN(n9400) );
  OAI22_X1 U9872 ( .A1(n8458), .A2(s_data_in_f[2]), .B1(\fmem_data[26][2] ), 
        .B2(n8457), .ZN(n8455) );
  INV_X1 U9873 ( .A(n8455), .ZN(n9401) );
  OAI22_X1 U9874 ( .A1(n8458), .A2(s_data_in_f[1]), .B1(\fmem_data[26][1] ), 
        .B2(n8457), .ZN(n8456) );
  INV_X1 U9875 ( .A(n8456), .ZN(n9402) );
  OAI22_X1 U9876 ( .A1(n8458), .A2(s_data_in_f[0]), .B1(\fmem_data[26][0] ), 
        .B2(n8457), .ZN(n8459) );
  INV_X1 U9877 ( .A(n8459), .ZN(n9403) );
  NAND3_X1 U9878 ( .A1(fmem_addr[0]), .A2(n8711), .A3(n8709), .ZN(n8643) );
  OAI22_X1 U9879 ( .A1(n8468), .A2(s_data_in_f[7]), .B1(\fmem_data[25][7] ), 
        .B2(n8467), .ZN(n8460) );
  INV_X1 U9880 ( .A(n8460), .ZN(n9404) );
  OAI22_X1 U9881 ( .A1(n8468), .A2(s_data_in_f[6]), .B1(\fmem_data[25][6] ), 
        .B2(n8467), .ZN(n8461) );
  INV_X1 U9882 ( .A(n8461), .ZN(n9405) );
  OAI22_X1 U9883 ( .A1(n8468), .A2(s_data_in_f[5]), .B1(\fmem_data[25][5] ), 
        .B2(n8467), .ZN(n8462) );
  INV_X1 U9884 ( .A(n8462), .ZN(n9406) );
  OAI22_X1 U9885 ( .A1(n8468), .A2(s_data_in_f[4]), .B1(\fmem_data[25][4] ), 
        .B2(n8467), .ZN(n8463) );
  INV_X1 U9886 ( .A(n8463), .ZN(n9407) );
  OAI22_X1 U9887 ( .A1(n8468), .A2(s_data_in_f[3]), .B1(\fmem_data[25][3] ), 
        .B2(n8467), .ZN(n8464) );
  INV_X1 U9888 ( .A(n8464), .ZN(n9408) );
  OAI22_X1 U9889 ( .A1(n8468), .A2(s_data_in_f[2]), .B1(\fmem_data[25][2] ), 
        .B2(n8467), .ZN(n8465) );
  INV_X1 U9890 ( .A(n8465), .ZN(n9409) );
  OAI22_X1 U9891 ( .A1(n8468), .A2(s_data_in_f[1]), .B1(\fmem_data[25][1] ), 
        .B2(n8467), .ZN(n8466) );
  INV_X1 U9892 ( .A(n8466), .ZN(n9410) );
  OAI22_X1 U9893 ( .A1(n8468), .A2(s_data_in_f[0]), .B1(\fmem_data[25][0] ), 
        .B2(n8467), .ZN(n8469) );
  INV_X1 U9894 ( .A(n8469), .ZN(n9411) );
  NAND3_X1 U9895 ( .A1(n8710), .A2(n8711), .A3(n8709), .ZN(n8655) );
  OAI22_X1 U9896 ( .A1(n8479), .A2(s_data_in_f[7]), .B1(\fmem_data[24][7] ), 
        .B2(n8478), .ZN(n8471) );
  INV_X1 U9897 ( .A(n8471), .ZN(n9412) );
  OAI22_X1 U9898 ( .A1(n8479), .A2(s_data_in_f[6]), .B1(\fmem_data[24][6] ), 
        .B2(n8478), .ZN(n8472) );
  INV_X1 U9899 ( .A(n8472), .ZN(n9413) );
  OAI22_X1 U9900 ( .A1(n8479), .A2(s_data_in_f[5]), .B1(\fmem_data[24][5] ), 
        .B2(n8478), .ZN(n8473) );
  INV_X1 U9901 ( .A(n8473), .ZN(n9414) );
  OAI22_X1 U9902 ( .A1(n8479), .A2(s_data_in_f[4]), .B1(\fmem_data[24][4] ), 
        .B2(n8478), .ZN(n8474) );
  INV_X1 U9903 ( .A(n8474), .ZN(n9415) );
  OAI22_X1 U9904 ( .A1(n8479), .A2(s_data_in_f[3]), .B1(\fmem_data[24][3] ), 
        .B2(n8478), .ZN(n8475) );
  INV_X1 U9905 ( .A(n8475), .ZN(n9416) );
  OAI22_X1 U9906 ( .A1(n8479), .A2(s_data_in_f[2]), .B1(\fmem_data[24][2] ), 
        .B2(n8478), .ZN(n8476) );
  INV_X1 U9907 ( .A(n8476), .ZN(n9417) );
  OAI22_X1 U9908 ( .A1(n8479), .A2(s_data_in_f[1]), .B1(\fmem_data[24][1] ), 
        .B2(n8478), .ZN(n8477) );
  INV_X1 U9909 ( .A(n8477), .ZN(n9418) );
  OAI22_X1 U9910 ( .A1(n8479), .A2(s_data_in_f[0]), .B1(\fmem_data[24][0] ), 
        .B2(n8478), .ZN(n8480) );
  INV_X1 U9911 ( .A(n8480), .ZN(n9419) );
  OAI22_X1 U9912 ( .A1(n8490), .A2(s_data_in_f[7]), .B1(\fmem_data[23][7] ), 
        .B2(n8489), .ZN(n8482) );
  INV_X1 U9913 ( .A(n8482), .ZN(n9420) );
  OAI22_X1 U9914 ( .A1(n8490), .A2(s_data_in_f[6]), .B1(\fmem_data[23][6] ), 
        .B2(n8489), .ZN(n8483) );
  INV_X1 U9915 ( .A(n8483), .ZN(n9421) );
  OAI22_X1 U9916 ( .A1(n8490), .A2(s_data_in_f[5]), .B1(\fmem_data[23][5] ), 
        .B2(n8489), .ZN(n8484) );
  INV_X1 U9917 ( .A(n8484), .ZN(n9422) );
  OAI22_X1 U9918 ( .A1(n8490), .A2(s_data_in_f[4]), .B1(\fmem_data[23][4] ), 
        .B2(n8489), .ZN(n8485) );
  INV_X1 U9919 ( .A(n8485), .ZN(n9423) );
  OAI22_X1 U9920 ( .A1(n8490), .A2(s_data_in_f[3]), .B1(\fmem_data[23][3] ), 
        .B2(n8489), .ZN(n8486) );
  INV_X1 U9921 ( .A(n8486), .ZN(n9424) );
  OAI22_X1 U9922 ( .A1(n8490), .A2(s_data_in_f[2]), .B1(\fmem_data[23][2] ), 
        .B2(n8489), .ZN(n8487) );
  INV_X1 U9923 ( .A(n8487), .ZN(n9425) );
  OAI22_X1 U9924 ( .A1(n8490), .A2(s_data_in_f[1]), .B1(\fmem_data[23][1] ), 
        .B2(n8489), .ZN(n8488) );
  INV_X1 U9925 ( .A(n8488), .ZN(n9426) );
  OAI22_X1 U9926 ( .A1(n8490), .A2(s_data_in_f[0]), .B1(\fmem_data[23][0] ), 
        .B2(n8489), .ZN(n8491) );
  INV_X1 U9927 ( .A(n8491), .ZN(n9427) );
  OAI22_X1 U9928 ( .A1(n8500), .A2(s_data_in_f[7]), .B1(\fmem_data[22][7] ), 
        .B2(n8499), .ZN(n8492) );
  INV_X1 U9929 ( .A(n8492), .ZN(n9428) );
  OAI22_X1 U9930 ( .A1(n8500), .A2(s_data_in_f[6]), .B1(\fmem_data[22][6] ), 
        .B2(n8499), .ZN(n8493) );
  INV_X1 U9931 ( .A(n8493), .ZN(n9429) );
  OAI22_X1 U9932 ( .A1(n8500), .A2(s_data_in_f[5]), .B1(\fmem_data[22][5] ), 
        .B2(n8499), .ZN(n8494) );
  INV_X1 U9933 ( .A(n8494), .ZN(n9430) );
  OAI22_X1 U9934 ( .A1(n8500), .A2(s_data_in_f[4]), .B1(\fmem_data[22][4] ), 
        .B2(n8499), .ZN(n8495) );
  INV_X1 U9935 ( .A(n8495), .ZN(n9431) );
  OAI22_X1 U9936 ( .A1(n8500), .A2(s_data_in_f[3]), .B1(\fmem_data[22][3] ), 
        .B2(n8499), .ZN(n8496) );
  INV_X1 U9937 ( .A(n8496), .ZN(n9432) );
  OAI22_X1 U9938 ( .A1(n8500), .A2(s_data_in_f[2]), .B1(\fmem_data[22][2] ), 
        .B2(n8499), .ZN(n8497) );
  INV_X1 U9939 ( .A(n8497), .ZN(n9433) );
  OAI22_X1 U9940 ( .A1(n8500), .A2(s_data_in_f[1]), .B1(\fmem_data[22][1] ), 
        .B2(n8499), .ZN(n8498) );
  INV_X1 U9941 ( .A(n8498), .ZN(n9434) );
  OAI22_X1 U9942 ( .A1(n8500), .A2(s_data_in_f[0]), .B1(\fmem_data[22][0] ), 
        .B2(n8499), .ZN(n8501) );
  INV_X1 U9943 ( .A(n8501), .ZN(n9435) );
  OAI22_X1 U9944 ( .A1(n8510), .A2(s_data_in_f[7]), .B1(\fmem_data[21][7] ), 
        .B2(n8509), .ZN(n8502) );
  INV_X1 U9945 ( .A(n8502), .ZN(n9436) );
  OAI22_X1 U9946 ( .A1(n8510), .A2(s_data_in_f[6]), .B1(\fmem_data[21][6] ), 
        .B2(n8509), .ZN(n8503) );
  INV_X1 U9947 ( .A(n8503), .ZN(n9437) );
  OAI22_X1 U9948 ( .A1(n8510), .A2(s_data_in_f[5]), .B1(\fmem_data[21][5] ), 
        .B2(n8509), .ZN(n8504) );
  INV_X1 U9949 ( .A(n8504), .ZN(n9438) );
  OAI22_X1 U9950 ( .A1(n8510), .A2(s_data_in_f[4]), .B1(\fmem_data[21][4] ), 
        .B2(n8509), .ZN(n8505) );
  INV_X1 U9951 ( .A(n8505), .ZN(n9439) );
  OAI22_X1 U9952 ( .A1(n8510), .A2(s_data_in_f[3]), .B1(\fmem_data[21][3] ), 
        .B2(n8509), .ZN(n8506) );
  INV_X1 U9953 ( .A(n8506), .ZN(n9440) );
  OAI22_X1 U9954 ( .A1(n8510), .A2(s_data_in_f[2]), .B1(\fmem_data[21][2] ), 
        .B2(n8509), .ZN(n8507) );
  INV_X1 U9955 ( .A(n8507), .ZN(n9441) );
  OAI22_X1 U9956 ( .A1(n8510), .A2(s_data_in_f[1]), .B1(\fmem_data[21][1] ), 
        .B2(n8509), .ZN(n8508) );
  INV_X1 U9957 ( .A(n8508), .ZN(n9442) );
  OAI22_X1 U9958 ( .A1(n8510), .A2(s_data_in_f[0]), .B1(\fmem_data[21][0] ), 
        .B2(n8509), .ZN(n8511) );
  INV_X1 U9959 ( .A(n8511), .ZN(n9443) );
  OAI22_X1 U9960 ( .A1(n8520), .A2(s_data_in_f[7]), .B1(\fmem_data[20][7] ), 
        .B2(n8519), .ZN(n8512) );
  INV_X1 U9961 ( .A(n8512), .ZN(n9444) );
  OAI22_X1 U9962 ( .A1(n8520), .A2(s_data_in_f[6]), .B1(\fmem_data[20][6] ), 
        .B2(n8519), .ZN(n8513) );
  INV_X1 U9963 ( .A(n8513), .ZN(n9445) );
  OAI22_X1 U9964 ( .A1(n8520), .A2(s_data_in_f[5]), .B1(\fmem_data[20][5] ), 
        .B2(n8519), .ZN(n8514) );
  INV_X1 U9965 ( .A(n8514), .ZN(n9446) );
  OAI22_X1 U9966 ( .A1(n8520), .A2(s_data_in_f[4]), .B1(\fmem_data[20][4] ), 
        .B2(n8519), .ZN(n8515) );
  INV_X1 U9967 ( .A(n8515), .ZN(n9447) );
  OAI22_X1 U9968 ( .A1(n8520), .A2(s_data_in_f[3]), .B1(\fmem_data[20][3] ), 
        .B2(n8519), .ZN(n8516) );
  INV_X1 U9969 ( .A(n8516), .ZN(n9448) );
  OAI22_X1 U9970 ( .A1(n8520), .A2(s_data_in_f[2]), .B1(\fmem_data[20][2] ), 
        .B2(n8519), .ZN(n8517) );
  INV_X1 U9971 ( .A(n8517), .ZN(n9449) );
  OAI22_X1 U9972 ( .A1(n8520), .A2(s_data_in_f[1]), .B1(\fmem_data[20][1] ), 
        .B2(n8519), .ZN(n8518) );
  INV_X1 U9973 ( .A(n8518), .ZN(n9450) );
  OAI22_X1 U9974 ( .A1(n8520), .A2(s_data_in_f[0]), .B1(\fmem_data[20][0] ), 
        .B2(n8519), .ZN(n8521) );
  INV_X1 U9975 ( .A(n8521), .ZN(n9451) );
  OAI22_X1 U9976 ( .A1(n8530), .A2(s_data_in_f[7]), .B1(\fmem_data[19][7] ), 
        .B2(n8529), .ZN(n8522) );
  INV_X1 U9977 ( .A(n8522), .ZN(n9452) );
  OAI22_X1 U9978 ( .A1(n8530), .A2(s_data_in_f[6]), .B1(\fmem_data[19][6] ), 
        .B2(n8529), .ZN(n8523) );
  INV_X1 U9979 ( .A(n8523), .ZN(n9453) );
  OAI22_X1 U9980 ( .A1(n8530), .A2(s_data_in_f[5]), .B1(\fmem_data[19][5] ), 
        .B2(n8529), .ZN(n8524) );
  INV_X1 U9981 ( .A(n8524), .ZN(n9454) );
  OAI22_X1 U9982 ( .A1(n8530), .A2(s_data_in_f[4]), .B1(\fmem_data[19][4] ), 
        .B2(n8529), .ZN(n8525) );
  INV_X1 U9983 ( .A(n8525), .ZN(n9455) );
  OAI22_X1 U9984 ( .A1(n8530), .A2(s_data_in_f[3]), .B1(\fmem_data[19][3] ), 
        .B2(n8529), .ZN(n8526) );
  INV_X1 U9985 ( .A(n8526), .ZN(n9456) );
  OAI22_X1 U9986 ( .A1(n8530), .A2(s_data_in_f[2]), .B1(\fmem_data[19][2] ), 
        .B2(n8529), .ZN(n8527) );
  INV_X1 U9987 ( .A(n8527), .ZN(n9457) );
  OAI22_X1 U9988 ( .A1(n8530), .A2(s_data_in_f[1]), .B1(\fmem_data[19][1] ), 
        .B2(n8529), .ZN(n8528) );
  INV_X1 U9989 ( .A(n8528), .ZN(n9458) );
  OAI22_X1 U9990 ( .A1(n8530), .A2(s_data_in_f[0]), .B1(\fmem_data[19][0] ), 
        .B2(n8529), .ZN(n8531) );
  INV_X1 U9991 ( .A(n8531), .ZN(n9459) );
  OAI22_X1 U9992 ( .A1(n8540), .A2(s_data_in_f[7]), .B1(\fmem_data[18][7] ), 
        .B2(n8539), .ZN(n8532) );
  INV_X1 U9993 ( .A(n8532), .ZN(n9460) );
  OAI22_X1 U9994 ( .A1(n8540), .A2(s_data_in_f[6]), .B1(\fmem_data[18][6] ), 
        .B2(n8539), .ZN(n8533) );
  INV_X1 U9995 ( .A(n8533), .ZN(n9461) );
  OAI22_X1 U9996 ( .A1(n8540), .A2(s_data_in_f[5]), .B1(\fmem_data[18][5] ), 
        .B2(n8539), .ZN(n8534) );
  INV_X1 U9997 ( .A(n8534), .ZN(n9462) );
  OAI22_X1 U9998 ( .A1(n8540), .A2(s_data_in_f[4]), .B1(\fmem_data[18][4] ), 
        .B2(n8539), .ZN(n8535) );
  INV_X1 U9999 ( .A(n8535), .ZN(n9463) );
  OAI22_X1 U10000 ( .A1(n8540), .A2(s_data_in_f[3]), .B1(\fmem_data[18][3] ), 
        .B2(n8539), .ZN(n8536) );
  INV_X1 U10001 ( .A(n8536), .ZN(n9464) );
  OAI22_X1 U10002 ( .A1(n8540), .A2(s_data_in_f[2]), .B1(\fmem_data[18][2] ), 
        .B2(n8539), .ZN(n8537) );
  INV_X1 U10003 ( .A(n8537), .ZN(n9465) );
  OAI22_X1 U10004 ( .A1(n8540), .A2(s_data_in_f[1]), .B1(\fmem_data[18][1] ), 
        .B2(n8539), .ZN(n8538) );
  INV_X1 U10005 ( .A(n8538), .ZN(n9466) );
  OAI22_X1 U10006 ( .A1(n8540), .A2(s_data_in_f[0]), .B1(\fmem_data[18][0] ), 
        .B2(n8539), .ZN(n8541) );
  INV_X1 U10007 ( .A(n8541), .ZN(n9467) );
  OAI22_X1 U10008 ( .A1(n8550), .A2(s_data_in_f[7]), .B1(\fmem_data[17][7] ), 
        .B2(n8549), .ZN(n8542) );
  INV_X1 U10009 ( .A(n8542), .ZN(n9468) );
  OAI22_X1 U10010 ( .A1(n8550), .A2(s_data_in_f[6]), .B1(\fmem_data[17][6] ), 
        .B2(n8549), .ZN(n8543) );
  INV_X1 U10011 ( .A(n8543), .ZN(n9469) );
  OAI22_X1 U10012 ( .A1(n8550), .A2(s_data_in_f[5]), .B1(\fmem_data[17][5] ), 
        .B2(n8549), .ZN(n8544) );
  INV_X1 U10013 ( .A(n8544), .ZN(n9470) );
  OAI22_X1 U10014 ( .A1(n8550), .A2(s_data_in_f[4]), .B1(\fmem_data[17][4] ), 
        .B2(n8549), .ZN(n8545) );
  INV_X1 U10015 ( .A(n8545), .ZN(n9471) );
  OAI22_X1 U10016 ( .A1(n8550), .A2(s_data_in_f[3]), .B1(\fmem_data[17][3] ), 
        .B2(n8549), .ZN(n8546) );
  INV_X1 U10017 ( .A(n8546), .ZN(n9472) );
  OAI22_X1 U10018 ( .A1(n8550), .A2(s_data_in_f[2]), .B1(\fmem_data[17][2] ), 
        .B2(n8549), .ZN(n8547) );
  INV_X1 U10019 ( .A(n8547), .ZN(n9473) );
  OAI22_X1 U10020 ( .A1(n8550), .A2(s_data_in_f[1]), .B1(\fmem_data[17][1] ), 
        .B2(n8549), .ZN(n8548) );
  INV_X1 U10021 ( .A(n8548), .ZN(n9474) );
  OAI22_X1 U10022 ( .A1(n8550), .A2(s_data_in_f[0]), .B1(\fmem_data[17][0] ), 
        .B2(n8549), .ZN(n8551) );
  INV_X1 U10023 ( .A(n8551), .ZN(n9475) );
  OAI22_X1 U10024 ( .A1(n8561), .A2(s_data_in_f[7]), .B1(\fmem_data[16][7] ), 
        .B2(n8560), .ZN(n8553) );
  INV_X1 U10025 ( .A(n8553), .ZN(n9476) );
  OAI22_X1 U10026 ( .A1(n8561), .A2(s_data_in_f[6]), .B1(\fmem_data[16][6] ), 
        .B2(n8560), .ZN(n8554) );
  INV_X1 U10027 ( .A(n8554), .ZN(n9477) );
  OAI22_X1 U10028 ( .A1(n8561), .A2(s_data_in_f[5]), .B1(\fmem_data[16][5] ), 
        .B2(n8560), .ZN(n8555) );
  INV_X1 U10029 ( .A(n8555), .ZN(n9478) );
  OAI22_X1 U10030 ( .A1(n8561), .A2(s_data_in_f[4]), .B1(\fmem_data[16][4] ), 
        .B2(n8560), .ZN(n8556) );
  INV_X1 U10031 ( .A(n8556), .ZN(n9479) );
  OAI22_X1 U10032 ( .A1(n8561), .A2(s_data_in_f[3]), .B1(\fmem_data[16][3] ), 
        .B2(n8560), .ZN(n8557) );
  INV_X1 U10033 ( .A(n8557), .ZN(n9480) );
  OAI22_X1 U10034 ( .A1(n8561), .A2(s_data_in_f[2]), .B1(\fmem_data[16][2] ), 
        .B2(n8560), .ZN(n8558) );
  INV_X1 U10035 ( .A(n8558), .ZN(n9481) );
  OAI22_X1 U10036 ( .A1(n8561), .A2(s_data_in_f[1]), .B1(\fmem_data[16][1] ), 
        .B2(n8560), .ZN(n8559) );
  INV_X1 U10037 ( .A(n8559), .ZN(n9482) );
  OAI22_X1 U10038 ( .A1(n8561), .A2(s_data_in_f[0]), .B1(\fmem_data[16][0] ), 
        .B2(n8560), .ZN(n8562) );
  INV_X1 U10039 ( .A(n8562), .ZN(n9483) );
  OAI22_X1 U10040 ( .A1(n8678), .A2(s_data_in_f[7]), .B1(\fmem_data[15][7] ), 
        .B2(n8563), .ZN(n8846) );
  OAI22_X1 U10041 ( .A1(n8678), .A2(s_data_in_f[6]), .B1(\fmem_data[15][6] ), 
        .B2(n8563), .ZN(n8847) );
  OAI22_X1 U10042 ( .A1(n8678), .A2(s_data_in_f[5]), .B1(\fmem_data[15][5] ), 
        .B2(n8563), .ZN(n8848) );
  OAI22_X1 U10043 ( .A1(n8678), .A2(s_data_in_f[4]), .B1(\fmem_data[15][4] ), 
        .B2(n8563), .ZN(n8849) );
  OAI22_X1 U10044 ( .A1(n8678), .A2(s_data_in_f[3]), .B1(\fmem_data[15][3] ), 
        .B2(n8563), .ZN(n8850) );
  OAI22_X1 U10045 ( .A1(n8678), .A2(s_data_in_f[2]), .B1(\fmem_data[15][2] ), 
        .B2(n8563), .ZN(n8851) );
  OAI22_X1 U10046 ( .A1(n8678), .A2(s_data_in_f[1]), .B1(\fmem_data[15][1] ), 
        .B2(n8563), .ZN(n8852) );
  OAI22_X1 U10047 ( .A1(n8678), .A2(s_data_in_f[0]), .B1(\fmem_data[15][0] ), 
        .B2(n8563), .ZN(n8853) );
  OAI22_X1 U10048 ( .A1(n8565), .A2(s_data_in_f[7]), .B1(\fmem_data[14][7] ), 
        .B2(n8564), .ZN(n8854) );
  OAI22_X1 U10049 ( .A1(n8565), .A2(s_data_in_f[6]), .B1(\fmem_data[14][6] ), 
        .B2(n8564), .ZN(n8855) );
  OAI22_X1 U10050 ( .A1(n8565), .A2(s_data_in_f[5]), .B1(\fmem_data[14][5] ), 
        .B2(n8564), .ZN(n8856) );
  OAI22_X1 U10051 ( .A1(n8565), .A2(s_data_in_f[4]), .B1(\fmem_data[14][4] ), 
        .B2(n8564), .ZN(n8857) );
  OAI22_X1 U10052 ( .A1(n8565), .A2(s_data_in_f[3]), .B1(\fmem_data[14][3] ), 
        .B2(n8564), .ZN(n8858) );
  OAI22_X1 U10053 ( .A1(n8565), .A2(s_data_in_f[2]), .B1(\fmem_data[14][2] ), 
        .B2(n8564), .ZN(n8859) );
  OAI22_X1 U10054 ( .A1(n8565), .A2(s_data_in_f[1]), .B1(\fmem_data[14][1] ), 
        .B2(n8564), .ZN(n8860) );
  OAI22_X1 U10055 ( .A1(n8565), .A2(s_data_in_f[0]), .B1(\fmem_data[14][0] ), 
        .B2(n8564), .ZN(n8861) );
  OAI22_X1 U10056 ( .A1(n8567), .A2(s_data_in_f[7]), .B1(\fmem_data[13][7] ), 
        .B2(n8566), .ZN(n8862) );
  OAI22_X1 U10057 ( .A1(n8567), .A2(s_data_in_f[6]), .B1(\fmem_data[13][6] ), 
        .B2(n8566), .ZN(n8863) );
  OAI22_X1 U10058 ( .A1(n8567), .A2(s_data_in_f[5]), .B1(\fmem_data[13][5] ), 
        .B2(n8566), .ZN(n8864) );
  OAI22_X1 U10059 ( .A1(n8567), .A2(s_data_in_f[4]), .B1(\fmem_data[13][4] ), 
        .B2(n8566), .ZN(n8865) );
  OAI22_X1 U10060 ( .A1(n8567), .A2(s_data_in_f[3]), .B1(\fmem_data[13][3] ), 
        .B2(n8566), .ZN(n8866) );
  OAI22_X1 U10061 ( .A1(n8567), .A2(s_data_in_f[2]), .B1(\fmem_data[13][2] ), 
        .B2(n8566), .ZN(n8867) );
  OAI22_X1 U10062 ( .A1(n8567), .A2(s_data_in_f[1]), .B1(\fmem_data[13][1] ), 
        .B2(n8566), .ZN(n8868) );
  OAI22_X1 U10063 ( .A1(n8567), .A2(s_data_in_f[0]), .B1(\fmem_data[13][0] ), 
        .B2(n8566), .ZN(n8869) );
  OAI22_X1 U10064 ( .A1(n8569), .A2(s_data_in_f[7]), .B1(\fmem_data[12][7] ), 
        .B2(n8568), .ZN(n8870) );
  OAI22_X1 U10065 ( .A1(n8569), .A2(s_data_in_f[6]), .B1(\fmem_data[12][6] ), 
        .B2(n8568), .ZN(n8871) );
  OAI22_X1 U10066 ( .A1(n8569), .A2(s_data_in_f[5]), .B1(\fmem_data[12][5] ), 
        .B2(n8568), .ZN(n8872) );
  OAI22_X1 U10067 ( .A1(n8569), .A2(s_data_in_f[4]), .B1(\fmem_data[12][4] ), 
        .B2(n8568), .ZN(n8873) );
  OAI22_X1 U10068 ( .A1(n8569), .A2(s_data_in_f[3]), .B1(\fmem_data[12][3] ), 
        .B2(n8568), .ZN(n8874) );
  OAI22_X1 U10069 ( .A1(n8569), .A2(s_data_in_f[2]), .B1(\fmem_data[12][2] ), 
        .B2(n8568), .ZN(n8875) );
  OAI22_X1 U10070 ( .A1(n8569), .A2(s_data_in_f[1]), .B1(\fmem_data[12][1] ), 
        .B2(n8568), .ZN(n8876) );
  OAI22_X1 U10071 ( .A1(n8569), .A2(s_data_in_f[0]), .B1(\fmem_data[12][0] ), 
        .B2(n8568), .ZN(n8877) );
  OAI22_X1 U10072 ( .A1(n8571), .A2(s_data_in_f[7]), .B1(\fmem_data[11][7] ), 
        .B2(n8570), .ZN(n8878) );
  OAI22_X1 U10073 ( .A1(n8571), .A2(s_data_in_f[6]), .B1(\fmem_data[11][6] ), 
        .B2(n8570), .ZN(n8879) );
  OAI22_X1 U10074 ( .A1(n8571), .A2(s_data_in_f[5]), .B1(\fmem_data[11][5] ), 
        .B2(n8570), .ZN(n8880) );
  OAI22_X1 U10075 ( .A1(n8571), .A2(s_data_in_f[4]), .B1(\fmem_data[11][4] ), 
        .B2(n8570), .ZN(n8881) );
  OAI22_X1 U10076 ( .A1(n8571), .A2(s_data_in_f[3]), .B1(\fmem_data[11][3] ), 
        .B2(n8570), .ZN(n8882) );
  OAI22_X1 U10077 ( .A1(n8571), .A2(s_data_in_f[2]), .B1(\fmem_data[11][2] ), 
        .B2(n8570), .ZN(n8883) );
  OAI22_X1 U10078 ( .A1(n8571), .A2(s_data_in_f[1]), .B1(\fmem_data[11][1] ), 
        .B2(n8570), .ZN(n8884) );
  OAI22_X1 U10079 ( .A1(n8571), .A2(s_data_in_f[0]), .B1(\fmem_data[11][0] ), 
        .B2(n8570), .ZN(n8885) );
  OAI22_X1 U10080 ( .A1(n8573), .A2(s_data_in_f[7]), .B1(\fmem_data[10][7] ), 
        .B2(n8572), .ZN(n8886) );
  OAI22_X1 U10081 ( .A1(n8573), .A2(s_data_in_f[6]), .B1(\fmem_data[10][6] ), 
        .B2(n8572), .ZN(n8887) );
  OAI22_X1 U10082 ( .A1(n8573), .A2(s_data_in_f[5]), .B1(\fmem_data[10][5] ), 
        .B2(n8572), .ZN(n8888) );
  OAI22_X1 U10083 ( .A1(n8573), .A2(s_data_in_f[4]), .B1(\fmem_data[10][4] ), 
        .B2(n8572), .ZN(n8889) );
  OAI22_X1 U10084 ( .A1(n8573), .A2(s_data_in_f[3]), .B1(\fmem_data[10][3] ), 
        .B2(n8572), .ZN(n8890) );
  OAI22_X1 U10085 ( .A1(n8573), .A2(s_data_in_f[2]), .B1(\fmem_data[10][2] ), 
        .B2(n8572), .ZN(n8891) );
  OAI22_X1 U10086 ( .A1(n8573), .A2(s_data_in_f[1]), .B1(\fmem_data[10][1] ), 
        .B2(n8572), .ZN(n8892) );
  OAI22_X1 U10087 ( .A1(n8573), .A2(s_data_in_f[0]), .B1(\fmem_data[10][0] ), 
        .B2(n8572), .ZN(n8893) );
  OAI22_X1 U10088 ( .A1(n8575), .A2(s_data_in_f[7]), .B1(\fmem_data[9][7] ), 
        .B2(n8574), .ZN(n8894) );
  OAI22_X1 U10089 ( .A1(n8575), .A2(s_data_in_f[6]), .B1(\fmem_data[9][6] ), 
        .B2(n8574), .ZN(n8895) );
  OAI22_X1 U10090 ( .A1(n8575), .A2(s_data_in_f[5]), .B1(\fmem_data[9][5] ), 
        .B2(n8574), .ZN(n8896) );
  OAI22_X1 U10091 ( .A1(n8575), .A2(s_data_in_f[4]), .B1(\fmem_data[9][4] ), 
        .B2(n8574), .ZN(n8897) );
  OAI22_X1 U10092 ( .A1(n8575), .A2(s_data_in_f[3]), .B1(\fmem_data[9][3] ), 
        .B2(n8574), .ZN(n8898) );
  OAI22_X1 U10093 ( .A1(n8575), .A2(s_data_in_f[2]), .B1(\fmem_data[9][2] ), 
        .B2(n8574), .ZN(n8899) );
  OAI22_X1 U10094 ( .A1(n8575), .A2(s_data_in_f[1]), .B1(\fmem_data[9][1] ), 
        .B2(n8574), .ZN(n8900) );
  OAI22_X1 U10095 ( .A1(n8575), .A2(s_data_in_f[0]), .B1(\fmem_data[9][0] ), 
        .B2(n8574), .ZN(n8901) );
  OAI22_X1 U10096 ( .A1(n8578), .A2(s_data_in_f[7]), .B1(\fmem_data[8][7] ), 
        .B2(n8577), .ZN(n8902) );
  OAI22_X1 U10097 ( .A1(n8578), .A2(s_data_in_f[6]), .B1(\fmem_data[8][6] ), 
        .B2(n8577), .ZN(n8903) );
  OAI22_X1 U10098 ( .A1(n8578), .A2(s_data_in_f[5]), .B1(\fmem_data[8][5] ), 
        .B2(n8577), .ZN(n8904) );
  OAI22_X1 U10099 ( .A1(n8578), .A2(s_data_in_f[4]), .B1(\fmem_data[8][4] ), 
        .B2(n8577), .ZN(n8905) );
  OAI22_X1 U10100 ( .A1(n8578), .A2(s_data_in_f[3]), .B1(\fmem_data[8][3] ), 
        .B2(n8577), .ZN(n8906) );
  OAI22_X1 U10101 ( .A1(n8578), .A2(s_data_in_f[2]), .B1(\fmem_data[8][2] ), 
        .B2(n8577), .ZN(n8907) );
  OAI22_X1 U10102 ( .A1(n8578), .A2(s_data_in_f[1]), .B1(\fmem_data[8][1] ), 
        .B2(n8577), .ZN(n8908) );
  OAI22_X1 U10103 ( .A1(n8578), .A2(s_data_in_f[0]), .B1(\fmem_data[8][0] ), 
        .B2(n8577), .ZN(n8909) );
  OAI22_X1 U10104 ( .A1(n8588), .A2(s_data_in_f[7]), .B1(\fmem_data[7][7] ), 
        .B2(n8587), .ZN(n8580) );
  INV_X1 U10105 ( .A(n8580), .ZN(n9484) );
  OAI22_X1 U10106 ( .A1(n8588), .A2(s_data_in_f[6]), .B1(\fmem_data[7][6] ), 
        .B2(n8587), .ZN(n8581) );
  INV_X1 U10107 ( .A(n8581), .ZN(n9485) );
  OAI22_X1 U10108 ( .A1(n8588), .A2(s_data_in_f[5]), .B1(\fmem_data[7][5] ), 
        .B2(n8587), .ZN(n8582) );
  INV_X1 U10109 ( .A(n8582), .ZN(n9486) );
  OAI22_X1 U10110 ( .A1(n8588), .A2(s_data_in_f[4]), .B1(\fmem_data[7][4] ), 
        .B2(n8587), .ZN(n8583) );
  INV_X1 U10111 ( .A(n8583), .ZN(n9487) );
  OAI22_X1 U10112 ( .A1(n8588), .A2(s_data_in_f[3]), .B1(\fmem_data[7][3] ), 
        .B2(n8587), .ZN(n8584) );
  INV_X1 U10113 ( .A(n8584), .ZN(n9488) );
  OAI22_X1 U10114 ( .A1(n8588), .A2(s_data_in_f[2]), .B1(\fmem_data[7][2] ), 
        .B2(n8587), .ZN(n8585) );
  INV_X1 U10115 ( .A(n8585), .ZN(n9489) );
  OAI22_X1 U10116 ( .A1(n8588), .A2(s_data_in_f[1]), .B1(\fmem_data[7][1] ), 
        .B2(n8587), .ZN(n8586) );
  INV_X1 U10117 ( .A(n8586), .ZN(n9490) );
  OAI22_X1 U10118 ( .A1(n8588), .A2(s_data_in_f[0]), .B1(\fmem_data[7][0] ), 
        .B2(n8587), .ZN(n8589) );
  INV_X1 U10119 ( .A(n8589), .ZN(n9491) );
  OAI22_X1 U10120 ( .A1(n8599), .A2(s_data_in_f[7]), .B1(\fmem_data[6][7] ), 
        .B2(n8598), .ZN(n8591) );
  INV_X1 U10121 ( .A(n8591), .ZN(n9492) );
  OAI22_X1 U10122 ( .A1(n8599), .A2(s_data_in_f[6]), .B1(\fmem_data[6][6] ), 
        .B2(n8598), .ZN(n8592) );
  INV_X1 U10123 ( .A(n8592), .ZN(n9493) );
  OAI22_X1 U10124 ( .A1(n8599), .A2(s_data_in_f[5]), .B1(\fmem_data[6][5] ), 
        .B2(n8598), .ZN(n8593) );
  INV_X1 U10125 ( .A(n8593), .ZN(n9494) );
  OAI22_X1 U10126 ( .A1(n8599), .A2(s_data_in_f[4]), .B1(\fmem_data[6][4] ), 
        .B2(n8598), .ZN(n8594) );
  INV_X1 U10127 ( .A(n8594), .ZN(n9495) );
  OAI22_X1 U10128 ( .A1(n8599), .A2(s_data_in_f[3]), .B1(\fmem_data[6][3] ), 
        .B2(n8598), .ZN(n8595) );
  INV_X1 U10129 ( .A(n8595), .ZN(n9496) );
  OAI22_X1 U10130 ( .A1(n8599), .A2(s_data_in_f[2]), .B1(\fmem_data[6][2] ), 
        .B2(n8598), .ZN(n8596) );
  INV_X1 U10131 ( .A(n8596), .ZN(n9497) );
  OAI22_X1 U10132 ( .A1(n8599), .A2(s_data_in_f[1]), .B1(\fmem_data[6][1] ), 
        .B2(n8598), .ZN(n8597) );
  INV_X1 U10133 ( .A(n8597), .ZN(n9498) );
  OAI22_X1 U10134 ( .A1(n8599), .A2(s_data_in_f[0]), .B1(\fmem_data[6][0] ), 
        .B2(n8598), .ZN(n8600) );
  INV_X1 U10135 ( .A(n8600), .ZN(n9499) );
  OAI22_X1 U10136 ( .A1(n8610), .A2(s_data_in_f[7]), .B1(\fmem_data[5][7] ), 
        .B2(n8609), .ZN(n8602) );
  INV_X1 U10137 ( .A(n8602), .ZN(n9500) );
  OAI22_X1 U10138 ( .A1(n8610), .A2(s_data_in_f[6]), .B1(\fmem_data[5][6] ), 
        .B2(n8609), .ZN(n8603) );
  INV_X1 U10139 ( .A(n8603), .ZN(n9501) );
  OAI22_X1 U10140 ( .A1(n8610), .A2(s_data_in_f[5]), .B1(\fmem_data[5][5] ), 
        .B2(n8609), .ZN(n8604) );
  INV_X1 U10141 ( .A(n8604), .ZN(n9502) );
  OAI22_X1 U10142 ( .A1(n8610), .A2(s_data_in_f[4]), .B1(\fmem_data[5][4] ), 
        .B2(n8609), .ZN(n8605) );
  INV_X1 U10143 ( .A(n8605), .ZN(n9503) );
  OAI22_X1 U10144 ( .A1(n8610), .A2(s_data_in_f[3]), .B1(\fmem_data[5][3] ), 
        .B2(n8609), .ZN(n8606) );
  INV_X1 U10145 ( .A(n8606), .ZN(n9504) );
  OAI22_X1 U10146 ( .A1(n8610), .A2(s_data_in_f[2]), .B1(\fmem_data[5][2] ), 
        .B2(n8609), .ZN(n8607) );
  INV_X1 U10147 ( .A(n8607), .ZN(n9505) );
  OAI22_X1 U10148 ( .A1(n8610), .A2(s_data_in_f[1]), .B1(\fmem_data[5][1] ), 
        .B2(n8609), .ZN(n8608) );
  INV_X1 U10149 ( .A(n8608), .ZN(n9506) );
  OAI22_X1 U10150 ( .A1(n8610), .A2(s_data_in_f[0]), .B1(\fmem_data[5][0] ), 
        .B2(n8609), .ZN(n8611) );
  INV_X1 U10151 ( .A(n8611), .ZN(n9507) );
  OAI22_X1 U10152 ( .A1(n8620), .A2(s_data_in_f[7]), .B1(\fmem_data[4][7] ), 
        .B2(n8619), .ZN(n8910) );
  OAI22_X1 U10153 ( .A1(n8620), .A2(s_data_in_f[6]), .B1(\fmem_data[4][6] ), 
        .B2(n8619), .ZN(n8613) );
  INV_X1 U10154 ( .A(n8613), .ZN(n9508) );
  OAI22_X1 U10155 ( .A1(n8620), .A2(s_data_in_f[5]), .B1(\fmem_data[4][5] ), 
        .B2(n8619), .ZN(n8614) );
  INV_X1 U10156 ( .A(n8614), .ZN(n9509) );
  OAI22_X1 U10157 ( .A1(n8620), .A2(s_data_in_f[4]), .B1(\fmem_data[4][4] ), 
        .B2(n8619), .ZN(n8615) );
  INV_X1 U10158 ( .A(n8615), .ZN(n9510) );
  OAI22_X1 U10159 ( .A1(n8620), .A2(s_data_in_f[3]), .B1(\fmem_data[4][3] ), 
        .B2(n8619), .ZN(n8616) );
  INV_X1 U10160 ( .A(n8616), .ZN(n9511) );
  OAI22_X1 U10161 ( .A1(n8620), .A2(s_data_in_f[2]), .B1(\fmem_data[4][2] ), 
        .B2(n8619), .ZN(n8617) );
  INV_X1 U10162 ( .A(n8617), .ZN(n9512) );
  OAI22_X1 U10163 ( .A1(n8620), .A2(s_data_in_f[1]), .B1(\fmem_data[4][1] ), 
        .B2(n8619), .ZN(n8618) );
  INV_X1 U10164 ( .A(n8618), .ZN(n9513) );
  OAI22_X1 U10165 ( .A1(n8620), .A2(s_data_in_f[0]), .B1(\fmem_data[4][0] ), 
        .B2(n8619), .ZN(n8621) );
  INV_X1 U10166 ( .A(n8621), .ZN(n9514) );
  OAI22_X1 U10167 ( .A1(n8630), .A2(s_data_in_f[7]), .B1(\fmem_data[3][7] ), 
        .B2(n8629), .ZN(n8622) );
  INV_X1 U10168 ( .A(n8622), .ZN(n9515) );
  OAI22_X1 U10169 ( .A1(n8630), .A2(s_data_in_f[6]), .B1(\fmem_data[3][6] ), 
        .B2(n8629), .ZN(n8623) );
  INV_X1 U10170 ( .A(n8623), .ZN(n9516) );
  OAI22_X1 U10171 ( .A1(n8630), .A2(s_data_in_f[5]), .B1(\fmem_data[3][5] ), 
        .B2(n8629), .ZN(n8624) );
  INV_X1 U10172 ( .A(n8624), .ZN(n9517) );
  OAI22_X1 U10173 ( .A1(n8630), .A2(s_data_in_f[4]), .B1(\fmem_data[3][4] ), 
        .B2(n8629), .ZN(n8625) );
  INV_X1 U10174 ( .A(n8625), .ZN(n9518) );
  OAI22_X1 U10175 ( .A1(n8630), .A2(s_data_in_f[3]), .B1(\fmem_data[3][3] ), 
        .B2(n8629), .ZN(n8626) );
  INV_X1 U10176 ( .A(n8626), .ZN(n9519) );
  OAI22_X1 U10177 ( .A1(n8630), .A2(s_data_in_f[2]), .B1(\fmem_data[3][2] ), 
        .B2(n8629), .ZN(n8627) );
  INV_X1 U10178 ( .A(n8627), .ZN(n9520) );
  OAI22_X1 U10179 ( .A1(n8630), .A2(s_data_in_f[1]), .B1(\fmem_data[3][1] ), 
        .B2(n8629), .ZN(n8628) );
  INV_X1 U10180 ( .A(n8628), .ZN(n9521) );
  OAI22_X1 U10181 ( .A1(n8630), .A2(s_data_in_f[0]), .B1(\fmem_data[3][0] ), 
        .B2(n8629), .ZN(n8631) );
  INV_X1 U10182 ( .A(n8631), .ZN(n9522) );
  OAI22_X1 U10183 ( .A1(n8641), .A2(s_data_in_f[7]), .B1(\fmem_data[2][7] ), 
        .B2(n8640), .ZN(n8633) );
  INV_X1 U10184 ( .A(n8633), .ZN(n9523) );
  OAI22_X1 U10185 ( .A1(n8641), .A2(s_data_in_f[6]), .B1(\fmem_data[2][6] ), 
        .B2(n8640), .ZN(n8634) );
  INV_X1 U10186 ( .A(n8634), .ZN(n9524) );
  OAI22_X1 U10187 ( .A1(n8641), .A2(s_data_in_f[5]), .B1(\fmem_data[2][5] ), 
        .B2(n8640), .ZN(n8635) );
  INV_X1 U10188 ( .A(n8635), .ZN(n9525) );
  OAI22_X1 U10189 ( .A1(n8641), .A2(s_data_in_f[4]), .B1(\fmem_data[2][4] ), 
        .B2(n8640), .ZN(n8636) );
  INV_X1 U10190 ( .A(n8636), .ZN(n9526) );
  OAI22_X1 U10191 ( .A1(n8641), .A2(s_data_in_f[3]), .B1(\fmem_data[2][3] ), 
        .B2(n8640), .ZN(n8637) );
  INV_X1 U10192 ( .A(n8637), .ZN(n9527) );
  OAI22_X1 U10193 ( .A1(n8641), .A2(s_data_in_f[2]), .B1(\fmem_data[2][2] ), 
        .B2(n8640), .ZN(n8638) );
  INV_X1 U10194 ( .A(n8638), .ZN(n9528) );
  OAI22_X1 U10195 ( .A1(n8641), .A2(s_data_in_f[1]), .B1(\fmem_data[2][1] ), 
        .B2(n8640), .ZN(n8639) );
  INV_X1 U10196 ( .A(n8639), .ZN(n9529) );
  OAI22_X1 U10197 ( .A1(n8641), .A2(s_data_in_f[0]), .B1(\fmem_data[2][0] ), 
        .B2(n8640), .ZN(n8642) );
  INV_X1 U10198 ( .A(n8642), .ZN(n9530) );
  OAI22_X1 U10199 ( .A1(n8652), .A2(s_data_in_f[7]), .B1(\fmem_data[1][7] ), 
        .B2(n8651), .ZN(n8644) );
  INV_X1 U10200 ( .A(n8644), .ZN(n9531) );
  OAI22_X1 U10201 ( .A1(n8652), .A2(s_data_in_f[6]), .B1(\fmem_data[1][6] ), 
        .B2(n8651), .ZN(n8645) );
  INV_X1 U10202 ( .A(n8645), .ZN(n9532) );
  OAI22_X1 U10203 ( .A1(n8652), .A2(s_data_in_f[5]), .B1(\fmem_data[1][5] ), 
        .B2(n8651), .ZN(n8646) );
  INV_X1 U10204 ( .A(n8646), .ZN(n9533) );
  OAI22_X1 U10205 ( .A1(n8652), .A2(s_data_in_f[4]), .B1(\fmem_data[1][4] ), 
        .B2(n8651), .ZN(n8647) );
  INV_X1 U10206 ( .A(n8647), .ZN(n9534) );
  OAI22_X1 U10207 ( .A1(n8652), .A2(s_data_in_f[3]), .B1(\fmem_data[1][3] ), 
        .B2(n8651), .ZN(n8648) );
  INV_X1 U10208 ( .A(n8648), .ZN(n9535) );
  OAI22_X1 U10209 ( .A1(n8652), .A2(s_data_in_f[2]), .B1(\fmem_data[1][2] ), 
        .B2(n8651), .ZN(n8649) );
  INV_X1 U10210 ( .A(n8649), .ZN(n9536) );
  OAI22_X1 U10211 ( .A1(n8652), .A2(s_data_in_f[1]), .B1(\fmem_data[1][1] ), 
        .B2(n8651), .ZN(n8650) );
  INV_X1 U10212 ( .A(n8650), .ZN(n9537) );
  OAI22_X1 U10213 ( .A1(n8652), .A2(s_data_in_f[0]), .B1(\fmem_data[1][0] ), 
        .B2(n8651), .ZN(n8653) );
  INV_X1 U10214 ( .A(n8653), .ZN(n9538) );
  OAI22_X1 U10215 ( .A1(n8664), .A2(s_data_in_f[7]), .B1(\fmem_data[0][7] ), 
        .B2(n8663), .ZN(n8656) );
  INV_X1 U10216 ( .A(n8656), .ZN(n9539) );
  OAI22_X1 U10217 ( .A1(n8664), .A2(s_data_in_f[6]), .B1(\fmem_data[0][6] ), 
        .B2(n8663), .ZN(n8657) );
  INV_X1 U10218 ( .A(n8657), .ZN(n9540) );
  OAI22_X1 U10219 ( .A1(n8664), .A2(s_data_in_f[5]), .B1(\fmem_data[0][5] ), 
        .B2(n8663), .ZN(n8658) );
  INV_X1 U10220 ( .A(n8658), .ZN(n9541) );
  OAI22_X1 U10221 ( .A1(n8664), .A2(s_data_in_f[4]), .B1(\fmem_data[0][4] ), 
        .B2(n8663), .ZN(n8659) );
  INV_X1 U10222 ( .A(n8659), .ZN(n9542) );
  OAI22_X1 U10223 ( .A1(n8664), .A2(s_data_in_f[3]), .B1(\fmem_data[0][3] ), 
        .B2(n8663), .ZN(n8660) );
  INV_X1 U10224 ( .A(n8660), .ZN(n9543) );
  OAI22_X1 U10225 ( .A1(n8664), .A2(s_data_in_f[2]), .B1(\fmem_data[0][2] ), 
        .B2(n8663), .ZN(n8661) );
  INV_X1 U10226 ( .A(n8661), .ZN(n9544) );
  OAI22_X1 U10227 ( .A1(n8664), .A2(s_data_in_f[1]), .B1(\fmem_data[0][1] ), 
        .B2(n8663), .ZN(n8662) );
  INV_X1 U10228 ( .A(n8662), .ZN(n9545) );
  OAI22_X1 U10229 ( .A1(n8664), .A2(s_data_in_f[0]), .B1(\fmem_data[0][0] ), 
        .B2(n8663), .ZN(n8665) );
  INV_X1 U10230 ( .A(n8665), .ZN(n9546) );
  NAND2_X1 U10231 ( .A1(\ctrl_inst/xmem_tracker [4]), .A2(n8688), .ZN(n8669)
         );
  NAND3_X1 U10232 ( .A1(\ctrl_inst/xmem_tracker [3]), .A2(
        \ctrl_inst/xmem_tracker [2]), .A3(n8674), .ZN(n8670) );
  AOI21_X1 U10233 ( .B1(n8669), .B2(n8670), .A(n8668), .ZN(n10318) );
  INV_X1 U10234 ( .A(n8670), .ZN(n8672) );
  AOI22_X1 U10235 ( .A1(\ctrl_inst/xmem_tracker [3]), .A2(n8688), .B1(
        \ctrl_inst/xmem_tracker [2]), .B2(n8674), .ZN(n8671) );
  NOR2_X1 U10236 ( .A1(n8672), .A2(n8671), .ZN(n10319) );
  AOI21_X1 U10237 ( .B1(n8688), .B2(\ctrl_inst/xmem_tracker [2]), .A(n8674), 
        .ZN(n8673) );
  AOI21_X1 U10238 ( .B1(n8674), .B2(\ctrl_inst/xmem_tracker [2]), .A(n8673), 
        .ZN(n10320) );
  NAND2_X1 U10239 ( .A1(n8688), .A2(n8675), .ZN(n8679) );
  AOI21_X1 U10240 ( .B1(n8746), .B2(n8678), .A(n8679), .ZN(n3397) );
  NAND2_X1 U10241 ( .A1(n8675), .A2(n3434), .ZN(n8686) );
  OAI22_X1 U10242 ( .A1(n8676), .A2(n8686), .B1(n8712), .B2(n8679), .ZN(n8677)
         );
  AND2_X1 U10243 ( .A1(n8678), .A2(n8677), .ZN(n3396) );
  OAI33_X1 U10244 ( .A1(n8681), .A2(n8710), .A3(n8680), .B1(n8682), .B2(n8679), 
        .B3(fmem_addr[0]), .ZN(n3395) );
  NAND2_X1 U10245 ( .A1(fmem_addr[0]), .A2(n8681), .ZN(n8684) );
  NAND2_X1 U10246 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n8683) );
  OAI21_X1 U10247 ( .B1(n8683), .B2(n8682), .A(n8688), .ZN(n8687) );
  AOI21_X1 U10248 ( .B1(n8711), .B2(n8684), .A(n8687), .ZN(n3394) );
  OAI22_X1 U10249 ( .A1(n8709), .A2(n8687), .B1(n8686), .B2(n8685), .ZN(n3393)
         );
  OAI21_X1 U10250 ( .B1(n8689), .B2(n8716), .A(n8688), .ZN(n3392) );
  OAI21_X1 U10251 ( .B1(n8691), .B2(n8713), .A(n8690), .ZN(n8692) );
  NAND2_X1 U10252 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  AOI22_X1 U10253 ( .A1(\ctrl_inst/pline_cntr [1]), .A2(n8695), .B1(n8694), 
        .B2(n8744), .ZN(n3120) );
endmodule

